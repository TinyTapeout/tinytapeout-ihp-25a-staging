module tt_um_dlmiles_tt08_poc_uart (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire clk_regs;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire rst_n_sync;
 wire sync_reset;
 wire \uart.resetCommandStrobe ;
 wire \uart.resetCommandUnit_1.async.area_io_q ;
 wire \uart.resetCommandUnit_1.async.area_io_r ;
 wire \uart.resetCommandUnit_1.ff ;
 wire \uart.resetCommandUnit_1.io_resetIn ;
 wire \uart.resetCommandUnit_1.reg1 ;
 wire \uart.uartArea_uart.busCtrl.io_regAddr[0] ;
 wire \uart.uartArea_uart.busCtrl.io_regAddr[1] ;
 wire \uart.uartArea_uart.busCtrl.io_regAddr[2] ;
 wire \uart.uartArea_uart.busCtrl.io_regAddr[3] ;
 wire \uart.uartArea_uart.busCtrl.io_regAddr[4] ;
 wire \uart.uartArea_uart.busCtrl.lastWasWrite ;
 wire \uart.uartArea_uart.busCtrl.oe ;
 wire \uart.uartArea_uart.commFilter.ctsFilter.io_b ;
 wire \uart.uartArea_uart.commFilter.ctsFilter.io_c ;
 wire \uart.uartArea_uart.commFilter.ctsFilter.io_o ;
 wire \uart.uartArea_uart.commFilter.dcdFilter.io_b ;
 wire \uart.uartArea_uart.commFilter.dcdFilter.io_c ;
 wire \uart.uartArea_uart.commFilter.dcdFilter.io_o ;
 wire \uart.uartArea_uart.commFilter.dsrFilter.io_b ;
 wire \uart.uartArea_uart.commFilter.dsrFilter.io_c ;
 wire \uart.uartArea_uart.commFilter.dsrFilter.io_o ;
 wire \uart.uartArea_uart.commFilter.io_ttl_ri ;
 wire \uart.uartArea_uart.commFilter.riFilter.io_b ;
 wire \uart.uartArea_uart.commFilter.riFilter.io_c ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptControl[0] ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptControl[1] ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptControl[2] ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptControl[3] ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptControl[4] ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptControl[5] ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptControl[6] ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptStatus[0] ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptStatus[1] ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptStatus[2] ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptStatus[3] ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptStatus[4] ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptStatus[5] ;
 wire \uart.uartArea_uart.regCtrl.io_regInterruptStatus[6] ;
 wire \uart.uartArea_uart.regCtrl.reg007[0] ;
 wire \uart.uartArea_uart.regCtrl.reg007[1] ;
 wire \uart.uartArea_uart.regCtrl.reg007[2] ;
 wire \uart.uartArea_uart.regCtrl.reg007[3] ;
 wire \uart.uartArea_uart.regCtrl.reg007[4] ;
 wire \uart.uartArea_uart.regCtrl.reg007[5] ;
 wire \uart.uartArea_uart.regCtrl.reg007[6] ;
 wire \uart.uartArea_uart.regCtrl.reg007[7] ;
 wire \uart.uartArea_uart.regCtrl.regFifoRxEnable ;
 wire \uart.uartArea_uart.regCtrl.regFifoTxEnable ;
 wire \uart.uartArea_uart.regCtrl.regModemCtrlChanged[0] ;
 wire \uart.uartArea_uart.regCtrl.regModemCtrlChanged[1] ;
 wire \uart.uartArea_uart.regCtrl.regModemCtrlChanged[2] ;
 wire \uart.uartArea_uart.regCtrl.regModemCtrlChanged[3] ;
 wire \uart.uartArea_uart.regCtrl.regModemCtrlHistory[0] ;
 wire \uart.uartArea_uart.regCtrl.regModemCtrlHistory[1] ;
 wire \uart.uartArea_uart.regCtrl.regModemCtrlHistory[3] ;
 wire \uart.uartArea_uart.regCtrl.riSignalNext ;
 wire \uart.uartArea_uart.regCtrl.txHolderBit9 ;
 wire \uart.uartArea_uart.regCtrl.txOverrun ;
 wire \uart.uartArea_uart.rxFifo.count[0] ;
 wire \uart.uartArea_uart.rxFifo.count[1] ;
 wire \uart.uartArea_uart.rxFifo.count[2] ;
 wire \uart.uartArea_uart.rxFifo.count[3] ;
 wire \uart.uartArea_uart.rxFifo.io_fifoRdAddr[0] ;
 wire \uart.uartArea_uart.rxFifo.io_fifoRdAddr[1] ;
 wire \uart.uartArea_uart.rxFifo.io_fifoRdAddr[2] ;
 wire \uart.uartArea_uart.rxFifo.io_fifoRdAddr[3] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_10[0] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_10[1] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_10[2] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_10[3] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_10[4] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_10[5] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_10[6] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_10[7] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_10[8] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_11[0] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_11[1] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_11[2] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_11[3] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_11[4] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_11[5] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_11[6] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_11[7] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_11[8] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_12[0] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_12[1] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_12[2] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_12[3] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_12[4] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_12[5] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_12[6] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_12[7] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_12[8] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_13[0] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_13[1] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_13[2] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_13[3] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_13[4] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_13[5] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_13[6] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_13[7] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_13[8] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_14[0] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_14[1] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_14[2] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_14[3] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_14[4] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_14[5] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_14[6] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_14[7] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_14[8] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_8[0] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_8[1] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_8[2] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_8[3] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_8[4] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_8[5] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_8[6] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_8[7] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_8[8] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_9[0] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_9[1] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_9[2] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_9[3] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_9[4] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_9[5] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_9[6] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_9[7] ;
 wire \uart.uartArea_uart.sharedFifo.fifoRegs_9[8] ;
 wire \uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[0] ;
 wire \uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[1] ;
 wire \uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[2] ;
 wire \uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[3] ;
 wire \uart.uartArea_uart.txFifo.count[0] ;
 wire \uart.uartArea_uart.txFifo.count[1] ;
 wire \uart.uartArea_uart.txFifo.count[2] ;
 wire \uart.uartArea_uart.txFifo.count[3] ;
 wire \uart.uartArea_uart.uartClocking_1.bitCtr[0] ;
 wire \uart.uartArea_uart.uartClocking_1.bitCtr[1] ;
 wire \uart.uartArea_uart.uartClocking_1.bitCtr[2] ;
 wire \uart.uartArea_uart.uartClocking_1.bitCtr[3] ;
 wire \uart.uartArea_uart.uartClocking_1.divisorCtr[0] ;
 wire \uart.uartArea_uart.uartClocking_1.divisorCtr[1] ;
 wire \uart.uartArea_uart.uartClocking_1.divisorCtr[2] ;
 wire \uart.uartArea_uart.uartClocking_1.divisorCtr[3] ;
 wire \uart.uartArea_uart.uartClocking_1.divisorCtr[4] ;
 wire \uart.uartArea_uart.uartClocking_1.divisorCtr[5] ;
 wire \uart.uartArea_uart.uartClocking_1.divisorCtr[6] ;
 wire \uart.uartArea_uart.uartClocking_1.divisorCtr[7] ;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire \async_reset_ctrl/_00_ ;
 wire \async_reset_ctrl/_01_ ;
 wire \async_reset_ctrl/_02_ ;
 wire net223;
 wire \async_reset_ctrl/_04_ ;
 wire net224;
 wire \async_reset_ctrl/_06_ ;
 wire \async_reset_ctrl/_07_ ;
 wire \async_reset_ctrl/_08_ ;
 wire \async_reset_ctrl/_09_ ;
 wire \async_reset_ctrl/_10_ ;
 wire net221;
 wire net222;
 wire \async_reset_ctrl/async_reset_in_triggered ;
 wire \async_reset_ctrl/dff3.d ;
 wire \async_reset_ctrl/dff3.q ;
 wire \async_reset_ctrl/dff_async_set1.q ;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire delaynet_0_clk;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;

 sg13g2_inv_1 _0732_ (.Y(_0150_),
    .A(\uart.uartArea_uart.rxFifo.count[3] ));
 sg13g2_inv_1 _0733_ (.Y(_0151_),
    .A(net330));
 sg13g2_inv_1 _0734_ (.Y(_0152_),
    .A(\uart.uartArea_uart.commFilter.dcdFilter.io_o ));
 sg13g2_inv_1 _0735_ (.Y(_0153_),
    .A(net301));
 sg13g2_inv_1 _0736_ (.Y(_0154_),
    .A(net377));
 sg13g2_inv_1 _0737_ (.Y(_0155_),
    .A(net367));
 sg13g2_inv_1 _0738_ (.Y(_0156_),
    .A(net379));
 sg13g2_inv_1 _0739_ (.Y(_0157_),
    .A(net415));
 sg13g2_inv_1 _0740_ (.Y(_0158_),
    .A(net233));
 sg13g2_inv_1 _0741_ (.Y(_0159_),
    .A(net230));
 sg13g2_inv_1 _0742_ (.Y(_0160_),
    .A(\uart.uartArea_uart.uartClocking_1.bitCtr[0] ));
 sg13g2_inv_1 _0743_ (.Y(_0161_),
    .A(net179));
 sg13g2_inv_1 _0744_ (.Y(_0162_),
    .A(net180));
 sg13g2_inv_1 _0745_ (.Y(_0163_),
    .A(net181));
 sg13g2_inv_2 _0746_ (.Y(_0164_),
    .A(net182));
 sg13g2_inv_1 _0747_ (.Y(_0165_),
    .A(net183));
 sg13g2_inv_1 _0748_ (.Y(_0166_),
    .A(net9));
 sg13g2_inv_1 _0749_ (.Y(_0167_),
    .A(net8));
 sg13g2_inv_1 _0750_ (.Y(_0168_),
    .A(net187));
 sg13g2_inv_1 _0751_ (.Y(_0169_),
    .A(net176));
 sg13g2_inv_1 _0752_ (.Y(_0170_),
    .A(net177));
 sg13g2_inv_2 _0753_ (.Y(_0171_),
    .A(_0000_));
 sg13g2_inv_1 _0754_ (.Y(_0172_),
    .A(net250));
 sg13g2_inv_1 _0755_ (.Y(_0173_),
    .A(\uart.uartArea_uart.regCtrl.riSignalNext ));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_and2_1 _0757_ (.A(\uart.uartArea_uart.busCtrl.io_regAddr[3] ),
    .B(\uart.uartArea_uart.busCtrl.io_regAddr[2] ),
    .X(_0174_));
 sg13g2_nand2_1 _0758_ (.Y(_0175_),
    .A(net409),
    .B(\uart.uartArea_uart.busCtrl.io_regAddr[2] ));
 sg13g2_nand2b_1 _0759_ (.Y(_0176_),
    .B(\uart.uartArea_uart.busCtrl.io_regAddr[0] ),
    .A_N(\uart.uartArea_uart.busCtrl.io_regAddr[4] ));
 sg13g2_nand3b_1 _0760_ (.B(\uart.uartArea_uart.busCtrl.io_regAddr[1] ),
    .C(\uart.uartArea_uart.busCtrl.io_regAddr[0] ),
    .Y(_0177_),
    .A_N(\uart.uartArea_uart.busCtrl.io_regAddr[4] ));
 sg13g2_or2_1 _0761_ (.X(_0178_),
    .B(_0177_),
    .A(_0175_));
 sg13g2_and2_1 _0762_ (.A(net3),
    .B(net2),
    .X(_0049_));
 sg13g2_nor2b_1 _0763_ (.A(\uart.uartArea_uart.busCtrl.lastWasWrite ),
    .B_N(_0049_),
    .Y(_0179_));
 sg13g2_nand3b_1 _0764_ (.B(net2),
    .C(net3),
    .Y(_0180_),
    .A_N(\uart.uartArea_uart.busCtrl.lastWasWrite ));
 sg13g2_nand2_2 _0765_ (.Y(_0181_),
    .A(net179),
    .B(net174));
 sg13g2_nor2_1 _0766_ (.A(_0178_),
    .B(_0181_),
    .Y(\uart.resetCommandStrobe ));
 sg13g2_nand2b_1 _0767_ (.Y(_0182_),
    .B(rst_n_sync),
    .A_N(\uart.resetCommandUnit_1.async.area_io_r ));
 sg13g2_nor4_1 _0768_ (.A(\uart.resetCommandUnit_1.ff ),
    .B(_0178_),
    .C(_0181_),
    .D(_0182_),
    .Y(_0050_));
 sg13g2_nand2b_1 _0769_ (.Y(_0183_),
    .B(net177),
    .A_N(net176));
 sg13g2_xor2_1 _0770_ (.B(net177),
    .A(net176),
    .X(_0184_));
 sg13g2_nor2_1 _0771_ (.A(net176),
    .B(net177),
    .Y(_0185_));
 sg13g2_nor2b_1 _0772_ (.A(\uart.uartArea_uart.busCtrl.io_regAddr[2] ),
    .B_N(\uart.uartArea_uart.busCtrl.io_regAddr[3] ),
    .Y(_0186_));
 sg13g2_a22oi_1 _0773_ (.Y(_0187_),
    .B1(_0185_),
    .B2(_0186_),
    .A2(_0184_),
    .A1(_0174_));
 sg13g2_o21ai_1 _0774_ (.B1(_0178_),
    .Y(_0188_),
    .A1(_0171_),
    .A2(_0187_));
 sg13g2_nand3_1 _0775_ (.B(net174),
    .C(_0188_),
    .A(net187),
    .Y(_0189_));
 sg13g2_nor2_1 _0776_ (.A(\uart.uartArea_uart.busCtrl.io_regAddr[3] ),
    .B(\uart.uartArea_uart.busCtrl.io_regAddr[2] ),
    .Y(_0190_));
 sg13g2_or2_1 _0777_ (.X(_0191_),
    .B(\uart.uartArea_uart.busCtrl.io_regAddr[2] ),
    .A(\uart.uartArea_uart.busCtrl.io_regAddr[3] ));
 sg13g2_nand2_1 _0778_ (.Y(_0192_),
    .A(_0000_),
    .B(_0190_));
 sg13g2_nor3_2 _0779_ (.A(net176),
    .B(net177),
    .C(_0192_),
    .Y(_0193_));
 sg13g2_nand3_1 _0780_ (.B(_0185_),
    .C(_0190_),
    .A(_0000_),
    .Y(_0194_));
 sg13g2_nor2b_1 _0781_ (.A(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[2] ),
    .B_N(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[3] ),
    .Y(_0195_));
 sg13g2_nand2b_1 _0782_ (.Y(_0196_),
    .B(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[3] ),
    .A_N(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[2] ));
 sg13g2_nand2_1 _0783_ (.Y(_0197_),
    .A(net373),
    .B(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[0] ));
 sg13g2_nor2_1 _0784_ (.A(_0196_),
    .B(_0197_),
    .Y(_0198_));
 sg13g2_nand2b_1 _0785_ (.Y(_0199_),
    .B(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[1] ),
    .A_N(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[0] ));
 sg13g2_nor2_2 _0786_ (.A(_0196_),
    .B(_0199_),
    .Y(_0200_));
 sg13g2_nand2b_1 _0787_ (.Y(_0201_),
    .B(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[0] ),
    .A_N(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[1] ));
 sg13g2_nor2_1 _0788_ (.A(_0196_),
    .B(_0201_),
    .Y(_0202_));
 sg13g2_and2_1 _0789_ (.A(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[3] ),
    .B(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[2] ),
    .X(_0203_));
 sg13g2_nand2_1 _0790_ (.Y(_0204_),
    .A(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[3] ),
    .B(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[2] ));
 sg13g2_nor2_1 _0791_ (.A(_0201_),
    .B(_0204_),
    .Y(_0205_));
 sg13g2_or2_1 _0792_ (.X(_0206_),
    .B(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[0] ),
    .A(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[1] ));
 sg13g2_a22oi_1 _0793_ (.Y(_0207_),
    .B1(_0206_),
    .B2(_0195_),
    .A2(_0203_),
    .A1(_0197_));
 sg13g2_nor2_1 _0794_ (.A(_0204_),
    .B(_0206_),
    .Y(_0208_));
 sg13g2_nor2_1 _0795_ (.A(_0199_),
    .B(_0204_),
    .Y(_0209_));
 sg13g2_nand2_1 _0796_ (.Y(_0210_),
    .A(\uart.uartArea_uart.sharedFifo.fifoRegs_14[8] ),
    .B(net158));
 sg13g2_a22oi_1 _0797_ (.Y(_0211_),
    .B1(net161),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_13[8] ),
    .A2(net163),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_10[8] ));
 sg13g2_inv_1 _0798_ (.Y(_0212_),
    .A(_0211_));
 sg13g2_a22oi_1 _0799_ (.Y(_0213_),
    .B1(net159),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_12[8] ),
    .A2(net162),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_9[8] ));
 sg13g2_a22oi_1 _0800_ (.Y(_0214_),
    .B1(net160),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_8[8] ),
    .A2(net164),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_11[8] ));
 sg13g2_nand3_1 _0801_ (.B(_0213_),
    .C(_0214_),
    .A(_0210_),
    .Y(_0215_));
 sg13g2_o21ai_1 _0802_ (.B1(_0193_),
    .Y(_0216_),
    .A1(_0212_),
    .A2(_0215_));
 sg13g2_nand2b_2 _0803_ (.Y(_0217_),
    .B(\uart.uartArea_uart.busCtrl.io_regAddr[2] ),
    .A_N(\uart.uartArea_uart.busCtrl.io_regAddr[3] ));
 sg13g2_nor4_2 _0804_ (.A(net176),
    .B(net177),
    .C(_0171_),
    .Y(_0218_),
    .D(_0217_));
 sg13g2_nor3_1 _0805_ (.A(\uart.uartArea_uart.txFifo.count[2] ),
    .B(\uart.uartArea_uart.txFifo.count[1] ),
    .C(\uart.uartArea_uart.txFifo.count[0] ),
    .Y(_0219_));
 sg13g2_nand2_2 _0806_ (.Y(_0220_),
    .A(\uart.uartArea_uart.txFifo.count[3] ),
    .B(_0219_));
 sg13g2_inv_1 _0807_ (.Y(_0221_),
    .A(_0220_));
 sg13g2_nor4_2 _0808_ (.A(_0169_),
    .B(net177),
    .C(\uart.uartArea_uart.busCtrl.io_regAddr[2] ),
    .Y(_0222_),
    .D(_0171_));
 sg13g2_a22oi_1 _0809_ (.Y(_0223_),
    .B1(_0222_),
    .B2(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[0] ),
    .A2(_0220_),
    .A1(_0218_));
 sg13g2_nor2_2 _0810_ (.A(_0177_),
    .B(_0217_),
    .Y(_0224_));
 sg13g2_nor3_2 _0811_ (.A(net176),
    .B(_0176_),
    .C(_0217_),
    .Y(_0225_));
 sg13g2_a22oi_1 _0812_ (.Y(_0226_),
    .B1(_0225_),
    .B2(\uart.uartArea_uart.regCtrl.regModemCtrlChanged[0] ),
    .A2(_0224_),
    .A1(\uart.uartArea_uart.regCtrl.reg007[0] ));
 sg13g2_o21ai_1 _0813_ (.B1(net177),
    .Y(_0227_),
    .A1(\uart.uartArea_uart.busCtrl.io_regAddr[1] ),
    .A2(_0175_));
 sg13g2_a21oi_1 _0814_ (.A1(_0169_),
    .A2(_0217_),
    .Y(_0228_),
    .B1(_0176_));
 sg13g2_a21oi_1 _0815_ (.A1(_0000_),
    .A2(_0227_),
    .Y(_0229_),
    .B1(_0228_));
 sg13g2_a21o_2 _0816_ (.A2(_0227_),
    .A1(_0000_),
    .B1(_0228_),
    .X(_0230_));
 sg13g2_nor2_2 _0817_ (.A(_0177_),
    .B(_0191_),
    .Y(_0231_));
 sg13g2_a21oi_1 _0818_ (.A1(\uart.uartArea_uart.regCtrl.io_regInterruptControl[0] ),
    .A2(_0231_),
    .Y(_0232_),
    .B1(net152));
 sg13g2_and4_1 _0819_ (.A(_0189_),
    .B(_0223_),
    .C(_0226_),
    .D(_0232_),
    .X(_0233_));
 sg13g2_a22oi_1 _0820_ (.Y(_0234_),
    .B1(net161),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_13[0] ),
    .A2(net163),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_10[0] ));
 sg13g2_a22oi_1 _0821_ (.Y(_0235_),
    .B1(net158),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_14[0] ),
    .A2(net164),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_11[0] ));
 sg13g2_a22oi_1 _0822_ (.Y(_0236_),
    .B1(net159),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_12[0] ),
    .A2(net162),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_9[0] ));
 sg13g2_nand2_1 _0823_ (.Y(_0237_),
    .A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[0] ),
    .B(net160));
 sg13g2_and4_1 _0824_ (.A(_0234_),
    .B(_0235_),
    .C(_0236_),
    .D(_0237_),
    .X(_0238_));
 sg13g2_a22oi_1 _0825_ (.Y(uio_out[0]),
    .B1(_0238_),
    .B2(net151),
    .A2(_0233_),
    .A1(_0216_));
 sg13g2_nand3_1 _0826_ (.B(net174),
    .C(_0188_),
    .A(net185),
    .Y(_0239_));
 sg13g2_nor3_1 _0827_ (.A(net348),
    .B(\uart.uartArea_uart.rxFifo.count[1] ),
    .C(\uart.uartArea_uart.rxFifo.count[0] ),
    .Y(_0240_));
 sg13g2_nand3_1 _0828_ (.B(_0193_),
    .C(_0240_),
    .A(\uart.uartArea_uart.rxFifo.count[3] ),
    .Y(_0241_));
 sg13g2_and2_1 _0829_ (.A(\uart.uartArea_uart.txFifo.count[1] ),
    .B(\uart.uartArea_uart.txFifo.count[0] ),
    .X(_0242_));
 sg13g2_nand4_1 _0830_ (.B(\uart.uartArea_uart.txFifo.count[2] ),
    .C(_0218_),
    .A(_0157_),
    .Y(_0243_),
    .D(_0242_));
 sg13g2_a221oi_1 _0831_ (.B2(\uart.uartArea_uart.regCtrl.regModemCtrlChanged[1] ),
    .C1(net152),
    .B1(net157),
    .A1(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[1] ),
    .Y(_0244_),
    .A2(_0222_));
 sg13g2_a22oi_1 _0832_ (.Y(_0245_),
    .B1(_0231_),
    .B2(\uart.uartArea_uart.regCtrl.io_regInterruptControl[1] ),
    .A2(_0224_),
    .A1(\uart.uartArea_uart.regCtrl.reg007[1] ));
 sg13g2_and4_1 _0833_ (.A(_0241_),
    .B(_0243_),
    .C(_0244_),
    .D(_0245_),
    .X(_0246_));
 sg13g2_nand2_1 _0834_ (.Y(_0247_),
    .A(\uart.uartArea_uart.sharedFifo.fifoRegs_14[1] ),
    .B(net158));
 sg13g2_a22oi_1 _0835_ (.Y(_0248_),
    .B1(net161),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_13[1] ),
    .A2(net164),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_11[1] ));
 sg13g2_a22oi_1 _0836_ (.Y(_0249_),
    .B1(net160),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_8[1] ),
    .A2(net162),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_9[1] ));
 sg13g2_a22oi_1 _0837_ (.Y(_0250_),
    .B1(net159),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_12[1] ),
    .A2(net163),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_10[1] ));
 sg13g2_and4_1 _0838_ (.A(_0247_),
    .B(_0248_),
    .C(_0249_),
    .D(_0250_),
    .X(_0251_));
 sg13g2_a22oi_1 _0839_ (.Y(uio_out[1]),
    .B1(_0251_),
    .B2(net151),
    .A2(_0246_),
    .A1(_0239_));
 sg13g2_nand3_1 _0840_ (.B(_0179_),
    .C(_0188_),
    .A(net184),
    .Y(_0252_));
 sg13g2_and4_1 _0841_ (.A(_0150_),
    .B(\uart.uartArea_uart.rxFifo.count[2] ),
    .C(\uart.uartArea_uart.rxFifo.count[1] ),
    .D(\uart.uartArea_uart.rxFifo.count[0] ),
    .X(_0253_));
 sg13g2_and2_1 _0842_ (.A(_0157_),
    .B(_0219_),
    .X(_0254_));
 sg13g2_a22oi_1 _0843_ (.Y(_0255_),
    .B1(net157),
    .B2(\uart.uartArea_uart.regCtrl.regModemCtrlChanged[2] ),
    .A2(_0222_),
    .A1(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[2] ));
 sg13g2_a22oi_1 _0844_ (.Y(_0256_),
    .B1(_0231_),
    .B2(\uart.uartArea_uart.regCtrl.io_regInterruptControl[2] ),
    .A2(_0224_),
    .A1(\uart.uartArea_uart.regCtrl.reg007[2] ));
 sg13g2_a22oi_1 _0845_ (.Y(_0257_),
    .B1(_0254_),
    .B2(_0218_),
    .A2(_0253_),
    .A1(_0193_));
 sg13g2_and4_1 _0846_ (.A(_0230_),
    .B(_0255_),
    .C(_0256_),
    .D(_0257_),
    .X(_0258_));
 sg13g2_a22oi_1 _0847_ (.Y(_0259_),
    .B1(_0209_),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_14[2] ),
    .A2(net161),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_13[2] ));
 sg13g2_nand2_1 _0848_ (.Y(_0260_),
    .A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[2] ),
    .B(_0207_));
 sg13g2_a22oi_1 _0849_ (.Y(_0261_),
    .B1(_0208_),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_12[2] ),
    .A2(net162),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_9[2] ));
 sg13g2_a22oi_1 _0850_ (.Y(_0262_),
    .B1(net163),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_10[2] ),
    .A2(_0198_),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_11[2] ));
 sg13g2_and4_2 _0851_ (.A(_0259_),
    .B(_0260_),
    .C(_0261_),
    .D(_0262_),
    .X(_0263_));
 sg13g2_a22oi_1 _0852_ (.Y(uio_out[2]),
    .B1(_0263_),
    .B2(net151),
    .A2(_0258_),
    .A1(_0252_));
 sg13g2_nand3_1 _0853_ (.B(net174),
    .C(_0188_),
    .A(net10),
    .Y(_0264_));
 sg13g2_nor2b_2 _0854_ (.A(\uart.uartArea_uart.rxFifo.count[3] ),
    .B_N(_0240_),
    .Y(_0265_));
 sg13g2_a22oi_1 _0855_ (.Y(_0266_),
    .B1(_0265_),
    .B2(_0193_),
    .A2(net157),
    .A1(\uart.uartArea_uart.regCtrl.regModemCtrlChanged[3] ));
 sg13g2_a22oi_1 _0856_ (.Y(_0267_),
    .B1(_0224_),
    .B2(\uart.uartArea_uart.regCtrl.reg007[3] ),
    .A2(_0222_),
    .A1(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[3] ));
 sg13g2_a21oi_1 _0857_ (.A1(\uart.uartArea_uart.regCtrl.io_regInterruptControl[3] ),
    .A2(_0231_),
    .Y(_0268_),
    .B1(net152));
 sg13g2_and3_1 _0858_ (.X(_0269_),
    .A(_0266_),
    .B(_0267_),
    .C(_0268_));
 sg13g2_a22oi_1 _0859_ (.Y(_0270_),
    .B1(net159),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_12[3] ),
    .A2(net161),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_13[3] ));
 sg13g2_a22oi_1 _0860_ (.Y(_0271_),
    .B1(net158),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_14[3] ),
    .A2(net164),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_11[3] ));
 sg13g2_a22oi_1 _0861_ (.Y(_0272_),
    .B1(net162),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_9[3] ),
    .A2(net163),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_10[3] ));
 sg13g2_nand2_1 _0862_ (.Y(_0273_),
    .A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[3] ),
    .B(net160));
 sg13g2_and4_1 _0863_ (.A(_0270_),
    .B(_0271_),
    .C(_0272_),
    .D(_0273_),
    .X(_0274_));
 sg13g2_a22oi_1 _0864_ (.Y(uio_out[3]),
    .B1(_0274_),
    .B2(net151),
    .A2(_0269_),
    .A1(_0264_));
 sg13g2_nand3_1 _0865_ (.B(_0179_),
    .C(_0188_),
    .A(net11),
    .Y(_0275_));
 sg13g2_a22oi_1 _0866_ (.Y(_0276_),
    .B1(_0224_),
    .B2(\uart.uartArea_uart.regCtrl.reg007[4] ),
    .A2(_0222_),
    .A1(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[4] ));
 sg13g2_a22oi_1 _0867_ (.Y(_0277_),
    .B1(_0231_),
    .B2(\uart.uartArea_uart.regCtrl.io_regInterruptControl[4] ),
    .A2(net157),
    .A1(\uart.uartArea_uart.commFilter.ctsFilter.io_o ));
 sg13g2_and3_1 _0868_ (.X(_0278_),
    .A(_0230_),
    .B(_0276_),
    .C(_0277_));
 sg13g2_a22oi_1 _0869_ (.Y(_0279_),
    .B1(_0205_),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_13[4] ),
    .A2(net164),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_11[4] ));
 sg13g2_a22oi_1 _0870_ (.Y(_0280_),
    .B1(net158),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_14[4] ),
    .A2(_0202_),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_9[4] ));
 sg13g2_a22oi_1 _0871_ (.Y(_0281_),
    .B1(net159),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_12[4] ),
    .A2(net163),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_10[4] ));
 sg13g2_nand2_1 _0872_ (.Y(_0282_),
    .A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[4] ),
    .B(net160));
 sg13g2_and4_1 _0873_ (.A(_0279_),
    .B(_0280_),
    .C(_0281_),
    .D(_0282_),
    .X(_0283_));
 sg13g2_a22oi_1 _0874_ (.Y(uio_out[4]),
    .B1(_0283_),
    .B2(net151),
    .A2(_0278_),
    .A1(_0275_));
 sg13g2_a22oi_1 _0875_ (.Y(_0284_),
    .B1(net159),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_12[5] ),
    .A2(net164),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_11[5] ));
 sg13g2_and2_1 _0876_ (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[5] ),
    .B(net160),
    .X(_0285_));
 sg13g2_a221oi_1 _0877_ (.B2(\uart.uartArea_uart.sharedFifo.fifoRegs_14[5] ),
    .C1(_0285_),
    .B1(net158),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_10[5] ),
    .Y(_0286_),
    .A2(_0200_));
 sg13g2_a22oi_1 _0878_ (.Y(_0287_),
    .B1(net161),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_13[5] ),
    .A2(net162),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_9[5] ));
 sg13g2_nand4_1 _0879_ (.B(_0284_),
    .C(_0286_),
    .A(net151),
    .Y(_0288_),
    .D(_0287_));
 sg13g2_nand3_1 _0880_ (.B(net174),
    .C(_0188_),
    .A(net12),
    .Y(_0289_));
 sg13g2_a22oi_1 _0881_ (.Y(_0290_),
    .B1(_0224_),
    .B2(\uart.uartArea_uart.regCtrl.reg007[5] ),
    .A2(_0222_),
    .A1(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[5] ));
 sg13g2_a22oi_1 _0882_ (.Y(_0291_),
    .B1(_0231_),
    .B2(\uart.uartArea_uart.regCtrl.io_regInterruptControl[5] ),
    .A2(net157),
    .A1(\uart.uartArea_uart.commFilter.dsrFilter.io_o ));
 sg13g2_nand4_1 _0883_ (.B(_0289_),
    .C(_0290_),
    .A(_0230_),
    .Y(_0292_),
    .D(_0291_));
 sg13g2_and2_2 _0884_ (.A(_0288_),
    .B(_0292_),
    .X(uio_out[5]));
 sg13g2_nand2_1 _0885_ (.Y(_0293_),
    .A(net13),
    .B(net174));
 sg13g2_nand2b_1 _0886_ (.Y(_0294_),
    .B(_0188_),
    .A_N(_0293_));
 sg13g2_nand2_1 _0887_ (.Y(_0295_),
    .A(\uart.uartArea_uart.regCtrl.riSignalNext ),
    .B(net157));
 sg13g2_nor2b_2 _0888_ (.A(_0177_),
    .B_N(_0186_),
    .Y(_0296_));
 sg13g2_a22oi_1 _0889_ (.Y(_0297_),
    .B1(_0231_),
    .B2(\uart.uartArea_uart.regCtrl.io_regInterruptControl[6] ),
    .A2(_0224_),
    .A1(\uart.uartArea_uart.regCtrl.reg007[6] ));
 sg13g2_a22oi_1 _0890_ (.Y(_0298_),
    .B1(_0296_),
    .B2(\uart.uartArea_uart.regCtrl.regFifoRxEnable ),
    .A2(_0222_),
    .A1(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[6] ));
 sg13g2_and4_1 _0891_ (.A(_0230_),
    .B(_0295_),
    .C(_0297_),
    .D(_0298_),
    .X(_0299_));
 sg13g2_nand2_1 _0892_ (.Y(_0300_),
    .A(\uart.uartArea_uart.sharedFifo.fifoRegs_13[6] ),
    .B(net161));
 sg13g2_a22oi_1 _0893_ (.Y(_0301_),
    .B1(net158),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_14[6] ),
    .A2(net163),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_10[6] ));
 sg13g2_a22oi_1 _0894_ (.Y(_0302_),
    .B1(net160),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_8[6] ),
    .A2(net164),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_11[6] ));
 sg13g2_a22oi_1 _0895_ (.Y(_0303_),
    .B1(net159),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_12[6] ),
    .A2(net162),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_9[6] ));
 sg13g2_and4_1 _0896_ (.A(_0300_),
    .B(_0301_),
    .C(_0302_),
    .D(_0303_),
    .X(_0304_));
 sg13g2_a22oi_1 _0897_ (.Y(uio_out[6]),
    .B1(_0304_),
    .B2(net151),
    .A2(_0299_),
    .A1(_0294_));
 sg13g2_nand2b_1 _0898_ (.Y(_0305_),
    .B(_0188_),
    .A_N(_0181_));
 sg13g2_a22oi_1 _0899_ (.Y(_0306_),
    .B1(_0224_),
    .B2(\uart.uartArea_uart.regCtrl.reg007[7] ),
    .A2(_0218_),
    .A1(\uart.uartArea_uart.regCtrl.txOverrun ));
 sg13g2_o21ai_1 _0900_ (.B1(_0306_),
    .Y(_0307_),
    .A1(_0194_),
    .A2(_0265_));
 sg13g2_a221oi_1 _0901_ (.B2(\uart.uartArea_uart.regCtrl.regFifoTxEnable ),
    .C1(net152),
    .B1(_0296_),
    .A1(\uart.uartArea_uart.commFilter.dcdFilter.io_o ),
    .Y(_0308_),
    .A2(net157));
 sg13g2_nor2b_1 _0902_ (.A(_0307_),
    .B_N(_0308_),
    .Y(_0309_));
 sg13g2_nand2_1 _0903_ (.Y(_0310_),
    .A(\uart.uartArea_uart.sharedFifo.fifoRegs_9[7] ),
    .B(net162));
 sg13g2_a22oi_1 _0904_ (.Y(_0311_),
    .B1(net159),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_12[7] ),
    .A2(net161),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_13[7] ));
 sg13g2_a22oi_1 _0905_ (.Y(_0312_),
    .B1(net160),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_8[7] ),
    .A2(net164),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_11[7] ));
 sg13g2_a22oi_1 _0906_ (.Y(_0313_),
    .B1(net158),
    .B2(\uart.uartArea_uart.sharedFifo.fifoRegs_14[7] ),
    .A2(net163),
    .A1(\uart.uartArea_uart.sharedFifo.fifoRegs_10[7] ));
 sg13g2_and4_1 _0907_ (.A(_0310_),
    .B(_0311_),
    .C(_0312_),
    .D(_0313_),
    .X(_0314_));
 sg13g2_a22oi_1 _0908_ (.Y(uio_out[7]),
    .B1(_0314_),
    .B2(net151),
    .A2(_0309_),
    .A1(_0305_));
 sg13g2_nor3_1 _0909_ (.A(net401),
    .B(\uart.uartArea_uart.uartClocking_1.divisorCtr[1] ),
    .C(net412),
    .Y(_0315_));
 sg13g2_or4_2 _0910_ (.A(\uart.uartArea_uart.uartClocking_1.divisorCtr[0] ),
    .B(\uart.uartArea_uart.uartClocking_1.divisorCtr[1] ),
    .C(\uart.uartArea_uart.uartClocking_1.divisorCtr[2] ),
    .D(net265),
    .X(_0316_));
 sg13g2_nor3_1 _0911_ (.A(net420),
    .B(net426),
    .C(_0316_),
    .Y(_0317_));
 sg13g2_nor4_2 _0912_ (.A(\uart.uartArea_uart.uartClocking_1.divisorCtr[4] ),
    .B(\uart.uartArea_uart.uartClocking_1.divisorCtr[5] ),
    .C(\uart.uartArea_uart.uartClocking_1.divisorCtr[6] ),
    .Y(_0318_),
    .D(_0316_));
 sg13g2_nand2_2 _0913_ (.Y(_0319_),
    .A(_0172_),
    .B(_0318_));
 sg13g2_nor2b_1 _0914_ (.A(net408),
    .B_N(\uart.resetCommandUnit_1.async.area_io_r ),
    .Y(_0320_));
 sg13g2_nand2b_1 _0915_ (.Y(_0321_),
    .B(\uart.resetCommandUnit_1.async.area_io_r ),
    .A_N(\uart.resetCommandUnit_1.io_resetIn ));
 sg13g2_nand2_2 _0916_ (.Y(_0322_),
    .A(_0319_),
    .B(net169));
 sg13g2_and3_1 _0917_ (.X(_0006_),
    .A(net231),
    .B(_0319_),
    .C(net169));
 sg13g2_xor2_1 _0918_ (.B(\uart.uartArea_uart.uartClocking_1.divisorCtr[1] ),
    .A(net401),
    .X(_0323_));
 sg13g2_nor2_1 _0919_ (.A(_0322_),
    .B(net402),
    .Y(_0007_));
 sg13g2_o21ai_1 _0920_ (.B1(net412),
    .Y(_0324_),
    .A1(net401),
    .A2(\uart.uartArea_uart.uartClocking_1.divisorCtr[1] ));
 sg13g2_nor2b_1 _0921_ (.A(net413),
    .B_N(_0324_),
    .Y(_0325_));
 sg13g2_nor2_1 _0922_ (.A(_0322_),
    .B(net414),
    .Y(_0008_));
 sg13g2_nand2b_1 _0923_ (.Y(_0326_),
    .B(net265),
    .A_N(_0315_));
 sg13g2_a21oi_1 _0924_ (.A1(_0316_),
    .A2(net266),
    .Y(_0009_),
    .B1(_0322_));
 sg13g2_xor2_1 _0925_ (.B(_0316_),
    .A(net420),
    .X(_0327_));
 sg13g2_nor2_1 _0926_ (.A(_0322_),
    .B(net421),
    .Y(_0010_));
 sg13g2_o21ai_1 _0927_ (.B1(net426),
    .Y(_0328_),
    .A1(net420),
    .A2(_0316_));
 sg13g2_nor2b_1 _0928_ (.A(net427),
    .B_N(_0328_),
    .Y(_0329_));
 sg13g2_nor2_1 _0929_ (.A(_0322_),
    .B(_0329_),
    .Y(_0011_));
 sg13g2_xnor2_1 _0930_ (.Y(_0330_),
    .A(net387),
    .B(_0317_));
 sg13g2_nor2_1 _0931_ (.A(_0322_),
    .B(net388),
    .Y(_0012_));
 sg13g2_nor3_1 _0932_ (.A(_0172_),
    .B(_0318_),
    .C(net170),
    .Y(_0013_));
 sg13g2_nand2_1 _0933_ (.Y(_0331_),
    .A(_0153_),
    .B(net377));
 sg13g2_a21oi_1 _0934_ (.A1(net301),
    .A2(_0154_),
    .Y(_0332_),
    .B1(\uart.uartArea_uart.regCtrl.regModemCtrlChanged[1] ));
 sg13g2_a21oi_1 _0935_ (.A1(_0331_),
    .A2(_0332_),
    .Y(_0014_),
    .B1(net171));
 sg13g2_a21oi_1 _0936_ (.A1(net230),
    .A2(_0173_),
    .Y(_0333_),
    .B1(net270));
 sg13g2_nor2_1 _0937_ (.A(net171),
    .B(net271),
    .Y(_0015_));
 sg13g2_nor4_2 _0938_ (.A(_0171_),
    .B(net172),
    .C(_0183_),
    .Y(_0334_),
    .D(_0191_));
 sg13g2_a21oi_1 _0939_ (.A1(_0221_),
    .A2(_0334_),
    .Y(_0335_),
    .B1(net243));
 sg13g2_nor2_1 _0940_ (.A(net170),
    .B(net244),
    .Y(_0016_));
 sg13g2_nor2_1 _0941_ (.A(net172),
    .B(_0194_),
    .Y(_0336_));
 sg13g2_mux2_1 _0942_ (.A0(net425),
    .A1(net186),
    .S(_0336_),
    .X(_0017_));
 sg13g2_a21oi_1 _0943_ (.A1(net174),
    .A2(_0296_),
    .Y(_0337_),
    .B1(net170));
 sg13g2_a21o_2 _0944_ (.A2(_0296_),
    .A1(net174),
    .B1(net170),
    .X(_0338_));
 sg13g2_nand2_1 _0945_ (.Y(_0339_),
    .A(net254),
    .B(net150));
 sg13g2_nand2_1 _0946_ (.Y(_0340_),
    .A(_0296_),
    .B(net167));
 sg13g2_o21ai_1 _0947_ (.B1(_0339_),
    .Y(_0018_),
    .A1(_0181_),
    .A2(_0340_));
 sg13g2_nand2_1 _0948_ (.Y(_0341_),
    .A(net249),
    .B(net150));
 sg13g2_o21ai_1 _0949_ (.B1(_0341_),
    .Y(_0019_),
    .A1(_0293_),
    .A2(_0340_));
 sg13g2_nand2_1 _0950_ (.Y(_0342_),
    .A(_0151_),
    .B(\uart.uartArea_uart.commFilter.dcdFilter.io_o ));
 sg13g2_a21oi_1 _0951_ (.A1(net330),
    .A2(_0152_),
    .Y(_0343_),
    .B1(net341));
 sg13g2_a21oi_1 _0952_ (.A1(_0342_),
    .A2(net342),
    .Y(_0020_),
    .B1(net170));
 sg13g2_nand2b_2 _0953_ (.Y(_0344_),
    .B(net3),
    .A_N(net2));
 sg13g2_nand4_1 _0954_ (.B(_0170_),
    .C(_0000_),
    .A(net176),
    .Y(_0345_),
    .D(_0190_));
 sg13g2_a21oi_2 _0955_ (.B1(_0345_),
    .Y(_0346_),
    .A2(_0344_),
    .A1(net172));
 sg13g2_o21ai_1 _0956_ (.B1(_0346_),
    .Y(_0347_),
    .A1(net187),
    .A2(net172));
 sg13g2_and3_1 _0957_ (.X(_0021_),
    .A(net242),
    .B(net165),
    .C(_0347_));
 sg13g2_o21ai_1 _0958_ (.B1(_0346_),
    .Y(_0348_),
    .A1(net8),
    .A2(net172));
 sg13g2_and3_1 _0959_ (.X(_0022_),
    .A(net252),
    .B(net165),
    .C(_0348_));
 sg13g2_o21ai_1 _0960_ (.B1(_0346_),
    .Y(_0349_),
    .A1(net9),
    .A2(net173));
 sg13g2_and3_1 _0961_ (.X(_0023_),
    .A(net237),
    .B(net166),
    .C(_0349_));
 sg13g2_o21ai_1 _0962_ (.B1(_0346_),
    .Y(_0350_),
    .A1(net10),
    .A2(net172));
 sg13g2_and3_1 _0963_ (.X(_0024_),
    .A(net240),
    .B(net165),
    .C(_0350_));
 sg13g2_o21ai_1 _0964_ (.B1(_0346_),
    .Y(_0351_),
    .A1(net11),
    .A2(net173));
 sg13g2_and3_1 _0965_ (.X(_0025_),
    .A(net239),
    .B(net166),
    .C(_0351_));
 sg13g2_o21ai_1 _0966_ (.B1(_0346_),
    .Y(_0352_),
    .A1(net12),
    .A2(net173));
 sg13g2_and3_1 _0967_ (.X(_0026_),
    .A(net238),
    .B(net166),
    .C(_0352_));
 sg13g2_o21ai_1 _0968_ (.B1(_0346_),
    .Y(_0353_),
    .A1(net13),
    .A2(net173));
 sg13g2_and3_1 _0969_ (.X(_0027_),
    .A(net241),
    .B(net166),
    .C(_0353_));
 sg13g2_nor3_1 _0970_ (.A(_0177_),
    .B(net172),
    .C(_0191_),
    .Y(_0354_));
 sg13g2_o21ai_1 _0971_ (.B1(net167),
    .Y(_0355_),
    .A1(net407),
    .A2(net155));
 sg13g2_a21oi_1 _0972_ (.A1(_0168_),
    .A2(net155),
    .Y(_0028_),
    .B1(_0355_));
 sg13g2_o21ai_1 _0973_ (.B1(net165),
    .Y(_0356_),
    .A1(net392),
    .A2(net156));
 sg13g2_a21oi_1 _0974_ (.A1(_0167_),
    .A2(net156),
    .Y(_0029_),
    .B1(_0356_));
 sg13g2_o21ai_1 _0975_ (.B1(net167),
    .Y(_0357_),
    .A1(net403),
    .A2(net155));
 sg13g2_a21oi_1 _0976_ (.A1(_0166_),
    .A2(net155),
    .Y(_0030_),
    .B1(_0357_));
 sg13g2_o21ai_1 _0977_ (.B1(net165),
    .Y(_0358_),
    .A1(net398),
    .A2(net156));
 sg13g2_a21oi_1 _0978_ (.A1(_0165_),
    .A2(net156),
    .Y(_0031_),
    .B1(_0358_));
 sg13g2_o21ai_1 _0979_ (.B1(net167),
    .Y(_0359_),
    .A1(net406),
    .A2(net155));
 sg13g2_a21oi_1 _0980_ (.A1(_0164_),
    .A2(net155),
    .Y(_0032_),
    .B1(_0359_));
 sg13g2_o21ai_1 _0981_ (.B1(net166),
    .Y(_0360_),
    .A1(net419),
    .A2(net155));
 sg13g2_a21oi_1 _0982_ (.A1(_0163_),
    .A2(net156),
    .Y(_0033_),
    .B1(_0360_));
 sg13g2_o21ai_1 _0983_ (.B1(net166),
    .Y(_0361_),
    .A1(net397),
    .A2(net156));
 sg13g2_a21oi_1 _0984_ (.A1(_0162_),
    .A2(net155),
    .Y(_0034_),
    .B1(_0361_));
 sg13g2_nor3_2 _0985_ (.A(_0177_),
    .B(net172),
    .C(_0217_),
    .Y(_0362_));
 sg13g2_o21ai_1 _0986_ (.B1(net167),
    .Y(_0363_),
    .A1(net376),
    .A2(net153));
 sg13g2_a21oi_1 _0987_ (.A1(_0168_),
    .A2(net153),
    .Y(_0035_),
    .B1(_0363_));
 sg13g2_o21ai_1 _0988_ (.B1(net165),
    .Y(_0364_),
    .A1(net394),
    .A2(net154));
 sg13g2_a21oi_1 _0989_ (.A1(_0167_),
    .A2(net154),
    .Y(_0036_),
    .B1(_0364_));
 sg13g2_o21ai_1 _0990_ (.B1(net167),
    .Y(_0365_),
    .A1(net375),
    .A2(net153));
 sg13g2_a21oi_1 _0991_ (.A1(_0166_),
    .A2(net153),
    .Y(_0037_),
    .B1(_0365_));
 sg13g2_o21ai_1 _0992_ (.B1(net165),
    .Y(_0366_),
    .A1(net396),
    .A2(net154));
 sg13g2_a21oi_1 _0993_ (.A1(_0165_),
    .A2(net154),
    .Y(_0038_),
    .B1(_0366_));
 sg13g2_o21ai_1 _0994_ (.B1(net167),
    .Y(_0367_),
    .A1(net399),
    .A2(net153));
 sg13g2_a21oi_1 _0995_ (.A1(_0164_),
    .A2(net153),
    .Y(_0039_),
    .B1(_0367_));
 sg13g2_o21ai_1 _0996_ (.B1(net166),
    .Y(_0368_),
    .A1(net400),
    .A2(net153));
 sg13g2_a21oi_1 _0997_ (.A1(_0163_),
    .A2(net154),
    .Y(_0040_),
    .B1(_0368_));
 sg13g2_o21ai_1 _0998_ (.B1(net166),
    .Y(_0369_),
    .A1(net405),
    .A2(net153));
 sg13g2_a21oi_1 _0999_ (.A1(_0162_),
    .A2(_0362_),
    .Y(_0041_),
    .B1(_0369_));
 sg13g2_o21ai_1 _1000_ (.B1(net165),
    .Y(_0370_),
    .A1(net393),
    .A2(net154));
 sg13g2_a21oi_1 _1001_ (.A1(_0161_),
    .A2(net154),
    .Y(_0042_),
    .B1(_0370_));
 sg13g2_or4_2 _1002_ (.A(net313),
    .B(net384),
    .C(net389),
    .D(_0319_),
    .X(_0371_));
 sg13g2_nor2_2 _1003_ (.A(net383),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_mux2_1 _1004_ (.A0(net344),
    .A1(net363),
    .S(_0372_),
    .X(_0043_));
 sg13g2_nand2b_1 _1005_ (.Y(_0373_),
    .B(net2),
    .A_N(net3));
 sg13g2_nor2_1 _1006_ (.A(net187),
    .B(net178),
    .Y(_0374_));
 sg13g2_a21oi_1 _1007_ (.A1(_0170_),
    .A2(net178),
    .Y(_0044_),
    .B1(_0374_));
 sg13g2_nor2_1 _1008_ (.A(net8),
    .B(net178),
    .Y(_0375_));
 sg13g2_a21oi_1 _1009_ (.A1(_0169_),
    .A2(net178),
    .Y(_0045_),
    .B1(_0375_));
 sg13g2_nand2_1 _1010_ (.Y(_0376_),
    .A(net424),
    .B(_0373_));
 sg13g2_o21ai_1 _1011_ (.B1(_0376_),
    .Y(_0046_),
    .A1(_0166_),
    .A2(_0373_));
 sg13g2_nand2_1 _1012_ (.Y(_0377_),
    .A(net409),
    .B(net178));
 sg13g2_o21ai_1 _1013_ (.B1(_0377_),
    .Y(_0047_),
    .A1(_0165_),
    .A2(net178));
 sg13g2_nand2_1 _1014_ (.Y(_0378_),
    .A(net281),
    .B(net178));
 sg13g2_o21ai_1 _1015_ (.B1(_0378_),
    .Y(_0048_),
    .A1(_0164_),
    .A2(net178));
 sg13g2_nor2_1 _1016_ (.A(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[3] ),
    .B(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[2] ),
    .Y(_0379_));
 sg13g2_or2_1 _1017_ (.X(_0380_),
    .B(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[2] ),
    .A(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[3] ));
 sg13g2_and2_2 _1018_ (.A(_0220_),
    .B(_0334_),
    .X(_0381_));
 sg13g2_nand2_1 _1019_ (.Y(_0382_),
    .A(_0220_),
    .B(_0334_));
 sg13g2_nor2_1 _1020_ (.A(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[1] ),
    .B(_0382_),
    .Y(_0383_));
 sg13g2_and4_1 _1021_ (.A(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[0] ),
    .B(net149),
    .C(_0379_),
    .D(_0383_),
    .X(_0384_));
 sg13g2_mux2_1 _1022_ (.A0(net287),
    .A1(net186),
    .S(net147),
    .X(_0051_));
 sg13g2_mux2_1 _1023_ (.A0(net283),
    .A1(net185),
    .S(net147),
    .X(_0052_));
 sg13g2_mux2_1 _1024_ (.A0(net299),
    .A1(net184),
    .S(net147),
    .X(_0053_));
 sg13g2_mux2_1 _1025_ (.A0(net310),
    .A1(net183),
    .S(net147),
    .X(_0054_));
 sg13g2_mux2_1 _1026_ (.A0(net365),
    .A1(net182),
    .S(_0384_),
    .X(_0055_));
 sg13g2_mux2_1 _1027_ (.A0(net327),
    .A1(net181),
    .S(net147),
    .X(_0056_));
 sg13g2_mux2_1 _1028_ (.A0(net309),
    .A1(net180),
    .S(net147),
    .X(_0057_));
 sg13g2_mux2_1 _1029_ (.A0(net328),
    .A1(net14),
    .S(net147),
    .X(_0058_));
 sg13g2_mux2_1 _1030_ (.A0(net278),
    .A1(\uart.uartArea_uart.regCtrl.txHolderBit9 ),
    .S(net147),
    .X(_0059_));
 sg13g2_o21ai_1 _1031_ (.B1(net169),
    .Y(_0385_),
    .A1(net246),
    .A2(_0319_));
 sg13g2_a21oi_1 _1032_ (.A1(_0160_),
    .A2(_0319_),
    .Y(_0060_),
    .B1(net247));
 sg13g2_or3_1 _1033_ (.A(net384),
    .B(\uart.uartArea_uart.uartClocking_1.bitCtr[0] ),
    .C(_0319_),
    .X(_0386_));
 sg13g2_o21ai_1 _1034_ (.B1(net384),
    .Y(_0387_),
    .A1(\uart.uartArea_uart.uartClocking_1.bitCtr[0] ),
    .A2(_0319_));
 sg13g2_a21oi_1 _1035_ (.A1(_0386_),
    .A2(net385),
    .Y(_0061_),
    .B1(net170));
 sg13g2_nand2_1 _1036_ (.Y(_0388_),
    .A(net313),
    .B(_0386_));
 sg13g2_a21oi_1 _1037_ (.A1(_0371_),
    .A2(net314),
    .Y(_0062_),
    .B1(net170));
 sg13g2_xor2_1 _1038_ (.B(_0371_),
    .A(net383),
    .X(_0389_));
 sg13g2_nor2_1 _1039_ (.A(net170),
    .B(_0389_),
    .Y(_0063_));
 sg13g2_nand3_1 _1040_ (.B(net7),
    .C(\uart.uartArea_uart.commFilter.riFilter.io_b ),
    .A(net344),
    .Y(_0390_));
 sg13g2_nor3_1 _1041_ (.A(net344),
    .B(net7),
    .C(\uart.uartArea_uart.commFilter.riFilter.io_b ),
    .Y(_0391_));
 sg13g2_a21oi_1 _1042_ (.A1(_0159_),
    .A2(net345),
    .Y(_0064_),
    .B1(_0391_));
 sg13g2_nand3_1 _1043_ (.B(net5),
    .C(\uart.uartArea_uart.commFilter.dcdFilter.io_b ),
    .A(net322),
    .Y(_0392_));
 sg13g2_nor3_1 _1044_ (.A(net322),
    .B(net5),
    .C(\uart.uartArea_uart.commFilter.dcdFilter.io_b ),
    .Y(_0393_));
 sg13g2_a21oi_1 _1045_ (.A1(_0152_),
    .A2(net323),
    .Y(_0065_),
    .B1(_0393_));
 sg13g2_nand3_1 _1046_ (.B(net4),
    .C(\uart.uartArea_uart.commFilter.dsrFilter.io_b ),
    .A(net316),
    .Y(_0394_));
 sg13g2_nor3_1 _1047_ (.A(net316),
    .B(net4),
    .C(\uart.uartArea_uart.commFilter.dsrFilter.io_b ),
    .Y(_0395_));
 sg13g2_a21oi_1 _1048_ (.A1(_0154_),
    .A2(net317),
    .Y(_0066_),
    .B1(_0395_));
 sg13g2_nand3_1 _1049_ (.B(net6),
    .C(\uart.uartArea_uart.commFilter.ctsFilter.io_b ),
    .A(net353),
    .Y(_0396_));
 sg13g2_nor3_1 _1050_ (.A(net353),
    .B(net6),
    .C(\uart.uartArea_uart.commFilter.ctsFilter.io_b ),
    .Y(_0397_));
 sg13g2_a21oi_1 _1051_ (.A1(_0156_),
    .A2(net354),
    .Y(_0067_),
    .B1(_0397_));
 sg13g2_mux2_1 _1052_ (.A0(net363),
    .A1(net7),
    .S(_0372_),
    .X(_0068_));
 sg13g2_mux2_1 _1053_ (.A0(net322),
    .A1(net369),
    .S(_0372_),
    .X(_0069_));
 sg13g2_mux2_1 _1054_ (.A0(net369),
    .A1(net5),
    .S(_0372_),
    .X(_0070_));
 sg13g2_mux2_1 _1055_ (.A0(net316),
    .A1(net351),
    .S(_0372_),
    .X(_0071_));
 sg13g2_mux2_1 _1056_ (.A0(net351),
    .A1(net4),
    .S(_0372_),
    .X(_0072_));
 sg13g2_mux2_1 _1057_ (.A0(net353),
    .A1(net362),
    .S(_0372_),
    .X(_0073_));
 sg13g2_mux2_1 _1058_ (.A0(net362),
    .A1(net6),
    .S(_0372_),
    .X(_0074_));
 sg13g2_nor2_1 _1059_ (.A(net171),
    .B(_0344_),
    .Y(_0075_));
 sg13g2_nor2b_1 _1060_ (.A(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[3] ),
    .B_N(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[2] ),
    .Y(_0398_));
 sg13g2_nand2_1 _1061_ (.Y(_0399_),
    .A(net149),
    .B(_0398_));
 sg13g2_nand2_1 _1062_ (.Y(_0400_),
    .A(net431),
    .B(_0381_));
 sg13g2_and3_1 _1063_ (.X(_0401_),
    .A(net390),
    .B(net175),
    .C(_0381_));
 sg13g2_nand3_1 _1064_ (.B(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[0] ),
    .C(_0381_),
    .A(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[1] ),
    .Y(_0402_));
 sg13g2_nor2_2 _1065_ (.A(_0399_),
    .B(_0402_),
    .Y(_0403_));
 sg13g2_mux2_1 _1066_ (.A0(net282),
    .A1(net186),
    .S(net146),
    .X(_0076_));
 sg13g2_mux2_1 _1067_ (.A0(net284),
    .A1(net185),
    .S(net146),
    .X(_0077_));
 sg13g2_mux2_1 _1068_ (.A0(net291),
    .A1(net184),
    .S(_0403_),
    .X(_0078_));
 sg13g2_mux2_1 _1069_ (.A0(net306),
    .A1(net183),
    .S(net146),
    .X(_0079_));
 sg13g2_mux2_1 _1070_ (.A0(net304),
    .A1(net182),
    .S(net146),
    .X(_0080_));
 sg13g2_mux2_1 _1071_ (.A0(net335),
    .A1(net181),
    .S(net146),
    .X(_0081_));
 sg13g2_mux2_1 _1072_ (.A0(net288),
    .A1(net180),
    .S(net146),
    .X(_0082_));
 sg13g2_mux2_1 _1073_ (.A0(net303),
    .A1(net179),
    .S(net146),
    .X(_0083_));
 sg13g2_mux2_1 _1074_ (.A0(net263),
    .A1(\uart.uartArea_uart.regCtrl.txHolderBit9 ),
    .S(net146),
    .X(_0084_));
 sg13g2_nor3_2 _1075_ (.A(net175),
    .B(_0399_),
    .C(_0400_),
    .Y(_0404_));
 sg13g2_mux2_1 _1076_ (.A0(net275),
    .A1(net186),
    .S(net145),
    .X(_0085_));
 sg13g2_mux2_1 _1077_ (.A0(net253),
    .A1(net185),
    .S(net145),
    .X(_0086_));
 sg13g2_mux2_1 _1078_ (.A0(net273),
    .A1(net184),
    .S(_0404_),
    .X(_0087_));
 sg13g2_mux2_1 _1079_ (.A0(net274),
    .A1(net183),
    .S(net145),
    .X(_0088_));
 sg13g2_mux2_1 _1080_ (.A0(net290),
    .A1(net182),
    .S(net145),
    .X(_0089_));
 sg13g2_mux2_1 _1081_ (.A0(net268),
    .A1(net181),
    .S(net145),
    .X(_0090_));
 sg13g2_mux2_1 _1082_ (.A0(net298),
    .A1(net180),
    .S(net145),
    .X(_0091_));
 sg13g2_mux2_1 _1083_ (.A0(net286),
    .A1(net179),
    .S(net145),
    .X(_0092_));
 sg13g2_mux2_1 _1084_ (.A0(net296),
    .A1(\uart.uartArea_uart.regCtrl.txHolderBit9 ),
    .S(net145),
    .X(_0093_));
 sg13g2_and4_1 _1085_ (.A(net175),
    .B(net149),
    .C(_0383_),
    .D(_0398_),
    .X(_0405_));
 sg13g2_mux2_1 _1086_ (.A0(net329),
    .A1(net186),
    .S(net144),
    .X(_0094_));
 sg13g2_mux2_1 _1087_ (.A0(net289),
    .A1(net185),
    .S(net144),
    .X(_0095_));
 sg13g2_mux2_1 _1088_ (.A0(net319),
    .A1(net184),
    .S(_0405_),
    .X(_0096_));
 sg13g2_mux2_1 _1089_ (.A0(net259),
    .A1(net183),
    .S(net144),
    .X(_0097_));
 sg13g2_mux2_1 _1090_ (.A0(net285),
    .A1(net182),
    .S(net144),
    .X(_0098_));
 sg13g2_mux2_1 _1091_ (.A0(net332),
    .A1(net181),
    .S(net144),
    .X(_0099_));
 sg13g2_mux2_1 _1092_ (.A0(net258),
    .A1(net180),
    .S(net144),
    .X(_0100_));
 sg13g2_mux2_1 _1093_ (.A0(net269),
    .A1(net179),
    .S(net144),
    .X(_0101_));
 sg13g2_mux2_1 _1094_ (.A0(net260),
    .A1(\uart.uartArea_uart.regCtrl.txHolderBit9 ),
    .S(net144),
    .X(_0102_));
 sg13g2_or4_1 _1095_ (.A(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[1] ),
    .B(net175),
    .C(_0382_),
    .D(_0399_),
    .X(_0406_));
 sg13g2_mux2_1 _1096_ (.A0(net186),
    .A1(net352),
    .S(net143),
    .X(_0103_));
 sg13g2_mux2_1 _1097_ (.A0(net185),
    .A1(net359),
    .S(net143),
    .X(_0104_));
 sg13g2_mux2_1 _1098_ (.A0(net184),
    .A1(net337),
    .S(_0406_),
    .X(_0105_));
 sg13g2_mux2_1 _1099_ (.A0(net183),
    .A1(net347),
    .S(net143),
    .X(_0106_));
 sg13g2_mux2_1 _1100_ (.A0(net182),
    .A1(net358),
    .S(net143),
    .X(_0107_));
 sg13g2_mux2_1 _1101_ (.A0(net181),
    .A1(net357),
    .S(net143),
    .X(_0108_));
 sg13g2_mux2_1 _1102_ (.A0(net180),
    .A1(net356),
    .S(net143),
    .X(_0109_));
 sg13g2_mux2_1 _1103_ (.A0(net179),
    .A1(net364),
    .S(net143),
    .X(_0110_));
 sg13g2_mux2_1 _1104_ (.A0(\uart.uartArea_uart.regCtrl.txHolderBit9 ),
    .A1(net360),
    .S(net143),
    .X(_0111_));
 sg13g2_nor3_2 _1105_ (.A(net148),
    .B(_0380_),
    .C(_0402_),
    .Y(_0407_));
 sg13g2_mux2_1 _1106_ (.A0(net325),
    .A1(net186),
    .S(net142),
    .X(_0112_));
 sg13g2_mux2_1 _1107_ (.A0(net280),
    .A1(net185),
    .S(net142),
    .X(_0113_));
 sg13g2_mux2_1 _1108_ (.A0(net276),
    .A1(net184),
    .S(_0407_),
    .X(_0114_));
 sg13g2_mux2_1 _1109_ (.A0(net295),
    .A1(net183),
    .S(net142),
    .X(_0115_));
 sg13g2_mux2_1 _1110_ (.A0(net294),
    .A1(net182),
    .S(net142),
    .X(_0116_));
 sg13g2_mux2_1 _1111_ (.A0(net336),
    .A1(net181),
    .S(net142),
    .X(_0117_));
 sg13g2_mux2_1 _1112_ (.A0(net305),
    .A1(net180),
    .S(net142),
    .X(_0118_));
 sg13g2_mux2_1 _1113_ (.A0(net311),
    .A1(net179),
    .S(net142),
    .X(_0119_));
 sg13g2_mux2_1 _1114_ (.A0(net338),
    .A1(\uart.uartArea_uart.regCtrl.txHolderBit9 ),
    .S(net142),
    .X(_0120_));
 sg13g2_nor4_2 _1115_ (.A(net175),
    .B(net148),
    .C(_0380_),
    .Y(_0408_),
    .D(_0400_));
 sg13g2_mux2_1 _1116_ (.A0(net321),
    .A1(net186),
    .S(net141),
    .X(_0121_));
 sg13g2_mux2_1 _1117_ (.A0(net293),
    .A1(net185),
    .S(net141),
    .X(_0122_));
 sg13g2_mux2_1 _1118_ (.A0(net262),
    .A1(net184),
    .S(net141),
    .X(_0123_));
 sg13g2_mux2_1 _1119_ (.A0(net300),
    .A1(net183),
    .S(net141),
    .X(_0124_));
 sg13g2_mux2_1 _1120_ (.A0(net340),
    .A1(net182),
    .S(_0408_),
    .X(_0125_));
 sg13g2_mux2_1 _1121_ (.A0(net312),
    .A1(net181),
    .S(net141),
    .X(_0126_));
 sg13g2_mux2_1 _1122_ (.A0(net320),
    .A1(net180),
    .S(net141),
    .X(_0127_));
 sg13g2_mux2_1 _1123_ (.A0(net255),
    .A1(net179),
    .S(net141),
    .X(_0128_));
 sg13g2_mux2_1 _1124_ (.A0(net333),
    .A1(\uart.uartArea_uart.regCtrl.txHolderBit9 ),
    .S(net141),
    .X(_0129_));
 sg13g2_o21ai_1 _1125_ (.B1(net149),
    .Y(_0409_),
    .A1(net175),
    .A2(_0381_));
 sg13g2_a21oi_1 _1126_ (.A1(net175),
    .A2(_0381_),
    .Y(_0130_),
    .B1(_0409_));
 sg13g2_a21oi_1 _1127_ (.A1(net175),
    .A2(_0381_),
    .Y(_0410_),
    .B1(net390));
 sg13g2_nor3_1 _1128_ (.A(net148),
    .B(_0401_),
    .C(net391),
    .Y(_0131_));
 sg13g2_a21oi_1 _1129_ (.A1(net395),
    .A2(_0401_),
    .Y(_0411_),
    .B1(net148));
 sg13g2_nor2_1 _1130_ (.A(net395),
    .B(_0401_),
    .Y(_0412_));
 sg13g2_nor2b_1 _1131_ (.A(_0412_),
    .B_N(_0411_),
    .Y(_0132_));
 sg13g2_and2_1 _1132_ (.A(net256),
    .B(_0411_),
    .X(_0133_));
 sg13g2_o21ai_1 _1133_ (.B1(net149),
    .Y(_0413_),
    .A1(\uart.uartArea_uart.txFifo.count[0] ),
    .A2(_0381_));
 sg13g2_a21oi_1 _1134_ (.A1(_0158_),
    .A2(_0381_),
    .Y(_0134_),
    .B1(_0413_));
 sg13g2_a21oi_1 _1135_ (.A1(\uart.uartArea_uart.txFifo.count[0] ),
    .A2(_0334_),
    .Y(_0414_),
    .B1(net370));
 sg13g2_and3_1 _1136_ (.X(_0415_),
    .A(net370),
    .B(\uart.uartArea_uart.txFifo.count[0] ),
    .C(_0334_));
 sg13g2_nor3_1 _1137_ (.A(_0338_),
    .B(net371),
    .C(_0415_),
    .Y(_0135_));
 sg13g2_nand2_1 _1138_ (.Y(_0416_),
    .A(net422),
    .B(_0415_));
 sg13g2_o21ai_1 _1139_ (.B1(net149),
    .Y(_0417_),
    .A1(net422),
    .A2(_0415_));
 sg13g2_nor2b_1 _1140_ (.A(net423),
    .B_N(_0416_),
    .Y(_0136_));
 sg13g2_o21ai_1 _1141_ (.B1(net149),
    .Y(_0418_),
    .A1(_0157_),
    .A2(_0416_));
 sg13g2_a21oi_1 _1142_ (.A1(_0157_),
    .A2(_0416_),
    .Y(_0137_),
    .B1(_0418_));
 sg13g2_nand3b_1 _1143_ (.B(net157),
    .C(net3),
    .Y(_0419_),
    .A_N(net2));
 sg13g2_o21ai_1 _1144_ (.B1(net168),
    .Y(_0420_),
    .A1(\uart.uartArea_uart.commFilter.ctsFilter.io_o ),
    .A2(_0419_));
 sg13g2_a21oi_1 _1145_ (.A1(_0155_),
    .A2(_0419_),
    .Y(_0138_),
    .B1(_0420_));
 sg13g2_o21ai_1 _1146_ (.B1(net168),
    .Y(_0421_),
    .A1(\uart.uartArea_uart.commFilter.dsrFilter.io_o ),
    .A2(_0419_));
 sg13g2_a21oi_1 _1147_ (.A1(_0153_),
    .A2(_0419_),
    .Y(_0139_),
    .B1(_0421_));
 sg13g2_o21ai_1 _1148_ (.B1(net168),
    .Y(_0422_),
    .A1(\uart.uartArea_uart.commFilter.dcdFilter.io_o ),
    .A2(_0419_));
 sg13g2_a21oi_1 _1149_ (.A1(_0151_),
    .A2(_0419_),
    .Y(_0140_),
    .B1(_0422_));
 sg13g2_nor4_2 _1150_ (.A(_0183_),
    .B(_0192_),
    .C(_0265_),
    .Y(_0423_),
    .D(_0344_));
 sg13g2_o21ai_1 _1151_ (.B1(net149),
    .Y(_0424_),
    .A1(net404),
    .A2(_0423_));
 sg13g2_a21oi_1 _1152_ (.A1(net404),
    .A2(_0423_),
    .Y(_0141_),
    .B1(_0424_));
 sg13g2_a21oi_1 _1153_ (.A1(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[0] ),
    .A2(_0423_),
    .Y(_0425_),
    .B1(net373));
 sg13g2_nor2b_1 _1154_ (.A(_0197_),
    .B_N(_0423_),
    .Y(_0426_));
 sg13g2_nor3_1 _1155_ (.A(net148),
    .B(net374),
    .C(_0426_),
    .Y(_0142_));
 sg13g2_a21oi_1 _1156_ (.A1(net417),
    .A2(_0426_),
    .Y(_0427_),
    .B1(net148));
 sg13g2_nor2_1 _1157_ (.A(net417),
    .B(_0426_),
    .Y(_0428_));
 sg13g2_nor2b_1 _1158_ (.A(net418),
    .B_N(_0427_),
    .Y(_0143_));
 sg13g2_and2_1 _1159_ (.A(net307),
    .B(_0427_),
    .X(_0144_));
 sg13g2_nor2_1 _1160_ (.A(\uart.uartArea_uart.rxFifo.count[0] ),
    .B(_0423_),
    .Y(_0429_));
 sg13g2_nor2b_1 _1161_ (.A(net235),
    .B_N(_0423_),
    .Y(_0430_));
 sg13g2_nor3_1 _1162_ (.A(_0338_),
    .B(_0429_),
    .C(_0430_),
    .Y(_0145_));
 sg13g2_nand2b_1 _1163_ (.Y(_0431_),
    .B(_0423_),
    .A_N(\uart.uartArea_uart.rxFifo.count[0] ));
 sg13g2_xor2_1 _1164_ (.B(_0431_),
    .A(net410),
    .X(_0432_));
 sg13g2_nor2_1 _1165_ (.A(net148),
    .B(net411),
    .Y(_0146_));
 sg13g2_o21ai_1 _1166_ (.B1(net348),
    .Y(_0433_),
    .A1(\uart.uartArea_uart.rxFifo.count[1] ),
    .A2(_0431_));
 sg13g2_nand2_1 _1167_ (.Y(_0434_),
    .A(_0240_),
    .B(_0423_));
 sg13g2_a21oi_1 _1168_ (.A1(net349),
    .A2(_0434_),
    .Y(_0147_),
    .B1(net148));
 sg13g2_and3_1 _1169_ (.X(_0148_),
    .A(net326),
    .B(net150),
    .C(_0434_));
 sg13g2_nand2_1 _1170_ (.Y(_0435_),
    .A(_0155_),
    .B(net379));
 sg13g2_a21oi_1 _1171_ (.A1(net367),
    .A2(_0156_),
    .Y(_0436_),
    .B1(\uart.uartArea_uart.regCtrl.regModemCtrlChanged[0] ));
 sg13g2_a21oi_1 _1172_ (.A1(_0435_),
    .A2(_0436_),
    .Y(_0149_),
    .B1(net171));
 sg13g2_dfrbp_1 _1173_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net34),
    .D(net1),
    .Q_N(_0576_),
    .Q(rst_n_sync));
 sg13g2_dfrbp_1 _1174_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net95),
    .D(net232),
    .Q_N(_0004_),
    .Q(\uart.uartArea_uart.uartClocking_1.divisorCtr[0] ));
 sg13g2_dfrbp_1 _1175_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net94),
    .D(_0007_),
    .Q_N(_0575_),
    .Q(\uart.uartArea_uart.uartClocking_1.divisorCtr[1] ));
 sg13g2_dfrbp_1 _1176_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net93),
    .D(_0008_),
    .Q_N(_0574_),
    .Q(\uart.uartArea_uart.uartClocking_1.divisorCtr[2] ));
 sg13g2_dfrbp_1 _1177_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net92),
    .D(net267),
    .Q_N(_0573_),
    .Q(\uart.uartArea_uart.uartClocking_1.divisorCtr[3] ));
 sg13g2_dfrbp_1 _1178_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net91),
    .D(_0010_),
    .Q_N(_0572_),
    .Q(\uart.uartArea_uart.uartClocking_1.divisorCtr[4] ));
 sg13g2_dfrbp_1 _1179_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net90),
    .D(_0011_),
    .Q_N(_0571_),
    .Q(\uart.uartArea_uart.uartClocking_1.divisorCtr[5] ));
 sg13g2_dfrbp_1 _1180_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net89),
    .D(_0012_),
    .Q_N(_0570_),
    .Q(\uart.uartArea_uart.uartClocking_1.divisorCtr[6] ));
 sg13g2_dfrbp_1 _1181_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net88),
    .D(net251),
    .Q_N(_0569_),
    .Q(\uart.uartArea_uart.uartClocking_1.divisorCtr[7] ));
 sg13g2_dfrbp_1 _1182_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net87),
    .D(net378),
    .Q_N(_0568_),
    .Q(\uart.uartArea_uart.regCtrl.regModemCtrlChanged[1] ));
 sg13g2_dfrbp_1 _1183_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net35),
    .D(net272),
    .Q_N(_0577_),
    .Q(\uart.uartArea_uart.regCtrl.regModemCtrlChanged[2] ));
 sg13g2_dfrbp_1 _1184_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net36),
    .D(\uart.resetCommandStrobe ),
    .Q_N(_0578_),
    .Q(\uart.resetCommandUnit_1.ff ));
 sg13g2_dfrbp_1 _1185_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net65),
    .D(\uart.resetCommandUnit_1.async.area_io_q ),
    .Q_N(_0579_),
    .Q(\uart.resetCommandUnit_1.reg1 ));
 sg13g2_dfrbp_1 _1186_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net85),
    .D(net228),
    .Q_N(_0567_),
    .Q(\uart.resetCommandUnit_1.async.area_io_r ));
 sg13g2_dfrbp_1 _1187_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net83),
    .D(net245),
    .Q_N(_0566_),
    .Q(\uart.uartArea_uart.regCtrl.txOverrun ));
 sg13g2_dfrbp_1 _1188_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net81),
    .D(_0017_),
    .Q_N(_0565_),
    .Q(\uart.uartArea_uart.regCtrl.txHolderBit9 ));
 sg13g2_dfrbp_1 _1189_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net80),
    .D(_0018_),
    .Q_N(_0564_),
    .Q(\uart.uartArea_uart.regCtrl.regFifoTxEnable ));
 sg13g2_dfrbp_1 _1190_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net78),
    .D(_0019_),
    .Q_N(_0563_),
    .Q(\uart.uartArea_uart.regCtrl.regFifoRxEnable ));
 sg13g2_dfrbp_1 _1191_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net76),
    .D(net343),
    .Q_N(_0562_),
    .Q(\uart.uartArea_uart.regCtrl.regModemCtrlChanged[3] ));
 sg13g2_dfrbp_1 _1192_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net74),
    .D(_0021_),
    .Q_N(_0561_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[0] ));
 sg13g2_dfrbp_1 _1193_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net72),
    .D(_0022_),
    .Q_N(_0560_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[1] ));
 sg13g2_dfrbp_1 _1194_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net70),
    .D(_0023_),
    .Q_N(_0559_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[2] ));
 sg13g2_dfrbp_1 _1195_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net68),
    .D(_0024_),
    .Q_N(_0558_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[3] ));
 sg13g2_dfrbp_1 _1196_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net66),
    .D(_0025_),
    .Q_N(_0557_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[4] ));
 sg13g2_dfrbp_1 _1197_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net63),
    .D(_0026_),
    .Q_N(_0556_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[5] ));
 sg13g2_dfrbp_1 _1198_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net61),
    .D(_0027_),
    .Q_N(_0555_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[6] ));
 sg13g2_dfrbp_1 _1199_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net59),
    .D(_0028_),
    .Q_N(_0554_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptControl[0] ));
 sg13g2_dfrbp_1 _1200_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net57),
    .D(_0029_),
    .Q_N(_0553_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptControl[1] ));
 sg13g2_dfrbp_1 _1201_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net55),
    .D(_0030_),
    .Q_N(_0552_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptControl[2] ));
 sg13g2_dfrbp_1 _1202_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net53),
    .D(_0031_),
    .Q_N(_0551_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptControl[3] ));
 sg13g2_dfrbp_1 _1203_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net51),
    .D(_0032_),
    .Q_N(_0550_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptControl[4] ));
 sg13g2_dfrbp_1 _1204_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net49),
    .D(_0033_),
    .Q_N(_0549_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptControl[5] ));
 sg13g2_dfrbp_1 _1205_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net47),
    .D(_0034_),
    .Q_N(_0548_),
    .Q(\uart.uartArea_uart.regCtrl.io_regInterruptControl[6] ));
 sg13g2_dfrbp_1 _1206_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net45),
    .D(_0035_),
    .Q_N(_0547_),
    .Q(\uart.uartArea_uart.regCtrl.reg007[0] ));
 sg13g2_dfrbp_1 _1207_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net43),
    .D(_0036_),
    .Q_N(_0546_),
    .Q(\uart.uartArea_uart.regCtrl.reg007[1] ));
 sg13g2_dfrbp_1 _1208_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net41),
    .D(_0037_),
    .Q_N(_0545_),
    .Q(\uart.uartArea_uart.regCtrl.reg007[2] ));
 sg13g2_dfrbp_1 _1209_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net39),
    .D(_0038_),
    .Q_N(_0544_),
    .Q(\uart.uartArea_uart.regCtrl.reg007[3] ));
 sg13g2_dfrbp_1 _1210_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net37),
    .D(_0039_),
    .Q_N(_0543_),
    .Q(\uart.uartArea_uart.regCtrl.reg007[4] ));
 sg13g2_dfrbp_1 _1211_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net32),
    .D(_0040_),
    .Q_N(_0542_),
    .Q(\uart.uartArea_uart.regCtrl.reg007[5] ));
 sg13g2_dfrbp_1 _1212_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net30),
    .D(_0041_),
    .Q_N(_0541_),
    .Q(\uart.uartArea_uart.regCtrl.reg007[6] ));
 sg13g2_dfrbp_1 _1213_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net28),
    .D(_0042_),
    .Q_N(_0540_),
    .Q(\uart.uartArea_uart.regCtrl.reg007[7] ));
 sg13g2_dfrbp_1 _1214_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net219),
    .D(_0043_),
    .Q_N(_0580_),
    .Q(\uart.uartArea_uart.commFilter.riFilter.io_c ));
 sg13g2_dfrbp_1 _1215_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net26),
    .D(net230),
    .Q_N(_0539_),
    .Q(\uart.uartArea_uart.regCtrl.riSignalNext ));
 sg13g2_dfrbp_1 _1216_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net25),
    .D(_0044_),
    .Q_N(_0538_),
    .Q(\uart.uartArea_uart.busCtrl.io_regAddr[0] ));
 sg13g2_dfrbp_1 _1217_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net24),
    .D(_0045_),
    .Q_N(_0537_),
    .Q(\uart.uartArea_uart.busCtrl.io_regAddr[1] ));
 sg13g2_dfrbp_1 _1218_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net23),
    .D(_0046_),
    .Q_N(_0536_),
    .Q(\uart.uartArea_uart.busCtrl.io_regAddr[2] ));
 sg13g2_dfrbp_1 _1219_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net218),
    .D(_0047_),
    .Q_N(_0535_),
    .Q(\uart.uartArea_uart.busCtrl.io_regAddr[3] ));
 sg13g2_dfrbp_1 _1220_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net217),
    .D(_0048_),
    .Q_N(_0000_),
    .Q(\uart.uartArea_uart.busCtrl.io_regAddr[4] ));
 sg13g2_dfrbp_1 _1221_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net216),
    .D(_0049_),
    .Q_N(_0534_),
    .Q(\uart.uartArea_uart.busCtrl.lastWasWrite ));
 sg13g2_dfrbp_1 _1222_ (.CLK(net224),
    .RESET_B(net215),
    .D(_0050_),
    .Q_N(_0533_),
    .Q(\uart.resetCommandUnit_1.async.area_io_q ));
 sg13g2_dfrbp_1 _1223_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net213),
    .D(_0051_),
    .Q_N(_0532_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_14[0] ));
 sg13g2_dfrbp_1 _1224_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net212),
    .D(_0052_),
    .Q_N(_0531_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_14[1] ));
 sg13g2_dfrbp_1 _1225_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net211),
    .D(_0053_),
    .Q_N(_0530_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_14[2] ));
 sg13g2_dfrbp_1 _1226_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net210),
    .D(_0054_),
    .Q_N(_0529_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_14[3] ));
 sg13g2_dfrbp_1 _1227_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net209),
    .D(net366),
    .Q_N(_0528_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_14[4] ));
 sg13g2_dfrbp_1 _1228_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net208),
    .D(_0056_),
    .Q_N(_0527_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_14[5] ));
 sg13g2_dfrbp_1 _1229_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net207),
    .D(_0057_),
    .Q_N(_0526_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_14[6] ));
 sg13g2_dfrbp_1 _1230_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net206),
    .D(_0058_),
    .Q_N(_0525_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_14[7] ));
 sg13g2_dfrbp_1 _1231_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net205),
    .D(net279),
    .Q_N(_0524_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_14[8] ));
 sg13g2_dfrbp_1 _1232_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net204),
    .D(net248),
    .Q_N(_0003_),
    .Q(\uart.uartArea_uart.uartClocking_1.bitCtr[0] ));
 sg13g2_dfrbp_1 _1233_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net202),
    .D(net386),
    .Q_N(_0523_),
    .Q(\uart.uartArea_uart.uartClocking_1.bitCtr[1] ));
 sg13g2_dfrbp_1 _1234_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net200),
    .D(net315),
    .Q_N(_0522_),
    .Q(\uart.uartArea_uart.uartClocking_1.bitCtr[2] ));
 sg13g2_dfrbp_1 _1235_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net198),
    .D(_0063_),
    .Q_N(_0521_),
    .Q(\uart.uartArea_uart.uartClocking_1.bitCtr[3] ));
 sg13g2_dfrbp_1 _1236_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net196),
    .D(net346),
    .Q_N(_0520_),
    .Q(\uart.uartArea_uart.commFilter.io_ttl_ri ));
 sg13g2_dfrbp_1 _1237_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net194),
    .D(net324),
    .Q_N(_0519_),
    .Q(\uart.uartArea_uart.commFilter.dcdFilter.io_o ));
 sg13g2_dfrbp_1 _1238_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net192),
    .D(net318),
    .Q_N(_0518_),
    .Q(\uart.uartArea_uart.commFilter.dsrFilter.io_o ));
 sg13g2_dfrbp_1 _1239_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net190),
    .D(net355),
    .Q_N(_0517_),
    .Q(\uart.uartArea_uart.commFilter.ctsFilter.io_o ));
 sg13g2_dfrbp_1 _1240_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net188),
    .D(_0068_),
    .Q_N(_0516_),
    .Q(\uart.uartArea_uart.commFilter.riFilter.io_b ));
 sg13g2_dfrbp_1 _1241_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net140),
    .D(_0069_),
    .Q_N(_0515_),
    .Q(\uart.uartArea_uart.commFilter.dcdFilter.io_c ));
 sg13g2_dfrbp_1 _1242_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net139),
    .D(_0070_),
    .Q_N(_0514_),
    .Q(\uart.uartArea_uart.commFilter.dcdFilter.io_b ));
 sg13g2_dfrbp_1 _1243_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net138),
    .D(_0071_),
    .Q_N(_0513_),
    .Q(\uart.uartArea_uart.commFilter.dsrFilter.io_c ));
 sg13g2_dfrbp_1 _1244_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net137),
    .D(_0072_),
    .Q_N(_0512_),
    .Q(\uart.uartArea_uart.commFilter.dsrFilter.io_b ));
 sg13g2_dfrbp_1 _1245_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net136),
    .D(_0073_),
    .Q_N(_0511_),
    .Q(\uart.uartArea_uart.commFilter.ctsFilter.io_c ));
 sg13g2_dfrbp_1 _1246_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net135),
    .D(_0074_),
    .Q_N(_0510_),
    .Q(\uart.uartArea_uart.commFilter.ctsFilter.io_b ));
 sg13g2_dfrbp_1 _1247_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net134),
    .D(_0075_),
    .Q_N(_0509_),
    .Q(\uart.uartArea_uart.busCtrl.oe ));
 sg13g2_dfrbp_1 _1248_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net133),
    .D(_0076_),
    .Q_N(_0508_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_8[0] ));
 sg13g2_dfrbp_1 _1249_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net132),
    .D(_0077_),
    .Q_N(_0507_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_8[1] ));
 sg13g2_dfrbp_1 _1250_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net131),
    .D(net292),
    .Q_N(_0506_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_8[2] ));
 sg13g2_dfrbp_1 _1251_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net130),
    .D(_0079_),
    .Q_N(_0505_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_8[3] ));
 sg13g2_dfrbp_1 _1252_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net129),
    .D(_0080_),
    .Q_N(_0504_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_8[4] ));
 sg13g2_dfrbp_1 _1253_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net128),
    .D(_0081_),
    .Q_N(_0503_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_8[5] ));
 sg13g2_dfrbp_1 _1254_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net127),
    .D(_0082_),
    .Q_N(_0502_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_8[6] ));
 sg13g2_dfrbp_1 _1255_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net126),
    .D(_0083_),
    .Q_N(_0501_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_8[7] ));
 sg13g2_dfrbp_1 _1256_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net125),
    .D(net264),
    .Q_N(_0500_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_8[8] ));
 sg13g2_dfrbp_1 _1257_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net124),
    .D(_0085_),
    .Q_N(_0499_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_9[0] ));
 sg13g2_dfrbp_1 _1258_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net123),
    .D(_0086_),
    .Q_N(_0498_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_9[1] ));
 sg13g2_dfrbp_1 _1259_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net122),
    .D(_0087_),
    .Q_N(_0497_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_9[2] ));
 sg13g2_dfrbp_1 _1260_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net121),
    .D(_0088_),
    .Q_N(_0496_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_9[3] ));
 sg13g2_dfrbp_1 _1261_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net120),
    .D(_0089_),
    .Q_N(_0495_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_9[4] ));
 sg13g2_dfrbp_1 _1262_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net119),
    .D(_0090_),
    .Q_N(_0494_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_9[5] ));
 sg13g2_dfrbp_1 _1263_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net118),
    .D(_0091_),
    .Q_N(_0493_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_9[6] ));
 sg13g2_dfrbp_1 _1264_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net117),
    .D(_0092_),
    .Q_N(_0492_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_9[7] ));
 sg13g2_dfrbp_1 _1265_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net116),
    .D(net297),
    .Q_N(_0491_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_9[8] ));
 sg13g2_dfrbp_1 _1266_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net115),
    .D(_0094_),
    .Q_N(_0490_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_10[0] ));
 sg13g2_dfrbp_1 _1267_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net114),
    .D(_0095_),
    .Q_N(_0489_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_10[1] ));
 sg13g2_dfrbp_1 _1268_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net113),
    .D(_0096_),
    .Q_N(_0488_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_10[2] ));
 sg13g2_dfrbp_1 _1269_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net112),
    .D(_0097_),
    .Q_N(_0487_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_10[3] ));
 sg13g2_dfrbp_1 _1270_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net111),
    .D(_0098_),
    .Q_N(_0486_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_10[4] ));
 sg13g2_dfrbp_1 _1271_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net110),
    .D(_0099_),
    .Q_N(_0485_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_10[5] ));
 sg13g2_dfrbp_1 _1272_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net109),
    .D(_0100_),
    .Q_N(_0484_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_10[6] ));
 sg13g2_dfrbp_1 _1273_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net108),
    .D(_0101_),
    .Q_N(_0483_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_10[7] ));
 sg13g2_dfrbp_1 _1274_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net107),
    .D(net261),
    .Q_N(_0482_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_10[8] ));
 sg13g2_dfrbp_1 _1275_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net106),
    .D(_0103_),
    .Q_N(_0481_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_11[0] ));
 sg13g2_dfrbp_1 _1276_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net105),
    .D(_0104_),
    .Q_N(_0480_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_11[1] ));
 sg13g2_dfrbp_1 _1277_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net104),
    .D(_0105_),
    .Q_N(_0479_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_11[2] ));
 sg13g2_dfrbp_1 _1278_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net103),
    .D(_0106_),
    .Q_N(_0478_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_11[3] ));
 sg13g2_dfrbp_1 _1279_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net102),
    .D(_0107_),
    .Q_N(_0477_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_11[4] ));
 sg13g2_dfrbp_1 _1280_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net101),
    .D(_0108_),
    .Q_N(_0476_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_11[5] ));
 sg13g2_dfrbp_1 _1281_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net100),
    .D(_0109_),
    .Q_N(_0475_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_11[6] ));
 sg13g2_dfrbp_1 _1282_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net99),
    .D(_0110_),
    .Q_N(_0474_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_11[7] ));
 sg13g2_dfrbp_1 _1283_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net98),
    .D(net361),
    .Q_N(_0473_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_11[8] ));
 sg13g2_dfrbp_1 _1284_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net97),
    .D(_0112_),
    .Q_N(_0472_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_12[0] ));
 sg13g2_dfrbp_1 _1285_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net96),
    .D(_0113_),
    .Q_N(_0471_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_12[1] ));
 sg13g2_dfrbp_1 _1286_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net86),
    .D(net277),
    .Q_N(_0470_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_12[2] ));
 sg13g2_dfrbp_1 _1287_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net84),
    .D(_0115_),
    .Q_N(_0469_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_12[3] ));
 sg13g2_dfrbp_1 _1288_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net82),
    .D(_0116_),
    .Q_N(_0468_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_12[4] ));
 sg13g2_dfrbp_1 _1289_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net79),
    .D(_0117_),
    .Q_N(_0467_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_12[5] ));
 sg13g2_dfrbp_1 _1290_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net77),
    .D(_0118_),
    .Q_N(_0466_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_12[6] ));
 sg13g2_dfrbp_1 _1291_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net75),
    .D(_0119_),
    .Q_N(_0465_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_12[7] ));
 sg13g2_dfrbp_1 _1292_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net73),
    .D(net339),
    .Q_N(_0464_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_12[8] ));
 sg13g2_dfrbp_1 _1293_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net71),
    .D(_0121_),
    .Q_N(_0463_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_13[0] ));
 sg13g2_dfrbp_1 _1294_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net69),
    .D(_0122_),
    .Q_N(_0462_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_13[1] ));
 sg13g2_dfrbp_1 _1295_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net67),
    .D(_0123_),
    .Q_N(_0461_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_13[2] ));
 sg13g2_dfrbp_1 _1296_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net64),
    .D(_0124_),
    .Q_N(_0460_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_13[3] ));
 sg13g2_dfrbp_1 _1297_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net62),
    .D(_0125_),
    .Q_N(_0459_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_13[4] ));
 sg13g2_dfrbp_1 _1298_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net60),
    .D(_0126_),
    .Q_N(_0458_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_13[5] ));
 sg13g2_dfrbp_1 _1299_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net58),
    .D(_0127_),
    .Q_N(_0457_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_13[6] ));
 sg13g2_dfrbp_1 _1300_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net56),
    .D(_0128_),
    .Q_N(_0456_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_13[7] ));
 sg13g2_dfrbp_1 _1301_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net54),
    .D(net334),
    .Q_N(_0455_),
    .Q(\uart.uartArea_uart.sharedFifo.fifoRegs_13[8] ));
 sg13g2_dfrbp_1 _1302_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net52),
    .D(_0130_),
    .Q_N(_0454_),
    .Q(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[0] ));
 sg13g2_dfrbp_1 _1303_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net48),
    .D(_0131_),
    .Q_N(_0453_),
    .Q(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[1] ));
 sg13g2_dfrbp_1 _1304_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net44),
    .D(_0132_),
    .Q_N(_0452_),
    .Q(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[2] ));
 sg13g2_dfrbp_1 _1305_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net40),
    .D(net257),
    .Q_N(_0451_),
    .Q(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[3] ));
 sg13g2_dfrbp_1 _1306_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net33),
    .D(net234),
    .Q_N(_0002_),
    .Q(\uart.uartArea_uart.txFifo.count[0] ));
 sg13g2_dfrbp_1 _1307_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net29),
    .D(net372),
    .Q_N(_0450_),
    .Q(\uart.uartArea_uart.txFifo.count[1] ));
 sg13g2_dfrbp_1 _1308_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net214),
    .D(_0136_),
    .Q_N(_0449_),
    .Q(\uart.uartArea_uart.txFifo.count[2] ));
 sg13g2_dfrbp_1 _1309_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net201),
    .D(net416),
    .Q_N(_0448_),
    .Q(\uart.uartArea_uart.txFifo.count[3] ));
 sg13g2_dfrbp_1 _1310_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net197),
    .D(net368),
    .Q_N(_0447_),
    .Q(\uart.uartArea_uart.regCtrl.regModemCtrlHistory[0] ));
 sg13g2_dfrbp_1 _1311_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net193),
    .D(net302),
    .Q_N(_0446_),
    .Q(\uart.uartArea_uart.regCtrl.regModemCtrlHistory[1] ));
 sg13g2_dfrbp_1 _1312_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net189),
    .D(net331),
    .Q_N(_0445_),
    .Q(\uart.uartArea_uart.regCtrl.regModemCtrlHistory[3] ));
 sg13g2_dfrbp_1 _1313_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net46),
    .D(_0141_),
    .Q_N(_0444_),
    .Q(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[0] ));
 sg13g2_dfrbp_1 _1314_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net38),
    .D(_0142_),
    .Q_N(_0443_),
    .Q(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[1] ));
 sg13g2_dfrbp_1 _1315_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net27),
    .D(_0143_),
    .Q_N(_0442_),
    .Q(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[2] ));
 sg13g2_dfrbp_1 _1316_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net199),
    .D(net308),
    .Q_N(_0441_),
    .Q(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[3] ));
 sg13g2_dfrbp_1 _1317_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net191),
    .D(net236),
    .Q_N(_0001_),
    .Q(\uart.uartArea_uart.rxFifo.count[0] ));
 sg13g2_dfrbp_1 _1318_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net42),
    .D(_0146_),
    .Q_N(_0440_),
    .Q(\uart.uartArea_uart.rxFifo.count[1] ));
 sg13g2_dfrbp_1 _1319_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net203),
    .D(net350),
    .Q_N(_0439_),
    .Q(\uart.uartArea_uart.rxFifo.count[2] ));
 sg13g2_dfrbp_1 _1320_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net50),
    .D(_0148_),
    .Q_N(_0438_),
    .Q(\uart.uartArea_uart.rxFifo.count[3] ));
 sg13g2_dfrbp_1 _1321_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net31),
    .D(net380),
    .Q_N(_0581_),
    .Q(\uart.uartArea_uart.regCtrl.regModemCtrlChanged[0] ));
 sg13g2_dfrbp_1 _1322_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net195),
    .D(net229),
    .Q_N(_0437_),
    .Q(\uart.resetCommandUnit_1.io_resetIn ));
 sg13g2_tiehi _1217__24 (.L_HI(net24));
 sg13g2_tiehi _1216__25 (.L_HI(net25));
 sg13g2_tiehi _1215__26 (.L_HI(net26));
 sg13g2_tiehi _1315__27 (.L_HI(net27));
 sg13g2_tiehi _1213__28 (.L_HI(net28));
 sg13g2_tiehi _1307__29 (.L_HI(net29));
 sg13g2_tiehi _1212__30 (.L_HI(net30));
 sg13g2_tiehi _1321__31 (.L_HI(net31));
 sg13g2_tiehi _1211__32 (.L_HI(net32));
 sg13g2_tiehi _1306__33 (.L_HI(net33));
 sg13g2_tiehi _1173__34 (.L_HI(net34));
 sg13g2_tiehi _1183__35 (.L_HI(net35));
 sg13g2_tiehi _1184__36 (.L_HI(net36));
 sg13g2_tiehi _1210__37 (.L_HI(net37));
 sg13g2_tiehi _1314__38 (.L_HI(net38));
 sg13g2_tiehi _1209__39 (.L_HI(net39));
 sg13g2_tiehi _1305__40 (.L_HI(net40));
 sg13g2_tiehi _1208__41 (.L_HI(net41));
 sg13g2_tiehi _1318__42 (.L_HI(net42));
 sg13g2_tiehi _1207__43 (.L_HI(net43));
 sg13g2_tiehi _1304__44 (.L_HI(net44));
 sg13g2_tiehi _1206__45 (.L_HI(net45));
 sg13g2_tiehi _1313__46 (.L_HI(net46));
 sg13g2_tiehi _1205__47 (.L_HI(net47));
 sg13g2_tiehi _1303__48 (.L_HI(net48));
 sg13g2_tiehi _1204__49 (.L_HI(net49));
 sg13g2_tiehi _1320__50 (.L_HI(net50));
 sg13g2_tiehi _1203__51 (.L_HI(net51));
 sg13g2_tiehi _1302__52 (.L_HI(net52));
 sg13g2_tiehi _1202__53 (.L_HI(net53));
 sg13g2_tiehi _1301__54 (.L_HI(net54));
 sg13g2_tiehi _1201__55 (.L_HI(net55));
 sg13g2_tiehi _1300__56 (.L_HI(net56));
 sg13g2_tiehi _1200__57 (.L_HI(net57));
 sg13g2_tiehi _1299__58 (.L_HI(net58));
 sg13g2_tiehi _1199__59 (.L_HI(net59));
 sg13g2_tiehi _1298__60 (.L_HI(net60));
 sg13g2_tiehi _1198__61 (.L_HI(net61));
 sg13g2_tiehi _1297__62 (.L_HI(net62));
 sg13g2_tiehi _1197__63 (.L_HI(net63));
 sg13g2_tiehi _1296__64 (.L_HI(net64));
 sg13g2_tiehi _1185__65 (.L_HI(net65));
 sg13g2_tiehi _1196__66 (.L_HI(net66));
 sg13g2_tiehi _1295__67 (.L_HI(net67));
 sg13g2_tiehi _1195__68 (.L_HI(net68));
 sg13g2_tiehi _1294__69 (.L_HI(net69));
 sg13g2_tiehi _1194__70 (.L_HI(net70));
 sg13g2_tiehi _1293__71 (.L_HI(net71));
 sg13g2_tiehi _1193__72 (.L_HI(net72));
 sg13g2_tiehi _1292__73 (.L_HI(net73));
 sg13g2_tiehi _1192__74 (.L_HI(net74));
 sg13g2_tiehi _1291__75 (.L_HI(net75));
 sg13g2_tiehi _1191__76 (.L_HI(net76));
 sg13g2_tiehi _1290__77 (.L_HI(net77));
 sg13g2_tiehi _1190__78 (.L_HI(net78));
 sg13g2_tiehi _1289__79 (.L_HI(net79));
 sg13g2_tiehi _1189__80 (.L_HI(net80));
 sg13g2_tiehi _1188__81 (.L_HI(net81));
 sg13g2_tiehi _1288__82 (.L_HI(net82));
 sg13g2_tiehi _1187__83 (.L_HI(net83));
 sg13g2_tiehi _1287__84 (.L_HI(net84));
 sg13g2_tiehi _1186__85 (.L_HI(net85));
 sg13g2_tiehi _1286__86 (.L_HI(net86));
 sg13g2_tiehi _1182__87 (.L_HI(net87));
 sg13g2_tiehi _1181__88 (.L_HI(net88));
 sg13g2_tiehi _1180__89 (.L_HI(net89));
 sg13g2_tiehi _1179__90 (.L_HI(net90));
 sg13g2_tiehi _1178__91 (.L_HI(net91));
 sg13g2_tiehi _1177__92 (.L_HI(net92));
 sg13g2_tiehi _1176__93 (.L_HI(net93));
 sg13g2_tiehi _1175__94 (.L_HI(net94));
 sg13g2_tiehi _1174__95 (.L_HI(net95));
 sg13g2_tiehi _1285__96 (.L_HI(net96));
 sg13g2_tiehi _1284__97 (.L_HI(net97));
 sg13g2_tiehi _1283__98 (.L_HI(net98));
 sg13g2_tiehi _1282__99 (.L_HI(net99));
 sg13g2_tiehi _1281__100 (.L_HI(net100));
 sg13g2_tiehi _1280__101 (.L_HI(net101));
 sg13g2_tiehi _1279__102 (.L_HI(net102));
 sg13g2_tiehi _1278__103 (.L_HI(net103));
 sg13g2_tiehi _1277__104 (.L_HI(net104));
 sg13g2_tiehi _1276__105 (.L_HI(net105));
 sg13g2_tiehi _1275__106 (.L_HI(net106));
 sg13g2_tiehi _1274__107 (.L_HI(net107));
 sg13g2_tiehi _1273__108 (.L_HI(net108));
 sg13g2_tiehi _1272__109 (.L_HI(net109));
 sg13g2_tiehi _1271__110 (.L_HI(net110));
 sg13g2_tiehi _1270__111 (.L_HI(net111));
 sg13g2_tiehi _1269__112 (.L_HI(net112));
 sg13g2_tiehi _1268__113 (.L_HI(net113));
 sg13g2_tiehi _1267__114 (.L_HI(net114));
 sg13g2_tiehi _1266__115 (.L_HI(net115));
 sg13g2_tiehi _1265__116 (.L_HI(net116));
 sg13g2_tiehi _1264__117 (.L_HI(net117));
 sg13g2_tiehi _1263__118 (.L_HI(net118));
 sg13g2_tiehi _1262__119 (.L_HI(net119));
 sg13g2_tiehi _1261__120 (.L_HI(net120));
 sg13g2_tiehi _1260__121 (.L_HI(net121));
 sg13g2_tiehi _1259__122 (.L_HI(net122));
 sg13g2_tiehi _1258__123 (.L_HI(net123));
 sg13g2_tiehi _1257__124 (.L_HI(net124));
 sg13g2_tiehi _1256__125 (.L_HI(net125));
 sg13g2_tiehi _1255__126 (.L_HI(net126));
 sg13g2_tiehi _1254__127 (.L_HI(net127));
 sg13g2_tiehi _1253__128 (.L_HI(net128));
 sg13g2_tiehi _1252__129 (.L_HI(net129));
 sg13g2_tiehi _1251__130 (.L_HI(net130));
 sg13g2_tiehi _1250__131 (.L_HI(net131));
 sg13g2_tiehi _1249__132 (.L_HI(net132));
 sg13g2_tiehi _1248__133 (.L_HI(net133));
 sg13g2_tiehi _1247__134 (.L_HI(net134));
 sg13g2_tiehi _1246__135 (.L_HI(net135));
 sg13g2_tiehi _1245__136 (.L_HI(net136));
 sg13g2_tiehi _1244__137 (.L_HI(net137));
 sg13g2_tiehi _1243__138 (.L_HI(net138));
 sg13g2_tiehi _1242__139 (.L_HI(net139));
 sg13g2_tiehi _1241__140 (.L_HI(net140));
 sg13g2_tiehi _1240__141 (.L_HI(net188));
 sg13g2_tiehi _1312__142 (.L_HI(net189));
 sg13g2_tiehi _1239__143 (.L_HI(net190));
 sg13g2_tiehi _1317__144 (.L_HI(net191));
 sg13g2_tiehi _1238__145 (.L_HI(net192));
 sg13g2_tiehi _1311__146 (.L_HI(net193));
 sg13g2_tiehi _1237__147 (.L_HI(net194));
 sg13g2_tiehi _1322__148 (.L_HI(net195));
 sg13g2_tiehi _1236__149 (.L_HI(net196));
 sg13g2_tiehi _1310__150 (.L_HI(net197));
 sg13g2_tiehi _1235__151 (.L_HI(net198));
 sg13g2_tiehi _1316__152 (.L_HI(net199));
 sg13g2_tiehi _1234__153 (.L_HI(net200));
 sg13g2_tiehi _1309__154 (.L_HI(net201));
 sg13g2_tiehi _1233__155 (.L_HI(net202));
 sg13g2_tiehi _1319__156 (.L_HI(net203));
 sg13g2_tiehi _1232__157 (.L_HI(net204));
 sg13g2_tiehi _1231__158 (.L_HI(net205));
 sg13g2_tiehi _1230__159 (.L_HI(net206));
 sg13g2_tiehi _1229__160 (.L_HI(net207));
 sg13g2_tiehi _1228__161 (.L_HI(net208));
 sg13g2_tiehi _1227__162 (.L_HI(net209));
 sg13g2_tiehi _1226__163 (.L_HI(net210));
 sg13g2_tiehi _1225__164 (.L_HI(net211));
 sg13g2_tiehi _1224__165 (.L_HI(net212));
 sg13g2_tiehi _1223__166 (.L_HI(net213));
 sg13g2_tiehi _1308__167 (.L_HI(net214));
 sg13g2_tiehi _1222__168 (.L_HI(net215));
 sg13g2_tiehi _1221__169 (.L_HI(net216));
 sg13g2_tiehi _1220__170 (.L_HI(net217));
 sg13g2_tiehi _1219__171 (.L_HI(net218));
 sg13g2_tiehi _1214__172 (.L_HI(net219));
 sg13g2_tiehi \async_reset_ctrl/_18__173  (.L_HI(net220));
 sg13g2_tielo tt_um_dlmiles_tt08_poc_uart_16 (.L_LO(net16));
 sg13g2_tielo tt_um_dlmiles_tt08_poc_uart_17 (.L_LO(net17));
 sg13g2_tielo tt_um_dlmiles_tt08_poc_uart_18 (.L_LO(net18));
 sg13g2_tielo tt_um_dlmiles_tt08_poc_uart_19 (.L_LO(net19));
 sg13g2_tielo tt_um_dlmiles_tt08_poc_uart_20 (.L_LO(net20));
 sg13g2_tielo tt_um_dlmiles_tt08_poc_uart_21 (.L_LO(net21));
 sg13g2_tielo tt_um_dlmiles_tt08_poc_uart_22 (.L_LO(net22));
 sg13g2_tiehi _1218__23 (.L_HI(net23));
 sg13g2_buf_1 _1481_ (.A(\uart.uartArea_uart.busCtrl.oe ),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1482_ (.A(\uart.uartArea_uart.busCtrl.oe ),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1483_ (.A(\uart.uartArea_uart.busCtrl.oe ),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1484_ (.A(\uart.uartArea_uart.busCtrl.oe ),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1485_ (.A(\uart.uartArea_uart.busCtrl.oe ),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1486_ (.A(\uart.uartArea_uart.busCtrl.oe ),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1487_ (.A(\uart.uartArea_uart.busCtrl.oe ),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1488_ (.A(\uart.uartArea_uart.busCtrl.oe ),
    .X(uio_oe[7]));
 sg13g2_inv_1 \async_reset_ctrl/_13_  (.Y(\async_reset_ctrl/_07_ ),
    .A(net226));
 sg13g2_nand2b_1 \async_reset_ctrl/_14_  (.Y(\async_reset_ctrl/_08_ ),
    .B(net381),
    .A_N(sync_reset));
 sg13g2_or2_1 \async_reset_ctrl/_15_  (.X(\async_reset_ctrl/_04_ ),
    .B(net382),
    .A(net225));
 sg13g2_nand2b_1 \async_reset_ctrl/_16_  (.Y(\async_reset_ctrl/_06_ ),
    .B(net1),
    .A_N(net381));
 sg13g2_dfrbp_1 \async_reset_ctrl/_17_  (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net221),
    .D(net225),
    .Q_N(\async_reset_ctrl/_10_ ),
    .Q(\async_reset_ctrl/dff3.q ));
 sg13g2_dfrbp_1 \async_reset_ctrl/_18_  (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net220),
    .D(net227),
    .Q_N(\async_reset_ctrl/_09_ ),
    .Q(sync_reset));
 sg13g2_dfrbp_1 \async_reset_ctrl/_19_  (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(\async_reset_ctrl/_04_ ),
    .D(net222),
    .Q_N(\async_reset_ctrl/dff_async_set1.q ),
    .Q(\async_reset_ctrl/_00_ ));
 sg13g2_dfrbp_1 \async_reset_ctrl/_20_  (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(\async_reset_ctrl/_06_ ),
    .D(net223),
    .Q_N(\async_reset_ctrl/async_reset_in_triggered ),
    .Q(\async_reset_ctrl/_01_ ));
 sg13g2_dfrbp_1 \async_reset_ctrl/_21_  (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net382),
    .D(\async_reset_ctrl/_07_ ),
    .Q_N(\async_reset_ctrl/dff3.d ),
    .Q(\async_reset_ctrl/_02_ ));
 sg13g2_tiehi \async_reset_ctrl/_17__174  (.L_HI(net221));
 sg13g2_tiehi \async_reset_ctrl/_19__175  (.L_HI(net222));
 sg13g2_tiehi \async_reset_ctrl/_20__176  (.L_HI(net223));
 sg13g2_inv_1 _0756__1 (.Y(net224),
    .A(clknet_1_0__leaf_clk));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(_0408_));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(_0407_));
 sg13g2_buf_4 fanout143 (.X(net143),
    .A(_0406_));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(_0405_));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(_0404_));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(_0403_));
 sg13g2_buf_4 fanout147 (.X(net147),
    .A(_0384_));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(_0338_));
 sg13g2_buf_2 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_0337_),
    .X(net150));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(_0229_));
 sg13g2_buf_1 fanout152 (.A(_0229_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_4 fanout154 (.X(net154),
    .A(_0362_));
 sg13g2_buf_2 fanout155 (.A(net156),
    .X(net155));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(_0354_));
 sg13g2_buf_2 fanout157 (.A(_0225_),
    .X(net157));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(_0209_));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(_0208_));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(_0207_));
 sg13g2_buf_4 fanout161 (.X(net161),
    .A(_0205_));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(_0202_));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(_0200_));
 sg13g2_buf_4 fanout164 (.X(net164),
    .A(_0198_));
 sg13g2_buf_2 fanout165 (.A(net169),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(net168),
    .X(net167));
 sg13g2_buf_1 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_0321_),
    .X(net169));
 sg13g2_buf_4 fanout170 (.X(net170),
    .A(_0320_));
 sg13g2_buf_2 fanout171 (.A(_0320_),
    .X(net171));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(_0180_));
 sg13g2_buf_1 fanout173 (.A(_0180_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_0179_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(net428),
    .X(net175));
 sg13g2_buf_4 fanout176 (.X(net176),
    .A(net430));
 sg13g2_buf_4 fanout177 (.X(net177),
    .A(net429));
 sg13g2_buf_2 fanout178 (.A(_0373_),
    .X(net178));
 sg13g2_buf_4 fanout179 (.X(net179),
    .A(net14));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(net13));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(net12));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(net11));
 sg13g2_buf_2 fanout183 (.A(net10),
    .X(net183));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(net9));
 sg13g2_buf_2 fanout185 (.A(net8),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(net187),
    .X(net186));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(uio_in[0]));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[6]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[7]),
    .X(net14));
 sg13g2_tielo tt_um_dlmiles_tt08_poc_uart_15 (.L_LO(net15));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_inv_1 clkload0 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_5_15__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_5_23__leaf_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\async_reset_ctrl/dff3.d ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold2 (.A(\async_reset_ctrl/dff_async_set1.q ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold3 (.A(\async_reset_ctrl/dff3.q ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold4 (.A(\uart.resetCommandUnit_1.reg1 ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold5 (.A(rst_n_sync),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold6 (.A(\uart.uartArea_uart.commFilter.io_ttl_ri ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0004_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0006_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0002_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0134_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0001_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0145_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold13 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[2] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold14 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[5] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold15 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[4] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold16 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[3] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold17 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[6] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold18 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[0] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold19 (.A(\uart.uartArea_uart.regCtrl.txOverrun ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0335_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0016_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0003_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0385_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0060_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold25 (.A(\uart.uartArea_uart.regCtrl.regFifoRxEnable ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold26 (.A(\uart.uartArea_uart.uartClocking_1.divisorCtr[7] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0013_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold28 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptStatus[1] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold29 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_9[1] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold30 (.A(\uart.uartArea_uart.regCtrl.regFifoTxEnable ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold31 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_13[7] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold32 (.A(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[3] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0133_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold34 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_10[6] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold35 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_10[3] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold36 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_10[8] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0102_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold38 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_13[2] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold39 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[8] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0084_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold41 (.A(\uart.uartArea_uart.uartClocking_1.divisorCtr[3] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0326_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0009_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold44 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_9[5] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold45 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_10[7] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold46 (.A(\uart.uartArea_uart.regCtrl.regModemCtrlChanged[2] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0333_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0015_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold49 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_9[2] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold50 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_9[3] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold51 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_9[0] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold52 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_12[2] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0114_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold54 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_14[8] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0059_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold56 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_12[1] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold57 (.A(\uart.uartArea_uart.busCtrl.io_regAddr[4] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold58 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[0] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold59 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_14[1] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold60 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[1] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold61 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_10[4] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold62 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_9[7] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold63 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_14[0] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold64 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[6] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold65 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_10[1] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold66 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_9[4] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold67 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[2] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0078_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold69 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_13[1] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold70 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_12[4] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold71 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_12[3] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold72 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_9[8] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0093_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold74 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_9[6] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold75 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_14[2] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold76 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_13[3] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold77 (.A(\uart.uartArea_uart.regCtrl.regModemCtrlHistory[1] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0139_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold79 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[7] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold80 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[4] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold81 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_12[6] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold82 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[3] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold83 (.A(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[3] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0144_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold85 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_14[6] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold86 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_14[3] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold87 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_12[7] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold88 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_13[5] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold89 (.A(\uart.uartArea_uart.uartClocking_1.bitCtr[2] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0388_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0062_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold92 (.A(\uart.uartArea_uart.commFilter.dsrFilter.io_c ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0394_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0066_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold95 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_10[2] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold96 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_13[6] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold97 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_13[0] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold98 (.A(\uart.uartArea_uart.commFilter.dcdFilter.io_c ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0392_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0065_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold101 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_12[0] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold102 (.A(\uart.uartArea_uart.rxFifo.count[3] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold103 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_14[5] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold104 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_14[7] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold105 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_10[0] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold106 (.A(\uart.uartArea_uart.regCtrl.regModemCtrlHistory[3] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0140_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold108 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_10[5] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold109 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_13[8] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0129_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold111 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_8[5] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold112 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_12[5] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold113 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_11[2] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold114 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_12[8] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0120_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold116 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_13[4] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold117 (.A(\uart.uartArea_uart.regCtrl.regModemCtrlChanged[3] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0343_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0020_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold120 (.A(\uart.uartArea_uart.commFilter.riFilter.io_c ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0390_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0064_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold123 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_11[3] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold124 (.A(\uart.uartArea_uart.rxFifo.count[2] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0433_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0147_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold127 (.A(\uart.uartArea_uart.commFilter.dsrFilter.io_b ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold128 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_11[0] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold129 (.A(\uart.uartArea_uart.commFilter.ctsFilter.io_c ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0396_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0067_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold132 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_11[6] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold133 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_11[5] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold134 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_11[4] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold135 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_11[1] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold136 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_11[8] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0111_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold138 (.A(\uart.uartArea_uart.commFilter.ctsFilter.io_b ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold139 (.A(\uart.uartArea_uart.commFilter.riFilter.io_b ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold140 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_11[7] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold141 (.A(\uart.uartArea_uart.sharedFifo.fifoRegs_14[4] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0055_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold143 (.A(\uart.uartArea_uart.regCtrl.regModemCtrlHistory[0] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0138_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold145 (.A(\uart.uartArea_uart.commFilter.dcdFilter.io_b ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold146 (.A(\uart.uartArea_uart.txFifo.count[1] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0414_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0135_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold149 (.A(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[1] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0425_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold151 (.A(\uart.uartArea_uart.regCtrl.reg007[2] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold152 (.A(\uart.uartArea_uart.regCtrl.reg007[0] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold153 (.A(\uart.uartArea_uart.commFilter.dsrFilter.io_o ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0014_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold155 (.A(\uart.uartArea_uart.commFilter.ctsFilter.io_o ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0149_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold157 (.A(\async_reset_ctrl/async_reset_in_triggered ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold158 (.A(\async_reset_ctrl/_08_ ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold159 (.A(\uart.uartArea_uart.uartClocking_1.bitCtr[3] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold160 (.A(\uart.uartArea_uart.uartClocking_1.bitCtr[1] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0387_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0061_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold163 (.A(\uart.uartArea_uart.uartClocking_1.divisorCtr[6] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0330_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold165 (.A(\uart.uartArea_uart.uartClocking_1.bitCtr[0] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold166 (.A(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[1] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0410_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold168 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptControl[1] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold169 (.A(\uart.uartArea_uart.regCtrl.reg007[7] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold170 (.A(\uart.uartArea_uart.regCtrl.reg007[1] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold171 (.A(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[2] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold172 (.A(\uart.uartArea_uart.regCtrl.reg007[3] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold173 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptControl[6] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold174 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptControl[3] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold175 (.A(\uart.uartArea_uart.regCtrl.reg007[4] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold176 (.A(\uart.uartArea_uart.regCtrl.reg007[5] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold177 (.A(\uart.uartArea_uart.uartClocking_1.divisorCtr[0] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0323_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold179 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptControl[2] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold180 (.A(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[0] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold181 (.A(\uart.uartArea_uart.regCtrl.reg007[6] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold182 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptControl[4] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold183 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptControl[0] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold184 (.A(\uart.resetCommandUnit_1.io_resetIn ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold185 (.A(\uart.uartArea_uart.busCtrl.io_regAddr[3] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold186 (.A(\uart.uartArea_uart.rxFifo.count[1] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0432_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold188 (.A(\uart.uartArea_uart.uartClocking_1.divisorCtr[2] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0315_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0325_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold191 (.A(\uart.uartArea_uart.txFifo.count[3] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0137_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold193 (.A(\uart.uartArea_uart.rxFifo.io_fifoRdAddr[2] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0428_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold195 (.A(\uart.uartArea_uart.regCtrl.io_regInterruptControl[5] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold196 (.A(\uart.uartArea_uart.uartClocking_1.divisorCtr[4] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0327_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold198 (.A(\uart.uartArea_uart.txFifo.count[2] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0417_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold200 (.A(\uart.uartArea_uart.busCtrl.io_regAddr[2] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold201 (.A(\uart.uartArea_uart.regCtrl.txHolderBit9 ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold202 (.A(\uart.uartArea_uart.uartClocking_1.divisorCtr[5] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0317_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold204 (.A(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[0] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold205 (.A(\uart.uartArea_uart.busCtrl.io_regAddr[0] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold206 (.A(\uart.uartArea_uart.busCtrl.io_regAddr[1] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold207 (.A(\uart.uartArea_uart.sharedFifo.io_txFifoWrAddr[1] ),
    .X(net431));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_4 FILLER_22_189 ();
 sg13g2_fill_2 FILLER_22_193 ();
 sg13g2_fill_2 FILLER_22_200 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_decap_8 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_214 ();
 sg13g2_decap_8 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_235 ();
 sg13g2_decap_8 FILLER_22_242 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_256 ();
 sg13g2_decap_8 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_4 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_186 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_4 FILLER_24_175 ();
 sg13g2_fill_1 FILLER_24_179 ();
 sg13g2_fill_2 FILLER_24_210 ();
 sg13g2_decap_4 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_247 ();
 sg13g2_decap_8 FILLER_24_254 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_268 ();
 sg13g2_decap_8 FILLER_24_275 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_decap_8 FILLER_24_289 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_310 ();
 sg13g2_decap_8 FILLER_24_317 ();
 sg13g2_decap_8 FILLER_24_324 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_4 FILLER_25_182 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_221 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_decap_8 FILLER_25_265 ();
 sg13g2_decap_8 FILLER_25_272 ();
 sg13g2_decap_8 FILLER_25_279 ();
 sg13g2_decap_8 FILLER_25_286 ();
 sg13g2_decap_8 FILLER_25_293 ();
 sg13g2_decap_8 FILLER_25_300 ();
 sg13g2_decap_8 FILLER_25_307 ();
 sg13g2_decap_8 FILLER_25_314 ();
 sg13g2_decap_8 FILLER_25_321 ();
 sg13g2_decap_8 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_decap_8 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_349 ();
 sg13g2_decap_8 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_fill_2 FILLER_26_189 ();
 sg13g2_fill_2 FILLER_26_200 ();
 sg13g2_fill_1 FILLER_26_202 ();
 sg13g2_fill_1 FILLER_26_208 ();
 sg13g2_fill_1 FILLER_26_232 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_4 FILLER_27_154 ();
 sg13g2_fill_1 FILLER_27_158 ();
 sg13g2_decap_4 FILLER_27_168 ();
 sg13g2_fill_1 FILLER_27_198 ();
 sg13g2_fill_1 FILLER_27_213 ();
 sg13g2_fill_1 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_254 ();
 sg13g2_decap_8 FILLER_27_267 ();
 sg13g2_decap_8 FILLER_27_274 ();
 sg13g2_decap_8 FILLER_27_281 ();
 sg13g2_decap_8 FILLER_27_288 ();
 sg13g2_decap_8 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_decap_8 FILLER_27_309 ();
 sg13g2_decap_8 FILLER_27_316 ();
 sg13g2_decap_8 FILLER_27_323 ();
 sg13g2_decap_8 FILLER_27_330 ();
 sg13g2_decap_8 FILLER_27_337 ();
 sg13g2_decap_8 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_4 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_137 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_decap_4 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_225 ();
 sg13g2_decap_8 FILLER_28_244 ();
 sg13g2_fill_2 FILLER_28_251 ();
 sg13g2_fill_2 FILLER_28_257 ();
 sg13g2_decap_8 FILLER_28_268 ();
 sg13g2_decap_8 FILLER_28_275 ();
 sg13g2_decap_8 FILLER_28_282 ();
 sg13g2_decap_8 FILLER_28_289 ();
 sg13g2_decap_8 FILLER_28_296 ();
 sg13g2_decap_8 FILLER_28_303 ();
 sg13g2_decap_8 FILLER_28_310 ();
 sg13g2_decap_8 FILLER_28_317 ();
 sg13g2_decap_8 FILLER_28_324 ();
 sg13g2_decap_8 FILLER_28_331 ();
 sg13g2_decap_8 FILLER_28_338 ();
 sg13g2_decap_8 FILLER_28_345 ();
 sg13g2_decap_8 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_28_359 ();
 sg13g2_decap_8 FILLER_28_366 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_4 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_fill_2 FILLER_29_207 ();
 sg13g2_fill_1 FILLER_29_209 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_264 ();
 sg13g2_decap_8 FILLER_29_274 ();
 sg13g2_decap_8 FILLER_29_281 ();
 sg13g2_decap_8 FILLER_29_288 ();
 sg13g2_decap_8 FILLER_29_295 ();
 sg13g2_decap_8 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_309 ();
 sg13g2_decap_8 FILLER_29_316 ();
 sg13g2_decap_8 FILLER_29_323 ();
 sg13g2_decap_8 FILLER_29_330 ();
 sg13g2_decap_8 FILLER_29_337 ();
 sg13g2_decap_8 FILLER_29_344 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_4 FILLER_30_140 ();
 sg13g2_fill_2 FILLER_30_144 ();
 sg13g2_fill_2 FILLER_30_170 ();
 sg13g2_fill_2 FILLER_30_215 ();
 sg13g2_fill_1 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_222 ();
 sg13g2_decap_4 FILLER_30_229 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_fill_2 FILLER_30_239 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_decap_8 FILLER_30_278 ();
 sg13g2_decap_8 FILLER_30_285 ();
 sg13g2_decap_8 FILLER_30_292 ();
 sg13g2_decap_8 FILLER_30_299 ();
 sg13g2_decap_8 FILLER_30_306 ();
 sg13g2_decap_8 FILLER_30_313 ();
 sg13g2_decap_8 FILLER_30_320 ();
 sg13g2_decap_8 FILLER_30_327 ();
 sg13g2_decap_8 FILLER_30_334 ();
 sg13g2_decap_8 FILLER_30_341 ();
 sg13g2_decap_8 FILLER_30_348 ();
 sg13g2_decap_8 FILLER_30_355 ();
 sg13g2_decap_8 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_30_369 ();
 sg13g2_decap_8 FILLER_30_376 ();
 sg13g2_decap_8 FILLER_30_383 ();
 sg13g2_decap_8 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_fill_2 FILLER_31_147 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_fill_2 FILLER_31_196 ();
 sg13g2_fill_1 FILLER_31_198 ();
 sg13g2_fill_2 FILLER_31_212 ();
 sg13g2_fill_1 FILLER_31_214 ();
 sg13g2_decap_8 FILLER_31_293 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_decap_8 FILLER_31_307 ();
 sg13g2_decap_8 FILLER_31_314 ();
 sg13g2_decap_8 FILLER_31_321 ();
 sg13g2_decap_8 FILLER_31_328 ();
 sg13g2_decap_8 FILLER_31_335 ();
 sg13g2_decap_8 FILLER_31_342 ();
 sg13g2_decap_8 FILLER_31_349 ();
 sg13g2_decap_8 FILLER_31_356 ();
 sg13g2_decap_8 FILLER_31_363 ();
 sg13g2_decap_8 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_31_384 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_4 FILLER_32_119 ();
 sg13g2_fill_2 FILLER_32_123 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_decap_4 FILLER_32_194 ();
 sg13g2_fill_2 FILLER_32_198 ();
 sg13g2_decap_8 FILLER_32_285 ();
 sg13g2_decap_8 FILLER_32_292 ();
 sg13g2_decap_8 FILLER_32_299 ();
 sg13g2_decap_8 FILLER_32_306 ();
 sg13g2_decap_8 FILLER_32_313 ();
 sg13g2_decap_8 FILLER_32_320 ();
 sg13g2_decap_8 FILLER_32_327 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_341 ();
 sg13g2_decap_8 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_362 ();
 sg13g2_decap_8 FILLER_32_369 ();
 sg13g2_decap_8 FILLER_32_376 ();
 sg13g2_decap_8 FILLER_32_383 ();
 sg13g2_decap_8 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_397 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_126 ();
 sg13g2_fill_2 FILLER_33_167 ();
 sg13g2_fill_2 FILLER_33_198 ();
 sg13g2_fill_2 FILLER_33_208 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_277 ();
 sg13g2_fill_1 FILLER_33_279 ();
 sg13g2_decap_8 FILLER_33_289 ();
 sg13g2_decap_8 FILLER_33_296 ();
 sg13g2_decap_8 FILLER_33_303 ();
 sg13g2_decap_8 FILLER_33_310 ();
 sg13g2_decap_8 FILLER_33_317 ();
 sg13g2_decap_8 FILLER_33_324 ();
 sg13g2_decap_8 FILLER_33_331 ();
 sg13g2_decap_8 FILLER_33_338 ();
 sg13g2_decap_8 FILLER_33_345 ();
 sg13g2_decap_8 FILLER_33_352 ();
 sg13g2_decap_8 FILLER_33_359 ();
 sg13g2_decap_8 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_380 ();
 sg13g2_decap_8 FILLER_33_387 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_fill_2 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_213 ();
 sg13g2_fill_2 FILLER_34_226 ();
 sg13g2_fill_2 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_242 ();
 sg13g2_fill_1 FILLER_34_255 ();
 sg13g2_decap_4 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_265 ();
 sg13g2_decap_8 FILLER_34_269 ();
 sg13g2_decap_8 FILLER_34_276 ();
 sg13g2_decap_8 FILLER_34_283 ();
 sg13g2_decap_8 FILLER_34_290 ();
 sg13g2_decap_8 FILLER_34_297 ();
 sg13g2_decap_8 FILLER_34_304 ();
 sg13g2_decap_8 FILLER_34_311 ();
 sg13g2_decap_8 FILLER_34_318 ();
 sg13g2_decap_8 FILLER_34_325 ();
 sg13g2_decap_8 FILLER_34_332 ();
 sg13g2_decap_8 FILLER_34_339 ();
 sg13g2_decap_8 FILLER_34_346 ();
 sg13g2_decap_8 FILLER_34_353 ();
 sg13g2_decap_8 FILLER_34_360 ();
 sg13g2_decap_8 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_34_374 ();
 sg13g2_decap_8 FILLER_34_381 ();
 sg13g2_decap_8 FILLER_34_388 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_4 FILLER_35_119 ();
 sg13g2_fill_2 FILLER_35_123 ();
 sg13g2_decap_8 FILLER_35_288 ();
 sg13g2_decap_8 FILLER_35_295 ();
 sg13g2_decap_8 FILLER_35_302 ();
 sg13g2_decap_8 FILLER_35_309 ();
 sg13g2_decap_8 FILLER_35_316 ();
 sg13g2_decap_8 FILLER_35_323 ();
 sg13g2_decap_8 FILLER_35_330 ();
 sg13g2_decap_8 FILLER_35_337 ();
 sg13g2_decap_8 FILLER_35_344 ();
 sg13g2_decap_8 FILLER_35_351 ();
 sg13g2_decap_8 FILLER_35_358 ();
 sg13g2_decap_8 FILLER_35_365 ();
 sg13g2_decap_8 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_248 ();
 sg13g2_decap_8 FILLER_36_302 ();
 sg13g2_decap_8 FILLER_36_309 ();
 sg13g2_decap_8 FILLER_36_316 ();
 sg13g2_decap_8 FILLER_36_323 ();
 sg13g2_decap_8 FILLER_36_330 ();
 sg13g2_decap_8 FILLER_36_337 ();
 sg13g2_decap_8 FILLER_36_344 ();
 sg13g2_decap_8 FILLER_36_351 ();
 sg13g2_decap_8 FILLER_36_358 ();
 sg13g2_decap_8 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_2 FILLER_37_176 ();
 sg13g2_fill_2 FILLER_37_201 ();
 sg13g2_fill_1 FILLER_37_203 ();
 sg13g2_fill_1 FILLER_37_215 ();
 sg13g2_fill_2 FILLER_37_239 ();
 sg13g2_fill_1 FILLER_37_241 ();
 sg13g2_decap_8 FILLER_37_305 ();
 sg13g2_decap_8 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_decap_8 FILLER_37_333 ();
 sg13g2_decap_8 FILLER_37_340 ();
 sg13g2_decap_8 FILLER_37_347 ();
 sg13g2_decap_8 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_37_361 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_4 FILLER_38_126 ();
 sg13g2_fill_1 FILLER_38_181 ();
 sg13g2_fill_2 FILLER_38_187 ();
 sg13g2_fill_2 FILLER_38_233 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_decap_8 FILLER_38_299 ();
 sg13g2_decap_8 FILLER_38_306 ();
 sg13g2_decap_8 FILLER_38_313 ();
 sg13g2_decap_8 FILLER_38_320 ();
 sg13g2_decap_8 FILLER_38_327 ();
 sg13g2_decap_8 FILLER_38_334 ();
 sg13g2_decap_8 FILLER_38_341 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_decap_8 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_362 ();
 sg13g2_decap_8 FILLER_38_369 ();
 sg13g2_decap_8 FILLER_38_376 ();
 sg13g2_decap_8 FILLER_38_383 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_4 FILLER_39_119 ();
 sg13g2_fill_2 FILLER_39_123 ();
 sg13g2_fill_2 FILLER_39_197 ();
 sg13g2_fill_1 FILLER_39_211 ();
 sg13g2_fill_2 FILLER_39_239 ();
 sg13g2_fill_1 FILLER_39_246 ();
 sg13g2_fill_1 FILLER_39_263 ();
 sg13g2_decap_8 FILLER_39_290 ();
 sg13g2_decap_8 FILLER_39_297 ();
 sg13g2_decap_8 FILLER_39_304 ();
 sg13g2_decap_8 FILLER_39_311 ();
 sg13g2_decap_8 FILLER_39_318 ();
 sg13g2_decap_8 FILLER_39_325 ();
 sg13g2_decap_8 FILLER_39_332 ();
 sg13g2_decap_8 FILLER_39_339 ();
 sg13g2_decap_8 FILLER_39_346 ();
 sg13g2_decap_8 FILLER_39_353 ();
 sg13g2_decap_8 FILLER_39_360 ();
 sg13g2_decap_8 FILLER_39_367 ();
 sg13g2_decap_8 FILLER_39_374 ();
 sg13g2_decap_8 FILLER_39_381 ();
 sg13g2_decap_8 FILLER_39_388 ();
 sg13g2_decap_8 FILLER_39_395 ();
 sg13g2_decap_8 FILLER_39_402 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_fill_2 FILLER_40_168 ();
 sg13g2_fill_1 FILLER_40_170 ();
 sg13g2_fill_2 FILLER_40_197 ();
 sg13g2_fill_1 FILLER_40_199 ();
 sg13g2_fill_2 FILLER_40_244 ();
 sg13g2_fill_1 FILLER_40_246 ();
 sg13g2_fill_2 FILLER_40_252 ();
 sg13g2_fill_1 FILLER_40_254 ();
 sg13g2_decap_8 FILLER_40_281 ();
 sg13g2_decap_8 FILLER_40_288 ();
 sg13g2_decap_8 FILLER_40_295 ();
 sg13g2_decap_8 FILLER_40_302 ();
 sg13g2_decap_8 FILLER_40_309 ();
 sg13g2_decap_8 FILLER_40_316 ();
 sg13g2_decap_8 FILLER_40_323 ();
 sg13g2_decap_8 FILLER_40_330 ();
 sg13g2_decap_8 FILLER_40_337 ();
 sg13g2_decap_8 FILLER_40_344 ();
 sg13g2_decap_8 FILLER_40_351 ();
 sg13g2_decap_8 FILLER_40_358 ();
 sg13g2_decap_8 FILLER_40_365 ();
 sg13g2_decap_8 FILLER_40_372 ();
 sg13g2_decap_8 FILLER_40_379 ();
 sg13g2_decap_8 FILLER_40_386 ();
 sg13g2_decap_8 FILLER_40_393 ();
 sg13g2_decap_8 FILLER_40_400 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_fill_1 FILLER_41_151 ();
 sg13g2_fill_2 FILLER_41_167 ();
 sg13g2_fill_2 FILLER_41_175 ();
 sg13g2_fill_1 FILLER_41_177 ();
 sg13g2_fill_1 FILLER_41_188 ();
 sg13g2_decap_8 FILLER_41_241 ();
 sg13g2_fill_2 FILLER_41_248 ();
 sg13g2_fill_1 FILLER_41_250 ();
 sg13g2_decap_8 FILLER_41_267 ();
 sg13g2_decap_8 FILLER_41_278 ();
 sg13g2_decap_8 FILLER_41_285 ();
 sg13g2_decap_8 FILLER_41_292 ();
 sg13g2_decap_8 FILLER_41_299 ();
 sg13g2_decap_8 FILLER_41_306 ();
 sg13g2_decap_8 FILLER_41_313 ();
 sg13g2_decap_8 FILLER_41_320 ();
 sg13g2_decap_8 FILLER_41_327 ();
 sg13g2_decap_8 FILLER_41_334 ();
 sg13g2_decap_8 FILLER_41_341 ();
 sg13g2_decap_8 FILLER_41_348 ();
 sg13g2_decap_8 FILLER_41_355 ();
 sg13g2_decap_8 FILLER_41_362 ();
 sg13g2_decap_8 FILLER_41_369 ();
 sg13g2_decap_8 FILLER_41_376 ();
 sg13g2_decap_8 FILLER_41_383 ();
 sg13g2_decap_8 FILLER_41_390 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_fill_1 FILLER_42_126 ();
 sg13g2_decap_4 FILLER_42_153 ();
 sg13g2_fill_1 FILLER_42_157 ();
 sg13g2_decap_8 FILLER_42_194 ();
 sg13g2_decap_8 FILLER_42_201 ();
 sg13g2_decap_8 FILLER_42_208 ();
 sg13g2_fill_1 FILLER_42_215 ();
 sg13g2_decap_4 FILLER_42_220 ();
 sg13g2_fill_1 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_242 ();
 sg13g2_decap_4 FILLER_42_249 ();
 sg13g2_fill_1 FILLER_42_253 ();
 sg13g2_decap_8 FILLER_42_290 ();
 sg13g2_decap_8 FILLER_42_297 ();
 sg13g2_decap_8 FILLER_42_304 ();
 sg13g2_decap_8 FILLER_42_311 ();
 sg13g2_decap_8 FILLER_42_318 ();
 sg13g2_decap_8 FILLER_42_325 ();
 sg13g2_decap_8 FILLER_42_332 ();
 sg13g2_decap_8 FILLER_42_339 ();
 sg13g2_decap_8 FILLER_42_346 ();
 sg13g2_decap_8 FILLER_42_353 ();
 sg13g2_decap_8 FILLER_42_360 ();
 sg13g2_decap_8 FILLER_42_367 ();
 sg13g2_decap_8 FILLER_42_374 ();
 sg13g2_decap_8 FILLER_42_381 ();
 sg13g2_decap_8 FILLER_42_388 ();
 sg13g2_decap_8 FILLER_42_395 ();
 sg13g2_decap_8 FILLER_42_402 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_4 FILLER_43_152 ();
 sg13g2_fill_1 FILLER_43_156 ();
 sg13g2_decap_8 FILLER_43_183 ();
 sg13g2_fill_1 FILLER_43_190 ();
 sg13g2_fill_1 FILLER_43_207 ();
 sg13g2_decap_8 FILLER_43_223 ();
 sg13g2_decap_4 FILLER_43_230 ();
 sg13g2_decap_8 FILLER_43_289 ();
 sg13g2_decap_8 FILLER_43_296 ();
 sg13g2_decap_8 FILLER_43_303 ();
 sg13g2_decap_8 FILLER_43_310 ();
 sg13g2_decap_8 FILLER_43_317 ();
 sg13g2_decap_8 FILLER_43_324 ();
 sg13g2_decap_8 FILLER_43_331 ();
 sg13g2_decap_8 FILLER_43_338 ();
 sg13g2_decap_4 FILLER_43_345 ();
 sg13g2_fill_1 FILLER_43_349 ();
 sg13g2_decap_8 FILLER_43_376 ();
 sg13g2_decap_8 FILLER_43_383 ();
 sg13g2_decap_8 FILLER_43_390 ();
 sg13g2_decap_8 FILLER_43_397 ();
 sg13g2_decap_4 FILLER_43_404 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_fill_2 FILLER_44_119 ();
 sg13g2_decap_4 FILLER_44_184 ();
 sg13g2_fill_2 FILLER_44_232 ();
 sg13g2_fill_1 FILLER_44_234 ();
 sg13g2_decap_8 FILLER_44_299 ();
 sg13g2_decap_8 FILLER_44_306 ();
 sg13g2_decap_8 FILLER_44_313 ();
 sg13g2_decap_8 FILLER_44_320 ();
 sg13g2_decap_8 FILLER_44_327 ();
 sg13g2_fill_2 FILLER_44_334 ();
 sg13g2_fill_1 FILLER_44_336 ();
 sg13g2_decap_4 FILLER_44_342 ();
 sg13g2_fill_2 FILLER_44_346 ();
 sg13g2_decap_8 FILLER_44_387 ();
 sg13g2_decap_8 FILLER_44_394 ();
 sg13g2_decap_8 FILLER_44_401 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_4 FILLER_45_126 ();
 sg13g2_fill_2 FILLER_45_130 ();
 sg13g2_decap_4 FILLER_45_155 ();
 sg13g2_fill_2 FILLER_45_204 ();
 sg13g2_fill_1 FILLER_45_215 ();
 sg13g2_decap_8 FILLER_45_292 ();
 sg13g2_decap_8 FILLER_45_299 ();
 sg13g2_decap_8 FILLER_45_306 ();
 sg13g2_decap_8 FILLER_45_313 ();
 sg13g2_decap_8 FILLER_45_320 ();
 sg13g2_decap_4 FILLER_45_341 ();
 sg13g2_decap_8 FILLER_45_397 ();
 sg13g2_decap_4 FILLER_45_404 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_4 FILLER_46_133 ();
 sg13g2_fill_2 FILLER_46_137 ();
 sg13g2_decap_8 FILLER_46_143 ();
 sg13g2_fill_1 FILLER_46_150 ();
 sg13g2_decap_4 FILLER_46_160 ();
 sg13g2_fill_1 FILLER_46_164 ();
 sg13g2_fill_2 FILLER_46_178 ();
 sg13g2_decap_4 FILLER_46_227 ();
 sg13g2_fill_1 FILLER_46_231 ();
 sg13g2_fill_2 FILLER_46_251 ();
 sg13g2_fill_2 FILLER_46_264 ();
 sg13g2_fill_1 FILLER_46_266 ();
 sg13g2_fill_1 FILLER_46_274 ();
 sg13g2_decap_8 FILLER_46_306 ();
 sg13g2_decap_8 FILLER_46_313 ();
 sg13g2_decap_8 FILLER_46_320 ();
 sg13g2_fill_2 FILLER_46_327 ();
 sg13g2_decap_8 FILLER_46_394 ();
 sg13g2_decap_8 FILLER_46_401 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_fill_2 FILLER_47_126 ();
 sg13g2_decap_4 FILLER_47_164 ();
 sg13g2_fill_2 FILLER_47_173 ();
 sg13g2_fill_1 FILLER_47_185 ();
 sg13g2_decap_8 FILLER_47_222 ();
 sg13g2_decap_8 FILLER_47_229 ();
 sg13g2_fill_2 FILLER_47_236 ();
 sg13g2_fill_1 FILLER_47_238 ();
 sg13g2_fill_1 FILLER_47_256 ();
 sg13g2_decap_8 FILLER_47_310 ();
 sg13g2_decap_8 FILLER_47_317 ();
 sg13g2_decap_8 FILLER_47_324 ();
 sg13g2_decap_8 FILLER_47_331 ();
 sg13g2_fill_2 FILLER_47_338 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_fill_2 FILLER_47_406 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_fill_2 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_fill_1 FILLER_48_161 ();
 sg13g2_decap_4 FILLER_48_219 ();
 sg13g2_fill_1 FILLER_48_254 ();
 sg13g2_decap_8 FILLER_48_298 ();
 sg13g2_decap_8 FILLER_48_305 ();
 sg13g2_decap_8 FILLER_48_312 ();
 sg13g2_decap_8 FILLER_48_319 ();
 sg13g2_decap_4 FILLER_48_326 ();
 sg13g2_decap_8 FILLER_48_339 ();
 sg13g2_decap_4 FILLER_48_346 ();
 sg13g2_fill_2 FILLER_48_367 ();
 sg13g2_decap_8 FILLER_48_381 ();
 sg13g2_decap_8 FILLER_48_388 ();
 sg13g2_decap_8 FILLER_48_395 ();
 sg13g2_decap_8 FILLER_48_402 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_fill_2 FILLER_49_133 ();
 sg13g2_fill_1 FILLER_49_135 ();
 sg13g2_fill_2 FILLER_49_162 ();
 sg13g2_fill_1 FILLER_49_190 ();
 sg13g2_decap_4 FILLER_49_209 ();
 sg13g2_fill_2 FILLER_49_287 ();
 sg13g2_fill_1 FILLER_49_297 ();
 sg13g2_decap_4 FILLER_49_307 ();
 sg13g2_fill_2 FILLER_49_353 ();
 sg13g2_fill_1 FILLER_49_355 ();
 sg13g2_decap_8 FILLER_49_391 ();
 sg13g2_decap_8 FILLER_49_398 ();
 sg13g2_decap_4 FILLER_49_405 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_fill_2 FILLER_50_133 ();
 sg13g2_fill_1 FILLER_50_135 ();
 sg13g2_decap_4 FILLER_50_140 ();
 sg13g2_fill_2 FILLER_50_174 ();
 sg13g2_fill_1 FILLER_50_238 ();
 sg13g2_fill_2 FILLER_50_254 ();
 sg13g2_fill_1 FILLER_50_256 ();
 sg13g2_fill_1 FILLER_50_271 ();
 sg13g2_fill_1 FILLER_50_290 ();
 sg13g2_decap_4 FILLER_50_296 ();
 sg13g2_fill_1 FILLER_50_359 ();
 sg13g2_decap_8 FILLER_50_396 ();
 sg13g2_decap_4 FILLER_50_403 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_4 FILLER_51_119 ();
 sg13g2_fill_2 FILLER_51_123 ();
 sg13g2_fill_2 FILLER_51_151 ();
 sg13g2_fill_1 FILLER_51_172 ();
 sg13g2_decap_8 FILLER_51_186 ();
 sg13g2_decap_8 FILLER_51_193 ();
 sg13g2_fill_2 FILLER_51_200 ();
 sg13g2_fill_1 FILLER_51_202 ();
 sg13g2_fill_2 FILLER_51_216 ();
 sg13g2_decap_8 FILLER_51_249 ();
 sg13g2_fill_2 FILLER_51_256 ();
 sg13g2_decap_8 FILLER_51_263 ();
 sg13g2_fill_2 FILLER_51_270 ();
 sg13g2_fill_1 FILLER_51_276 ();
 sg13g2_decap_8 FILLER_51_296 ();
 sg13g2_fill_1 FILLER_51_303 ();
 sg13g2_decap_8 FILLER_51_400 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_decap_4 FILLER_52_133 ();
 sg13g2_fill_2 FILLER_52_137 ();
 sg13g2_fill_1 FILLER_52_178 ();
 sg13g2_fill_2 FILLER_52_224 ();
 sg13g2_fill_1 FILLER_52_246 ();
 sg13g2_fill_1 FILLER_52_275 ();
 sg13g2_fill_1 FILLER_52_294 ();
 sg13g2_fill_2 FILLER_52_300 ();
 sg13g2_fill_1 FILLER_52_356 ();
 sg13g2_decap_8 FILLER_52_400 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_4 FILLER_53_126 ();
 sg13g2_decap_4 FILLER_53_172 ();
 sg13g2_fill_1 FILLER_53_176 ();
 sg13g2_fill_1 FILLER_53_210 ();
 sg13g2_fill_1 FILLER_53_268 ();
 sg13g2_fill_1 FILLER_53_312 ();
 sg13g2_fill_2 FILLER_53_322 ();
 sg13g2_fill_1 FILLER_53_356 ();
 sg13g2_decap_8 FILLER_53_392 ();
 sg13g2_decap_8 FILLER_53_399 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_fill_2 FILLER_54_126 ();
 sg13g2_fill_1 FILLER_54_157 ();
 sg13g2_fill_1 FILLER_54_210 ();
 sg13g2_fill_2 FILLER_54_225 ();
 sg13g2_fill_2 FILLER_54_255 ();
 sg13g2_fill_2 FILLER_54_270 ();
 sg13g2_fill_1 FILLER_54_358 ();
 sg13g2_decap_8 FILLER_54_392 ();
 sg13g2_decap_8 FILLER_54_399 ();
 sg13g2_fill_2 FILLER_54_406 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_fill_2 FILLER_55_126 ();
 sg13g2_fill_2 FILLER_55_164 ();
 sg13g2_fill_1 FILLER_55_166 ();
 sg13g2_fill_1 FILLER_55_181 ();
 sg13g2_fill_2 FILLER_55_191 ();
 sg13g2_decap_4 FILLER_55_207 ();
 sg13g2_fill_2 FILLER_55_211 ();
 sg13g2_decap_4 FILLER_55_248 ();
 sg13g2_fill_2 FILLER_55_252 ();
 sg13g2_fill_1 FILLER_55_283 ();
 sg13g2_fill_2 FILLER_55_296 ();
 sg13g2_decap_8 FILLER_55_382 ();
 sg13g2_decap_8 FILLER_55_389 ();
 sg13g2_decap_8 FILLER_55_396 ();
 sg13g2_decap_4 FILLER_55_403 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_fill_2 FILLER_56_162 ();
 sg13g2_fill_1 FILLER_56_164 ();
 sg13g2_fill_2 FILLER_56_190 ();
 sg13g2_fill_1 FILLER_56_192 ();
 sg13g2_decap_4 FILLER_56_244 ();
 sg13g2_fill_2 FILLER_56_268 ();
 sg13g2_fill_2 FILLER_56_296 ();
 sg13g2_fill_2 FILLER_56_361 ();
 sg13g2_fill_1 FILLER_56_363 ();
 sg13g2_decap_8 FILLER_56_373 ();
 sg13g2_decap_8 FILLER_56_380 ();
 sg13g2_decap_8 FILLER_56_387 ();
 sg13g2_decap_8 FILLER_56_394 ();
 sg13g2_decap_8 FILLER_56_401 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_fill_2 FILLER_57_119 ();
 sg13g2_decap_4 FILLER_57_156 ();
 sg13g2_fill_1 FILLER_57_160 ();
 sg13g2_fill_1 FILLER_57_187 ();
 sg13g2_decap_8 FILLER_57_224 ();
 sg13g2_decap_8 FILLER_57_231 ();
 sg13g2_decap_4 FILLER_57_251 ();
 sg13g2_fill_2 FILLER_57_255 ();
 sg13g2_decap_4 FILLER_57_262 ();
 sg13g2_fill_2 FILLER_57_266 ();
 sg13g2_fill_2 FILLER_57_276 ();
 sg13g2_fill_1 FILLER_57_278 ();
 sg13g2_decap_8 FILLER_57_283 ();
 sg13g2_decap_4 FILLER_57_290 ();
 sg13g2_fill_2 FILLER_57_355 ();
 sg13g2_fill_1 FILLER_57_357 ();
 sg13g2_decap_8 FILLER_57_371 ();
 sg13g2_decap_8 FILLER_57_378 ();
 sg13g2_decap_8 FILLER_57_385 ();
 sg13g2_decap_8 FILLER_57_392 ();
 sg13g2_decap_8 FILLER_57_399 ();
 sg13g2_fill_2 FILLER_57_406 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_fill_2 FILLER_58_159 ();
 sg13g2_decap_8 FILLER_58_200 ();
 sg13g2_fill_1 FILLER_58_207 ();
 sg13g2_decap_8 FILLER_58_225 ();
 sg13g2_decap_8 FILLER_58_232 ();
 sg13g2_decap_8 FILLER_58_239 ();
 sg13g2_decap_8 FILLER_58_246 ();
 sg13g2_fill_1 FILLER_58_258 ();
 sg13g2_fill_2 FILLER_58_324 ();
 sg13g2_fill_1 FILLER_58_326 ();
 sg13g2_decap_8 FILLER_58_367 ();
 sg13g2_decap_8 FILLER_58_374 ();
 sg13g2_decap_8 FILLER_58_381 ();
 sg13g2_decap_8 FILLER_58_388 ();
 sg13g2_decap_8 FILLER_58_395 ();
 sg13g2_decap_8 FILLER_58_402 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_4 FILLER_59_133 ();
 sg13g2_fill_2 FILLER_59_137 ();
 sg13g2_fill_2 FILLER_59_185 ();
 sg13g2_fill_1 FILLER_59_187 ();
 sg13g2_decap_8 FILLER_59_211 ();
 sg13g2_decap_8 FILLER_59_218 ();
 sg13g2_fill_2 FILLER_59_225 ();
 sg13g2_fill_1 FILLER_59_239 ();
 sg13g2_decap_4 FILLER_59_263 ();
 sg13g2_fill_2 FILLER_59_267 ();
 sg13g2_decap_4 FILLER_59_274 ();
 sg13g2_decap_4 FILLER_59_282 ();
 sg13g2_fill_1 FILLER_59_292 ();
 sg13g2_decap_8 FILLER_59_356 ();
 sg13g2_decap_8 FILLER_59_363 ();
 sg13g2_decap_8 FILLER_59_370 ();
 sg13g2_decap_8 FILLER_59_377 ();
 sg13g2_decap_8 FILLER_59_384 ();
 sg13g2_decap_8 FILLER_59_391 ();
 sg13g2_decap_8 FILLER_59_398 ();
 sg13g2_decap_4 FILLER_59_405 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_decap_8 FILLER_60_133 ();
 sg13g2_decap_8 FILLER_60_140 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_decap_8 FILLER_60_154 ();
 sg13g2_decap_8 FILLER_60_161 ();
 sg13g2_decap_8 FILLER_60_168 ();
 sg13g2_fill_2 FILLER_60_175 ();
 sg13g2_fill_1 FILLER_60_177 ();
 sg13g2_fill_2 FILLER_60_186 ();
 sg13g2_fill_1 FILLER_60_188 ();
 sg13g2_decap_4 FILLER_60_215 ();
 sg13g2_fill_1 FILLER_60_219 ();
 sg13g2_decap_4 FILLER_60_277 ();
 sg13g2_decap_8 FILLER_60_285 ();
 sg13g2_fill_2 FILLER_60_292 ();
 sg13g2_decap_8 FILLER_60_365 ();
 sg13g2_decap_8 FILLER_60_372 ();
 sg13g2_decap_8 FILLER_60_379 ();
 sg13g2_decap_8 FILLER_60_386 ();
 sg13g2_decap_8 FILLER_60_393 ();
 sg13g2_decap_8 FILLER_60_400 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_decap_8 FILLER_61_133 ();
 sg13g2_decap_8 FILLER_61_140 ();
 sg13g2_fill_1 FILLER_61_147 ();
 sg13g2_fill_1 FILLER_61_177 ();
 sg13g2_fill_2 FILLER_61_223 ();
 sg13g2_fill_2 FILLER_61_237 ();
 sg13g2_fill_1 FILLER_61_239 ();
 sg13g2_fill_1 FILLER_61_343 ();
 sg13g2_decap_8 FILLER_61_375 ();
 sg13g2_decap_8 FILLER_61_382 ();
 sg13g2_decap_8 FILLER_61_389 ();
 sg13g2_decap_8 FILLER_61_396 ();
 sg13g2_decap_4 FILLER_61_403 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_fill_1 FILLER_62_133 ();
 sg13g2_decap_4 FILLER_62_164 ();
 sg13g2_fill_2 FILLER_62_178 ();
 sg13g2_fill_1 FILLER_62_194 ();
 sg13g2_decap_4 FILLER_62_214 ();
 sg13g2_decap_4 FILLER_62_240 ();
 sg13g2_fill_2 FILLER_62_264 ();
 sg13g2_fill_1 FILLER_62_266 ();
 sg13g2_fill_2 FILLER_62_297 ();
 sg13g2_fill_1 FILLER_62_359 ();
 sg13g2_decap_8 FILLER_62_373 ();
 sg13g2_decap_8 FILLER_62_380 ();
 sg13g2_decap_8 FILLER_62_387 ();
 sg13g2_decap_8 FILLER_62_394 ();
 sg13g2_decap_8 FILLER_62_401 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_fill_2 FILLER_63_126 ();
 sg13g2_fill_2 FILLER_63_214 ();
 sg13g2_fill_1 FILLER_63_216 ();
 sg13g2_decap_8 FILLER_63_226 ();
 sg13g2_fill_2 FILLER_63_233 ();
 sg13g2_decap_4 FILLER_63_247 ();
 sg13g2_decap_4 FILLER_63_273 ();
 sg13g2_fill_2 FILLER_63_281 ();
 sg13g2_fill_2 FILLER_63_292 ();
 sg13g2_fill_1 FILLER_63_308 ();
 sg13g2_decap_8 FILLER_63_367 ();
 sg13g2_decap_8 FILLER_63_374 ();
 sg13g2_decap_8 FILLER_63_381 ();
 sg13g2_decap_8 FILLER_63_388 ();
 sg13g2_decap_8 FILLER_63_395 ();
 sg13g2_decap_8 FILLER_63_402 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_fill_1 FILLER_64_126 ();
 sg13g2_fill_1 FILLER_64_198 ();
 sg13g2_fill_2 FILLER_64_225 ();
 sg13g2_fill_1 FILLER_64_227 ();
 sg13g2_fill_1 FILLER_64_236 ();
 sg13g2_fill_2 FILLER_64_242 ();
 sg13g2_fill_1 FILLER_64_254 ();
 sg13g2_decap_4 FILLER_64_259 ();
 sg13g2_fill_1 FILLER_64_263 ();
 sg13g2_fill_2 FILLER_64_276 ();
 sg13g2_fill_1 FILLER_64_317 ();
 sg13g2_decap_8 FILLER_64_363 ();
 sg13g2_decap_8 FILLER_64_370 ();
 sg13g2_decap_8 FILLER_64_377 ();
 sg13g2_decap_8 FILLER_64_384 ();
 sg13g2_decap_8 FILLER_64_391 ();
 sg13g2_decap_8 FILLER_64_398 ();
 sg13g2_decap_4 FILLER_64_405 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_4 FILLER_65_133 ();
 sg13g2_fill_2 FILLER_65_164 ();
 sg13g2_fill_1 FILLER_65_166 ();
 sg13g2_fill_1 FILLER_65_198 ();
 sg13g2_fill_2 FILLER_65_223 ();
 sg13g2_fill_2 FILLER_65_238 ();
 sg13g2_fill_1 FILLER_65_240 ();
 sg13g2_fill_1 FILLER_65_252 ();
 sg13g2_fill_1 FILLER_65_259 ();
 sg13g2_fill_1 FILLER_65_291 ();
 sg13g2_fill_1 FILLER_65_337 ();
 sg13g2_decap_8 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_371 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_decap_8 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_399 ();
 sg13g2_fill_2 FILLER_65_406 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_fill_2 FILLER_66_140 ();
 sg13g2_fill_1 FILLER_66_142 ();
 sg13g2_fill_1 FILLER_66_153 ();
 sg13g2_decap_8 FILLER_66_182 ();
 sg13g2_decap_4 FILLER_66_189 ();
 sg13g2_fill_2 FILLER_66_193 ();
 sg13g2_fill_2 FILLER_66_199 ();
 sg13g2_fill_1 FILLER_66_201 ();
 sg13g2_fill_1 FILLER_66_208 ();
 sg13g2_fill_2 FILLER_66_222 ();
 sg13g2_fill_1 FILLER_66_244 ();
 sg13g2_fill_1 FILLER_66_305 ();
 sg13g2_decap_8 FILLER_66_372 ();
 sg13g2_decap_8 FILLER_66_379 ();
 sg13g2_decap_8 FILLER_66_386 ();
 sg13g2_decap_8 FILLER_66_393 ();
 sg13g2_decap_8 FILLER_66_400 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_4 FILLER_67_140 ();
 sg13g2_fill_2 FILLER_67_144 ();
 sg13g2_fill_2 FILLER_67_167 ();
 sg13g2_fill_1 FILLER_67_169 ();
 sg13g2_decap_4 FILLER_67_193 ();
 sg13g2_fill_2 FILLER_67_197 ();
 sg13g2_fill_2 FILLER_67_225 ();
 sg13g2_fill_1 FILLER_67_253 ();
 sg13g2_fill_1 FILLER_67_347 ();
 sg13g2_decap_8 FILLER_67_374 ();
 sg13g2_decap_8 FILLER_67_381 ();
 sg13g2_decap_8 FILLER_67_388 ();
 sg13g2_decap_8 FILLER_67_395 ();
 sg13g2_decap_8 FILLER_67_402 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_4 FILLER_68_126 ();
 sg13g2_fill_2 FILLER_68_191 ();
 sg13g2_fill_1 FILLER_68_227 ();
 sg13g2_fill_1 FILLER_68_266 ();
 sg13g2_decap_8 FILLER_68_395 ();
 sg13g2_decap_8 FILLER_68_402 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_fill_2 FILLER_69_133 ();
 sg13g2_fill_2 FILLER_69_251 ();
 sg13g2_fill_1 FILLER_69_253 ();
 sg13g2_fill_1 FILLER_69_262 ();
 sg13g2_decap_8 FILLER_69_267 ();
 sg13g2_fill_2 FILLER_69_274 ();
 sg13g2_fill_1 FILLER_69_276 ();
 sg13g2_decap_4 FILLER_69_281 ();
 sg13g2_fill_2 FILLER_69_329 ();
 sg13g2_fill_1 FILLER_69_331 ();
 sg13g2_fill_1 FILLER_69_371 ();
 sg13g2_decap_8 FILLER_69_385 ();
 sg13g2_decap_8 FILLER_69_392 ();
 sg13g2_decap_8 FILLER_69_399 ();
 sg13g2_fill_2 FILLER_69_406 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_4 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_199 ();
 sg13g2_decap_4 FILLER_70_206 ();
 sg13g2_fill_2 FILLER_70_253 ();
 sg13g2_fill_1 FILLER_70_255 ();
 sg13g2_decap_8 FILLER_70_276 ();
 sg13g2_fill_1 FILLER_70_331 ();
 sg13g2_fill_1 FILLER_70_336 ();
 sg13g2_decap_8 FILLER_70_341 ();
 sg13g2_fill_2 FILLER_70_348 ();
 sg13g2_fill_2 FILLER_70_355 ();
 sg13g2_decap_8 FILLER_70_370 ();
 sg13g2_decap_8 FILLER_70_377 ();
 sg13g2_decap_8 FILLER_70_384 ();
 sg13g2_decap_8 FILLER_70_391 ();
 sg13g2_decap_8 FILLER_70_398 ();
 sg13g2_decap_4 FILLER_70_405 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_fill_1 FILLER_71_147 ();
 sg13g2_fill_1 FILLER_71_158 ();
 sg13g2_fill_2 FILLER_71_168 ();
 sg13g2_fill_1 FILLER_71_170 ();
 sg13g2_decap_8 FILLER_71_186 ();
 sg13g2_decap_8 FILLER_71_203 ();
 sg13g2_decap_8 FILLER_71_210 ();
 sg13g2_decap_4 FILLER_71_217 ();
 sg13g2_fill_1 FILLER_71_266 ();
 sg13g2_decap_8 FILLER_71_329 ();
 sg13g2_decap_8 FILLER_71_336 ();
 sg13g2_decap_8 FILLER_71_343 ();
 sg13g2_decap_4 FILLER_71_350 ();
 sg13g2_fill_1 FILLER_71_354 ();
 sg13g2_decap_8 FILLER_71_358 ();
 sg13g2_decap_8 FILLER_71_365 ();
 sg13g2_decap_8 FILLER_71_372 ();
 sg13g2_decap_8 FILLER_71_379 ();
 sg13g2_decap_8 FILLER_71_386 ();
 sg13g2_decap_8 FILLER_71_393 ();
 sg13g2_decap_8 FILLER_71_400 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_fill_2 FILLER_72_166 ();
 sg13g2_fill_2 FILLER_72_210 ();
 sg13g2_fill_2 FILLER_72_260 ();
 sg13g2_decap_8 FILLER_72_345 ();
 sg13g2_decap_8 FILLER_72_352 ();
 sg13g2_decap_8 FILLER_72_359 ();
 sg13g2_decap_8 FILLER_72_366 ();
 sg13g2_decap_8 FILLER_72_373 ();
 sg13g2_decap_8 FILLER_72_380 ();
 sg13g2_decap_8 FILLER_72_387 ();
 sg13g2_decap_8 FILLER_72_394 ();
 sg13g2_decap_8 FILLER_72_401 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_fill_1 FILLER_73_166 ();
 sg13g2_fill_1 FILLER_73_193 ();
 sg13g2_fill_1 FILLER_73_262 ();
 sg13g2_fill_2 FILLER_73_278 ();
 sg13g2_fill_2 FILLER_73_302 ();
 sg13g2_decap_8 FILLER_73_344 ();
 sg13g2_decap_8 FILLER_73_351 ();
 sg13g2_decap_8 FILLER_73_358 ();
 sg13g2_decap_8 FILLER_73_365 ();
 sg13g2_decap_8 FILLER_73_372 ();
 sg13g2_decap_8 FILLER_73_379 ();
 sg13g2_decap_8 FILLER_73_386 ();
 sg13g2_decap_8 FILLER_73_393 ();
 sg13g2_decap_8 FILLER_73_400 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_4 FILLER_74_140 ();
 sg13g2_fill_1 FILLER_74_144 ();
 sg13g2_fill_1 FILLER_74_159 ();
 sg13g2_fill_2 FILLER_74_169 ();
 sg13g2_fill_1 FILLER_74_171 ();
 sg13g2_fill_1 FILLER_74_182 ();
 sg13g2_fill_2 FILLER_74_223 ();
 sg13g2_fill_2 FILLER_74_239 ();
 sg13g2_decap_8 FILLER_74_337 ();
 sg13g2_decap_8 FILLER_74_344 ();
 sg13g2_decap_8 FILLER_74_351 ();
 sg13g2_decap_8 FILLER_74_358 ();
 sg13g2_decap_8 FILLER_74_365 ();
 sg13g2_decap_8 FILLER_74_372 ();
 sg13g2_decap_8 FILLER_74_379 ();
 sg13g2_decap_8 FILLER_74_386 ();
 sg13g2_decap_8 FILLER_74_393 ();
 sg13g2_decap_8 FILLER_74_400 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_4 FILLER_75_154 ();
 sg13g2_fill_1 FILLER_75_158 ();
 sg13g2_decap_8 FILLER_75_163 ();
 sg13g2_fill_2 FILLER_75_170 ();
 sg13g2_fill_2 FILLER_75_181 ();
 sg13g2_fill_1 FILLER_75_183 ();
 sg13g2_decap_4 FILLER_75_192 ();
 sg13g2_fill_1 FILLER_75_196 ();
 sg13g2_fill_2 FILLER_75_210 ();
 sg13g2_fill_1 FILLER_75_287 ();
 sg13g2_fill_2 FILLER_75_314 ();
 sg13g2_decap_8 FILLER_75_328 ();
 sg13g2_decap_8 FILLER_75_335 ();
 sg13g2_decap_8 FILLER_75_342 ();
 sg13g2_decap_8 FILLER_75_349 ();
 sg13g2_decap_8 FILLER_75_356 ();
 sg13g2_decap_8 FILLER_75_363 ();
 sg13g2_decap_8 FILLER_75_370 ();
 sg13g2_decap_8 FILLER_75_377 ();
 sg13g2_decap_8 FILLER_75_384 ();
 sg13g2_decap_8 FILLER_75_391 ();
 sg13g2_decap_8 FILLER_75_398 ();
 sg13g2_decap_4 FILLER_75_405 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_fill_2 FILLER_76_175 ();
 sg13g2_fill_1 FILLER_76_177 ();
 sg13g2_decap_8 FILLER_76_186 ();
 sg13g2_decap_8 FILLER_76_193 ();
 sg13g2_decap_8 FILLER_76_200 ();
 sg13g2_decap_8 FILLER_76_207 ();
 sg13g2_decap_8 FILLER_76_214 ();
 sg13g2_fill_2 FILLER_76_221 ();
 sg13g2_fill_1 FILLER_76_227 ();
 sg13g2_fill_2 FILLER_76_243 ();
 sg13g2_fill_2 FILLER_76_285 ();
 sg13g2_decap_8 FILLER_76_339 ();
 sg13g2_decap_8 FILLER_76_346 ();
 sg13g2_decap_8 FILLER_76_353 ();
 sg13g2_decap_8 FILLER_76_360 ();
 sg13g2_decap_8 FILLER_76_367 ();
 sg13g2_decap_8 FILLER_76_374 ();
 sg13g2_decap_8 FILLER_76_381 ();
 sg13g2_decap_8 FILLER_76_388 ();
 sg13g2_decap_8 FILLER_76_395 ();
 sg13g2_decap_8 FILLER_76_402 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_fill_2 FILLER_77_217 ();
 sg13g2_fill_1 FILLER_77_250 ();
 sg13g2_decap_8 FILLER_77_351 ();
 sg13g2_decap_8 FILLER_77_358 ();
 sg13g2_decap_8 FILLER_77_365 ();
 sg13g2_decap_8 FILLER_77_372 ();
 sg13g2_decap_8 FILLER_77_379 ();
 sg13g2_decap_8 FILLER_77_386 ();
 sg13g2_decap_8 FILLER_77_393 ();
 sg13g2_decap_8 FILLER_77_400 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_fill_2 FILLER_78_224 ();
 sg13g2_fill_2 FILLER_78_234 ();
 sg13g2_fill_1 FILLER_78_236 ();
 sg13g2_fill_1 FILLER_78_277 ();
 sg13g2_decap_8 FILLER_78_282 ();
 sg13g2_fill_2 FILLER_78_289 ();
 sg13g2_fill_1 FILLER_78_291 ();
 sg13g2_fill_1 FILLER_78_296 ();
 sg13g2_decap_8 FILLER_78_340 ();
 sg13g2_decap_8 FILLER_78_347 ();
 sg13g2_decap_8 FILLER_78_354 ();
 sg13g2_decap_8 FILLER_78_361 ();
 sg13g2_decap_8 FILLER_78_368 ();
 sg13g2_decap_8 FILLER_78_375 ();
 sg13g2_decap_8 FILLER_78_382 ();
 sg13g2_decap_8 FILLER_78_389 ();
 sg13g2_decap_8 FILLER_78_396 ();
 sg13g2_decap_4 FILLER_78_403 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_4 FILLER_79_224 ();
 sg13g2_fill_2 FILLER_79_228 ();
 sg13g2_fill_2 FILLER_79_265 ();
 sg13g2_fill_2 FILLER_79_293 ();
 sg13g2_fill_1 FILLER_79_295 ();
 sg13g2_fill_1 FILLER_79_312 ();
 sg13g2_fill_2 FILLER_79_332 ();
 sg13g2_fill_1 FILLER_79_334 ();
 sg13g2_decap_8 FILLER_79_344 ();
 sg13g2_decap_8 FILLER_79_351 ();
 sg13g2_decap_8 FILLER_79_358 ();
 sg13g2_decap_8 FILLER_79_365 ();
 sg13g2_decap_8 FILLER_79_372 ();
 sg13g2_decap_8 FILLER_79_379 ();
 sg13g2_decap_8 FILLER_79_386 ();
 sg13g2_decap_8 FILLER_79_393 ();
 sg13g2_decap_8 FILLER_79_400 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_decap_8 FILLER_80_77 ();
 sg13g2_decap_8 FILLER_80_84 ();
 sg13g2_decap_8 FILLER_80_91 ();
 sg13g2_decap_8 FILLER_80_98 ();
 sg13g2_decap_8 FILLER_80_105 ();
 sg13g2_decap_8 FILLER_80_112 ();
 sg13g2_decap_8 FILLER_80_119 ();
 sg13g2_decap_8 FILLER_80_126 ();
 sg13g2_decap_8 FILLER_80_133 ();
 sg13g2_decap_8 FILLER_80_140 ();
 sg13g2_decap_8 FILLER_80_147 ();
 sg13g2_decap_8 FILLER_80_154 ();
 sg13g2_decap_8 FILLER_80_161 ();
 sg13g2_decap_8 FILLER_80_168 ();
 sg13g2_decap_8 FILLER_80_175 ();
 sg13g2_fill_2 FILLER_80_182 ();
 sg13g2_decap_4 FILLER_80_188 ();
 sg13g2_decap_4 FILLER_80_196 ();
 sg13g2_decap_4 FILLER_80_204 ();
 sg13g2_decap_4 FILLER_80_212 ();
 sg13g2_decap_4 FILLER_80_220 ();
 sg13g2_decap_4 FILLER_80_228 ();
 sg13g2_decap_4 FILLER_80_236 ();
 sg13g2_decap_4 FILLER_80_244 ();
 sg13g2_fill_2 FILLER_80_261 ();
 sg13g2_fill_1 FILLER_80_263 ();
 sg13g2_fill_2 FILLER_80_269 ();
 sg13g2_fill_1 FILLER_80_271 ();
 sg13g2_fill_2 FILLER_80_277 ();
 sg13g2_fill_1 FILLER_80_279 ();
 sg13g2_fill_2 FILLER_80_285 ();
 sg13g2_fill_1 FILLER_80_287 ();
 sg13g2_fill_2 FILLER_80_293 ();
 sg13g2_fill_1 FILLER_80_295 ();
 sg13g2_fill_1 FILLER_80_305 ();
 sg13g2_fill_2 FILLER_80_322 ();
 sg13g2_decap_8 FILLER_80_341 ();
 sg13g2_decap_4 FILLER_80_348 ();
 sg13g2_fill_2 FILLER_80_357 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_decap_8 FILLER_80_365 ();
 sg13g2_decap_4 FILLER_80_372 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uo_out[0] = net15;
 assign uo_out[1] = net16;
 assign uo_out[2] = net17;
 assign uo_out[3] = net18;
 assign uo_out[4] = net19;
 assign uo_out[5] = net20;
 assign uo_out[6] = net21;
 assign uo_out[7] = net22;
endmodule

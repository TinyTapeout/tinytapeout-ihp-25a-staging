module tt_um_jamesrosssharp_1bitam (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire COMP_OUT;
 wire PWM_OUT;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire clknet_leaf_0_clk;
 wire \am_sdr0.I_out[0] ;
 wire \am_sdr0.I_out[1] ;
 wire \am_sdr0.I_out[2] ;
 wire \am_sdr0.I_out[3] ;
 wire \am_sdr0.I_out[4] ;
 wire \am_sdr0.I_out[5] ;
 wire \am_sdr0.I_out[6] ;
 wire \am_sdr0.I_out[7] ;
 wire \am_sdr0.Q_out[0] ;
 wire \am_sdr0.Q_out[1] ;
 wire \am_sdr0.Q_out[2] ;
 wire \am_sdr0.Q_out[3] ;
 wire \am_sdr0.Q_out[4] ;
 wire \am_sdr0.Q_out[5] ;
 wire \am_sdr0.Q_out[6] ;
 wire \am_sdr0.Q_out[7] ;
 wire \am_sdr0.am0.I_in[0] ;
 wire \am_sdr0.am0.I_in[1] ;
 wire \am_sdr0.am0.I_in[2] ;
 wire \am_sdr0.am0.I_in[3] ;
 wire \am_sdr0.am0.I_in[4] ;
 wire \am_sdr0.am0.I_in[5] ;
 wire \am_sdr0.am0.I_in[6] ;
 wire \am_sdr0.am0.I_in[7] ;
 wire \am_sdr0.am0.Q_in[0] ;
 wire \am_sdr0.am0.Q_in[1] ;
 wire \am_sdr0.am0.Q_in[2] ;
 wire \am_sdr0.am0.Q_in[3] ;
 wire \am_sdr0.am0.Q_in[4] ;
 wire \am_sdr0.am0.Q_in[5] ;
 wire \am_sdr0.am0.Q_in[6] ;
 wire \am_sdr0.am0.Q_in[7] ;
 wire \am_sdr0.am0.a[0] ;
 wire \am_sdr0.am0.a[10] ;
 wire \am_sdr0.am0.a[11] ;
 wire \am_sdr0.am0.a[12] ;
 wire \am_sdr0.am0.a[13] ;
 wire \am_sdr0.am0.a[14] ;
 wire \am_sdr0.am0.a[15] ;
 wire \am_sdr0.am0.a[1] ;
 wire \am_sdr0.am0.a[2] ;
 wire \am_sdr0.am0.a[3] ;
 wire \am_sdr0.am0.a[4] ;
 wire \am_sdr0.am0.a[5] ;
 wire \am_sdr0.am0.a[6] ;
 wire \am_sdr0.am0.a[7] ;
 wire \am_sdr0.am0.a[8] ;
 wire \am_sdr0.am0.a[9] ;
 wire \am_sdr0.am0.count2[0] ;
 wire \am_sdr0.am0.count2[1] ;
 wire \am_sdr0.am0.count2[2] ;
 wire \am_sdr0.am0.count2[3] ;
 wire \am_sdr0.am0.count[0] ;
 wire \am_sdr0.am0.count[1] ;
 wire \am_sdr0.am0.demod_out[10] ;
 wire \am_sdr0.am0.demod_out[11] ;
 wire \am_sdr0.am0.demod_out[12] ;
 wire \am_sdr0.am0.demod_out[13] ;
 wire \am_sdr0.am0.demod_out[14] ;
 wire \am_sdr0.am0.demod_out[15] ;
 wire \am_sdr0.am0.demod_out[8] ;
 wire \am_sdr0.am0.demod_out[9] ;
 wire \am_sdr0.am0.left[0] ;
 wire \am_sdr0.am0.left[1] ;
 wire \am_sdr0.am0.left[2] ;
 wire \am_sdr0.am0.left[3] ;
 wire \am_sdr0.am0.left[4] ;
 wire \am_sdr0.am0.left[5] ;
 wire \am_sdr0.am0.left[6] ;
 wire \am_sdr0.am0.left[7] ;
 wire \am_sdr0.am0.left[8] ;
 wire \am_sdr0.am0.left[9] ;
 wire \am_sdr0.am0.load_tick ;
 wire \am_sdr0.am0.m_count[0] ;
 wire \am_sdr0.am0.m_count[1] ;
 wire \am_sdr0.am0.m_count[2] ;
 wire \am_sdr0.am0.m_count[3] ;
 wire \am_sdr0.am0.multA[0] ;
 wire \am_sdr0.am0.multA[10] ;
 wire \am_sdr0.am0.multA[11] ;
 wire \am_sdr0.am0.multA[12] ;
 wire \am_sdr0.am0.multA[13] ;
 wire \am_sdr0.am0.multA[14] ;
 wire \am_sdr0.am0.multA[15] ;
 wire \am_sdr0.am0.multA[16] ;
 wire \am_sdr0.am0.multA[1] ;
 wire \am_sdr0.am0.multA[2] ;
 wire \am_sdr0.am0.multA[3] ;
 wire \am_sdr0.am0.multA[4] ;
 wire \am_sdr0.am0.multA[5] ;
 wire \am_sdr0.am0.multA[6] ;
 wire \am_sdr0.am0.multA[7] ;
 wire \am_sdr0.am0.multA[8] ;
 wire \am_sdr0.am0.multA[9] ;
 wire \am_sdr0.am0.multB[0] ;
 wire \am_sdr0.am0.multB[1] ;
 wire \am_sdr0.am0.multB[2] ;
 wire \am_sdr0.am0.multB[3] ;
 wire \am_sdr0.am0.multB[4] ;
 wire \am_sdr0.am0.multB[5] ;
 wire \am_sdr0.am0.multB[6] ;
 wire \am_sdr0.am0.multB[7] ;
 wire \am_sdr0.am0.q[0] ;
 wire \am_sdr0.am0.q[1] ;
 wire \am_sdr0.am0.q[2] ;
 wire \am_sdr0.am0.q[3] ;
 wire \am_sdr0.am0.q[4] ;
 wire \am_sdr0.am0.q[5] ;
 wire \am_sdr0.am0.q[6] ;
 wire \am_sdr0.am0.q[7] ;
 wire \am_sdr0.am0.r[0] ;
 wire \am_sdr0.am0.r[1] ;
 wire \am_sdr0.am0.r[2] ;
 wire \am_sdr0.am0.r[3] ;
 wire \am_sdr0.am0.r[4] ;
 wire \am_sdr0.am0.r[5] ;
 wire \am_sdr0.am0.r[6] ;
 wire \am_sdr0.am0.r[7] ;
 wire \am_sdr0.am0.r[9] ;
 wire \am_sdr0.am0.right[0] ;
 wire \am_sdr0.am0.right[1] ;
 wire \am_sdr0.am0.right[2] ;
 wire \am_sdr0.am0.right[3] ;
 wire \am_sdr0.am0.right[4] ;
 wire \am_sdr0.am0.right[5] ;
 wire \am_sdr0.am0.right[6] ;
 wire \am_sdr0.am0.right[7] ;
 wire \am_sdr0.am0.right[8] ;
 wire \am_sdr0.am0.right[9] ;
 wire \am_sdr0.am0.sqrt_done ;
 wire \am_sdr0.am0.sqrt_state[0] ;
 wire \am_sdr0.am0.sqrt_state[1] ;
 wire \am_sdr0.am0.state[0] ;
 wire \am_sdr0.am0.state[1] ;
 wire \am_sdr0.am0.state[2] ;
 wire \am_sdr0.am0.state[3] ;
 wire \am_sdr0.am0.state[4] ;
 wire \am_sdr0.am0.state[5] ;
 wire \am_sdr0.am0.state[6] ;
 wire \am_sdr0.am0.sum[0] ;
 wire \am_sdr0.am0.sum[10] ;
 wire \am_sdr0.am0.sum[11] ;
 wire \am_sdr0.am0.sum[12] ;
 wire \am_sdr0.am0.sum[13] ;
 wire \am_sdr0.am0.sum[14] ;
 wire \am_sdr0.am0.sum[15] ;
 wire \am_sdr0.am0.sum[16] ;
 wire \am_sdr0.am0.sum[1] ;
 wire \am_sdr0.am0.sum[2] ;
 wire \am_sdr0.am0.sum[3] ;
 wire \am_sdr0.am0.sum[4] ;
 wire \am_sdr0.am0.sum[5] ;
 wire \am_sdr0.am0.sum[6] ;
 wire \am_sdr0.am0.sum[7] ;
 wire \am_sdr0.am0.sum[8] ;
 wire \am_sdr0.am0.sum[9] ;
 wire \am_sdr0.cic0.comb1[0] ;
 wire \am_sdr0.cic0.comb1[10] ;
 wire \am_sdr0.cic0.comb1[11] ;
 wire \am_sdr0.cic0.comb1[12] ;
 wire \am_sdr0.cic0.comb1[13] ;
 wire \am_sdr0.cic0.comb1[14] ;
 wire \am_sdr0.cic0.comb1[15] ;
 wire \am_sdr0.cic0.comb1[16] ;
 wire \am_sdr0.cic0.comb1[17] ;
 wire \am_sdr0.cic0.comb1[18] ;
 wire \am_sdr0.cic0.comb1[19] ;
 wire \am_sdr0.cic0.comb1[1] ;
 wire \am_sdr0.cic0.comb1[2] ;
 wire \am_sdr0.cic0.comb1[3] ;
 wire \am_sdr0.cic0.comb1[4] ;
 wire \am_sdr0.cic0.comb1[5] ;
 wire \am_sdr0.cic0.comb1[6] ;
 wire \am_sdr0.cic0.comb1[7] ;
 wire \am_sdr0.cic0.comb1[8] ;
 wire \am_sdr0.cic0.comb1[9] ;
 wire \am_sdr0.cic0.comb1_in_del[0] ;
 wire \am_sdr0.cic0.comb1_in_del[10] ;
 wire \am_sdr0.cic0.comb1_in_del[11] ;
 wire \am_sdr0.cic0.comb1_in_del[12] ;
 wire \am_sdr0.cic0.comb1_in_del[13] ;
 wire \am_sdr0.cic0.comb1_in_del[14] ;
 wire \am_sdr0.cic0.comb1_in_del[15] ;
 wire \am_sdr0.cic0.comb1_in_del[16] ;
 wire \am_sdr0.cic0.comb1_in_del[17] ;
 wire \am_sdr0.cic0.comb1_in_del[18] ;
 wire \am_sdr0.cic0.comb1_in_del[19] ;
 wire \am_sdr0.cic0.comb1_in_del[1] ;
 wire \am_sdr0.cic0.comb1_in_del[2] ;
 wire \am_sdr0.cic0.comb1_in_del[3] ;
 wire \am_sdr0.cic0.comb1_in_del[4] ;
 wire \am_sdr0.cic0.comb1_in_del[5] ;
 wire \am_sdr0.cic0.comb1_in_del[6] ;
 wire \am_sdr0.cic0.comb1_in_del[7] ;
 wire \am_sdr0.cic0.comb1_in_del[8] ;
 wire \am_sdr0.cic0.comb1_in_del[9] ;
 wire \am_sdr0.cic0.comb2[0] ;
 wire \am_sdr0.cic0.comb2[10] ;
 wire \am_sdr0.cic0.comb2[11] ;
 wire \am_sdr0.cic0.comb2[12] ;
 wire \am_sdr0.cic0.comb2[13] ;
 wire \am_sdr0.cic0.comb2[14] ;
 wire \am_sdr0.cic0.comb2[15] ;
 wire \am_sdr0.cic0.comb2[16] ;
 wire \am_sdr0.cic0.comb2[17] ;
 wire \am_sdr0.cic0.comb2[18] ;
 wire \am_sdr0.cic0.comb2[19] ;
 wire \am_sdr0.cic0.comb2[1] ;
 wire \am_sdr0.cic0.comb2[2] ;
 wire \am_sdr0.cic0.comb2[3] ;
 wire \am_sdr0.cic0.comb2[4] ;
 wire \am_sdr0.cic0.comb2[5] ;
 wire \am_sdr0.cic0.comb2[6] ;
 wire \am_sdr0.cic0.comb2[7] ;
 wire \am_sdr0.cic0.comb2[8] ;
 wire \am_sdr0.cic0.comb2[9] ;
 wire \am_sdr0.cic0.comb2_in_del[0] ;
 wire \am_sdr0.cic0.comb2_in_del[10] ;
 wire \am_sdr0.cic0.comb2_in_del[11] ;
 wire \am_sdr0.cic0.comb2_in_del[12] ;
 wire \am_sdr0.cic0.comb2_in_del[13] ;
 wire \am_sdr0.cic0.comb2_in_del[14] ;
 wire \am_sdr0.cic0.comb2_in_del[15] ;
 wire \am_sdr0.cic0.comb2_in_del[16] ;
 wire \am_sdr0.cic0.comb2_in_del[17] ;
 wire \am_sdr0.cic0.comb2_in_del[18] ;
 wire \am_sdr0.cic0.comb2_in_del[19] ;
 wire \am_sdr0.cic0.comb2_in_del[1] ;
 wire \am_sdr0.cic0.comb2_in_del[2] ;
 wire \am_sdr0.cic0.comb2_in_del[3] ;
 wire \am_sdr0.cic0.comb2_in_del[4] ;
 wire \am_sdr0.cic0.comb2_in_del[5] ;
 wire \am_sdr0.cic0.comb2_in_del[6] ;
 wire \am_sdr0.cic0.comb2_in_del[7] ;
 wire \am_sdr0.cic0.comb2_in_del[8] ;
 wire \am_sdr0.cic0.comb2_in_del[9] ;
 wire \am_sdr0.cic0.comb3[12] ;
 wire \am_sdr0.cic0.comb3[13] ;
 wire \am_sdr0.cic0.comb3[14] ;
 wire \am_sdr0.cic0.comb3[15] ;
 wire \am_sdr0.cic0.comb3[16] ;
 wire \am_sdr0.cic0.comb3[17] ;
 wire \am_sdr0.cic0.comb3[18] ;
 wire \am_sdr0.cic0.comb3[19] ;
 wire \am_sdr0.cic0.comb3_in_del[0] ;
 wire \am_sdr0.cic0.comb3_in_del[10] ;
 wire \am_sdr0.cic0.comb3_in_del[11] ;
 wire \am_sdr0.cic0.comb3_in_del[12] ;
 wire \am_sdr0.cic0.comb3_in_del[13] ;
 wire \am_sdr0.cic0.comb3_in_del[14] ;
 wire \am_sdr0.cic0.comb3_in_del[15] ;
 wire \am_sdr0.cic0.comb3_in_del[16] ;
 wire \am_sdr0.cic0.comb3_in_del[17] ;
 wire \am_sdr0.cic0.comb3_in_del[18] ;
 wire \am_sdr0.cic0.comb3_in_del[19] ;
 wire \am_sdr0.cic0.comb3_in_del[1] ;
 wire \am_sdr0.cic0.comb3_in_del[2] ;
 wire \am_sdr0.cic0.comb3_in_del[3] ;
 wire \am_sdr0.cic0.comb3_in_del[4] ;
 wire \am_sdr0.cic0.comb3_in_del[5] ;
 wire \am_sdr0.cic0.comb3_in_del[6] ;
 wire \am_sdr0.cic0.comb3_in_del[7] ;
 wire \am_sdr0.cic0.comb3_in_del[8] ;
 wire \am_sdr0.cic0.comb3_in_del[9] ;
 wire \am_sdr0.cic0.count[0] ;
 wire \am_sdr0.cic0.count[1] ;
 wire \am_sdr0.cic0.count[2] ;
 wire \am_sdr0.cic0.count[3] ;
 wire \am_sdr0.cic0.count[4] ;
 wire \am_sdr0.cic0.count[5] ;
 wire \am_sdr0.cic0.count[6] ;
 wire \am_sdr0.cic0.count[7] ;
 wire \am_sdr0.cic0.integ1[0] ;
 wire \am_sdr0.cic0.integ1[10] ;
 wire \am_sdr0.cic0.integ1[11] ;
 wire \am_sdr0.cic0.integ1[12] ;
 wire \am_sdr0.cic0.integ1[13] ;
 wire \am_sdr0.cic0.integ1[14] ;
 wire \am_sdr0.cic0.integ1[15] ;
 wire \am_sdr0.cic0.integ1[16] ;
 wire \am_sdr0.cic0.integ1[17] ;
 wire \am_sdr0.cic0.integ1[18] ;
 wire \am_sdr0.cic0.integ1[19] ;
 wire \am_sdr0.cic0.integ1[1] ;
 wire \am_sdr0.cic0.integ1[20] ;
 wire \am_sdr0.cic0.integ1[21] ;
 wire \am_sdr0.cic0.integ1[22] ;
 wire \am_sdr0.cic0.integ1[23] ;
 wire \am_sdr0.cic0.integ1[24] ;
 wire \am_sdr0.cic0.integ1[25] ;
 wire \am_sdr0.cic0.integ1[2] ;
 wire \am_sdr0.cic0.integ1[3] ;
 wire \am_sdr0.cic0.integ1[4] ;
 wire \am_sdr0.cic0.integ1[5] ;
 wire \am_sdr0.cic0.integ1[6] ;
 wire \am_sdr0.cic0.integ1[7] ;
 wire \am_sdr0.cic0.integ1[8] ;
 wire \am_sdr0.cic0.integ1[9] ;
 wire \am_sdr0.cic0.integ2[0] ;
 wire \am_sdr0.cic0.integ2[10] ;
 wire \am_sdr0.cic0.integ2[11] ;
 wire \am_sdr0.cic0.integ2[12] ;
 wire \am_sdr0.cic0.integ2[13] ;
 wire \am_sdr0.cic0.integ2[14] ;
 wire \am_sdr0.cic0.integ2[15] ;
 wire \am_sdr0.cic0.integ2[16] ;
 wire \am_sdr0.cic0.integ2[17] ;
 wire \am_sdr0.cic0.integ2[18] ;
 wire \am_sdr0.cic0.integ2[19] ;
 wire \am_sdr0.cic0.integ2[1] ;
 wire \am_sdr0.cic0.integ2[20] ;
 wire \am_sdr0.cic0.integ2[21] ;
 wire \am_sdr0.cic0.integ2[22] ;
 wire \am_sdr0.cic0.integ2[2] ;
 wire \am_sdr0.cic0.integ2[3] ;
 wire \am_sdr0.cic0.integ2[4] ;
 wire \am_sdr0.cic0.integ2[5] ;
 wire \am_sdr0.cic0.integ2[6] ;
 wire \am_sdr0.cic0.integ2[7] ;
 wire \am_sdr0.cic0.integ2[8] ;
 wire \am_sdr0.cic0.integ2[9] ;
 wire \am_sdr0.cic0.integ3[0] ;
 wire \am_sdr0.cic0.integ3[10] ;
 wire \am_sdr0.cic0.integ3[11] ;
 wire \am_sdr0.cic0.integ3[12] ;
 wire \am_sdr0.cic0.integ3[13] ;
 wire \am_sdr0.cic0.integ3[14] ;
 wire \am_sdr0.cic0.integ3[15] ;
 wire \am_sdr0.cic0.integ3[16] ;
 wire \am_sdr0.cic0.integ3[17] ;
 wire \am_sdr0.cic0.integ3[18] ;
 wire \am_sdr0.cic0.integ3[19] ;
 wire \am_sdr0.cic0.integ3[1] ;
 wire \am_sdr0.cic0.integ3[2] ;
 wire \am_sdr0.cic0.integ3[3] ;
 wire \am_sdr0.cic0.integ3[4] ;
 wire \am_sdr0.cic0.integ3[5] ;
 wire \am_sdr0.cic0.integ3[6] ;
 wire \am_sdr0.cic0.integ3[7] ;
 wire \am_sdr0.cic0.integ3[8] ;
 wire \am_sdr0.cic0.integ3[9] ;
 wire \am_sdr0.cic0.integ_sample[0] ;
 wire \am_sdr0.cic0.integ_sample[10] ;
 wire \am_sdr0.cic0.integ_sample[11] ;
 wire \am_sdr0.cic0.integ_sample[12] ;
 wire \am_sdr0.cic0.integ_sample[13] ;
 wire \am_sdr0.cic0.integ_sample[14] ;
 wire \am_sdr0.cic0.integ_sample[15] ;
 wire \am_sdr0.cic0.integ_sample[16] ;
 wire \am_sdr0.cic0.integ_sample[17] ;
 wire \am_sdr0.cic0.integ_sample[18] ;
 wire \am_sdr0.cic0.integ_sample[19] ;
 wire \am_sdr0.cic0.integ_sample[1] ;
 wire \am_sdr0.cic0.integ_sample[2] ;
 wire \am_sdr0.cic0.integ_sample[3] ;
 wire \am_sdr0.cic0.integ_sample[4] ;
 wire \am_sdr0.cic0.integ_sample[5] ;
 wire \am_sdr0.cic0.integ_sample[6] ;
 wire \am_sdr0.cic0.integ_sample[7] ;
 wire \am_sdr0.cic0.integ_sample[8] ;
 wire \am_sdr0.cic0.integ_sample[9] ;
 wire \am_sdr0.cic0.out_tick ;
 wire \am_sdr0.cic0.sample ;
 wire \am_sdr0.cic0.x_out[10] ;
 wire \am_sdr0.cic0.x_out[11] ;
 wire \am_sdr0.cic0.x_out[12] ;
 wire \am_sdr0.cic0.x_out[13] ;
 wire \am_sdr0.cic0.x_out[14] ;
 wire \am_sdr0.cic0.x_out[15] ;
 wire \am_sdr0.cic0.x_out[8] ;
 wire \am_sdr0.cic0.x_out[9] ;
 wire \am_sdr0.cic1.comb1[0] ;
 wire \am_sdr0.cic1.comb1[10] ;
 wire \am_sdr0.cic1.comb1[11] ;
 wire \am_sdr0.cic1.comb1[12] ;
 wire \am_sdr0.cic1.comb1[13] ;
 wire \am_sdr0.cic1.comb1[14] ;
 wire \am_sdr0.cic1.comb1[15] ;
 wire \am_sdr0.cic1.comb1[16] ;
 wire \am_sdr0.cic1.comb1[17] ;
 wire \am_sdr0.cic1.comb1[18] ;
 wire \am_sdr0.cic1.comb1[19] ;
 wire \am_sdr0.cic1.comb1[1] ;
 wire \am_sdr0.cic1.comb1[2] ;
 wire \am_sdr0.cic1.comb1[3] ;
 wire \am_sdr0.cic1.comb1[4] ;
 wire \am_sdr0.cic1.comb1[5] ;
 wire \am_sdr0.cic1.comb1[6] ;
 wire \am_sdr0.cic1.comb1[7] ;
 wire \am_sdr0.cic1.comb1[8] ;
 wire \am_sdr0.cic1.comb1[9] ;
 wire \am_sdr0.cic1.comb1_in_del[0] ;
 wire \am_sdr0.cic1.comb1_in_del[10] ;
 wire \am_sdr0.cic1.comb1_in_del[11] ;
 wire \am_sdr0.cic1.comb1_in_del[12] ;
 wire \am_sdr0.cic1.comb1_in_del[13] ;
 wire \am_sdr0.cic1.comb1_in_del[14] ;
 wire \am_sdr0.cic1.comb1_in_del[15] ;
 wire \am_sdr0.cic1.comb1_in_del[16] ;
 wire \am_sdr0.cic1.comb1_in_del[17] ;
 wire \am_sdr0.cic1.comb1_in_del[18] ;
 wire \am_sdr0.cic1.comb1_in_del[19] ;
 wire \am_sdr0.cic1.comb1_in_del[1] ;
 wire \am_sdr0.cic1.comb1_in_del[2] ;
 wire \am_sdr0.cic1.comb1_in_del[3] ;
 wire \am_sdr0.cic1.comb1_in_del[4] ;
 wire \am_sdr0.cic1.comb1_in_del[5] ;
 wire \am_sdr0.cic1.comb1_in_del[6] ;
 wire \am_sdr0.cic1.comb1_in_del[7] ;
 wire \am_sdr0.cic1.comb1_in_del[8] ;
 wire \am_sdr0.cic1.comb1_in_del[9] ;
 wire \am_sdr0.cic1.comb2[0] ;
 wire \am_sdr0.cic1.comb2[10] ;
 wire \am_sdr0.cic1.comb2[11] ;
 wire \am_sdr0.cic1.comb2[12] ;
 wire \am_sdr0.cic1.comb2[13] ;
 wire \am_sdr0.cic1.comb2[14] ;
 wire \am_sdr0.cic1.comb2[15] ;
 wire \am_sdr0.cic1.comb2[16] ;
 wire \am_sdr0.cic1.comb2[17] ;
 wire \am_sdr0.cic1.comb2[18] ;
 wire \am_sdr0.cic1.comb2[19] ;
 wire \am_sdr0.cic1.comb2[1] ;
 wire \am_sdr0.cic1.comb2[2] ;
 wire \am_sdr0.cic1.comb2[3] ;
 wire \am_sdr0.cic1.comb2[4] ;
 wire \am_sdr0.cic1.comb2[5] ;
 wire \am_sdr0.cic1.comb2[6] ;
 wire \am_sdr0.cic1.comb2[7] ;
 wire \am_sdr0.cic1.comb2[8] ;
 wire \am_sdr0.cic1.comb2[9] ;
 wire \am_sdr0.cic1.comb2_in_del[0] ;
 wire \am_sdr0.cic1.comb2_in_del[10] ;
 wire \am_sdr0.cic1.comb2_in_del[11] ;
 wire \am_sdr0.cic1.comb2_in_del[12] ;
 wire \am_sdr0.cic1.comb2_in_del[13] ;
 wire \am_sdr0.cic1.comb2_in_del[14] ;
 wire \am_sdr0.cic1.comb2_in_del[15] ;
 wire \am_sdr0.cic1.comb2_in_del[16] ;
 wire \am_sdr0.cic1.comb2_in_del[17] ;
 wire \am_sdr0.cic1.comb2_in_del[18] ;
 wire \am_sdr0.cic1.comb2_in_del[19] ;
 wire \am_sdr0.cic1.comb2_in_del[1] ;
 wire \am_sdr0.cic1.comb2_in_del[2] ;
 wire \am_sdr0.cic1.comb2_in_del[3] ;
 wire \am_sdr0.cic1.comb2_in_del[4] ;
 wire \am_sdr0.cic1.comb2_in_del[5] ;
 wire \am_sdr0.cic1.comb2_in_del[6] ;
 wire \am_sdr0.cic1.comb2_in_del[7] ;
 wire \am_sdr0.cic1.comb2_in_del[8] ;
 wire \am_sdr0.cic1.comb2_in_del[9] ;
 wire \am_sdr0.cic1.comb3[12] ;
 wire \am_sdr0.cic1.comb3[13] ;
 wire \am_sdr0.cic1.comb3[14] ;
 wire \am_sdr0.cic1.comb3[15] ;
 wire \am_sdr0.cic1.comb3[16] ;
 wire \am_sdr0.cic1.comb3[17] ;
 wire \am_sdr0.cic1.comb3[18] ;
 wire \am_sdr0.cic1.comb3[19] ;
 wire \am_sdr0.cic1.comb3_in_del[0] ;
 wire \am_sdr0.cic1.comb3_in_del[10] ;
 wire \am_sdr0.cic1.comb3_in_del[11] ;
 wire \am_sdr0.cic1.comb3_in_del[12] ;
 wire \am_sdr0.cic1.comb3_in_del[13] ;
 wire \am_sdr0.cic1.comb3_in_del[14] ;
 wire \am_sdr0.cic1.comb3_in_del[15] ;
 wire \am_sdr0.cic1.comb3_in_del[16] ;
 wire \am_sdr0.cic1.comb3_in_del[17] ;
 wire \am_sdr0.cic1.comb3_in_del[18] ;
 wire \am_sdr0.cic1.comb3_in_del[19] ;
 wire \am_sdr0.cic1.comb3_in_del[1] ;
 wire \am_sdr0.cic1.comb3_in_del[2] ;
 wire \am_sdr0.cic1.comb3_in_del[3] ;
 wire \am_sdr0.cic1.comb3_in_del[4] ;
 wire \am_sdr0.cic1.comb3_in_del[5] ;
 wire \am_sdr0.cic1.comb3_in_del[6] ;
 wire \am_sdr0.cic1.comb3_in_del[7] ;
 wire \am_sdr0.cic1.comb3_in_del[8] ;
 wire \am_sdr0.cic1.comb3_in_del[9] ;
 wire \am_sdr0.cic1.count[0] ;
 wire \am_sdr0.cic1.count[1] ;
 wire \am_sdr0.cic1.count[2] ;
 wire \am_sdr0.cic1.count[3] ;
 wire \am_sdr0.cic1.count[4] ;
 wire \am_sdr0.cic1.count[5] ;
 wire \am_sdr0.cic1.count[6] ;
 wire \am_sdr0.cic1.count[7] ;
 wire \am_sdr0.cic1.integ1[0] ;
 wire \am_sdr0.cic1.integ1[10] ;
 wire \am_sdr0.cic1.integ1[11] ;
 wire \am_sdr0.cic1.integ1[12] ;
 wire \am_sdr0.cic1.integ1[13] ;
 wire \am_sdr0.cic1.integ1[14] ;
 wire \am_sdr0.cic1.integ1[15] ;
 wire \am_sdr0.cic1.integ1[16] ;
 wire \am_sdr0.cic1.integ1[17] ;
 wire \am_sdr0.cic1.integ1[18] ;
 wire \am_sdr0.cic1.integ1[19] ;
 wire \am_sdr0.cic1.integ1[1] ;
 wire \am_sdr0.cic1.integ1[20] ;
 wire \am_sdr0.cic1.integ1[21] ;
 wire \am_sdr0.cic1.integ1[22] ;
 wire \am_sdr0.cic1.integ1[23] ;
 wire \am_sdr0.cic1.integ1[24] ;
 wire \am_sdr0.cic1.integ1[25] ;
 wire \am_sdr0.cic1.integ1[2] ;
 wire \am_sdr0.cic1.integ1[3] ;
 wire \am_sdr0.cic1.integ1[4] ;
 wire \am_sdr0.cic1.integ1[5] ;
 wire \am_sdr0.cic1.integ1[6] ;
 wire \am_sdr0.cic1.integ1[7] ;
 wire \am_sdr0.cic1.integ1[8] ;
 wire \am_sdr0.cic1.integ1[9] ;
 wire \am_sdr0.cic1.integ2[0] ;
 wire \am_sdr0.cic1.integ2[10] ;
 wire \am_sdr0.cic1.integ2[11] ;
 wire \am_sdr0.cic1.integ2[12] ;
 wire \am_sdr0.cic1.integ2[13] ;
 wire \am_sdr0.cic1.integ2[14] ;
 wire \am_sdr0.cic1.integ2[15] ;
 wire \am_sdr0.cic1.integ2[16] ;
 wire \am_sdr0.cic1.integ2[17] ;
 wire \am_sdr0.cic1.integ2[18] ;
 wire \am_sdr0.cic1.integ2[19] ;
 wire \am_sdr0.cic1.integ2[1] ;
 wire \am_sdr0.cic1.integ2[20] ;
 wire \am_sdr0.cic1.integ2[21] ;
 wire \am_sdr0.cic1.integ2[22] ;
 wire \am_sdr0.cic1.integ2[2] ;
 wire \am_sdr0.cic1.integ2[3] ;
 wire \am_sdr0.cic1.integ2[4] ;
 wire \am_sdr0.cic1.integ2[5] ;
 wire \am_sdr0.cic1.integ2[6] ;
 wire \am_sdr0.cic1.integ2[7] ;
 wire \am_sdr0.cic1.integ2[8] ;
 wire \am_sdr0.cic1.integ2[9] ;
 wire \am_sdr0.cic1.integ3[0] ;
 wire \am_sdr0.cic1.integ3[10] ;
 wire \am_sdr0.cic1.integ3[11] ;
 wire \am_sdr0.cic1.integ3[12] ;
 wire \am_sdr0.cic1.integ3[13] ;
 wire \am_sdr0.cic1.integ3[14] ;
 wire \am_sdr0.cic1.integ3[15] ;
 wire \am_sdr0.cic1.integ3[16] ;
 wire \am_sdr0.cic1.integ3[17] ;
 wire \am_sdr0.cic1.integ3[18] ;
 wire \am_sdr0.cic1.integ3[19] ;
 wire \am_sdr0.cic1.integ3[1] ;
 wire \am_sdr0.cic1.integ3[2] ;
 wire \am_sdr0.cic1.integ3[3] ;
 wire \am_sdr0.cic1.integ3[4] ;
 wire \am_sdr0.cic1.integ3[5] ;
 wire \am_sdr0.cic1.integ3[6] ;
 wire \am_sdr0.cic1.integ3[7] ;
 wire \am_sdr0.cic1.integ3[8] ;
 wire \am_sdr0.cic1.integ3[9] ;
 wire \am_sdr0.cic1.integ_sample[0] ;
 wire \am_sdr0.cic1.integ_sample[10] ;
 wire \am_sdr0.cic1.integ_sample[11] ;
 wire \am_sdr0.cic1.integ_sample[12] ;
 wire \am_sdr0.cic1.integ_sample[13] ;
 wire \am_sdr0.cic1.integ_sample[14] ;
 wire \am_sdr0.cic1.integ_sample[15] ;
 wire \am_sdr0.cic1.integ_sample[16] ;
 wire \am_sdr0.cic1.integ_sample[17] ;
 wire \am_sdr0.cic1.integ_sample[18] ;
 wire \am_sdr0.cic1.integ_sample[19] ;
 wire \am_sdr0.cic1.integ_sample[1] ;
 wire \am_sdr0.cic1.integ_sample[2] ;
 wire \am_sdr0.cic1.integ_sample[3] ;
 wire \am_sdr0.cic1.integ_sample[4] ;
 wire \am_sdr0.cic1.integ_sample[5] ;
 wire \am_sdr0.cic1.integ_sample[6] ;
 wire \am_sdr0.cic1.integ_sample[7] ;
 wire \am_sdr0.cic1.integ_sample[8] ;
 wire \am_sdr0.cic1.integ_sample[9] ;
 wire \am_sdr0.cic1.out_tick ;
 wire \am_sdr0.cic1.sample ;
 wire \am_sdr0.cic1.x_out[10] ;
 wire \am_sdr0.cic1.x_out[11] ;
 wire \am_sdr0.cic1.x_out[12] ;
 wire \am_sdr0.cic1.x_out[13] ;
 wire \am_sdr0.cic1.x_out[14] ;
 wire \am_sdr0.cic1.x_out[15] ;
 wire \am_sdr0.cic1.x_out[8] ;
 wire \am_sdr0.cic1.x_out[9] ;
 wire \am_sdr0.cic2.comb1[0] ;
 wire \am_sdr0.cic2.comb1[10] ;
 wire \am_sdr0.cic2.comb1[11] ;
 wire \am_sdr0.cic2.comb1[12] ;
 wire \am_sdr0.cic2.comb1[13] ;
 wire \am_sdr0.cic2.comb1[14] ;
 wire \am_sdr0.cic2.comb1[15] ;
 wire \am_sdr0.cic2.comb1[16] ;
 wire \am_sdr0.cic2.comb1[17] ;
 wire \am_sdr0.cic2.comb1[18] ;
 wire \am_sdr0.cic2.comb1[19] ;
 wire \am_sdr0.cic2.comb1[1] ;
 wire \am_sdr0.cic2.comb1[2] ;
 wire \am_sdr0.cic2.comb1[3] ;
 wire \am_sdr0.cic2.comb1[4] ;
 wire \am_sdr0.cic2.comb1[5] ;
 wire \am_sdr0.cic2.comb1[6] ;
 wire \am_sdr0.cic2.comb1[7] ;
 wire \am_sdr0.cic2.comb1[8] ;
 wire \am_sdr0.cic2.comb1[9] ;
 wire \am_sdr0.cic2.comb1_in_del[0] ;
 wire \am_sdr0.cic2.comb1_in_del[10] ;
 wire \am_sdr0.cic2.comb1_in_del[11] ;
 wire \am_sdr0.cic2.comb1_in_del[12] ;
 wire \am_sdr0.cic2.comb1_in_del[13] ;
 wire \am_sdr0.cic2.comb1_in_del[14] ;
 wire \am_sdr0.cic2.comb1_in_del[15] ;
 wire \am_sdr0.cic2.comb1_in_del[16] ;
 wire \am_sdr0.cic2.comb1_in_del[17] ;
 wire \am_sdr0.cic2.comb1_in_del[18] ;
 wire \am_sdr0.cic2.comb1_in_del[19] ;
 wire \am_sdr0.cic2.comb1_in_del[1] ;
 wire \am_sdr0.cic2.comb1_in_del[2] ;
 wire \am_sdr0.cic2.comb1_in_del[3] ;
 wire \am_sdr0.cic2.comb1_in_del[4] ;
 wire \am_sdr0.cic2.comb1_in_del[5] ;
 wire \am_sdr0.cic2.comb1_in_del[6] ;
 wire \am_sdr0.cic2.comb1_in_del[7] ;
 wire \am_sdr0.cic2.comb1_in_del[8] ;
 wire \am_sdr0.cic2.comb1_in_del[9] ;
 wire \am_sdr0.cic2.comb2[0] ;
 wire \am_sdr0.cic2.comb2[10] ;
 wire \am_sdr0.cic2.comb2[11] ;
 wire \am_sdr0.cic2.comb2[12] ;
 wire \am_sdr0.cic2.comb2[13] ;
 wire \am_sdr0.cic2.comb2[14] ;
 wire \am_sdr0.cic2.comb2[15] ;
 wire \am_sdr0.cic2.comb2[16] ;
 wire \am_sdr0.cic2.comb2[17] ;
 wire \am_sdr0.cic2.comb2[18] ;
 wire \am_sdr0.cic2.comb2[19] ;
 wire \am_sdr0.cic2.comb2[1] ;
 wire \am_sdr0.cic2.comb2[2] ;
 wire \am_sdr0.cic2.comb2[3] ;
 wire \am_sdr0.cic2.comb2[4] ;
 wire \am_sdr0.cic2.comb2[5] ;
 wire \am_sdr0.cic2.comb2[6] ;
 wire \am_sdr0.cic2.comb2[7] ;
 wire \am_sdr0.cic2.comb2[8] ;
 wire \am_sdr0.cic2.comb2[9] ;
 wire \am_sdr0.cic2.comb2_in_del[0] ;
 wire \am_sdr0.cic2.comb2_in_del[10] ;
 wire \am_sdr0.cic2.comb2_in_del[11] ;
 wire \am_sdr0.cic2.comb2_in_del[12] ;
 wire \am_sdr0.cic2.comb2_in_del[13] ;
 wire \am_sdr0.cic2.comb2_in_del[14] ;
 wire \am_sdr0.cic2.comb2_in_del[15] ;
 wire \am_sdr0.cic2.comb2_in_del[16] ;
 wire \am_sdr0.cic2.comb2_in_del[17] ;
 wire \am_sdr0.cic2.comb2_in_del[18] ;
 wire \am_sdr0.cic2.comb2_in_del[19] ;
 wire \am_sdr0.cic2.comb2_in_del[1] ;
 wire \am_sdr0.cic2.comb2_in_del[2] ;
 wire \am_sdr0.cic2.comb2_in_del[3] ;
 wire \am_sdr0.cic2.comb2_in_del[4] ;
 wire \am_sdr0.cic2.comb2_in_del[5] ;
 wire \am_sdr0.cic2.comb2_in_del[6] ;
 wire \am_sdr0.cic2.comb2_in_del[7] ;
 wire \am_sdr0.cic2.comb2_in_del[8] ;
 wire \am_sdr0.cic2.comb2_in_del[9] ;
 wire \am_sdr0.cic2.comb3[12] ;
 wire \am_sdr0.cic2.comb3[13] ;
 wire \am_sdr0.cic2.comb3[14] ;
 wire \am_sdr0.cic2.comb3[15] ;
 wire \am_sdr0.cic2.comb3[16] ;
 wire \am_sdr0.cic2.comb3[17] ;
 wire \am_sdr0.cic2.comb3[18] ;
 wire \am_sdr0.cic2.comb3[19] ;
 wire \am_sdr0.cic2.comb3_in_del[0] ;
 wire \am_sdr0.cic2.comb3_in_del[10] ;
 wire \am_sdr0.cic2.comb3_in_del[11] ;
 wire \am_sdr0.cic2.comb3_in_del[12] ;
 wire \am_sdr0.cic2.comb3_in_del[13] ;
 wire \am_sdr0.cic2.comb3_in_del[14] ;
 wire \am_sdr0.cic2.comb3_in_del[15] ;
 wire \am_sdr0.cic2.comb3_in_del[16] ;
 wire \am_sdr0.cic2.comb3_in_del[17] ;
 wire \am_sdr0.cic2.comb3_in_del[18] ;
 wire \am_sdr0.cic2.comb3_in_del[19] ;
 wire \am_sdr0.cic2.comb3_in_del[1] ;
 wire \am_sdr0.cic2.comb3_in_del[2] ;
 wire \am_sdr0.cic2.comb3_in_del[3] ;
 wire \am_sdr0.cic2.comb3_in_del[4] ;
 wire \am_sdr0.cic2.comb3_in_del[5] ;
 wire \am_sdr0.cic2.comb3_in_del[6] ;
 wire \am_sdr0.cic2.comb3_in_del[7] ;
 wire \am_sdr0.cic2.comb3_in_del[8] ;
 wire \am_sdr0.cic2.comb3_in_del[9] ;
 wire \am_sdr0.cic2.count[0] ;
 wire \am_sdr0.cic2.count[1] ;
 wire \am_sdr0.cic2.count[2] ;
 wire \am_sdr0.cic2.count[3] ;
 wire \am_sdr0.cic2.count[4] ;
 wire \am_sdr0.cic2.count[5] ;
 wire \am_sdr0.cic2.count[6] ;
 wire \am_sdr0.cic2.count[7] ;
 wire \am_sdr0.cic2.integ1[0] ;
 wire \am_sdr0.cic2.integ1[10] ;
 wire \am_sdr0.cic2.integ1[11] ;
 wire \am_sdr0.cic2.integ1[12] ;
 wire \am_sdr0.cic2.integ1[13] ;
 wire \am_sdr0.cic2.integ1[14] ;
 wire \am_sdr0.cic2.integ1[15] ;
 wire \am_sdr0.cic2.integ1[16] ;
 wire \am_sdr0.cic2.integ1[17] ;
 wire \am_sdr0.cic2.integ1[18] ;
 wire \am_sdr0.cic2.integ1[19] ;
 wire \am_sdr0.cic2.integ1[1] ;
 wire \am_sdr0.cic2.integ1[20] ;
 wire \am_sdr0.cic2.integ1[21] ;
 wire \am_sdr0.cic2.integ1[22] ;
 wire \am_sdr0.cic2.integ1[23] ;
 wire \am_sdr0.cic2.integ1[24] ;
 wire \am_sdr0.cic2.integ1[25] ;
 wire \am_sdr0.cic2.integ1[2] ;
 wire \am_sdr0.cic2.integ1[3] ;
 wire \am_sdr0.cic2.integ1[4] ;
 wire \am_sdr0.cic2.integ1[5] ;
 wire \am_sdr0.cic2.integ1[6] ;
 wire \am_sdr0.cic2.integ1[7] ;
 wire \am_sdr0.cic2.integ1[8] ;
 wire \am_sdr0.cic2.integ1[9] ;
 wire \am_sdr0.cic2.integ2[0] ;
 wire \am_sdr0.cic2.integ2[10] ;
 wire \am_sdr0.cic2.integ2[11] ;
 wire \am_sdr0.cic2.integ2[12] ;
 wire \am_sdr0.cic2.integ2[13] ;
 wire \am_sdr0.cic2.integ2[14] ;
 wire \am_sdr0.cic2.integ2[15] ;
 wire \am_sdr0.cic2.integ2[16] ;
 wire \am_sdr0.cic2.integ2[17] ;
 wire \am_sdr0.cic2.integ2[18] ;
 wire \am_sdr0.cic2.integ2[19] ;
 wire \am_sdr0.cic2.integ2[1] ;
 wire \am_sdr0.cic2.integ2[20] ;
 wire \am_sdr0.cic2.integ2[21] ;
 wire \am_sdr0.cic2.integ2[22] ;
 wire \am_sdr0.cic2.integ2[2] ;
 wire \am_sdr0.cic2.integ2[3] ;
 wire \am_sdr0.cic2.integ2[4] ;
 wire \am_sdr0.cic2.integ2[5] ;
 wire \am_sdr0.cic2.integ2[6] ;
 wire \am_sdr0.cic2.integ2[7] ;
 wire \am_sdr0.cic2.integ2[8] ;
 wire \am_sdr0.cic2.integ2[9] ;
 wire \am_sdr0.cic2.integ3[0] ;
 wire \am_sdr0.cic2.integ3[10] ;
 wire \am_sdr0.cic2.integ3[11] ;
 wire \am_sdr0.cic2.integ3[12] ;
 wire \am_sdr0.cic2.integ3[13] ;
 wire \am_sdr0.cic2.integ3[14] ;
 wire \am_sdr0.cic2.integ3[15] ;
 wire \am_sdr0.cic2.integ3[16] ;
 wire \am_sdr0.cic2.integ3[17] ;
 wire \am_sdr0.cic2.integ3[18] ;
 wire \am_sdr0.cic2.integ3[19] ;
 wire \am_sdr0.cic2.integ3[1] ;
 wire \am_sdr0.cic2.integ3[2] ;
 wire \am_sdr0.cic2.integ3[3] ;
 wire \am_sdr0.cic2.integ3[4] ;
 wire \am_sdr0.cic2.integ3[5] ;
 wire \am_sdr0.cic2.integ3[6] ;
 wire \am_sdr0.cic2.integ3[7] ;
 wire \am_sdr0.cic2.integ3[8] ;
 wire \am_sdr0.cic2.integ3[9] ;
 wire \am_sdr0.cic2.integ_sample[0] ;
 wire \am_sdr0.cic2.integ_sample[10] ;
 wire \am_sdr0.cic2.integ_sample[11] ;
 wire \am_sdr0.cic2.integ_sample[12] ;
 wire \am_sdr0.cic2.integ_sample[13] ;
 wire \am_sdr0.cic2.integ_sample[14] ;
 wire \am_sdr0.cic2.integ_sample[15] ;
 wire \am_sdr0.cic2.integ_sample[16] ;
 wire \am_sdr0.cic2.integ_sample[17] ;
 wire \am_sdr0.cic2.integ_sample[18] ;
 wire \am_sdr0.cic2.integ_sample[19] ;
 wire \am_sdr0.cic2.integ_sample[1] ;
 wire \am_sdr0.cic2.integ_sample[2] ;
 wire \am_sdr0.cic2.integ_sample[3] ;
 wire \am_sdr0.cic2.integ_sample[4] ;
 wire \am_sdr0.cic2.integ_sample[5] ;
 wire \am_sdr0.cic2.integ_sample[6] ;
 wire \am_sdr0.cic2.integ_sample[7] ;
 wire \am_sdr0.cic2.integ_sample[8] ;
 wire \am_sdr0.cic2.integ_sample[9] ;
 wire \am_sdr0.cic2.sample ;
 wire \am_sdr0.cic3.comb1[0] ;
 wire \am_sdr0.cic3.comb1[10] ;
 wire \am_sdr0.cic3.comb1[11] ;
 wire \am_sdr0.cic3.comb1[12] ;
 wire \am_sdr0.cic3.comb1[13] ;
 wire \am_sdr0.cic3.comb1[14] ;
 wire \am_sdr0.cic3.comb1[15] ;
 wire \am_sdr0.cic3.comb1[16] ;
 wire \am_sdr0.cic3.comb1[17] ;
 wire \am_sdr0.cic3.comb1[18] ;
 wire \am_sdr0.cic3.comb1[19] ;
 wire \am_sdr0.cic3.comb1[1] ;
 wire \am_sdr0.cic3.comb1[2] ;
 wire \am_sdr0.cic3.comb1[3] ;
 wire \am_sdr0.cic3.comb1[4] ;
 wire \am_sdr0.cic3.comb1[5] ;
 wire \am_sdr0.cic3.comb1[6] ;
 wire \am_sdr0.cic3.comb1[7] ;
 wire \am_sdr0.cic3.comb1[8] ;
 wire \am_sdr0.cic3.comb1[9] ;
 wire \am_sdr0.cic3.comb1_in_del[0] ;
 wire \am_sdr0.cic3.comb1_in_del[10] ;
 wire \am_sdr0.cic3.comb1_in_del[11] ;
 wire \am_sdr0.cic3.comb1_in_del[12] ;
 wire \am_sdr0.cic3.comb1_in_del[13] ;
 wire \am_sdr0.cic3.comb1_in_del[14] ;
 wire \am_sdr0.cic3.comb1_in_del[15] ;
 wire \am_sdr0.cic3.comb1_in_del[16] ;
 wire \am_sdr0.cic3.comb1_in_del[17] ;
 wire \am_sdr0.cic3.comb1_in_del[18] ;
 wire \am_sdr0.cic3.comb1_in_del[19] ;
 wire \am_sdr0.cic3.comb1_in_del[1] ;
 wire \am_sdr0.cic3.comb1_in_del[2] ;
 wire \am_sdr0.cic3.comb1_in_del[3] ;
 wire \am_sdr0.cic3.comb1_in_del[4] ;
 wire \am_sdr0.cic3.comb1_in_del[5] ;
 wire \am_sdr0.cic3.comb1_in_del[6] ;
 wire \am_sdr0.cic3.comb1_in_del[7] ;
 wire \am_sdr0.cic3.comb1_in_del[8] ;
 wire \am_sdr0.cic3.comb1_in_del[9] ;
 wire \am_sdr0.cic3.comb2[0] ;
 wire \am_sdr0.cic3.comb2[10] ;
 wire \am_sdr0.cic3.comb2[11] ;
 wire \am_sdr0.cic3.comb2[12] ;
 wire \am_sdr0.cic3.comb2[13] ;
 wire \am_sdr0.cic3.comb2[14] ;
 wire \am_sdr0.cic3.comb2[15] ;
 wire \am_sdr0.cic3.comb2[16] ;
 wire \am_sdr0.cic3.comb2[17] ;
 wire \am_sdr0.cic3.comb2[18] ;
 wire \am_sdr0.cic3.comb2[19] ;
 wire \am_sdr0.cic3.comb2[1] ;
 wire \am_sdr0.cic3.comb2[2] ;
 wire \am_sdr0.cic3.comb2[3] ;
 wire \am_sdr0.cic3.comb2[4] ;
 wire \am_sdr0.cic3.comb2[5] ;
 wire \am_sdr0.cic3.comb2[6] ;
 wire \am_sdr0.cic3.comb2[7] ;
 wire \am_sdr0.cic3.comb2[8] ;
 wire \am_sdr0.cic3.comb2[9] ;
 wire \am_sdr0.cic3.comb2_in_del[0] ;
 wire \am_sdr0.cic3.comb2_in_del[10] ;
 wire \am_sdr0.cic3.comb2_in_del[11] ;
 wire \am_sdr0.cic3.comb2_in_del[12] ;
 wire \am_sdr0.cic3.comb2_in_del[13] ;
 wire \am_sdr0.cic3.comb2_in_del[14] ;
 wire \am_sdr0.cic3.comb2_in_del[15] ;
 wire \am_sdr0.cic3.comb2_in_del[16] ;
 wire \am_sdr0.cic3.comb2_in_del[17] ;
 wire \am_sdr0.cic3.comb2_in_del[18] ;
 wire \am_sdr0.cic3.comb2_in_del[19] ;
 wire \am_sdr0.cic3.comb2_in_del[1] ;
 wire \am_sdr0.cic3.comb2_in_del[2] ;
 wire \am_sdr0.cic3.comb2_in_del[3] ;
 wire \am_sdr0.cic3.comb2_in_del[4] ;
 wire \am_sdr0.cic3.comb2_in_del[5] ;
 wire \am_sdr0.cic3.comb2_in_del[6] ;
 wire \am_sdr0.cic3.comb2_in_del[7] ;
 wire \am_sdr0.cic3.comb2_in_del[8] ;
 wire \am_sdr0.cic3.comb2_in_del[9] ;
 wire \am_sdr0.cic3.comb3[12] ;
 wire \am_sdr0.cic3.comb3[13] ;
 wire \am_sdr0.cic3.comb3[14] ;
 wire \am_sdr0.cic3.comb3[15] ;
 wire \am_sdr0.cic3.comb3[16] ;
 wire \am_sdr0.cic3.comb3[17] ;
 wire \am_sdr0.cic3.comb3[18] ;
 wire \am_sdr0.cic3.comb3[19] ;
 wire \am_sdr0.cic3.comb3_in_del[0] ;
 wire \am_sdr0.cic3.comb3_in_del[10] ;
 wire \am_sdr0.cic3.comb3_in_del[11] ;
 wire \am_sdr0.cic3.comb3_in_del[12] ;
 wire \am_sdr0.cic3.comb3_in_del[13] ;
 wire \am_sdr0.cic3.comb3_in_del[14] ;
 wire \am_sdr0.cic3.comb3_in_del[15] ;
 wire \am_sdr0.cic3.comb3_in_del[16] ;
 wire \am_sdr0.cic3.comb3_in_del[17] ;
 wire \am_sdr0.cic3.comb3_in_del[18] ;
 wire \am_sdr0.cic3.comb3_in_del[19] ;
 wire \am_sdr0.cic3.comb3_in_del[1] ;
 wire \am_sdr0.cic3.comb3_in_del[2] ;
 wire \am_sdr0.cic3.comb3_in_del[3] ;
 wire \am_sdr0.cic3.comb3_in_del[4] ;
 wire \am_sdr0.cic3.comb3_in_del[5] ;
 wire \am_sdr0.cic3.comb3_in_del[6] ;
 wire \am_sdr0.cic3.comb3_in_del[7] ;
 wire \am_sdr0.cic3.comb3_in_del[8] ;
 wire \am_sdr0.cic3.comb3_in_del[9] ;
 wire \am_sdr0.cic3.count[0] ;
 wire \am_sdr0.cic3.count[1] ;
 wire \am_sdr0.cic3.count[2] ;
 wire \am_sdr0.cic3.count[3] ;
 wire \am_sdr0.cic3.count[4] ;
 wire \am_sdr0.cic3.count[5] ;
 wire \am_sdr0.cic3.count[6] ;
 wire \am_sdr0.cic3.count[7] ;
 wire \am_sdr0.cic3.integ1[0] ;
 wire \am_sdr0.cic3.integ1[10] ;
 wire \am_sdr0.cic3.integ1[11] ;
 wire \am_sdr0.cic3.integ1[12] ;
 wire \am_sdr0.cic3.integ1[13] ;
 wire \am_sdr0.cic3.integ1[14] ;
 wire \am_sdr0.cic3.integ1[15] ;
 wire \am_sdr0.cic3.integ1[16] ;
 wire \am_sdr0.cic3.integ1[17] ;
 wire \am_sdr0.cic3.integ1[18] ;
 wire \am_sdr0.cic3.integ1[19] ;
 wire \am_sdr0.cic3.integ1[1] ;
 wire \am_sdr0.cic3.integ1[20] ;
 wire \am_sdr0.cic3.integ1[21] ;
 wire \am_sdr0.cic3.integ1[22] ;
 wire \am_sdr0.cic3.integ1[23] ;
 wire \am_sdr0.cic3.integ1[24] ;
 wire \am_sdr0.cic3.integ1[25] ;
 wire \am_sdr0.cic3.integ1[2] ;
 wire \am_sdr0.cic3.integ1[3] ;
 wire \am_sdr0.cic3.integ1[4] ;
 wire \am_sdr0.cic3.integ1[5] ;
 wire \am_sdr0.cic3.integ1[6] ;
 wire \am_sdr0.cic3.integ1[7] ;
 wire \am_sdr0.cic3.integ1[8] ;
 wire \am_sdr0.cic3.integ1[9] ;
 wire \am_sdr0.cic3.integ2[0] ;
 wire \am_sdr0.cic3.integ2[10] ;
 wire \am_sdr0.cic3.integ2[11] ;
 wire \am_sdr0.cic3.integ2[12] ;
 wire \am_sdr0.cic3.integ2[13] ;
 wire \am_sdr0.cic3.integ2[14] ;
 wire \am_sdr0.cic3.integ2[15] ;
 wire \am_sdr0.cic3.integ2[16] ;
 wire \am_sdr0.cic3.integ2[17] ;
 wire \am_sdr0.cic3.integ2[18] ;
 wire \am_sdr0.cic3.integ2[19] ;
 wire \am_sdr0.cic3.integ2[1] ;
 wire \am_sdr0.cic3.integ2[20] ;
 wire \am_sdr0.cic3.integ2[21] ;
 wire \am_sdr0.cic3.integ2[22] ;
 wire \am_sdr0.cic3.integ2[2] ;
 wire \am_sdr0.cic3.integ2[3] ;
 wire \am_sdr0.cic3.integ2[4] ;
 wire \am_sdr0.cic3.integ2[5] ;
 wire \am_sdr0.cic3.integ2[6] ;
 wire \am_sdr0.cic3.integ2[7] ;
 wire \am_sdr0.cic3.integ2[8] ;
 wire \am_sdr0.cic3.integ2[9] ;
 wire \am_sdr0.cic3.integ3[0] ;
 wire \am_sdr0.cic3.integ3[10] ;
 wire \am_sdr0.cic3.integ3[11] ;
 wire \am_sdr0.cic3.integ3[12] ;
 wire \am_sdr0.cic3.integ3[13] ;
 wire \am_sdr0.cic3.integ3[14] ;
 wire \am_sdr0.cic3.integ3[15] ;
 wire \am_sdr0.cic3.integ3[16] ;
 wire \am_sdr0.cic3.integ3[17] ;
 wire \am_sdr0.cic3.integ3[18] ;
 wire \am_sdr0.cic3.integ3[19] ;
 wire \am_sdr0.cic3.integ3[1] ;
 wire \am_sdr0.cic3.integ3[2] ;
 wire \am_sdr0.cic3.integ3[3] ;
 wire \am_sdr0.cic3.integ3[4] ;
 wire \am_sdr0.cic3.integ3[5] ;
 wire \am_sdr0.cic3.integ3[6] ;
 wire \am_sdr0.cic3.integ3[7] ;
 wire \am_sdr0.cic3.integ3[8] ;
 wire \am_sdr0.cic3.integ3[9] ;
 wire \am_sdr0.cic3.integ_sample[0] ;
 wire \am_sdr0.cic3.integ_sample[10] ;
 wire \am_sdr0.cic3.integ_sample[11] ;
 wire \am_sdr0.cic3.integ_sample[12] ;
 wire \am_sdr0.cic3.integ_sample[13] ;
 wire \am_sdr0.cic3.integ_sample[14] ;
 wire \am_sdr0.cic3.integ_sample[15] ;
 wire \am_sdr0.cic3.integ_sample[16] ;
 wire \am_sdr0.cic3.integ_sample[17] ;
 wire \am_sdr0.cic3.integ_sample[18] ;
 wire \am_sdr0.cic3.integ_sample[19] ;
 wire \am_sdr0.cic3.integ_sample[1] ;
 wire \am_sdr0.cic3.integ_sample[2] ;
 wire \am_sdr0.cic3.integ_sample[3] ;
 wire \am_sdr0.cic3.integ_sample[4] ;
 wire \am_sdr0.cic3.integ_sample[5] ;
 wire \am_sdr0.cic3.integ_sample[6] ;
 wire \am_sdr0.cic3.integ_sample[7] ;
 wire \am_sdr0.cic3.integ_sample[8] ;
 wire \am_sdr0.cic3.integ_sample[9] ;
 wire \am_sdr0.cic3.sample ;
 wire \am_sdr0.cos[0] ;
 wire \am_sdr0.cos[1] ;
 wire \am_sdr0.cos[2] ;
 wire \am_sdr0.cos[3] ;
 wire \am_sdr0.cos[4] ;
 wire \am_sdr0.cos[5] ;
 wire \am_sdr0.cos[6] ;
 wire \am_sdr0.cos[7] ;
 wire \am_sdr0.count[0] ;
 wire \am_sdr0.count[1] ;
 wire \am_sdr0.count[2] ;
 wire \am_sdr0.count[3] ;
 wire \am_sdr0.count[4] ;
 wire \am_sdr0.count[5] ;
 wire \am_sdr0.count[6] ;
 wire \am_sdr0.count[7] ;
 wire \am_sdr0.gain_spi[0] ;
 wire \am_sdr0.gain_spi[1] ;
 wire \am_sdr0.gain_spi[2] ;
 wire \am_sdr0.mix0.RF_in_q ;
 wire \am_sdr0.mix0.RF_in_qq ;
 wire \am_sdr0.mix0.cos_q[0] ;
 wire \am_sdr0.mix0.cos_q[1] ;
 wire \am_sdr0.mix0.cos_q[2] ;
 wire \am_sdr0.mix0.cos_q[3] ;
 wire \am_sdr0.mix0.cos_q[4] ;
 wire \am_sdr0.mix0.cos_q[5] ;
 wire \am_sdr0.mix0.cos_q[6] ;
 wire \am_sdr0.mix0.cos_q[7] ;
 wire \am_sdr0.mix0.sin_in[0] ;
 wire \am_sdr0.mix0.sin_in[1] ;
 wire \am_sdr0.mix0.sin_in[2] ;
 wire \am_sdr0.mix0.sin_in[3] ;
 wire \am_sdr0.mix0.sin_in[4] ;
 wire \am_sdr0.mix0.sin_in[5] ;
 wire \am_sdr0.mix0.sin_in[6] ;
 wire \am_sdr0.mix0.sin_in[7] ;
 wire \am_sdr0.mix0.sin_q[0] ;
 wire \am_sdr0.mix0.sin_q[1] ;
 wire \am_sdr0.mix0.sin_q[2] ;
 wire \am_sdr0.mix0.sin_q[3] ;
 wire \am_sdr0.mix0.sin_q[4] ;
 wire \am_sdr0.mix0.sin_q[5] ;
 wire \am_sdr0.mix0.sin_q[6] ;
 wire \am_sdr0.mix0.sin_q[7] ;
 wire \am_sdr0.nco0.phase[0] ;
 wire \am_sdr0.nco0.phase[10] ;
 wire \am_sdr0.nco0.phase[11] ;
 wire \am_sdr0.nco0.phase[12] ;
 wire \am_sdr0.nco0.phase[13] ;
 wire \am_sdr0.nco0.phase[14] ;
 wire \am_sdr0.nco0.phase[15] ;
 wire \am_sdr0.nco0.phase[16] ;
 wire \am_sdr0.nco0.phase[17] ;
 wire \am_sdr0.nco0.phase[18] ;
 wire \am_sdr0.nco0.phase[19] ;
 wire \am_sdr0.nco0.phase[1] ;
 wire \am_sdr0.nco0.phase[20] ;
 wire \am_sdr0.nco0.phase[21] ;
 wire \am_sdr0.nco0.phase[22] ;
 wire \am_sdr0.nco0.phase[23] ;
 wire \am_sdr0.nco0.phase[24] ;
 wire \am_sdr0.nco0.phase[25] ;
 wire \am_sdr0.nco0.phase[2] ;
 wire \am_sdr0.nco0.phase[3] ;
 wire \am_sdr0.nco0.phase[4] ;
 wire \am_sdr0.nco0.phase[5] ;
 wire \am_sdr0.nco0.phase[6] ;
 wire \am_sdr0.nco0.phase[7] ;
 wire \am_sdr0.nco0.phase[8] ;
 wire \am_sdr0.nco0.phase[9] ;
 wire \am_sdr0.nco0.phase_inc[0] ;
 wire \am_sdr0.nco0.phase_inc[10] ;
 wire \am_sdr0.nco0.phase_inc[11] ;
 wire \am_sdr0.nco0.phase_inc[12] ;
 wire \am_sdr0.nco0.phase_inc[13] ;
 wire \am_sdr0.nco0.phase_inc[14] ;
 wire \am_sdr0.nco0.phase_inc[15] ;
 wire \am_sdr0.nco0.phase_inc[16] ;
 wire \am_sdr0.nco0.phase_inc[17] ;
 wire \am_sdr0.nco0.phase_inc[18] ;
 wire \am_sdr0.nco0.phase_inc[19] ;
 wire \am_sdr0.nco0.phase_inc[1] ;
 wire \am_sdr0.nco0.phase_inc[20] ;
 wire \am_sdr0.nco0.phase_inc[21] ;
 wire \am_sdr0.nco0.phase_inc[22] ;
 wire \am_sdr0.nco0.phase_inc[23] ;
 wire \am_sdr0.nco0.phase_inc[24] ;
 wire \am_sdr0.nco0.phase_inc[25] ;
 wire \am_sdr0.nco0.phase_inc[2] ;
 wire \am_sdr0.nco0.phase_inc[3] ;
 wire \am_sdr0.nco0.phase_inc[4] ;
 wire \am_sdr0.nco0.phase_inc[5] ;
 wire \am_sdr0.nco0.phase_inc[6] ;
 wire \am_sdr0.nco0.phase_inc[7] ;
 wire \am_sdr0.nco0.phase_inc[8] ;
 wire \am_sdr0.nco0.phase_inc[9] ;
 wire \am_sdr0.spi0.CS_q ;
 wire \am_sdr0.spi0.CS_qq ;
 wire \am_sdr0.spi0.CS_qqq ;
 wire \am_sdr0.spi0.MOSI_q ;
 wire \am_sdr0.spi0.MOSI_qq ;
 wire \am_sdr0.spi0.SCK_q ;
 wire \am_sdr0.spi0.SCK_qq ;
 wire \am_sdr0.spi0.SCK_qqq ;
 wire \am_sdr0.spi0.shift_reg[0] ;
 wire \am_sdr0.spi0.shift_reg[10] ;
 wire \am_sdr0.spi0.shift_reg[11] ;
 wire \am_sdr0.spi0.shift_reg[12] ;
 wire \am_sdr0.spi0.shift_reg[13] ;
 wire \am_sdr0.spi0.shift_reg[14] ;
 wire \am_sdr0.spi0.shift_reg[15] ;
 wire \am_sdr0.spi0.shift_reg[16] ;
 wire \am_sdr0.spi0.shift_reg[17] ;
 wire \am_sdr0.spi0.shift_reg[18] ;
 wire \am_sdr0.spi0.shift_reg[19] ;
 wire \am_sdr0.spi0.shift_reg[1] ;
 wire \am_sdr0.spi0.shift_reg[20] ;
 wire \am_sdr0.spi0.shift_reg[21] ;
 wire \am_sdr0.spi0.shift_reg[22] ;
 wire \am_sdr0.spi0.shift_reg[23] ;
 wire \am_sdr0.spi0.shift_reg[24] ;
 wire \am_sdr0.spi0.shift_reg[25] ;
 wire \am_sdr0.spi0.shift_reg[26] ;
 wire \am_sdr0.spi0.shift_reg[27] ;
 wire \am_sdr0.spi0.shift_reg[28] ;
 wire \am_sdr0.spi0.shift_reg[2] ;
 wire \am_sdr0.spi0.shift_reg[3] ;
 wire \am_sdr0.spi0.shift_reg[4] ;
 wire \am_sdr0.spi0.shift_reg[5] ;
 wire \am_sdr0.spi0.shift_reg[6] ;
 wire \am_sdr0.spi0.shift_reg[7] ;
 wire \am_sdr0.spi0.shift_reg[8] ;
 wire \am_sdr0.spi0.shift_reg[9] ;
 wire \am_sdr0.spi0.state[0] ;
 wire \am_sdr0.spi0.state[1] ;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_145_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;

 sg13g2_inv_1 _07971_ (.Y(_01177_),
    .A(net1323));
 sg13g2_inv_1 _07972_ (.Y(_01178_),
    .A(net2047));
 sg13g2_inv_1 _07973_ (.Y(_01179_),
    .A(net1435));
 sg13g2_inv_1 _07974_ (.Y(_01180_),
    .A(\am_sdr0.am0.demod_out[13] ));
 sg13g2_inv_1 _07975_ (.Y(_01181_),
    .A(net1488));
 sg13g2_inv_1 _07976_ (.Y(_01182_),
    .A(\am_sdr0.am0.demod_out[12] ));
 sg13g2_inv_1 _07977_ (.Y(_01183_),
    .A(net2168));
 sg13g2_inv_1 _07978_ (.Y(_01184_),
    .A(\am_sdr0.am0.demod_out[11] ));
 sg13g2_inv_1 _07979_ (.Y(_01185_),
    .A(net1522));
 sg13g2_inv_2 _07980_ (.Y(_01186_),
    .A(\am_sdr0.am0.demod_out[10] ));
 sg13g2_inv_1 _07981_ (.Y(_01187_),
    .A(net2127));
 sg13g2_inv_1 _07982_ (.Y(_01188_),
    .A(net1647));
 sg13g2_inv_1 _07983_ (.Y(_01189_),
    .A(net2139));
 sg13g2_inv_1 _07984_ (.Y(_01190_),
    .A(\am_sdr0.am0.q[0] ));
 sg13g2_inv_1 _07985_ (.Y(_01191_),
    .A(net1235));
 sg13g2_inv_1 _07986_ (.Y(_01192_),
    .A(net2640));
 sg13g2_inv_1 _07987_ (.Y(_01193_),
    .A(net2415));
 sg13g2_inv_1 _07988_ (.Y(_01194_),
    .A(net1341));
 sg13g2_inv_1 _07989_ (.Y(_01195_),
    .A(net2161));
 sg13g2_inv_1 _07990_ (.Y(_01196_),
    .A(net1343));
 sg13g2_inv_1 _07991_ (.Y(_01197_),
    .A(net1415));
 sg13g2_inv_1 _07992_ (.Y(_01198_),
    .A(\am_sdr0.nco0.phase_inc[23] ));
 sg13g2_inv_1 _07993_ (.Y(_01199_),
    .A(net1455));
 sg13g2_inv_1 _07994_ (.Y(_01200_),
    .A(net1419));
 sg13g2_inv_1 _07995_ (.Y(_01201_),
    .A(net2557));
 sg13g2_inv_1 _07996_ (.Y(_01202_),
    .A(net1289));
 sg13g2_inv_1 _07997_ (.Y(_01203_),
    .A(net2043));
 sg13g2_inv_1 _07998_ (.Y(_01204_),
    .A(net2093));
 sg13g2_inv_1 _07999_ (.Y(_01205_),
    .A(net2498));
 sg13g2_inv_1 _08000_ (.Y(_01206_),
    .A(net1420));
 sg13g2_inv_1 _08001_ (.Y(_01207_),
    .A(net1345));
 sg13g2_inv_1 _08002_ (.Y(_01208_),
    .A(net1298));
 sg13g2_inv_1 _08003_ (.Y(_01209_),
    .A(net2439));
 sg13g2_inv_1 _08004_ (.Y(_01210_),
    .A(net1409));
 sg13g2_inv_1 _08005_ (.Y(_01211_),
    .A(net1315));
 sg13g2_inv_1 _08006_ (.Y(_01212_),
    .A(net2076));
 sg13g2_inv_1 _08007_ (.Y(_01213_),
    .A(net1422));
 sg13g2_inv_1 _08008_ (.Y(_01214_),
    .A(net2091));
 sg13g2_inv_1 _08009_ (.Y(_01215_),
    .A(net2244));
 sg13g2_inv_1 _08010_ (.Y(_01216_),
    .A(net2193));
 sg13g2_inv_1 _08011_ (.Y(_01217_),
    .A(net1291));
 sg13g2_inv_1 _08012_ (.Y(_01218_),
    .A(net2745));
 sg13g2_inv_1 _08013_ (.Y(_01219_),
    .A(net1271));
 sg13g2_inv_1 _08014_ (.Y(_01220_),
    .A(net2554));
 sg13g2_inv_1 _08015_ (.Y(_01221_),
    .A(net2054));
 sg13g2_inv_1 _08016_ (.Y(_01222_),
    .A(net2133));
 sg13g2_inv_1 _08017_ (.Y(_01223_),
    .A(net1721));
 sg13g2_inv_1 _08018_ (.Y(_01224_),
    .A(net2201));
 sg13g2_inv_1 _08019_ (.Y(_01225_),
    .A(net2550));
 sg13g2_inv_1 _08020_ (.Y(_01226_),
    .A(net2560));
 sg13g2_inv_1 _08021_ (.Y(_01227_),
    .A(net2633));
 sg13g2_inv_1 _08022_ (.Y(_01228_),
    .A(net2265));
 sg13g2_inv_1 _08023_ (.Y(_01229_),
    .A(net2092));
 sg13g2_inv_1 _08024_ (.Y(_01230_),
    .A(net2289));
 sg13g2_inv_1 _08025_ (.Y(_01231_),
    .A(\am_sdr0.cic0.comb3_in_del[11] ));
 sg13g2_inv_1 _08026_ (.Y(_01232_),
    .A(\am_sdr0.cic0.comb2[11] ));
 sg13g2_inv_1 _08027_ (.Y(_01233_),
    .A(net2212));
 sg13g2_inv_1 _08028_ (.Y(_01234_),
    .A(net2224));
 sg13g2_inv_1 _08029_ (.Y(_01235_),
    .A(\am_sdr0.cic0.comb3_in_del[8] ));
 sg13g2_inv_1 _08030_ (.Y(_01236_),
    .A(net2319));
 sg13g2_inv_1 _08031_ (.Y(_01237_),
    .A(\am_sdr0.cic0.comb3_in_del[7] ));
 sg13g2_inv_1 _08032_ (.Y(_01238_),
    .A(\am_sdr0.cic0.comb2[7] ));
 sg13g2_inv_1 _08033_ (.Y(_01239_),
    .A(\am_sdr0.cic0.comb3_in_del[6] ));
 sg13g2_inv_1 _08034_ (.Y(_01240_),
    .A(\am_sdr0.cic0.comb2[6] ));
 sg13g2_inv_1 _08035_ (.Y(_01241_),
    .A(\am_sdr0.cic0.comb3_in_del[5] ));
 sg13g2_inv_1 _08036_ (.Y(_01242_),
    .A(net2711));
 sg13g2_inv_1 _08037_ (.Y(_01243_),
    .A(\am_sdr0.cic0.comb3_in_del[4] ));
 sg13g2_inv_1 _08038_ (.Y(_01244_),
    .A(net2399));
 sg13g2_inv_1 _08039_ (.Y(_01245_),
    .A(net2079));
 sg13g2_inv_1 _08040_ (.Y(_01246_),
    .A(net2131));
 sg13g2_inv_1 _08041_ (.Y(_01247_),
    .A(net2074));
 sg13g2_inv_1 _08042_ (.Y(_01248_),
    .A(net2170));
 sg13g2_inv_1 _08043_ (.Y(_01249_),
    .A(net1368));
 sg13g2_inv_1 _08044_ (.Y(_01250_),
    .A(net1293));
 sg13g2_inv_1 _08045_ (.Y(_01251_),
    .A(net1306));
 sg13g2_inv_1 _08046_ (.Y(_01252_),
    .A(net1269));
 sg13g2_inv_1 _08047_ (.Y(_01253_),
    .A(net1495));
 sg13g2_inv_1 _08048_ (.Y(_01254_),
    .A(net1478));
 sg13g2_inv_1 _08049_ (.Y(_01255_),
    .A(net1339));
 sg13g2_inv_1 _08050_ (.Y(_01256_),
    .A(net1503));
 sg13g2_inv_1 _08051_ (.Y(_01257_),
    .A(net2123));
 sg13g2_inv_1 _08052_ (.Y(_01258_),
    .A(net2589));
 sg13g2_inv_1 _08053_ (.Y(_01259_),
    .A(\am_sdr0.cic0.comb2_in_del[17] ));
 sg13g2_inv_1 _08054_ (.Y(_01260_),
    .A(net2748));
 sg13g2_inv_1 _08055_ (.Y(_01261_),
    .A(net2272));
 sg13g2_inv_1 _08056_ (.Y(_01262_),
    .A(\am_sdr0.cic0.comb2_in_del[15] ));
 sg13g2_inv_1 _08057_ (.Y(_01263_),
    .A(net2743));
 sg13g2_inv_1 _08058_ (.Y(_01264_),
    .A(net2472));
 sg13g2_inv_1 _08059_ (.Y(_01265_),
    .A(net2694));
 sg13g2_inv_1 _08060_ (.Y(_01266_),
    .A(net2577));
 sg13g2_inv_1 _08061_ (.Y(_01267_),
    .A(\am_sdr0.cic0.comb1[11] ));
 sg13g2_inv_1 _08062_ (.Y(_01268_),
    .A(net2401));
 sg13g2_inv_1 _08063_ (.Y(_01269_),
    .A(\am_sdr0.cic0.comb2_in_del[9] ));
 sg13g2_inv_1 _08064_ (.Y(_01270_),
    .A(net2894));
 sg13g2_inv_1 _08065_ (.Y(_01271_),
    .A(net2440));
 sg13g2_inv_1 _08066_ (.Y(_01272_),
    .A(net2107));
 sg13g2_inv_1 _08067_ (.Y(_01273_),
    .A(net2331));
 sg13g2_inv_1 _08068_ (.Y(_01274_),
    .A(net2431));
 sg13g2_inv_1 _08069_ (.Y(_01275_),
    .A(net2823));
 sg13g2_inv_1 _08070_ (.Y(_01276_),
    .A(net2221));
 sg13g2_inv_1 _08071_ (.Y(_01277_),
    .A(net2545));
 sg13g2_inv_1 _08072_ (.Y(_01278_),
    .A(\am_sdr0.cic0.comb1[1] ));
 sg13g2_inv_1 _08073_ (.Y(_01279_),
    .A(net2377));
 sg13g2_inv_1 _08074_ (.Y(_01280_),
    .A(net2547));
 sg13g2_inv_1 _08075_ (.Y(_01281_),
    .A(net2287));
 sg13g2_inv_1 _08076_ (.Y(_01282_),
    .A(net2661));
 sg13g2_inv_1 _08077_ (.Y(_01283_),
    .A(\am_sdr0.cic0.comb1_in_del[17] ));
 sg13g2_inv_1 _08078_ (.Y(_01284_),
    .A(net2597));
 sg13g2_inv_1 _08079_ (.Y(_01285_),
    .A(\am_sdr0.cic0.integ_sample[16] ));
 sg13g2_inv_1 _08080_ (.Y(_01286_),
    .A(net2709));
 sg13g2_inv_1 _08081_ (.Y(_01287_),
    .A(\am_sdr0.cic0.integ_sample[14] ));
 sg13g2_inv_1 _08082_ (.Y(_01288_),
    .A(\am_sdr0.cic0.integ_sample[13] ));
 sg13g2_inv_1 _08083_ (.Y(_01289_),
    .A(\am_sdr0.cic0.integ_sample[12] ));
 sg13g2_inv_1 _08084_ (.Y(_01290_),
    .A(net2292));
 sg13g2_inv_1 _08085_ (.Y(_01291_),
    .A(net2636));
 sg13g2_inv_1 _08086_ (.Y(_01292_),
    .A(\am_sdr0.cic0.comb1_in_del[9] ));
 sg13g2_inv_1 _08087_ (.Y(_01293_),
    .A(\am_sdr0.cic0.integ_sample[9] ));
 sg13g2_inv_1 _08088_ (.Y(_01294_),
    .A(net2703));
 sg13g2_inv_1 _08089_ (.Y(_01295_),
    .A(\am_sdr0.cic0.integ_sample[7] ));
 sg13g2_inv_1 _08090_ (.Y(_01296_),
    .A(\am_sdr0.cic0.integ_sample[6] ));
 sg13g2_inv_1 _08091_ (.Y(_01297_),
    .A(\am_sdr0.cic0.comb1_in_del[5] ));
 sg13g2_inv_1 _08092_ (.Y(_01298_),
    .A(net2626));
 sg13g2_inv_1 _08093_ (.Y(_01299_),
    .A(net2738));
 sg13g2_inv_1 _08094_ (.Y(_01300_),
    .A(net2464));
 sg13g2_inv_1 _08095_ (.Y(_01301_),
    .A(net2705));
 sg13g2_inv_1 _08096_ (.Y(_01302_),
    .A(\am_sdr0.cic0.integ_sample[1] ));
 sg13g2_inv_1 _08097_ (.Y(_01303_),
    .A(net2121));
 sg13g2_inv_2 _08098_ (.Y(_01304_),
    .A(net1698));
 sg13g2_inv_1 _08099_ (.Y(_01305_),
    .A(net2061));
 sg13g2_inv_1 _08100_ (.Y(_01306_),
    .A(net1795));
 sg13g2_inv_1 _08101_ (.Y(_01307_),
    .A(net2145));
 sg13g2_inv_1 _08102_ (.Y(_01308_),
    .A(net2256));
 sg13g2_inv_1 _08103_ (.Y(_01309_),
    .A(net2147));
 sg13g2_inv_1 _08104_ (.Y(_01310_),
    .A(net2376));
 sg13g2_inv_1 _08105_ (.Y(_01311_),
    .A(net2500));
 sg13g2_inv_1 _08106_ (.Y(_01312_),
    .A(net2335));
 sg13g2_inv_1 _08107_ (.Y(_01313_),
    .A(net2367));
 sg13g2_inv_1 _08108_ (.Y(_01314_),
    .A(\am_sdr0.cic1.comb3_in_del[11] ));
 sg13g2_inv_1 _08109_ (.Y(_01315_),
    .A(\am_sdr0.cic1.comb2[11] ));
 sg13g2_inv_1 _08110_ (.Y(_01316_),
    .A(net2087));
 sg13g2_inv_1 _08111_ (.Y(_01317_),
    .A(net2207));
 sg13g2_inv_1 _08112_ (.Y(_01318_),
    .A(\am_sdr0.cic1.comb3_in_del[8] ));
 sg13g2_inv_1 _08113_ (.Y(_01319_),
    .A(net2403));
 sg13g2_inv_1 _08114_ (.Y(_01320_),
    .A(\am_sdr0.cic1.comb3_in_del[7] ));
 sg13g2_inv_1 _08115_ (.Y(_01321_),
    .A(net2494));
 sg13g2_inv_1 _08116_ (.Y(_01322_),
    .A(\am_sdr0.cic1.comb3_in_del[6] ));
 sg13g2_inv_1 _08117_ (.Y(_01323_),
    .A(net2392));
 sg13g2_inv_1 _08118_ (.Y(_01324_),
    .A(net2102));
 sg13g2_inv_1 _08119_ (.Y(_01325_),
    .A(\am_sdr0.cic1.comb3_in_del[4] ));
 sg13g2_inv_1 _08120_ (.Y(_01326_),
    .A(net2370));
 sg13g2_inv_1 _08121_ (.Y(_01327_),
    .A(net2183));
 sg13g2_inv_1 _08122_ (.Y(_01328_),
    .A(net2189));
 sg13g2_inv_1 _08123_ (.Y(_01329_),
    .A(net2307));
 sg13g2_inv_1 _08124_ (.Y(_01330_),
    .A(net2166));
 sg13g2_inv_1 _08125_ (.Y(_01331_),
    .A(net1484));
 sg13g2_inv_1 _08126_ (.Y(_01332_),
    .A(net1264));
 sg13g2_inv_1 _08127_ (.Y(_01333_),
    .A(net1347));
 sg13g2_inv_1 _08128_ (.Y(_01334_),
    .A(net1366));
 sg13g2_inv_1 _08129_ (.Y(_01335_),
    .A(net1226));
 sg13g2_inv_1 _08130_ (.Y(_01336_),
    .A(net1241));
 sg13g2_inv_1 _08131_ (.Y(_01337_),
    .A(net1337));
 sg13g2_inv_1 _08132_ (.Y(_01338_),
    .A(net1283));
 sg13g2_inv_1 _08133_ (.Y(_01339_),
    .A(net2119));
 sg13g2_inv_1 _08134_ (.Y(_01340_),
    .A(net2760));
 sg13g2_inv_1 _08135_ (.Y(_01341_),
    .A(net2816));
 sg13g2_inv_1 _08136_ (.Y(_01342_),
    .A(net2773));
 sg13g2_inv_1 _08137_ (.Y(_01343_),
    .A(net2606));
 sg13g2_inv_1 _08138_ (.Y(_01344_),
    .A(net2398));
 sg13g2_inv_1 _08139_ (.Y(_01345_),
    .A(net2327));
 sg13g2_inv_1 _08140_ (.Y(_01346_),
    .A(\am_sdr0.cic1.comb1[12] ));
 sg13g2_inv_1 _08141_ (.Y(_01347_),
    .A(\am_sdr0.cic1.comb1[11] ));
 sg13g2_inv_1 _08142_ (.Y(_01348_),
    .A(net2329));
 sg13g2_inv_1 _08143_ (.Y(_01349_),
    .A(\am_sdr0.cic1.comb2_in_del[9] ));
 sg13g2_inv_1 _08144_ (.Y(_01350_),
    .A(\am_sdr0.cic1.comb1[9] ));
 sg13g2_inv_1 _08145_ (.Y(_01351_),
    .A(net2485));
 sg13g2_inv_1 _08146_ (.Y(_01352_),
    .A(net2442));
 sg13g2_inv_1 _08147_ (.Y(_01353_),
    .A(net2732));
 sg13g2_inv_1 _08148_ (.Y(_01354_),
    .A(net2583));
 sg13g2_inv_1 _08149_ (.Y(_01355_),
    .A(net2670));
 sg13g2_inv_1 _08150_ (.Y(_01356_),
    .A(net2263));
 sg13g2_inv_1 _08151_ (.Y(_01357_),
    .A(net2492));
 sg13g2_inv_1 _08152_ (.Y(_01358_),
    .A(net2468));
 sg13g2_inv_1 _08153_ (.Y(_01359_),
    .A(net2458));
 sg13g2_inv_1 _08154_ (.Y(_01360_),
    .A(net2388));
 sg13g2_inv_1 _08155_ (.Y(_01361_),
    .A(net2141));
 sg13g2_inv_1 _08156_ (.Y(_01362_),
    .A(\am_sdr0.cic1.integ_sample[18] ));
 sg13g2_inv_1 _08157_ (.Y(_01363_),
    .A(net2351));
 sg13g2_inv_1 _08158_ (.Y(_01364_),
    .A(\am_sdr0.cic1.integ_sample[16] ));
 sg13g2_inv_1 _08159_ (.Y(_01365_),
    .A(\am_sdr0.cic1.integ_sample[15] ));
 sg13g2_inv_1 _08160_ (.Y(_01366_),
    .A(net2579));
 sg13g2_inv_1 _08161_ (.Y(_01367_),
    .A(net2804));
 sg13g2_inv_1 _08162_ (.Y(_01368_),
    .A(net2713));
 sg13g2_inv_1 _08163_ (.Y(_01369_),
    .A(net2298));
 sg13g2_inv_1 _08164_ (.Y(_01370_),
    .A(\am_sdr0.cic1.integ_sample[10] ));
 sg13g2_inv_1 _08165_ (.Y(_01371_),
    .A(\am_sdr0.cic1.comb1_in_del[9] ));
 sg13g2_inv_1 _08166_ (.Y(_01372_),
    .A(net2903));
 sg13g2_inv_1 _08167_ (.Y(_01373_),
    .A(\am_sdr0.cic1.integ_sample[8] ));
 sg13g2_inv_1 _08168_ (.Y(_01374_),
    .A(net2569));
 sg13g2_inv_1 _08169_ (.Y(_01375_),
    .A(net2751));
 sg13g2_inv_1 _08170_ (.Y(_01376_),
    .A(\am_sdr0.cic1.comb1_in_del[5] ));
 sg13g2_inv_1 _08171_ (.Y(_01377_),
    .A(net2877));
 sg13g2_inv_1 _08172_ (.Y(_01378_),
    .A(\am_sdr0.cic1.integ_sample[4] ));
 sg13g2_inv_1 _08173_ (.Y(_01379_),
    .A(net2593));
 sg13g2_inv_1 _08174_ (.Y(_01380_),
    .A(net2561));
 sg13g2_inv_1 _08175_ (.Y(_01381_),
    .A(net2359));
 sg13g2_inv_1 _08176_ (.Y(_01382_),
    .A(net2035));
 sg13g2_inv_2 _08177_ (.Y(_01383_),
    .A(net1756));
 sg13g2_inv_2 _08178_ (.Y(_01384_),
    .A(net1691));
 sg13g2_inv_1 _08179_ (.Y(_01385_),
    .A(net2811));
 sg13g2_inv_1 _08180_ (.Y(_01386_),
    .A(net2634));
 sg13g2_inv_1 _08181_ (.Y(_01387_),
    .A(\am_sdr0.cic2.integ2[8] ));
 sg13g2_inv_1 _08182_ (.Y(_01388_),
    .A(net2834));
 sg13g2_inv_1 _08183_ (.Y(_01389_),
    .A(\am_sdr0.cic2.integ2[5] ));
 sg13g2_inv_1 _08184_ (.Y(_01390_),
    .A(net2915));
 sg13g2_inv_1 _08185_ (.Y(_01391_),
    .A(net2898));
 sg13g2_inv_1 _08186_ (.Y(_01392_),
    .A(\am_sdr0.cic2.integ1[8] ));
 sg13g2_inv_1 _08187_ (.Y(_01393_),
    .A(net2918));
 sg13g2_inv_1 _08188_ (.Y(_01394_),
    .A(net2057));
 sg13g2_inv_1 _08189_ (.Y(_01395_),
    .A(net1827));
 sg13g2_inv_1 _08190_ (.Y(_01396_),
    .A(net2339));
 sg13g2_inv_1 _08191_ (.Y(_01397_),
    .A(net2039));
 sg13g2_inv_1 _08192_ (.Y(_01398_),
    .A(net2344));
 sg13g2_inv_1 _08193_ (.Y(_01399_),
    .A(net2104));
 sg13g2_inv_1 _08194_ (.Y(_01400_),
    .A(net2314));
 sg13g2_inv_1 _08195_ (.Y(_01401_),
    .A(net2509));
 sg13g2_inv_1 _08196_ (.Y(_01402_),
    .A(net2368));
 sg13g2_inv_1 _08197_ (.Y(_01403_),
    .A(net2799));
 sg13g2_inv_1 _08198_ (.Y(_01404_),
    .A(net2333));
 sg13g2_inv_1 _08199_ (.Y(_01405_),
    .A(net2172));
 sg13g2_inv_1 _08200_ (.Y(_01406_),
    .A(net2325));
 sg13g2_inv_1 _08201_ (.Y(_01407_),
    .A(\am_sdr0.cic2.comb3_in_del[7] ));
 sg13g2_inv_1 _08202_ (.Y(_01408_),
    .A(\am_sdr0.cic2.comb2[7] ));
 sg13g2_inv_1 _08203_ (.Y(_01409_),
    .A(net2249));
 sg13g2_inv_1 _08204_ (.Y(_01410_),
    .A(\am_sdr0.cic2.comb3_in_del[5] ));
 sg13g2_inv_1 _08205_ (.Y(_01411_),
    .A(net2381));
 sg13g2_inv_1 _08206_ (.Y(_01412_),
    .A(\am_sdr0.cic2.comb3_in_del[4] ));
 sg13g2_inv_1 _08207_ (.Y(_01413_),
    .A(net2529));
 sg13g2_inv_1 _08208_ (.Y(_01414_),
    .A(net2125));
 sg13g2_inv_1 _08209_ (.Y(_01415_),
    .A(net2111));
 sg13g2_inv_1 _08210_ (.Y(_01416_),
    .A(net2083));
 sg13g2_inv_1 _08211_ (.Y(_01417_),
    .A(net1466));
 sg13g2_inv_1 _08212_ (.Y(_01418_),
    .A(net1287));
 sg13g2_inv_1 _08213_ (.Y(_01419_),
    .A(net1246));
 sg13g2_inv_1 _08214_ (.Y(_01420_),
    .A(net1285));
 sg13g2_inv_1 _08215_ (.Y(_01421_),
    .A(net1262));
 sg13g2_inv_1 _08216_ (.Y(_01422_),
    .A(net1450));
 sg13g2_inv_1 _08217_ (.Y(_01423_),
    .A(net1295));
 sg13g2_inv_1 _08218_ (.Y(_01424_),
    .A(net1369));
 sg13g2_inv_1 _08219_ (.Y(_01425_),
    .A(net1231));
 sg13g2_inv_1 _08220_ (.Y(_01426_),
    .A(net2315));
 sg13g2_inv_1 _08221_ (.Y(_01427_),
    .A(net2245));
 sg13g2_inv_1 _08222_ (.Y(_01428_),
    .A(net2659));
 sg13g2_inv_1 _08223_ (.Y(_01429_),
    .A(net2631));
 sg13g2_inv_1 _08224_ (.Y(_01430_),
    .A(net2855));
 sg13g2_inv_1 _08225_ (.Y(_01431_),
    .A(net2567));
 sg13g2_inv_1 _08226_ (.Y(_01432_),
    .A(\am_sdr0.cic2.comb2_in_del[13] ));
 sg13g2_inv_1 _08227_ (.Y(_01433_),
    .A(net2538));
 sg13g2_inv_1 _08228_ (.Y(_01434_),
    .A(\am_sdr0.cic2.comb2_in_del[12] ));
 sg13g2_inv_1 _08229_ (.Y(_01435_),
    .A(net2794));
 sg13g2_inv_1 _08230_ (.Y(_01436_),
    .A(net2251));
 sg13g2_inv_1 _08231_ (.Y(_01437_),
    .A(net2496));
 sg13g2_inv_1 _08232_ (.Y(_01438_),
    .A(net2281));
 sg13g2_inv_1 _08233_ (.Y(_01439_),
    .A(net2479));
 sg13g2_inv_1 _08234_ (.Y(_01440_),
    .A(net2520));
 sg13g2_inv_1 _08235_ (.Y(_01441_),
    .A(net2394));
 sg13g2_inv_1 _08236_ (.Y(_01442_),
    .A(net2386));
 sg13g2_inv_1 _08237_ (.Y(_01443_),
    .A(net2222));
 sg13g2_inv_1 _08238_ (.Y(_01444_),
    .A(\am_sdr0.cic2.comb1[3] ));
 sg13g2_inv_1 _08239_ (.Y(_01445_),
    .A(net2420));
 sg13g2_inv_1 _08240_ (.Y(_01446_),
    .A(net2312));
 sg13g2_inv_1 _08241_ (.Y(_01447_),
    .A(\am_sdr0.cic2.comb2_in_del[0] ));
 sg13g2_inv_1 _08242_ (.Y(_01448_),
    .A(net2383));
 sg13g2_inv_1 _08243_ (.Y(_01449_),
    .A(net1486));
 sg13g2_inv_1 _08244_ (.Y(_01450_),
    .A(net2342));
 sg13g2_inv_1 _08245_ (.Y(_01451_),
    .A(net2234));
 sg13g2_inv_1 _08246_ (.Y(_01452_),
    .A(net2296));
 sg13g2_inv_1 _08247_ (.Y(_01453_),
    .A(net2226));
 sg13g2_inv_1 _08248_ (.Y(_01454_),
    .A(net1384));
 sg13g2_inv_1 _08249_ (.Y(_01455_),
    .A(net2616));
 sg13g2_inv_1 _08250_ (.Y(_01456_),
    .A(net2356));
 sg13g2_inv_1 _08251_ (.Y(_01457_),
    .A(net2066));
 sg13g2_inv_1 _08252_ (.Y(_01458_),
    .A(net2077));
 sg13g2_inv_1 _08253_ (.Y(_01459_),
    .A(\am_sdr0.cic2.comb1_in_del[9] ));
 sg13g2_inv_1 _08254_ (.Y(_01460_),
    .A(net2361));
 sg13g2_inv_1 _08255_ (.Y(_01461_),
    .A(net2151));
 sg13g2_inv_1 _08256_ (.Y(_01462_),
    .A(net2396));
 sg13g2_inv_1 _08257_ (.Y(_01463_),
    .A(net2374));
 sg13g2_inv_1 _08258_ (.Y(_01464_),
    .A(net2654));
 sg13g2_inv_1 _08259_ (.Y(_01465_),
    .A(net2447));
 sg13g2_inv_1 _08260_ (.Y(_01466_),
    .A(net2137));
 sg13g2_inv_1 _08261_ (.Y(_01467_),
    .A(net2599));
 sg13g2_inv_1 _08262_ (.Y(_01468_),
    .A(net2453));
 sg13g2_inv_1 _08263_ (.Y(_01469_),
    .A(net2068));
 sg13g2_inv_2 _08264_ (.Y(_01470_),
    .A(net1739));
 sg13g2_inv_1 _08265_ (.Y(_01471_),
    .A(net2478));
 sg13g2_inv_1 _08266_ (.Y(_01472_),
    .A(\am_sdr0.cic3.integ3[5] ));
 sg13g2_inv_1 _08267_ (.Y(_01473_),
    .A(net2467));
 sg13g2_inv_1 _08268_ (.Y(_01474_),
    .A(\am_sdr0.cic3.integ2[8] ));
 sg13g2_inv_1 _08269_ (.Y(_01475_),
    .A(\am_sdr0.cic3.integ2[5] ));
 sg13g2_inv_1 _08270_ (.Y(_01476_),
    .A(net2879));
 sg13g2_inv_1 _08271_ (.Y(_01477_),
    .A(net2946));
 sg13g2_inv_1 _08272_ (.Y(_01478_),
    .A(\am_sdr0.cic3.integ1[8] ));
 sg13g2_inv_1 _08273_ (.Y(_01479_),
    .A(net2963));
 sg13g2_inv_1 _08274_ (.Y(_01480_),
    .A(net2191));
 sg13g2_inv_1 _08275_ (.Y(_01481_),
    .A(net1863));
 sg13g2_inv_1 _08276_ (.Y(_01482_),
    .A(net2423));
 sg13g2_inv_1 _08277_ (.Y(_01483_),
    .A(net2203));
 sg13g2_inv_1 _08278_ (.Y(_01484_),
    .A(net2490));
 sg13g2_inv_1 _08279_ (.Y(_01485_),
    .A(\am_sdr0.cic3.comb2[15] ));
 sg13g2_inv_1 _08280_ (.Y(_01486_),
    .A(net2300));
 sg13g2_inv_1 _08281_ (.Y(_01487_),
    .A(net2542));
 sg13g2_inv_1 _08282_ (.Y(_01488_),
    .A(net2270));
 sg13g2_inv_1 _08283_ (.Y(_01489_),
    .A(\am_sdr0.cic3.comb3_in_del[11] ));
 sg13g2_inv_1 _08284_ (.Y(_01490_),
    .A(net2213));
 sg13g2_inv_1 _08285_ (.Y(_01491_),
    .A(\am_sdr0.cic3.comb3_in_del[10] ));
 sg13g2_inv_1 _08286_ (.Y(_01492_),
    .A(\am_sdr0.cic3.comb2[10] ));
 sg13g2_inv_1 _08287_ (.Y(_01493_),
    .A(net2181));
 sg13g2_inv_1 _08288_ (.Y(_01494_),
    .A(net2210));
 sg13g2_inv_1 _08289_ (.Y(_01495_),
    .A(\am_sdr0.cic3.comb3_in_del[7] ));
 sg13g2_inv_1 _08290_ (.Y(_01496_),
    .A(net2264));
 sg13g2_inv_1 _08291_ (.Y(_01497_),
    .A(net2199));
 sg13g2_inv_1 _08292_ (.Y(_01498_),
    .A(\am_sdr0.cic3.comb3_in_del[5] ));
 sg13g2_inv_1 _08293_ (.Y(_01499_),
    .A(net2232));
 sg13g2_inv_1 _08294_ (.Y(_01500_),
    .A(\am_sdr0.cic3.comb3_in_del[4] ));
 sg13g2_inv_1 _08295_ (.Y(_01501_),
    .A(net2228));
 sg13g2_inv_1 _08296_ (.Y(_01502_),
    .A(\am_sdr0.cic3.comb3_in_del[3] ));
 sg13g2_inv_1 _08297_ (.Y(_01503_),
    .A(net2188));
 sg13g2_inv_1 _08298_ (.Y(_01504_),
    .A(net2089));
 sg13g2_inv_1 _08299_ (.Y(_01505_),
    .A(net2045));
 sg13g2_inv_1 _08300_ (.Y(_01506_),
    .A(net1528));
 sg13g2_inv_1 _08301_ (.Y(_01507_),
    .A(net1332));
 sg13g2_inv_1 _08302_ (.Y(_01508_),
    .A(net1355));
 sg13g2_inv_1 _08303_ (.Y(_01509_),
    .A(net1349));
 sg13g2_inv_1 _08304_ (.Y(_01510_),
    .A(net1319));
 sg13g2_inv_1 _08305_ (.Y(_01511_),
    .A(net1462));
 sg13g2_inv_1 _08306_ (.Y(_01512_),
    .A(net1452));
 sg13g2_inv_1 _08307_ (.Y(_01513_),
    .A(net2149));
 sg13g2_inv_1 _08308_ (.Y(_01514_),
    .A(net1516));
 sg13g2_inv_1 _08309_ (.Y(_01515_),
    .A(\am_sdr0.cic3.comb1[19] ));
 sg13g2_inv_1 _08310_ (.Y(_01516_),
    .A(net2363));
 sg13g2_inv_1 _08311_ (.Y(_01517_),
    .A(net2736));
 sg13g2_inv_1 _08312_ (.Y(_01518_),
    .A(net2365));
 sg13g2_inv_1 _08313_ (.Y(_01519_),
    .A(net2758));
 sg13g2_inv_1 _08314_ (.Y(_01520_),
    .A(net2321));
 sg13g2_inv_1 _08315_ (.Y(_01521_),
    .A(net2540));
 sg13g2_inv_1 _08316_ (.Y(_01522_),
    .A(net2522));
 sg13g2_inv_1 _08317_ (.Y(_01523_),
    .A(net2236));
 sg13g2_inv_1 _08318_ (.Y(_01524_),
    .A(net2379));
 sg13g2_inv_1 _08319_ (.Y(_01525_),
    .A(\am_sdr0.cic3.comb2_in_del[9] ));
 sg13g2_inv_1 _08320_ (.Y(_01526_),
    .A(net2776));
 sg13g2_inv_1 _08321_ (.Y(_01527_),
    .A(\am_sdr0.cic3.comb1[8] ));
 sg13g2_inv_1 _08322_ (.Y(_01528_),
    .A(net2575));
 sg13g2_inv_1 _08323_ (.Y(_01529_),
    .A(\am_sdr0.cic3.comb1[6] ));
 sg13g2_inv_1 _08324_ (.Y(_01530_),
    .A(\am_sdr0.cic3.comb2_in_del[5] ));
 sg13g2_inv_1 _08325_ (.Y(_01531_),
    .A(net2449));
 sg13g2_inv_1 _08326_ (.Y(_01532_),
    .A(net2595));
 sg13g2_inv_1 _08327_ (.Y(_01533_),
    .A(net2553));
 sg13g2_inv_1 _08328_ (.Y(_01534_),
    .A(net2238));
 sg13g2_inv_1 _08329_ (.Y(_01535_),
    .A(net2347));
 sg13g2_inv_1 _08330_ (.Y(_01536_),
    .A(net2358));
 sg13g2_inv_1 _08331_ (.Y(_01537_),
    .A(net2260));
 sg13g2_inv_1 _08332_ (.Y(_01538_),
    .A(net2194));
 sg13g2_inv_1 _08333_ (.Y(_01539_),
    .A(net2476));
 sg13g2_inv_1 _08334_ (.Y(_01540_),
    .A(\am_sdr0.cic3.integ_sample[17] ));
 sg13g2_inv_1 _08335_ (.Y(_01541_),
    .A(net2621));
 sg13g2_inv_1 _08336_ (.Y(_01542_),
    .A(\am_sdr0.cic3.comb1_in_del[15] ));
 sg13g2_inv_1 _08337_ (.Y(_01543_),
    .A(\am_sdr0.cic3.integ_sample[15] ));
 sg13g2_inv_1 _08338_ (.Y(_01544_),
    .A(net2680));
 sg13g2_inv_1 _08339_ (.Y(_01545_),
    .A(\am_sdr0.cic3.integ_sample[13] ));
 sg13g2_inv_1 _08340_ (.Y(_01546_),
    .A(net2725));
 sg13g2_inv_1 _08341_ (.Y(_01547_),
    .A(net2302));
 sg13g2_inv_1 _08342_ (.Y(_01548_),
    .A(net2425));
 sg13g2_inv_1 _08343_ (.Y(_01549_),
    .A(\am_sdr0.cic3.comb1_in_del[9] ));
 sg13g2_inv_1 _08344_ (.Y(_01550_),
    .A(net2921));
 sg13g2_inv_1 _08345_ (.Y(_01551_),
    .A(net2504));
 sg13g2_inv_1 _08346_ (.Y(_01552_),
    .A(net2507));
 sg13g2_inv_1 _08347_ (.Y(_01553_),
    .A(net2587));
 sg13g2_inv_1 _08348_ (.Y(_01554_),
    .A(\am_sdr0.cic3.comb1_in_del[5] ));
 sg13g2_inv_1 _08349_ (.Y(_01555_),
    .A(net2891));
 sg13g2_inv_1 _08350_ (.Y(_01556_),
    .A(net2513));
 sg13g2_inv_1 _08351_ (.Y(_01557_),
    .A(net2445));
 sg13g2_inv_1 _08352_ (.Y(_01558_),
    .A(net2483));
 sg13g2_inv_1 _08353_ (.Y(_01559_),
    .A(net2349));
 sg13g2_inv_1 _08354_ (.Y(_01560_),
    .A(net2413));
 sg13g2_inv_1 _08355_ (.Y(_01561_),
    .A(net2262));
 sg13g2_inv_1 _08356_ (.Y(_01562_),
    .A(\am_sdr0.am0.sqrt_state[1] ));
 sg13g2_inv_1 _08357_ (.Y(_01563_),
    .A(\am_sdr0.am0.sum[1] ));
 sg13g2_inv_1 _08358_ (.Y(_01564_),
    .A(net2455));
 sg13g2_inv_1 _08359_ (.Y(_01565_),
    .A(net1966));
 sg13g2_inv_1 _08360_ (.Y(_01566_),
    .A(\am_sdr0.am0.m_count[3] ));
 sg13g2_inv_1 _08361_ (.Y(_01567_),
    .A(\am_sdr0.am0.sqrt_done ));
 sg13g2_inv_1 _08362_ (.Y(_01568_),
    .A(net1258));
 sg13g2_inv_1 _08363_ (.Y(_01569_),
    .A(net2113));
 sg13g2_inv_1 _08364_ (.Y(_01570_),
    .A(\am_sdr0.am0.count2[0] ));
 sg13g2_inv_1 _08365_ (.Y(_01571_),
    .A(net2097));
 sg13g2_inv_1 _08366_ (.Y(_01572_),
    .A(net1254));
 sg13g2_inv_1 _08367_ (.Y(_01573_),
    .A(net1256));
 sg13g2_inv_1 _08368_ (.Y(_01574_),
    .A(\am_sdr0.am0.load_tick ));
 sg13g2_inv_2 _08369_ (.Y(_01575_),
    .A(net2947));
 sg13g2_inv_2 _08370_ (.Y(_01576_),
    .A(net1654));
 sg13g2_inv_1 _08371_ (.Y(_01577_),
    .A(net1651));
 sg13g2_inv_1 _08372_ (.Y(_01578_),
    .A(net1525));
 sg13g2_inv_2 _08373_ (.Y(_01579_),
    .A(net1648));
 sg13g2_inv_1 _08374_ (.Y(_01580_),
    .A(\am_sdr0.am0.multA[15] ));
 sg13g2_inv_1 _08375_ (.Y(_01581_),
    .A(net1427));
 sg13g2_inv_1 _08376_ (.Y(_01582_),
    .A(\am_sdr0.count[7] ));
 sg13g2_inv_2 _08377_ (.Y(_01583_),
    .A(net1870));
 sg13g2_inv_2 _08378_ (.Y(_01584_),
    .A(\am_sdr0.count[5] ));
 sg13g2_inv_2 _08379_ (.Y(_01585_),
    .A(\am_sdr0.count[4] ));
 sg13g2_inv_2 _08380_ (.Y(_01586_),
    .A(net3157));
 sg13g2_inv_1 _08381_ (.Y(_01587_),
    .A(\am_sdr0.count[2] ));
 sg13g2_inv_1 _08382_ (.Y(_01588_),
    .A(\am_sdr0.cic0.integ2[20] ));
 sg13g2_inv_1 _08383_ (.Y(_01589_),
    .A(\am_sdr0.cic0.integ3[17] ));
 sg13g2_inv_1 _08384_ (.Y(_01590_),
    .A(\am_sdr0.cic1.integ2[20] ));
 sg13g2_inv_1 _08385_ (.Y(_01591_),
    .A(\am_sdr0.cic1.integ3[17] ));
 sg13g2_inv_1 _08386_ (.Y(_01592_),
    .A(_00069_));
 sg13g2_inv_1 _08387_ (.Y(_01593_),
    .A(_00072_));
 sg13g2_inv_1 _08388_ (.Y(_01594_),
    .A(net1164));
 sg13g2_inv_1 _08389_ (.Y(_01595_),
    .A(net1163));
 sg13g2_and3_1 _08390_ (.X(_01596_),
    .A(\am_sdr0.am0.m_count[1] ),
    .B(\am_sdr0.am0.m_count[0] ),
    .C(\am_sdr0.am0.m_count[2] ));
 sg13g2_nand3_1 _08391_ (.B(\am_sdr0.am0.m_count[0] ),
    .C(\am_sdr0.am0.m_count[2] ),
    .A(\am_sdr0.am0.m_count[1] ),
    .Y(_01597_));
 sg13g2_nor2_1 _08392_ (.A(\am_sdr0.am0.m_count[3] ),
    .B(_01597_),
    .Y(_01598_));
 sg13g2_nand2_2 _08393_ (.Y(_01599_),
    .A(_01566_),
    .B(_01596_));
 sg13g2_a21oi_1 _08394_ (.A1(\am_sdr0.am0.state[2] ),
    .A2(net1608),
    .Y(_01600_),
    .B1(net1275));
 sg13g2_nor2_1 _08395_ (.A(net1893),
    .B(net1276),
    .Y(_00020_));
 sg13g2_a21oi_1 _08396_ (.A1(_01567_),
    .A2(net1258),
    .Y(_01601_),
    .B1(net1260));
 sg13g2_nor2_1 _08397_ (.A(net1893),
    .B(net1261),
    .Y(_00021_));
 sg13g2_a21oi_1 _08398_ (.A1(net2827),
    .A2(net1608),
    .Y(_01602_),
    .B1(net1873));
 sg13g2_nor2_1 _08399_ (.A(net1893),
    .B(_01602_),
    .Y(_00019_));
 sg13g2_a21oi_1 _08400_ (.A1(\am_sdr0.am0.state[0] ),
    .A2(_01574_),
    .Y(_01603_),
    .B1(net1892));
 sg13g2_o21ai_1 _08401_ (.B1(_01603_),
    .Y(_00018_),
    .A1(_01567_),
    .A2(_01568_));
 sg13g2_nand2_1 _08402_ (.Y(_01604_),
    .A(net1653),
    .B(net1652));
 sg13g2_nand2_2 _08403_ (.Y(_01605_),
    .A(_01575_),
    .B(_01576_));
 sg13g2_nor2_1 _08404_ (.A(net1651),
    .B(_01605_),
    .Y(_01606_));
 sg13g2_a21oi_1 _08405_ (.A1(net1653),
    .A2(net1652),
    .Y(_01607_),
    .B1(_01606_));
 sg13g2_nand2_1 _08406_ (.Y(_01608_),
    .A(net1525),
    .B(net1650));
 sg13g2_nand2_1 _08407_ (.Y(_01609_),
    .A(net1653),
    .B(net1654));
 sg13g2_nand4_1 _08408_ (.B(net1649),
    .C(_01605_),
    .A(net1525),
    .Y(_01610_),
    .D(_01609_));
 sg13g2_o21ai_1 _08409_ (.B1(_01610_),
    .Y(_00001_),
    .A1(net1648),
    .A2(_01607_));
 sg13g2_nand2_2 _08410_ (.Y(_01611_),
    .A(net1653),
    .B(_01576_));
 sg13g2_a21oi_1 _08411_ (.A1(net1653),
    .A2(_01576_),
    .Y(_01612_),
    .B1(_01577_));
 sg13g2_o21ai_1 _08412_ (.B1(_01579_),
    .Y(_01613_),
    .A1(net1651),
    .A2(net2603));
 sg13g2_nand2_1 _08413_ (.Y(_01614_),
    .A(_01577_),
    .B(_01611_));
 sg13g2_nand2_1 _08414_ (.Y(_01615_),
    .A(net1651),
    .B(_01609_));
 sg13g2_nand3_1 _08415_ (.B(_01614_),
    .C(_01615_),
    .A(net1649),
    .Y(_01616_));
 sg13g2_o21ai_1 _08416_ (.B1(_01616_),
    .Y(_00002_),
    .A1(_01612_),
    .A2(_01613_));
 sg13g2_nand2_1 _08417_ (.Y(_01617_),
    .A(_01575_),
    .B(net1654));
 sg13g2_nand2_1 _08418_ (.Y(_01618_),
    .A(_01577_),
    .B(_01617_));
 sg13g2_nand3b_1 _08419_ (.B(_01618_),
    .C(net1649),
    .Y(_01619_),
    .A_N(_01612_));
 sg13g2_o21ai_1 _08420_ (.B1(_01615_),
    .Y(_01620_),
    .A1(net1652),
    .A2(net2409));
 sg13g2_o21ai_1 _08421_ (.B1(_01619_),
    .Y(_00003_),
    .A1(net1649),
    .A2(_01620_));
 sg13g2_nor2_1 _08422_ (.A(net1525),
    .B(net1649),
    .Y(_01621_));
 sg13g2_nand2_1 _08423_ (.Y(_01622_),
    .A(_01578_),
    .B(_01579_));
 sg13g2_nor2_1 _08424_ (.A(_01575_),
    .B(net1651),
    .Y(_01623_));
 sg13g2_a21oi_2 _08425_ (.B1(_01579_),
    .Y(_01624_),
    .A2(_01623_),
    .A1(net1654));
 sg13g2_nand2_2 _08426_ (.Y(_01625_),
    .A(net1652),
    .B(_01605_));
 sg13g2_a22oi_1 _08427_ (.Y(_00004_),
    .B1(_01624_),
    .B2(_01625_),
    .A2(_01621_),
    .A1(_01617_));
 sg13g2_o21ai_1 _08428_ (.B1(_01614_),
    .Y(_01626_),
    .A1(net1654),
    .A2(_01604_));
 sg13g2_a21oi_1 _08429_ (.A1(net1649),
    .A2(_01605_),
    .Y(_01627_),
    .B1(_01626_));
 sg13g2_a21oi_1 _08430_ (.A1(net1650),
    .A2(_01626_),
    .Y(_00005_),
    .B1(_01627_));
 sg13g2_nor3_1 _08431_ (.A(_01576_),
    .B(net1649),
    .C(net2603),
    .Y(_01628_));
 sg13g2_a221oi_1 _08432_ (.B2(_01604_),
    .C1(_01628_),
    .B1(_01624_),
    .A1(_01576_),
    .Y(_00006_),
    .A2(_01621_));
 sg13g2_o21ai_1 _08433_ (.B1(net1526),
    .Y(_00007_),
    .A1(net1650),
    .A2(_01625_));
 sg13g2_a21oi_1 _08434_ (.A1(net1651),
    .A2(_01609_),
    .Y(_01629_),
    .B1(_01623_));
 sg13g2_inv_1 _08435_ (.Y(_00008_),
    .A(_01629_));
 sg13g2_nand2b_1 _08436_ (.Y(_01630_),
    .B(net1169),
    .A_N(net1655));
 sg13g2_xnor2_1 _08437_ (.Y(_00030_),
    .A(net1505),
    .B(_01630_));
 sg13g2_nor2_1 _08438_ (.A(net1169),
    .B(\am_sdr0.mix0.sin_q[1] ),
    .Y(_01631_));
 sg13g2_a21oi_1 _08439_ (.A1(_00040_),
    .A2(_01631_),
    .Y(_01632_),
    .B1(net1655));
 sg13g2_o21ai_1 _08440_ (.B1(_01632_),
    .Y(_01633_),
    .A1(_00040_),
    .A2(_01631_));
 sg13g2_nand2_1 _08441_ (.Y(_01634_),
    .A(net1655),
    .B(net1460));
 sg13g2_nand2_1 _08442_ (.Y(_00031_),
    .A(_01633_),
    .B(_01634_));
 sg13g2_xor2_1 _08443_ (.B(_01632_),
    .A(net1250),
    .X(_00032_));
 sg13g2_nor4_2 _08444_ (.A(net1169),
    .B(\am_sdr0.mix0.sin_q[1] ),
    .C(\am_sdr0.mix0.sin_q[2] ),
    .Y(_01635_),
    .D(net1250));
 sg13g2_inv_1 _08445_ (.Y(_01636_),
    .A(_01635_));
 sg13g2_a21oi_1 _08446_ (.A1(_00041_),
    .A2(_01635_),
    .Y(_01637_),
    .B1(net1655));
 sg13g2_o21ai_1 _08447_ (.B1(_01637_),
    .Y(_01638_),
    .A1(_00041_),
    .A2(_01635_));
 sg13g2_nand2_1 _08448_ (.Y(_01639_),
    .A(net1655),
    .B(net1326));
 sg13g2_nand2_1 _08449_ (.Y(_00033_),
    .A(_01638_),
    .B(_01639_));
 sg13g2_xor2_1 _08450_ (.B(_01637_),
    .A(net1198),
    .X(_00034_));
 sg13g2_nor3_1 _08451_ (.A(\am_sdr0.mix0.sin_q[4] ),
    .B(net1198),
    .C(_01636_),
    .Y(_01640_));
 sg13g2_a21o_1 _08452_ (.A2(_01640_),
    .A1(_00042_),
    .B1(net1655),
    .X(_01641_));
 sg13g2_nor2_1 _08453_ (.A(_00042_),
    .B(_01640_),
    .Y(_01642_));
 sg13g2_nand2_1 _08454_ (.Y(_01643_),
    .A(net1655),
    .B(net1206));
 sg13g2_o21ai_1 _08455_ (.B1(_01643_),
    .Y(_00035_),
    .A1(_01641_),
    .A2(_01642_));
 sg13g2_xnor2_1 _08456_ (.Y(_00036_),
    .A(net1196),
    .B(_01641_));
 sg13g2_nand2b_1 _08457_ (.Y(_01644_),
    .B(net1168),
    .A_N(net1656));
 sg13g2_xnor2_1 _08458_ (.Y(_00023_),
    .A(net2255),
    .B(_01644_));
 sg13g2_nor2_1 _08459_ (.A(net1168),
    .B(\am_sdr0.mix0.cos_q[1] ),
    .Y(_01645_));
 sg13g2_a21oi_1 _08460_ (.A1(_00043_),
    .A2(_01645_),
    .Y(_01646_),
    .B1(net1656));
 sg13g2_o21ai_1 _08461_ (.B1(_01646_),
    .Y(_01647_),
    .A1(_00043_),
    .A2(_01645_));
 sg13g2_nand2_1 _08462_ (.Y(_01648_),
    .A(net1656),
    .B(net1445));
 sg13g2_nand2_1 _08463_ (.Y(_00024_),
    .A(_01647_),
    .B(net1446));
 sg13g2_xor2_1 _08464_ (.B(_01646_),
    .A(net1311),
    .X(_00025_));
 sg13g2_nor4_2 _08465_ (.A(net1168),
    .B(\am_sdr0.mix0.cos_q[1] ),
    .C(\am_sdr0.mix0.cos_q[2] ),
    .Y(_01649_),
    .D(\am_sdr0.mix0.cos_q[3] ));
 sg13g2_inv_1 _08466_ (.Y(_01650_),
    .A(_01649_));
 sg13g2_a21oi_1 _08467_ (.A1(_00044_),
    .A2(_01649_),
    .Y(_01651_),
    .B1(net1656));
 sg13g2_o21ai_1 _08468_ (.B1(_01651_),
    .Y(_01652_),
    .A1(_00044_),
    .A2(_01649_));
 sg13g2_nand2_1 _08469_ (.Y(_01653_),
    .A(net1656),
    .B(net1266));
 sg13g2_nand2_1 _08470_ (.Y(_00026_),
    .A(_01652_),
    .B(net1267));
 sg13g2_xor2_1 _08471_ (.B(_01651_),
    .A(net1237),
    .X(_00027_));
 sg13g2_nor3_1 _08472_ (.A(net1266),
    .B(net1237),
    .C(_01650_),
    .Y(_01654_));
 sg13g2_a21o_1 _08473_ (.A2(_01654_),
    .A1(_00045_),
    .B1(net1656),
    .X(_01655_));
 sg13g2_nor2_1 _08474_ (.A(_00045_),
    .B(_01654_),
    .Y(_01656_));
 sg13g2_nand2_1 _08475_ (.Y(_01657_),
    .A(net1655),
    .B(net2050));
 sg13g2_o21ai_1 _08476_ (.B1(_01657_),
    .Y(_00028_),
    .A1(_01655_),
    .A2(_01656_));
 sg13g2_xnor2_1 _08477_ (.Y(_00029_),
    .A(net1215),
    .B(_01655_));
 sg13g2_nor2b_1 _08478_ (.A(_01625_),
    .B_N(_01609_),
    .Y(_01658_));
 sg13g2_o21ai_1 _08479_ (.B1(net1648),
    .Y(_01659_),
    .A1(_01623_),
    .A2(_01658_));
 sg13g2_o21ai_1 _08480_ (.B1(_01659_),
    .Y(_00009_),
    .A1(_01605_),
    .A2(_01622_));
 sg13g2_a21oi_1 _08481_ (.A1(net1653),
    .A2(net1654),
    .Y(_01660_),
    .B1(net1651));
 sg13g2_nor2_1 _08482_ (.A(_01577_),
    .B(net2603),
    .Y(_01661_));
 sg13g2_or3_1 _08483_ (.A(net1648),
    .B(_01660_),
    .C(_01661_),
    .X(_01662_));
 sg13g2_o21ai_1 _08484_ (.B1(_01662_),
    .Y(_00010_),
    .A1(_01579_),
    .A2(_01611_));
 sg13g2_nand3_1 _08485_ (.B(net1654),
    .C(net1652),
    .A(_01575_),
    .Y(_01663_));
 sg13g2_o21ai_1 _08486_ (.B1(_01614_),
    .Y(_01664_),
    .A1(_01577_),
    .A2(net2409));
 sg13g2_a22oi_1 _08487_ (.Y(_00011_),
    .B1(_01664_),
    .B2(_01579_),
    .A2(_01663_),
    .A1(_01624_));
 sg13g2_nand3_1 _08488_ (.B(_01615_),
    .C(_01618_),
    .A(net1648),
    .Y(_01665_));
 sg13g2_nor2_1 _08489_ (.A(_01578_),
    .B(_01605_),
    .Y(_01666_));
 sg13g2_o21ai_1 _08490_ (.B1(_01665_),
    .Y(_00012_),
    .A1(net1648),
    .A2(_01666_));
 sg13g2_xnor2_1 _08491_ (.Y(_01667_),
    .A(net1648),
    .B(_01611_));
 sg13g2_nor2_1 _08492_ (.A(_01606_),
    .B(_01667_),
    .Y(_00013_));
 sg13g2_o21ai_1 _08493_ (.B1(_01665_),
    .Y(_00014_),
    .A1(net1648),
    .A2(_01629_));
 sg13g2_a21o_1 _08494_ (.A2(net1651),
    .A1(net1653),
    .B1(_01660_),
    .X(_00000_));
 sg13g2_and3_1 _08495_ (.X(_00015_),
    .A(net2827),
    .B(net2024),
    .C(net1610));
 sg13g2_and3_1 _08496_ (.X(_00016_),
    .A(net2021),
    .B(net1273),
    .C(\am_sdr0.am0.load_tick ));
 sg13g2_and3_1 _08497_ (.X(_00017_),
    .A(net2801),
    .B(net2024),
    .C(net1610));
 sg13g2_nor2_2 _08498_ (.A(\am_sdr0.am0.state[2] ),
    .B(\am_sdr0.am0.state[1] ),
    .Y(_01668_));
 sg13g2_nor3_1 _08499_ (.A(\am_sdr0.am0.state[2] ),
    .B(\am_sdr0.am0.state[1] ),
    .C(net1873),
    .Y(_01669_));
 sg13g2_inv_1 _08500_ (.Y(_01670_),
    .A(net1620));
 sg13g2_o21ai_1 _08501_ (.B1(net2024),
    .Y(_01671_),
    .A1(\am_sdr0.am0.state[4] ),
    .A2(_01670_));
 sg13g2_inv_1 _08502_ (.Y(_01672_),
    .A(net1587));
 sg13g2_nor2_1 _08503_ (.A(net1892),
    .B(_01668_),
    .Y(_01673_));
 sg13g2_a22oi_1 _08504_ (.Y(_01674_),
    .B1(net1604),
    .B2(net1166),
    .A2(net1587),
    .A1(\am_sdr0.am0.m_count[0] ));
 sg13g2_inv_1 _08505_ (.Y(_00079_),
    .A(net1167));
 sg13g2_a21oi_1 _08506_ (.A1(\am_sdr0.am0.m_count[0] ),
    .A2(_01672_),
    .Y(_01675_),
    .B1(net2162));
 sg13g2_and3_1 _08507_ (.X(_01676_),
    .A(net2162),
    .B(\am_sdr0.am0.m_count[0] ),
    .C(_01672_));
 sg13g2_nor3_1 _08508_ (.A(\am_sdr0.am0.state[2] ),
    .B(\am_sdr0.am0.state[1] ),
    .C(net1587),
    .Y(_01677_));
 sg13g2_nor3_1 _08509_ (.A(net2163),
    .B(_01676_),
    .C(_01677_),
    .Y(_00080_));
 sg13g2_o21ai_1 _08510_ (.B1(_01672_),
    .Y(_01678_),
    .A1(_01596_),
    .A2(_01668_));
 sg13g2_o21ai_1 _08511_ (.B1(_01678_),
    .Y(_01679_),
    .A1(net2778),
    .A2(_01676_));
 sg13g2_inv_1 _08512_ (.Y(_00081_),
    .A(net2779));
 sg13g2_and2_1 _08513_ (.A(net3178),
    .B(_01678_),
    .X(_01680_));
 sg13g2_or3_1 _08514_ (.A(_00015_),
    .B(_00017_),
    .C(_01680_),
    .X(_00082_));
 sg13g2_a22oi_1 _08515_ (.Y(_01681_),
    .B1(_01669_),
    .B2(net3159),
    .A2(net2897),
    .A1(\am_sdr0.am0.Q_in[0] ));
 sg13g2_nor2_1 _08516_ (.A(net1585),
    .B(net3160),
    .Y(_01682_));
 sg13g2_a221oi_1 _08517_ (.B2(net2821),
    .C1(_01682_),
    .B1(net1605),
    .A1(\am_sdr0.am0.multB[0] ),
    .Y(_01683_),
    .A2(net1585));
 sg13g2_inv_1 _08518_ (.Y(_00083_),
    .A(net2822));
 sg13g2_nand2_1 _08519_ (.Y(_01684_),
    .A(net2048),
    .B(net1604));
 sg13g2_nand2_1 _08520_ (.Y(_01685_),
    .A(\am_sdr0.am0.multB[1] ),
    .B(net1585));
 sg13g2_a22oi_1 _08521_ (.Y(_01686_),
    .B1(net1620),
    .B2(\am_sdr0.am0.I_in[1] ),
    .A2(net2897),
    .A1(\am_sdr0.am0.Q_in[1] ));
 sg13g2_or2_1 _08522_ (.X(_01687_),
    .B(_01686_),
    .A(net1587));
 sg13g2_nand3_1 _08523_ (.B(_01685_),
    .C(_01687_),
    .A(_01684_),
    .Y(_00084_));
 sg13g2_nand2_1 _08524_ (.Y(_01688_),
    .A(net1493),
    .B(net1604));
 sg13g2_nand2_1 _08525_ (.Y(_01689_),
    .A(\am_sdr0.am0.multB[2] ),
    .B(net1586));
 sg13g2_a22oi_1 _08526_ (.Y(_01690_),
    .B1(net1620),
    .B2(\am_sdr0.am0.I_in[2] ),
    .A2(net1873),
    .A1(\am_sdr0.am0.Q_in[2] ));
 sg13g2_or2_1 _08527_ (.X(_01691_),
    .B(_01690_),
    .A(net1585));
 sg13g2_nand3_1 _08528_ (.B(_01689_),
    .C(_01691_),
    .A(_01688_),
    .Y(_00085_));
 sg13g2_nand2_1 _08529_ (.Y(_01692_),
    .A(net1520),
    .B(net1604));
 sg13g2_nand2_1 _08530_ (.Y(_01693_),
    .A(net1493),
    .B(net1585));
 sg13g2_a22oi_1 _08531_ (.Y(_01694_),
    .B1(net1620),
    .B2(\am_sdr0.am0.I_in[3] ),
    .A2(net1873),
    .A1(\am_sdr0.am0.Q_in[3] ));
 sg13g2_or2_1 _08532_ (.X(_01695_),
    .B(_01694_),
    .A(net1585));
 sg13g2_nand3_1 _08533_ (.B(_01693_),
    .C(_01695_),
    .A(_01692_),
    .Y(_00086_));
 sg13g2_nand2_1 _08534_ (.Y(_01696_),
    .A(net1510),
    .B(net1604));
 sg13g2_nand2_1 _08535_ (.Y(_01697_),
    .A(\am_sdr0.am0.multB[4] ),
    .B(net1586));
 sg13g2_a22oi_1 _08536_ (.Y(_01698_),
    .B1(net1620),
    .B2(\am_sdr0.am0.I_in[4] ),
    .A2(net1873),
    .A1(\am_sdr0.am0.Q_in[4] ));
 sg13g2_or2_1 _08537_ (.X(_01699_),
    .B(_01698_),
    .A(net1585));
 sg13g2_nand3_1 _08538_ (.B(_01697_),
    .C(_01699_),
    .A(_01696_),
    .Y(_00087_));
 sg13g2_nand2_1 _08539_ (.Y(_01700_),
    .A(net2037),
    .B(net1604));
 sg13g2_nand2_1 _08540_ (.Y(_01701_),
    .A(net1510),
    .B(net1588));
 sg13g2_a22oi_1 _08541_ (.Y(_01702_),
    .B1(net1620),
    .B2(\am_sdr0.am0.I_in[5] ),
    .A2(net1873),
    .A1(\am_sdr0.am0.Q_in[5] ));
 sg13g2_or2_1 _08542_ (.X(_01703_),
    .B(_01702_),
    .A(net1585));
 sg13g2_nand3_1 _08543_ (.B(_01701_),
    .C(_01703_),
    .A(_01700_),
    .Y(_00088_));
 sg13g2_nand2_1 _08544_ (.Y(_01704_),
    .A(net1427),
    .B(net1604));
 sg13g2_nand2_1 _08545_ (.Y(_01705_),
    .A(\am_sdr0.am0.multB[6] ),
    .B(net1588));
 sg13g2_a22oi_1 _08546_ (.Y(_01706_),
    .B1(net1620),
    .B2(\am_sdr0.am0.I_in[6] ),
    .A2(net1873),
    .A1(\am_sdr0.am0.Q_in[6] ));
 sg13g2_or2_1 _08547_ (.X(_01707_),
    .B(_01706_),
    .A(net1587));
 sg13g2_nand3_1 _08548_ (.B(_01705_),
    .C(_01707_),
    .A(_01704_),
    .Y(_00089_));
 sg13g2_a22oi_1 _08549_ (.Y(_01708_),
    .B1(net1620),
    .B2(\am_sdr0.am0.I_in[7] ),
    .A2(net1873),
    .A1(\am_sdr0.am0.Q_in[7] ));
 sg13g2_or2_1 _08550_ (.X(_01709_),
    .B(_01708_),
    .A(net1587));
 sg13g2_o21ai_1 _08551_ (.B1(net1568),
    .Y(_00090_),
    .A1(_01581_),
    .A2(_01672_));
 sg13g2_a21o_1 _08552_ (.A2(net1586),
    .A1(net3113),
    .B1(_01682_),
    .X(_00091_));
 sg13g2_nand2_1 _08553_ (.Y(_01710_),
    .A(net3113),
    .B(net1604));
 sg13g2_nand2_1 _08554_ (.Y(_01711_),
    .A(net2925),
    .B(net1587));
 sg13g2_nand3_1 _08555_ (.B(_01710_),
    .C(_01711_),
    .A(_01687_),
    .Y(_00092_));
 sg13g2_nand2_1 _08556_ (.Y(_01712_),
    .A(net2925),
    .B(net1605));
 sg13g2_nand2_1 _08557_ (.Y(_01713_),
    .A(net2829),
    .B(net1588));
 sg13g2_nand3_1 _08558_ (.B(_01712_),
    .C(_01713_),
    .A(_01691_),
    .Y(_00093_));
 sg13g2_nand2_1 _08559_ (.Y(_01714_),
    .A(net2829),
    .B(net1605));
 sg13g2_nand2_1 _08560_ (.Y(_01715_),
    .A(\am_sdr0.am0.multA[3] ),
    .B(net1588));
 sg13g2_nand3_1 _08561_ (.B(_01714_),
    .C(_01715_),
    .A(_01695_),
    .Y(_00094_));
 sg13g2_nand2_1 _08562_ (.Y(_01716_),
    .A(net2909),
    .B(net1605));
 sg13g2_nand2_1 _08563_ (.Y(_01717_),
    .A(net2905),
    .B(net1588));
 sg13g2_nand3_1 _08564_ (.B(_01716_),
    .C(_01717_),
    .A(_01699_),
    .Y(_00095_));
 sg13g2_nand2_1 _08565_ (.Y(_01718_),
    .A(net2905),
    .B(net1605));
 sg13g2_nand2_1 _08566_ (.Y(_01719_),
    .A(net2831),
    .B(net1588));
 sg13g2_nand3_1 _08567_ (.B(_01718_),
    .C(_01719_),
    .A(_01703_),
    .Y(_00096_));
 sg13g2_nand2_1 _08568_ (.Y(_01720_),
    .A(net2831),
    .B(net1605));
 sg13g2_nand2_1 _08569_ (.Y(_01721_),
    .A(\am_sdr0.am0.multA[6] ),
    .B(net1589));
 sg13g2_nand3_1 _08570_ (.B(_01720_),
    .C(_01721_),
    .A(_01707_),
    .Y(_00097_));
 sg13g2_nand2_1 _08571_ (.Y(_01722_),
    .A(\am_sdr0.am0.multA[6] ),
    .B(net1606));
 sg13g2_nand2_1 _08572_ (.Y(_01723_),
    .A(net2678),
    .B(net1589));
 sg13g2_nand3_1 _08573_ (.B(_01722_),
    .C(_01723_),
    .A(net1568),
    .Y(_00098_));
 sg13g2_nand2_1 _08574_ (.Y(_01724_),
    .A(net2678),
    .B(net1606));
 sg13g2_nand2_1 _08575_ (.Y(_01725_),
    .A(net2730),
    .B(net1589));
 sg13g2_nand3_1 _08576_ (.B(_01724_),
    .C(_01725_),
    .A(net1567),
    .Y(_00099_));
 sg13g2_a22oi_1 _08577_ (.Y(_01726_),
    .B1(net1606),
    .B2(net2730),
    .A2(net1589),
    .A1(net2819));
 sg13g2_nand2_1 _08578_ (.Y(_00100_),
    .A(net1567),
    .B(_01726_));
 sg13g2_a22oi_1 _08579_ (.Y(_01727_),
    .B1(net1607),
    .B2(net2819),
    .A2(net1590),
    .A1(\am_sdr0.am0.multA[10] ));
 sg13g2_nand2_1 _08580_ (.Y(_00101_),
    .A(net1568),
    .B(net2820));
 sg13g2_nand2_1 _08581_ (.Y(_01728_),
    .A(net2985),
    .B(net1606));
 sg13g2_nand2_1 _08582_ (.Y(_01729_),
    .A(\am_sdr0.am0.multA[11] ),
    .B(net1590));
 sg13g2_nand3_1 _08583_ (.B(_01728_),
    .C(_01729_),
    .A(net1567),
    .Y(_00102_));
 sg13g2_a22oi_1 _08584_ (.Y(_01730_),
    .B1(net1606),
    .B2(net3011),
    .A2(net1590),
    .A1(net2948));
 sg13g2_nand2_1 _08585_ (.Y(_00103_),
    .A(net1567),
    .B(_01730_));
 sg13g2_a22oi_1 _08586_ (.Y(_01731_),
    .B1(net1607),
    .B2(net2948),
    .A2(net1589),
    .A1(net2697));
 sg13g2_nand2_1 _08587_ (.Y(_00104_),
    .A(net1567),
    .B(_01731_));
 sg13g2_nand2_1 _08588_ (.Y(_01732_),
    .A(net2697),
    .B(net1606));
 sg13g2_nand2_1 _08589_ (.Y(_01733_),
    .A(\am_sdr0.am0.multA[14] ),
    .B(net1589));
 sg13g2_nand3_1 _08590_ (.B(_01732_),
    .C(_01733_),
    .A(net1567),
    .Y(_00105_));
 sg13g2_a22oi_1 _08591_ (.Y(_01734_),
    .B1(net1606),
    .B2(net2781),
    .A2(net1589),
    .A1(net2451));
 sg13g2_nand2_1 _08592_ (.Y(_00106_),
    .A(net1567),
    .B(_01734_));
 sg13g2_a22oi_1 _08593_ (.Y(_01735_),
    .B1(net1606),
    .B2(net2451),
    .A2(net1589),
    .A1(\am_sdr0.am0.multA[16] ));
 sg13g2_nand2_1 _08594_ (.Y(_00107_),
    .A(net1567),
    .B(net2452));
 sg13g2_nand3b_1 _08595_ (.B(\am_sdr0.am0.multB[0] ),
    .C(_01603_),
    .Y(_01736_),
    .A_N(_01668_));
 sg13g2_inv_1 _08596_ (.Y(_01737_),
    .A(_01736_));
 sg13g2_o21ai_1 _08597_ (.B1(_00016_),
    .Y(_01738_),
    .A1(\am_sdr0.am0.multB[0] ),
    .A2(_01668_));
 sg13g2_and2_1 _08598_ (.A(net1584),
    .B(_01738_),
    .X(_01739_));
 sg13g2_nand2_1 _08599_ (.Y(_01740_),
    .A(net1431),
    .B(net1565));
 sg13g2_nor2b_1 _08600_ (.A(net1431),
    .B_N(\am_sdr0.am0.multA[0] ),
    .Y(_01741_));
 sg13g2_inv_1 _08601_ (.Y(_01742_),
    .A(_01741_));
 sg13g2_xnor2_1 _08602_ (.Y(_01743_),
    .A(net1431),
    .B(\am_sdr0.am0.multA[0] ));
 sg13g2_o21ai_1 _08603_ (.B1(_01740_),
    .Y(_00108_),
    .A1(net1584),
    .A2(_01743_));
 sg13g2_xnor2_1 _08604_ (.Y(_01744_),
    .A(\am_sdr0.am0.multA[0] ),
    .B(\am_sdr0.am0.multA[1] ));
 sg13g2_nor3_1 _08605_ (.A(\am_sdr0.am0.m_count[3] ),
    .B(_00058_),
    .C(_01597_),
    .Y(_01745_));
 sg13g2_a21oi_1 _08606_ (.A1(_01566_),
    .A2(_01596_),
    .Y(_01746_),
    .B1(_01744_));
 sg13g2_nor3_1 _08607_ (.A(_01563_),
    .B(_01745_),
    .C(_01746_),
    .Y(_01747_));
 sg13g2_o21ai_1 _08608_ (.B1(_01563_),
    .Y(_01748_),
    .A1(_01745_),
    .A2(_01746_));
 sg13g2_nand2b_1 _08609_ (.Y(_01749_),
    .B(_01748_),
    .A_N(_01747_));
 sg13g2_o21ai_1 _08610_ (.B1(net1566),
    .Y(_01750_),
    .A1(_01741_),
    .A2(_01749_));
 sg13g2_a21oi_1 _08611_ (.A1(_01741_),
    .A2(_01749_),
    .Y(_01751_),
    .B1(_01750_));
 sg13g2_a21o_1 _08612_ (.A2(net1565),
    .A1(net2503),
    .B1(_01751_),
    .X(_00109_));
 sg13g2_a21o_1 _08613_ (.A2(_01748_),
    .A1(_01742_),
    .B1(_01747_),
    .X(_01752_));
 sg13g2_nor3_1 _08614_ (.A(\am_sdr0.am0.multA[0] ),
    .B(\am_sdr0.am0.multA[1] ),
    .C(\am_sdr0.am0.multA[2] ),
    .Y(_01753_));
 sg13g2_o21ai_1 _08615_ (.B1(\am_sdr0.am0.multA[2] ),
    .Y(_01754_),
    .A1(\am_sdr0.am0.multA[0] ),
    .A2(\am_sdr0.am0.multA[1] ));
 sg13g2_nand2b_1 _08616_ (.Y(_01755_),
    .B(_01754_),
    .A_N(_01753_));
 sg13g2_mux2_1 _08617_ (.A0(_00060_),
    .A1(_01755_),
    .S(net1608),
    .X(_01756_));
 sg13g2_xnor2_1 _08618_ (.Y(_01757_),
    .A(_00059_),
    .B(_01756_));
 sg13g2_o21ai_1 _08619_ (.B1(net1566),
    .Y(_01758_),
    .A1(_01752_),
    .A2(_01757_));
 sg13g2_a21oi_1 _08620_ (.A1(_01752_),
    .A2(_01757_),
    .Y(_01759_),
    .B1(_01758_));
 sg13g2_a21o_1 _08621_ (.A2(net1565),
    .A1(net2277),
    .B1(_01759_),
    .X(_00110_));
 sg13g2_and2_1 _08622_ (.A(\am_sdr0.am0.sum[2] ),
    .B(_01756_),
    .X(_01760_));
 sg13g2_a21o_1 _08623_ (.A2(_01757_),
    .A1(_01752_),
    .B1(_01760_),
    .X(_01761_));
 sg13g2_nand2_1 _08624_ (.Y(_01762_),
    .A(_00061_),
    .B(net1610));
 sg13g2_or4_2 _08625_ (.A(\am_sdr0.am0.multA[0] ),
    .B(\am_sdr0.am0.multA[1] ),
    .C(\am_sdr0.am0.multA[2] ),
    .D(\am_sdr0.am0.multA[3] ),
    .X(_01763_));
 sg13g2_xnor2_1 _08626_ (.Y(_01764_),
    .A(\am_sdr0.am0.multA[3] ),
    .B(_01753_));
 sg13g2_o21ai_1 _08627_ (.B1(_01762_),
    .Y(_01765_),
    .A1(net1610),
    .A2(_01764_));
 sg13g2_and2_1 _08628_ (.A(\am_sdr0.am0.sum[3] ),
    .B(_01765_),
    .X(_01766_));
 sg13g2_xor2_1 _08629_ (.B(_01765_),
    .A(\am_sdr0.am0.sum[3] ),
    .X(_01767_));
 sg13g2_o21ai_1 _08630_ (.B1(net1566),
    .Y(_01768_),
    .A1(_01761_),
    .A2(_01767_));
 sg13g2_a21oi_1 _08631_ (.A1(_01761_),
    .A2(_01767_),
    .Y(_01769_),
    .B1(_01768_));
 sg13g2_a21o_1 _08632_ (.A2(net1565),
    .A1(net2687),
    .B1(_01769_),
    .X(_00111_));
 sg13g2_a21oi_2 _08633_ (.B1(_01766_),
    .Y(_01770_),
    .A2(_01767_),
    .A1(_01761_));
 sg13g2_nand2_1 _08634_ (.Y(_01771_),
    .A(_00063_),
    .B(net1610));
 sg13g2_nor2_1 _08635_ (.A(\am_sdr0.am0.multA[4] ),
    .B(_01763_),
    .Y(_01772_));
 sg13g2_xor2_1 _08636_ (.B(_01763_),
    .A(\am_sdr0.am0.multA[4] ),
    .X(_01773_));
 sg13g2_o21ai_1 _08637_ (.B1(_01771_),
    .Y(_01774_),
    .A1(net1610),
    .A2(_01773_));
 sg13g2_xor2_1 _08638_ (.B(_01774_),
    .A(_00062_),
    .X(_01775_));
 sg13g2_or2_1 _08639_ (.X(_01776_),
    .B(_01775_),
    .A(_01770_));
 sg13g2_a21oi_1 _08640_ (.A1(_01770_),
    .A2(_01775_),
    .Y(_01777_),
    .B1(net1584));
 sg13g2_a22oi_1 _08641_ (.Y(_01778_),
    .B1(_01776_),
    .B2(_01777_),
    .A2(net1565),
    .A1(net2099));
 sg13g2_inv_1 _08642_ (.Y(_00112_),
    .A(net2100));
 sg13g2_nor2_1 _08643_ (.A(\am_sdr0.am0.multA[5] ),
    .B(net1608),
    .Y(_01779_));
 sg13g2_xnor2_1 _08644_ (.Y(_01780_),
    .A(_00064_),
    .B(_01772_));
 sg13g2_a21oi_1 _08645_ (.A1(net1608),
    .A2(_01780_),
    .Y(_01781_),
    .B1(_01779_));
 sg13g2_nor2b_1 _08646_ (.A(\am_sdr0.am0.sum[5] ),
    .B_N(_01781_),
    .Y(_01782_));
 sg13g2_nand2b_1 _08647_ (.Y(_01783_),
    .B(\am_sdr0.am0.sum[5] ),
    .A_N(_01781_));
 sg13g2_nand2b_1 _08648_ (.Y(_01784_),
    .B(_01783_),
    .A_N(_01782_));
 sg13g2_nand2_1 _08649_ (.Y(_01785_),
    .A(\am_sdr0.am0.sum[4] ),
    .B(_01774_));
 sg13g2_and2_1 _08650_ (.A(_01776_),
    .B(_01785_),
    .X(_01786_));
 sg13g2_o21ai_1 _08651_ (.B1(net1566),
    .Y(_01787_),
    .A1(_01784_),
    .A2(_01786_));
 sg13g2_a21oi_1 _08652_ (.A1(_01784_),
    .A2(_01786_),
    .Y(_01788_),
    .B1(_01787_));
 sg13g2_a21o_1 _08653_ (.A2(net1565),
    .A1(net2729),
    .B1(_01788_),
    .X(_00113_));
 sg13g2_nand2_1 _08654_ (.Y(_01789_),
    .A(_00065_),
    .B(net1610));
 sg13g2_or2_1 _08655_ (.X(_01790_),
    .B(\am_sdr0.am0.multA[5] ),
    .A(\am_sdr0.am0.multA[4] ));
 sg13g2_or2_1 _08656_ (.X(_01791_),
    .B(_01790_),
    .A(_01763_));
 sg13g2_nor3_1 _08657_ (.A(\am_sdr0.am0.multA[6] ),
    .B(_01763_),
    .C(_01790_),
    .Y(_01792_));
 sg13g2_xor2_1 _08658_ (.B(_01791_),
    .A(\am_sdr0.am0.multA[6] ),
    .X(_01793_));
 sg13g2_o21ai_1 _08659_ (.B1(_01789_),
    .Y(_01794_),
    .A1(net1610),
    .A2(_01793_));
 sg13g2_and2_1 _08660_ (.A(\am_sdr0.am0.sum[6] ),
    .B(_01794_),
    .X(_01795_));
 sg13g2_xor2_1 _08661_ (.B(_01794_),
    .A(\am_sdr0.am0.sum[6] ),
    .X(_01796_));
 sg13g2_nor3_2 _08662_ (.A(_01770_),
    .B(_01775_),
    .C(_01784_),
    .Y(_01797_));
 sg13g2_o21ai_1 _08663_ (.B1(_01783_),
    .Y(_01798_),
    .A1(_01782_),
    .A2(_01785_));
 sg13g2_nor2_1 _08664_ (.A(_01797_),
    .B(_01798_),
    .Y(_01799_));
 sg13g2_nor2b_1 _08665_ (.A(_01799_),
    .B_N(_01796_),
    .Y(_01800_));
 sg13g2_nor3_1 _08666_ (.A(_01796_),
    .B(_01797_),
    .C(_01798_),
    .Y(_01801_));
 sg13g2_nor3_1 _08667_ (.A(net1584),
    .B(_01800_),
    .C(_01801_),
    .Y(_01802_));
 sg13g2_a21o_1 _08668_ (.A2(net1565),
    .A1(net2740),
    .B1(_01802_),
    .X(_00114_));
 sg13g2_nand2b_1 _08669_ (.Y(_01803_),
    .B(net1609),
    .A_N(\am_sdr0.am0.multA[7] ));
 sg13g2_xor2_1 _08670_ (.B(_01792_),
    .A(_00066_),
    .X(_01804_));
 sg13g2_o21ai_1 _08671_ (.B1(_01803_),
    .Y(_01805_),
    .A1(net1609),
    .A2(_01804_));
 sg13g2_nand2_1 _08672_ (.Y(_01806_),
    .A(\am_sdr0.am0.sum[7] ),
    .B(_01805_));
 sg13g2_xor2_1 _08673_ (.B(_01805_),
    .A(\am_sdr0.am0.sum[7] ),
    .X(_01807_));
 sg13g2_or2_1 _08674_ (.X(_01808_),
    .B(_01800_),
    .A(_01795_));
 sg13g2_o21ai_1 _08675_ (.B1(net1566),
    .Y(_01809_),
    .A1(_01807_),
    .A2(_01808_));
 sg13g2_a21oi_1 _08676_ (.A1(_01807_),
    .A2(_01808_),
    .Y(_01810_),
    .B1(_01809_));
 sg13g2_a21o_1 _08677_ (.A2(net1565),
    .A1(net2835),
    .B1(_01810_),
    .X(_00115_));
 sg13g2_nand2_1 _08678_ (.Y(_01811_),
    .A(net2247),
    .B(net1564));
 sg13g2_or2_1 _08679_ (.X(_01812_),
    .B(\am_sdr0.am0.multA[7] ),
    .A(\am_sdr0.am0.multA[6] ));
 sg13g2_nor2_1 _08680_ (.A(_01791_),
    .B(_01812_),
    .Y(_01813_));
 sg13g2_nor4_2 _08681_ (.A(\am_sdr0.am0.multA[8] ),
    .B(_01763_),
    .C(_01790_),
    .Y(_01814_),
    .D(_01812_));
 sg13g2_nand2_1 _08682_ (.Y(_01815_),
    .A(_00067_),
    .B(net1609));
 sg13g2_xnor2_1 _08683_ (.Y(_01816_),
    .A(\am_sdr0.am0.multA[8] ),
    .B(_01813_));
 sg13g2_o21ai_1 _08684_ (.B1(_01815_),
    .Y(_01817_),
    .A1(net1609),
    .A2(_01816_));
 sg13g2_nand2_1 _08685_ (.Y(_01818_),
    .A(\am_sdr0.am0.sum[8] ),
    .B(_01817_));
 sg13g2_xnor2_1 _08686_ (.Y(_01819_),
    .A(\am_sdr0.am0.sum[8] ),
    .B(_01817_));
 sg13g2_o21ai_1 _08687_ (.B1(_01795_),
    .Y(_01820_),
    .A1(\am_sdr0.am0.sum[7] ),
    .A2(_01805_));
 sg13g2_nand3b_1 _08688_ (.B(_01806_),
    .C(_01820_),
    .Y(_01821_),
    .A_N(_01798_));
 sg13g2_nand2_1 _08689_ (.Y(_01822_),
    .A(_01796_),
    .B(_01807_));
 sg13g2_nand3_1 _08690_ (.B(_01820_),
    .C(_01822_),
    .A(_01806_),
    .Y(_01823_));
 sg13g2_o21ai_1 _08691_ (.B1(_01823_),
    .Y(_01824_),
    .A1(_01797_),
    .A2(_01821_));
 sg13g2_nor2_1 _08692_ (.A(_01819_),
    .B(_01824_),
    .Y(_01825_));
 sg13g2_a21o_1 _08693_ (.A2(_01824_),
    .A1(_01819_),
    .B1(_01736_),
    .X(_01826_));
 sg13g2_o21ai_1 _08694_ (.B1(_01811_),
    .Y(_00116_),
    .A1(_01825_),
    .A2(_01826_));
 sg13g2_o21ai_1 _08695_ (.B1(_01818_),
    .Y(_01827_),
    .A1(_01819_),
    .A2(_01824_));
 sg13g2_nand2b_2 _08696_ (.Y(_01828_),
    .B(_01814_),
    .A_N(\am_sdr0.am0.multA[9] ));
 sg13g2_nand2_1 _08697_ (.Y(_01829_),
    .A(_00068_),
    .B(net1609));
 sg13g2_xnor2_1 _08698_ (.Y(_01830_),
    .A(\am_sdr0.am0.multA[9] ),
    .B(_01814_));
 sg13g2_o21ai_1 _08699_ (.B1(_01829_),
    .Y(_01831_),
    .A1(net1609),
    .A2(_01830_));
 sg13g2_nand2_1 _08700_ (.Y(_01832_),
    .A(\am_sdr0.am0.sum[9] ),
    .B(_01831_));
 sg13g2_nor2_1 _08701_ (.A(\am_sdr0.am0.sum[9] ),
    .B(_01831_),
    .Y(_01833_));
 sg13g2_xnor2_1 _08702_ (.Y(_01834_),
    .A(\am_sdr0.am0.sum[9] ),
    .B(_01831_));
 sg13g2_nor2b_1 _08703_ (.A(_01827_),
    .B_N(_01834_),
    .Y(_01835_));
 sg13g2_nor2b_1 _08704_ (.A(_01834_),
    .B_N(_01827_),
    .Y(_01836_));
 sg13g2_nor3_1 _08705_ (.A(net1584),
    .B(_01835_),
    .C(_01836_),
    .Y(_01837_));
 sg13g2_a21o_1 _08706_ (.A2(net1564),
    .A1(net2955),
    .B1(_01837_),
    .X(_00117_));
 sg13g2_o21ai_1 _08707_ (.B1(_01832_),
    .Y(_01838_),
    .A1(_01818_),
    .A2(_01833_));
 sg13g2_inv_1 _08708_ (.Y(_01839_),
    .A(_01838_));
 sg13g2_nor2_1 _08709_ (.A(_01819_),
    .B(_01834_),
    .Y(_01840_));
 sg13g2_inv_1 _08710_ (.Y(_01841_),
    .A(_01840_));
 sg13g2_o21ai_1 _08711_ (.B1(_01839_),
    .Y(_01842_),
    .A1(_01824_),
    .A2(_01841_));
 sg13g2_xor2_1 _08712_ (.B(_01828_),
    .A(\am_sdr0.am0.multA[10] ),
    .X(_01843_));
 sg13g2_nand2_1 _08713_ (.Y(_01844_),
    .A(_00069_),
    .B(net1609));
 sg13g2_o21ai_1 _08714_ (.B1(_01844_),
    .Y(_01845_),
    .A1(net1611),
    .A2(_01843_));
 sg13g2_nand2_1 _08715_ (.Y(_01846_),
    .A(\am_sdr0.am0.sum[10] ),
    .B(_01845_));
 sg13g2_xor2_1 _08716_ (.B(_01845_),
    .A(\am_sdr0.am0.sum[10] ),
    .X(_01847_));
 sg13g2_xnor2_1 _08717_ (.Y(_01848_),
    .A(\am_sdr0.am0.sum[10] ),
    .B(_01845_));
 sg13g2_nand2_1 _08718_ (.Y(_01849_),
    .A(_01842_),
    .B(_01847_));
 sg13g2_nor2_1 _08719_ (.A(_01842_),
    .B(_01847_),
    .Y(_01850_));
 sg13g2_nor2_1 _08720_ (.A(net1584),
    .B(_01850_),
    .Y(_01851_));
 sg13g2_a22oi_1 _08721_ (.Y(_01852_),
    .B1(_01849_),
    .B2(_01851_),
    .A2(net1564),
    .A1(net2938));
 sg13g2_inv_1 _08722_ (.Y(_00118_),
    .A(_01852_));
 sg13g2_nand2_1 _08723_ (.Y(_01853_),
    .A(net2470),
    .B(net1564));
 sg13g2_o21ai_1 _08724_ (.B1(_01599_),
    .Y(_01854_),
    .A1(_01592_),
    .A2(_01828_));
 sg13g2_xor2_1 _08725_ (.B(_01854_),
    .A(\am_sdr0.am0.multA[11] ),
    .X(_01855_));
 sg13g2_nor2_1 _08726_ (.A(\am_sdr0.am0.sum[11] ),
    .B(_01855_),
    .Y(_01856_));
 sg13g2_xnor2_1 _08727_ (.Y(_01857_),
    .A(\am_sdr0.am0.sum[11] ),
    .B(_01855_));
 sg13g2_a21oi_1 _08728_ (.A1(_01846_),
    .A2(_01849_),
    .Y(_01858_),
    .B1(_01857_));
 sg13g2_nand3_1 _08729_ (.B(_01849_),
    .C(_01857_),
    .A(_01846_),
    .Y(_01859_));
 sg13g2_nand2_1 _08730_ (.Y(_01860_),
    .A(_01737_),
    .B(_01859_));
 sg13g2_o21ai_1 _08731_ (.B1(_01853_),
    .Y(_00119_),
    .A1(_01858_),
    .A2(_01860_));
 sg13g2_nand2_1 _08732_ (.Y(_01861_),
    .A(net1480),
    .B(_01739_));
 sg13g2_nor2_1 _08733_ (.A(_01848_),
    .B(_01857_),
    .Y(_01862_));
 sg13g2_nand2_1 _08734_ (.Y(_01863_),
    .A(_01840_),
    .B(_01862_));
 sg13g2_nor2_1 _08735_ (.A(_01846_),
    .B(_01856_),
    .Y(_01864_));
 sg13g2_a221oi_1 _08736_ (.B2(_01838_),
    .C1(_01864_),
    .B1(_01862_),
    .A1(\am_sdr0.am0.sum[11] ),
    .Y(_01865_),
    .A2(_01855_));
 sg13g2_o21ai_1 _08737_ (.B1(_01865_),
    .Y(_01866_),
    .A1(_01824_),
    .A2(_01863_));
 sg13g2_nor3_1 _08738_ (.A(\am_sdr0.am0.multA[10] ),
    .B(\am_sdr0.am0.multA[11] ),
    .C(_01828_),
    .Y(_01867_));
 sg13g2_nor2_1 _08739_ (.A(net1609),
    .B(_01867_),
    .Y(_01868_));
 sg13g2_xnor2_1 _08740_ (.Y(_01869_),
    .A(\am_sdr0.am0.multA[12] ),
    .B(_01868_));
 sg13g2_nand2_1 _08741_ (.Y(_01870_),
    .A(\am_sdr0.am0.sum[12] ),
    .B(_01869_));
 sg13g2_xor2_1 _08742_ (.B(_01869_),
    .A(net2702),
    .X(_01871_));
 sg13g2_inv_1 _08743_ (.Y(_01872_),
    .A(_01871_));
 sg13g2_and2_1 _08744_ (.A(_01866_),
    .B(_01871_),
    .X(_01873_));
 sg13g2_o21ai_1 _08745_ (.B1(net1566),
    .Y(_01874_),
    .A1(_01866_),
    .A2(_01871_));
 sg13g2_o21ai_1 _08746_ (.B1(_01861_),
    .Y(_00120_),
    .A1(_01873_),
    .A2(_01874_));
 sg13g2_nand2_1 _08747_ (.Y(_01875_),
    .A(net2618),
    .B(net1564));
 sg13g2_nor2_1 _08748_ (.A(_00070_),
    .B(_01599_),
    .Y(_01876_));
 sg13g2_nor4_2 _08749_ (.A(\am_sdr0.am0.multA[10] ),
    .B(\am_sdr0.am0.multA[11] ),
    .C(\am_sdr0.am0.multA[12] ),
    .Y(_01877_),
    .D(_01828_));
 sg13g2_nor2b_1 _08750_ (.A(\am_sdr0.am0.multA[13] ),
    .B_N(_01877_),
    .Y(_01878_));
 sg13g2_xnor2_1 _08751_ (.Y(_01879_),
    .A(\am_sdr0.am0.multA[13] ),
    .B(_01877_));
 sg13g2_a21oi_2 _08752_ (.B1(_01876_),
    .Y(_01880_),
    .A2(_01879_),
    .A1(net1608));
 sg13g2_nand2_1 _08753_ (.Y(_01881_),
    .A(\am_sdr0.am0.sum[13] ),
    .B(_01880_));
 sg13g2_nor2_1 _08754_ (.A(\am_sdr0.am0.sum[13] ),
    .B(_01880_),
    .Y(_01882_));
 sg13g2_xnor2_1 _08755_ (.Y(_01883_),
    .A(\am_sdr0.am0.sum[13] ),
    .B(_01880_));
 sg13g2_a21oi_1 _08756_ (.A1(net1480),
    .A2(_01869_),
    .Y(_01884_),
    .B1(_01873_));
 sg13g2_xnor2_1 _08757_ (.Y(_01885_),
    .A(_01883_),
    .B(_01884_));
 sg13g2_o21ai_1 _08758_ (.B1(_01875_),
    .Y(_00121_),
    .A1(net1584),
    .A2(_01885_));
 sg13g2_nor2_1 _08759_ (.A(_01872_),
    .B(_01883_),
    .Y(_01886_));
 sg13g2_o21ai_1 _08760_ (.B1(_01881_),
    .Y(_01887_),
    .A1(_01870_),
    .A2(_01882_));
 sg13g2_a21o_1 _08761_ (.A2(_01886_),
    .A1(_01866_),
    .B1(_01887_),
    .X(_01888_));
 sg13g2_nor2_1 _08762_ (.A(_00071_),
    .B(net1608),
    .Y(_01889_));
 sg13g2_nor2b_1 _08763_ (.A(\am_sdr0.am0.multA[14] ),
    .B_N(_01878_),
    .Y(_01890_));
 sg13g2_xnor2_1 _08764_ (.Y(_01891_),
    .A(\am_sdr0.am0.multA[14] ),
    .B(_01878_));
 sg13g2_a21oi_2 _08765_ (.B1(_01889_),
    .Y(_01892_),
    .A2(_01891_),
    .A1(net1608));
 sg13g2_nand2_1 _08766_ (.Y(_01893_),
    .A(\am_sdr0.am0.sum[14] ),
    .B(_01892_));
 sg13g2_inv_1 _08767_ (.Y(_01894_),
    .A(_01893_));
 sg13g2_xnor2_1 _08768_ (.Y(_01895_),
    .A(\am_sdr0.am0.sum[14] ),
    .B(_01892_));
 sg13g2_inv_1 _08769_ (.Y(_01896_),
    .A(_01895_));
 sg13g2_nand2b_1 _08770_ (.Y(_01897_),
    .B(_01895_),
    .A_N(_01888_));
 sg13g2_a21oi_1 _08771_ (.A1(_01888_),
    .A2(_01896_),
    .Y(_01898_),
    .B1(net1584));
 sg13g2_a22oi_1 _08772_ (.Y(_01899_),
    .B1(_01897_),
    .B2(_01898_),
    .A2(net1564),
    .A1(net2767));
 sg13g2_inv_1 _08773_ (.Y(_00122_),
    .A(_01899_));
 sg13g2_nand2_1 _08774_ (.Y(_01900_),
    .A(net2032),
    .B(net1564));
 sg13g2_nand2b_1 _08775_ (.Y(_01901_),
    .B(\am_sdr0.am0.multA[15] ),
    .A_N(_01890_));
 sg13g2_a21oi_1 _08776_ (.A1(_01580_),
    .A2(_01890_),
    .Y(_01902_),
    .B1(net1611));
 sg13g2_a22oi_1 _08777_ (.Y(_01903_),
    .B1(_01901_),
    .B2(_01902_),
    .A2(net1611),
    .A1(_01593_));
 sg13g2_nor2_1 _08778_ (.A(\am_sdr0.am0.sum[15] ),
    .B(_01903_),
    .Y(_01904_));
 sg13g2_xnor2_1 _08779_ (.Y(_01905_),
    .A(\am_sdr0.am0.sum[15] ),
    .B(_01903_));
 sg13g2_a21oi_1 _08780_ (.A1(_01888_),
    .A2(_01896_),
    .Y(_01906_),
    .B1(_01894_));
 sg13g2_and2_1 _08781_ (.A(_01905_),
    .B(_01906_),
    .X(_01907_));
 sg13g2_o21ai_1 _08782_ (.B1(net1566),
    .Y(_01908_),
    .A1(_01905_),
    .A2(_01906_));
 sg13g2_o21ai_1 _08783_ (.B1(_01900_),
    .Y(_00123_),
    .A1(_01907_),
    .A2(_01908_));
 sg13g2_nand2_1 _08784_ (.Y(_01909_),
    .A(net2209),
    .B(net1564));
 sg13g2_nor2_1 _08785_ (.A(_01895_),
    .B(_01905_),
    .Y(_01910_));
 sg13g2_nor2_1 _08786_ (.A(_01893_),
    .B(_01904_),
    .Y(_01911_));
 sg13g2_a221oi_1 _08787_ (.B2(_01888_),
    .C1(_01911_),
    .B1(_01910_),
    .A1(\am_sdr0.am0.sum[15] ),
    .Y(_01912_),
    .A2(_01903_));
 sg13g2_xnor2_1 _08788_ (.Y(_01913_),
    .A(\am_sdr0.am0.sum[16] ),
    .B(\am_sdr0.am0.multA[16] ));
 sg13g2_xnor2_1 _08789_ (.Y(_01914_),
    .A(_01902_),
    .B(_01913_));
 sg13g2_and2_1 _08790_ (.A(_01912_),
    .B(_01914_),
    .X(_01915_));
 sg13g2_o21ai_1 _08791_ (.B1(net1566),
    .Y(_01916_),
    .A1(_01912_),
    .A2(_01914_));
 sg13g2_o21ai_1 _08792_ (.B1(_01909_),
    .Y(_00124_),
    .A1(_01915_),
    .A2(_01916_));
 sg13g2_nor2_1 _08793_ (.A(net2118),
    .B(net1893),
    .Y(_01917_));
 sg13g2_nor2_1 _08794_ (.A(_01562_),
    .B(\am_sdr0.am0.sqrt_state[0] ),
    .Y(_01918_));
 sg13g2_nand2b_2 _08795_ (.Y(_01919_),
    .B(\am_sdr0.am0.sqrt_state[1] ),
    .A_N(\am_sdr0.am0.sqrt_state[0] ));
 sg13g2_a21oi_2 _08796_ (.B1(net1893),
    .Y(_01920_),
    .A2(\am_sdr0.am0.sqrt_state[0] ),
    .A1(\am_sdr0.am0.sqrt_state[1] ));
 sg13g2_nor2_1 _08797_ (.A(\am_sdr0.am0.sqrt_state[1] ),
    .B(\am_sdr0.am0.sqrt_state[0] ),
    .Y(_01921_));
 sg13g2_nand2b_2 _08798_ (.Y(_01922_),
    .B(_01920_),
    .A_N(_01921_));
 sg13g2_inv_1 _08799_ (.Y(_00173_),
    .A(_01922_));
 sg13g2_a21oi_2 _08800_ (.B1(net1618),
    .Y(_01923_),
    .A2(net1256),
    .A1(_01564_));
 sg13g2_nor2_1 _08801_ (.A(_01922_),
    .B(_01923_),
    .Y(_01924_));
 sg13g2_nand2b_1 _08802_ (.Y(_01925_),
    .B(_00173_),
    .A_N(_01923_));
 sg13g2_nand3_1 _08803_ (.B(net1602),
    .C(net1583),
    .A(net1170),
    .Y(_01926_));
 sg13g2_o21ai_1 _08804_ (.B1(_01926_),
    .Y(_00125_),
    .A1(_01570_),
    .A2(net1583));
 sg13g2_nand3_1 _08805_ (.B(\am_sdr0.am0.count2[0] ),
    .C(net1583),
    .A(net3004),
    .Y(_01927_));
 sg13g2_a21oi_1 _08806_ (.A1(\am_sdr0.am0.count2[0] ),
    .A2(net1583),
    .Y(_01928_),
    .B1(net3004));
 sg13g2_nor2_2 _08807_ (.A(net1602),
    .B(_01922_),
    .Y(_01929_));
 sg13g2_nor2_1 _08808_ (.A(net3005),
    .B(_01929_),
    .Y(_01930_));
 sg13g2_and2_1 _08809_ (.A(_01927_),
    .B(_01930_),
    .X(_00126_));
 sg13g2_nand3_1 _08810_ (.B(\am_sdr0.am0.count2[0] ),
    .C(net1254),
    .A(\am_sdr0.am0.count2[1] ),
    .Y(_01931_));
 sg13g2_a21oi_1 _08811_ (.A1(net1602),
    .A2(_01931_),
    .Y(_01932_),
    .B1(_01925_));
 sg13g2_a21oi_1 _08812_ (.A1(_01572_),
    .A2(_01927_),
    .Y(_00127_),
    .B1(_01932_));
 sg13g2_or4_1 _08813_ (.A(net2097),
    .B(net1618),
    .C(_01925_),
    .D(_01931_),
    .X(_01933_));
 sg13g2_o21ai_1 _08814_ (.B1(_01933_),
    .Y(_00128_),
    .A1(_01571_),
    .A2(_01932_));
 sg13g2_nor2_1 _08815_ (.A(_01564_),
    .B(net1256),
    .Y(_01934_));
 sg13g2_o21ai_1 _08816_ (.B1(_00173_),
    .Y(_01935_),
    .A1(net1619),
    .A2(_01934_));
 sg13g2_nand2_1 _08817_ (.Y(_01936_),
    .A(net1212),
    .B(_01935_));
 sg13g2_nand3_1 _08818_ (.B(net1602),
    .C(net1257),
    .A(net2015),
    .Y(_01937_));
 sg13g2_nand2_1 _08819_ (.Y(_01938_),
    .A(net1233),
    .B(\am_sdr0.am0.right[0] ));
 sg13g2_xnor2_1 _08820_ (.Y(_01939_),
    .A(net1233),
    .B(\am_sdr0.am0.right[0] ));
 sg13g2_o21ai_1 _08821_ (.B1(_01936_),
    .Y(_00129_),
    .A1(net1580),
    .A2(net1234));
 sg13g2_nand2_1 _08822_ (.Y(_01940_),
    .A(net1217),
    .B(net1563));
 sg13g2_nor2_1 _08823_ (.A(\am_sdr0.am0.right[0] ),
    .B(\am_sdr0.am0.right[1] ),
    .Y(_01941_));
 sg13g2_nor2_1 _08824_ (.A(net1872),
    .B(_01941_),
    .Y(_01942_));
 sg13g2_and2_1 _08825_ (.A(\am_sdr0.am0.right[0] ),
    .B(\am_sdr0.am0.right[1] ),
    .X(_01943_));
 sg13g2_nor3_1 _08826_ (.A(net1872),
    .B(_01941_),
    .C(_01943_),
    .Y(_01944_));
 sg13g2_nor2b_1 _08827_ (.A(_00047_),
    .B_N(net1872),
    .Y(_01945_));
 sg13g2_o21ai_1 _08828_ (.B1(\am_sdr0.am0.left[1] ),
    .Y(_01946_),
    .A1(_01944_),
    .A2(_01945_));
 sg13g2_nor3_1 _08829_ (.A(\am_sdr0.am0.left[1] ),
    .B(_01944_),
    .C(_01945_),
    .Y(_01947_));
 sg13g2_or3_1 _08830_ (.A(\am_sdr0.am0.left[1] ),
    .B(_01944_),
    .C(_01945_),
    .X(_01948_));
 sg13g2_nand2_1 _08831_ (.Y(_01949_),
    .A(_01946_),
    .B(_01948_));
 sg13g2_a21oi_1 _08832_ (.A1(_01938_),
    .A2(_01949_),
    .Y(_01950_),
    .B1(_01937_));
 sg13g2_o21ai_1 _08833_ (.B1(_01950_),
    .Y(_01951_),
    .A1(_01938_),
    .A2(_01949_));
 sg13g2_nand2_1 _08834_ (.Y(_00130_),
    .A(_01940_),
    .B(_01951_));
 sg13g2_nand2_1 _08835_ (.Y(_01952_),
    .A(net1210),
    .B(net1563));
 sg13g2_o21ai_1 _08836_ (.B1(_01946_),
    .Y(_01953_),
    .A1(_01938_),
    .A2(_01947_));
 sg13g2_xnor2_1 _08837_ (.Y(_01954_),
    .A(_00048_),
    .B(_01942_));
 sg13g2_and2_1 _08838_ (.A(\am_sdr0.am0.left[2] ),
    .B(_01954_),
    .X(_01955_));
 sg13g2_xor2_1 _08839_ (.B(_01954_),
    .A(\am_sdr0.am0.left[2] ),
    .X(_01956_));
 sg13g2_a21oi_1 _08840_ (.A1(_01953_),
    .A2(_01956_),
    .Y(_01957_),
    .B1(net1580));
 sg13g2_o21ai_1 _08841_ (.B1(_01957_),
    .Y(_01958_),
    .A1(_01953_),
    .A2(_01956_));
 sg13g2_nand2_1 _08842_ (.Y(_00131_),
    .A(_01952_),
    .B(_01958_));
 sg13g2_a21oi_1 _08843_ (.A1(_01953_),
    .A2(_01956_),
    .Y(_01959_),
    .B1(_01955_));
 sg13g2_nand2b_1 _08844_ (.Y(_01960_),
    .B(net1872),
    .A_N(_00049_));
 sg13g2_nand2_1 _08845_ (.Y(_01961_),
    .A(_00048_),
    .B(_01941_));
 sg13g2_xnor2_1 _08846_ (.Y(_01962_),
    .A(\am_sdr0.am0.right[3] ),
    .B(_01961_));
 sg13g2_o21ai_1 _08847_ (.B1(_01960_),
    .Y(_01963_),
    .A1(net1872),
    .A2(_01962_));
 sg13g2_nand2_1 _08848_ (.Y(_01964_),
    .A(\am_sdr0.am0.left[3] ),
    .B(_01963_));
 sg13g2_xnor2_1 _08849_ (.Y(_01965_),
    .A(\am_sdr0.am0.left[3] ),
    .B(_01963_));
 sg13g2_nor2_1 _08850_ (.A(_01959_),
    .B(_01965_),
    .Y(_01966_));
 sg13g2_and2_1 _08851_ (.A(_01959_),
    .B(_01965_),
    .X(_01967_));
 sg13g2_nor3_1 _08852_ (.A(net1580),
    .B(_01966_),
    .C(_01967_),
    .Y(_01968_));
 sg13g2_a21o_1 _08853_ (.A2(net1563),
    .A1(net1222),
    .B1(_01968_),
    .X(_00132_));
 sg13g2_o21ai_1 _08854_ (.B1(_01964_),
    .Y(_01969_),
    .A1(_01959_),
    .A2(_01965_));
 sg13g2_nor4_2 _08855_ (.A(\am_sdr0.am0.right[0] ),
    .B(\am_sdr0.am0.right[1] ),
    .C(\am_sdr0.am0.right[2] ),
    .Y(_01970_),
    .D(\am_sdr0.am0.right[3] ));
 sg13g2_nor2_1 _08856_ (.A(\am_sdr0.am0.r[9] ),
    .B(_01970_),
    .Y(_01971_));
 sg13g2_xnor2_1 _08857_ (.Y(_01972_),
    .A(_00050_),
    .B(_01971_));
 sg13g2_nand2_1 _08858_ (.Y(_01973_),
    .A(\am_sdr0.am0.left[4] ),
    .B(_01972_));
 sg13g2_inv_1 _08859_ (.Y(_01974_),
    .A(_01973_));
 sg13g2_xor2_1 _08860_ (.B(_01972_),
    .A(\am_sdr0.am0.left[4] ),
    .X(_01975_));
 sg13g2_nand2_1 _08861_ (.Y(_01976_),
    .A(_01969_),
    .B(_01975_));
 sg13g2_nor2_1 _08862_ (.A(_01969_),
    .B(_01975_),
    .Y(_01977_));
 sg13g2_nor2_1 _08863_ (.A(net1580),
    .B(_01977_),
    .Y(_01978_));
 sg13g2_a22oi_1 _08864_ (.Y(_01979_),
    .B1(_01976_),
    .B2(_01978_),
    .A2(net1563),
    .A1(net1224));
 sg13g2_inv_1 _08865_ (.Y(_00133_),
    .A(_01979_));
 sg13g2_a21oi_1 _08866_ (.A1(_01969_),
    .A2(_01975_),
    .Y(_01980_),
    .B1(_01974_));
 sg13g2_nand2_1 _08867_ (.Y(_01981_),
    .A(_00050_),
    .B(_01970_));
 sg13g2_xor2_1 _08868_ (.B(_01981_),
    .A(\am_sdr0.am0.right[5] ),
    .X(_01982_));
 sg13g2_nand2_1 _08869_ (.Y(_01983_),
    .A(net1872),
    .B(_00052_));
 sg13g2_o21ai_1 _08870_ (.B1(_01983_),
    .Y(_01984_),
    .A1(net1871),
    .A2(_01982_));
 sg13g2_xnor2_1 _08871_ (.Y(_01985_),
    .A(net1336),
    .B(_01984_));
 sg13g2_nor2_1 _08872_ (.A(_01980_),
    .B(_01985_),
    .Y(_01986_));
 sg13g2_nand2_1 _08873_ (.Y(_01987_),
    .A(_01980_),
    .B(_01985_));
 sg13g2_nor2_1 _08874_ (.A(net1580),
    .B(_01986_),
    .Y(_01988_));
 sg13g2_a22oi_1 _08875_ (.Y(_01989_),
    .B1(_01987_),
    .B2(_01988_),
    .A2(net1563),
    .A1(net1313));
 sg13g2_inv_1 _08876_ (.Y(_00134_),
    .A(_01989_));
 sg13g2_nand2b_1 _08877_ (.Y(_01990_),
    .B(\am_sdr0.am0.left[5] ),
    .A_N(_01984_));
 sg13g2_o21ai_1 _08878_ (.B1(_01990_),
    .Y(_01991_),
    .A1(_01980_),
    .A2(_01985_));
 sg13g2_nor2_1 _08879_ (.A(\am_sdr0.am0.right[4] ),
    .B(\am_sdr0.am0.right[5] ),
    .Y(_01992_));
 sg13g2_and2_1 _08880_ (.A(_01970_),
    .B(_01992_),
    .X(_01993_));
 sg13g2_nor2_1 _08881_ (.A(net1871),
    .B(_01993_),
    .Y(_01994_));
 sg13g2_xnor2_1 _08882_ (.Y(_01995_),
    .A(_00053_),
    .B(_01994_));
 sg13g2_nand2_1 _08883_ (.Y(_01996_),
    .A(net1392),
    .B(_01995_));
 sg13g2_xor2_1 _08884_ (.B(_01995_),
    .A(\am_sdr0.am0.left[6] ),
    .X(_01997_));
 sg13g2_nand2_1 _08885_ (.Y(_01998_),
    .A(_01991_),
    .B(_01997_));
 sg13g2_nor2_1 _08886_ (.A(_01991_),
    .B(_01997_),
    .Y(_01999_));
 sg13g2_nor2_1 _08887_ (.A(net1580),
    .B(_01999_),
    .Y(_02000_));
 sg13g2_a22oi_1 _08888_ (.Y(_02001_),
    .B1(_01998_),
    .B2(_02000_),
    .A2(net1563),
    .A1(net1200));
 sg13g2_inv_1 _08889_ (.Y(_00135_),
    .A(_02001_));
 sg13g2_nand2b_1 _08890_ (.Y(_02002_),
    .B(net1871),
    .A_N(_00054_));
 sg13g2_nand2_1 _08891_ (.Y(_02003_),
    .A(_00053_),
    .B(_01993_));
 sg13g2_xnor2_1 _08892_ (.Y(_02004_),
    .A(\am_sdr0.am0.right[7] ),
    .B(_02003_));
 sg13g2_o21ai_1 _08893_ (.B1(_02002_),
    .Y(_02005_),
    .A1(net1871),
    .A2(_02004_));
 sg13g2_nand2_1 _08894_ (.Y(_02006_),
    .A(\am_sdr0.am0.left[7] ),
    .B(_02005_));
 sg13g2_xnor2_1 _08895_ (.Y(_02007_),
    .A(\am_sdr0.am0.left[7] ),
    .B(_02005_));
 sg13g2_a21oi_1 _08896_ (.A1(_01996_),
    .A2(_01998_),
    .Y(_02008_),
    .B1(_02007_));
 sg13g2_nand3_1 _08897_ (.B(_01998_),
    .C(_02007_),
    .A(_01996_),
    .Y(_02009_));
 sg13g2_nor2_1 _08898_ (.A(net1580),
    .B(_02008_),
    .Y(_02010_));
 sg13g2_a22oi_1 _08899_ (.Y(_02011_),
    .B1(_02009_),
    .B2(_02010_),
    .A2(net1563),
    .A1(net1352));
 sg13g2_inv_1 _08900_ (.Y(_00136_),
    .A(_02011_));
 sg13g2_nand2_1 _08901_ (.Y(_02012_),
    .A(net1871),
    .B(net1563));
 sg13g2_nor2_1 _08902_ (.A(\am_sdr0.am0.right[6] ),
    .B(\am_sdr0.am0.right[7] ),
    .Y(_02013_));
 sg13g2_and2_1 _08903_ (.A(_01993_),
    .B(_02013_),
    .X(_02014_));
 sg13g2_nor2b_1 _08904_ (.A(\am_sdr0.am0.right[8] ),
    .B_N(_02014_),
    .Y(_02015_));
 sg13g2_xnor2_1 _08905_ (.Y(_02016_),
    .A(\am_sdr0.am0.right[8] ),
    .B(_02014_));
 sg13g2_nand2_1 _08906_ (.Y(_02017_),
    .A(net1871),
    .B(_00057_));
 sg13g2_o21ai_1 _08907_ (.B1(_02017_),
    .Y(_02018_),
    .A1(net1871),
    .A2(_02016_));
 sg13g2_nand2_1 _08908_ (.Y(_02019_),
    .A(net3270),
    .B(_02018_));
 sg13g2_o21ai_1 _08909_ (.B1(_02006_),
    .Y(_02020_),
    .A1(_00056_),
    .A2(_02018_));
 sg13g2_o21ai_1 _08910_ (.B1(_02019_),
    .Y(_02021_),
    .A1(_02008_),
    .A2(_02020_));
 sg13g2_xor2_1 _08911_ (.B(_02015_),
    .A(\am_sdr0.am0.right[9] ),
    .X(_02022_));
 sg13g2_mux2_1 _08912_ (.A0(_02022_),
    .A1(_00055_),
    .S(net1871),
    .X(_02023_));
 sg13g2_xnor2_1 _08913_ (.Y(_02024_),
    .A(\am_sdr0.am0.left[9] ),
    .B(_02023_));
 sg13g2_inv_1 _08914_ (.Y(_02025_),
    .A(_02024_));
 sg13g2_nor2_1 _08915_ (.A(_02021_),
    .B(_02025_),
    .Y(_02026_));
 sg13g2_a21o_1 _08916_ (.A2(_02025_),
    .A1(_02021_),
    .B1(net1580),
    .X(_02027_));
 sg13g2_o21ai_1 _08917_ (.B1(_02012_),
    .Y(_00137_),
    .A1(net3271),
    .A2(_02027_));
 sg13g2_nand2_1 _08918_ (.Y(_02028_),
    .A(_01564_),
    .B(_01573_));
 sg13g2_a21o_1 _08919_ (.A2(_02028_),
    .A1(net1602),
    .B1(_01922_),
    .X(_02029_));
 sg13g2_a21oi_2 _08920_ (.B1(_01922_),
    .Y(_02030_),
    .A2(_02028_),
    .A1(net1600));
 sg13g2_a22oi_1 _08921_ (.Y(_02031_),
    .B1(net1579),
    .B2(net1248),
    .A2(_01929_),
    .A1(\am_sdr0.am0.sum[1] ));
 sg13g2_inv_1 _08922_ (.Y(_00138_),
    .A(net1249));
 sg13g2_a22oi_1 _08923_ (.Y(_02032_),
    .B1(net1579),
    .B2(net1239),
    .A2(_01929_),
    .A1(\am_sdr0.am0.sum[2] ));
 sg13g2_inv_1 _08924_ (.Y(_00139_),
    .A(net1240));
 sg13g2_and2_1 _08925_ (.A(\am_sdr0.am0.sum[3] ),
    .B(net1618),
    .X(_02033_));
 sg13g2_a21oi_1 _08926_ (.A1(net1248),
    .A2(net1600),
    .Y(_02034_),
    .B1(_02033_));
 sg13g2_nor2_1 _08927_ (.A(net1386),
    .B(net1572),
    .Y(_02035_));
 sg13g2_a21oi_1 _08928_ (.A1(net1572),
    .A2(_02034_),
    .Y(_00140_),
    .B1(_02035_));
 sg13g2_and2_1 _08929_ (.A(\am_sdr0.am0.sum[4] ),
    .B(net1618),
    .X(_02036_));
 sg13g2_a21oi_1 _08930_ (.A1(net1239),
    .A2(net1600),
    .Y(_02037_),
    .B1(_02036_));
 sg13g2_nor2_1 _08931_ (.A(net1458),
    .B(net1572),
    .Y(_02038_));
 sg13g2_a21oi_1 _08932_ (.A1(net1572),
    .A2(_02037_),
    .Y(_00141_),
    .B1(_02038_));
 sg13g2_and2_1 _08933_ (.A(\am_sdr0.am0.sum[5] ),
    .B(net1618),
    .X(_02039_));
 sg13g2_a21oi_1 _08934_ (.A1(net1386),
    .A2(net1600),
    .Y(_02040_),
    .B1(_02039_));
 sg13g2_nor2_1 _08935_ (.A(net2027),
    .B(net1572),
    .Y(_02041_));
 sg13g2_a21oi_1 _08936_ (.A1(net1572),
    .A2(_02040_),
    .Y(_00142_),
    .B1(_02041_));
 sg13g2_and2_1 _08937_ (.A(\am_sdr0.am0.sum[6] ),
    .B(net1618),
    .X(_02042_));
 sg13g2_a21oi_1 _08938_ (.A1(\am_sdr0.am0.a[3] ),
    .A2(net1600),
    .Y(_02043_),
    .B1(_02042_));
 sg13g2_nor2_1 _08939_ (.A(net1456),
    .B(net1573),
    .Y(_02044_));
 sg13g2_a21oi_1 _08940_ (.A1(net1572),
    .A2(_02043_),
    .Y(_00143_),
    .B1(_02044_));
 sg13g2_and2_1 _08941_ (.A(\am_sdr0.am0.sum[7] ),
    .B(net1619),
    .X(_02045_));
 sg13g2_a21oi_1 _08942_ (.A1(\am_sdr0.am0.a[4] ),
    .A2(net1600),
    .Y(_02046_),
    .B1(_02045_));
 sg13g2_nor2_1 _08943_ (.A(net1508),
    .B(net1573),
    .Y(_02047_));
 sg13g2_a21oi_1 _08944_ (.A1(net1572),
    .A2(_02046_),
    .Y(_00144_),
    .B1(_02047_));
 sg13g2_and2_1 _08945_ (.A(\am_sdr0.am0.sum[8] ),
    .B(net1619),
    .X(_02048_));
 sg13g2_a21oi_1 _08946_ (.A1(net1456),
    .A2(net1600),
    .Y(_02049_),
    .B1(_02048_));
 sg13g2_nor2_1 _08947_ (.A(net1491),
    .B(net1576),
    .Y(_02050_));
 sg13g2_a21oi_1 _08948_ (.A1(net1576),
    .A2(_02049_),
    .Y(_00145_),
    .B1(_02050_));
 sg13g2_and2_1 _08949_ (.A(\am_sdr0.am0.sum[9] ),
    .B(net1618),
    .X(_02051_));
 sg13g2_a21oi_1 _08950_ (.A1(\am_sdr0.am0.a[6] ),
    .A2(net1600),
    .Y(_02052_),
    .B1(_02051_));
 sg13g2_nor2_1 _08951_ (.A(net1413),
    .B(net1573),
    .Y(_02053_));
 sg13g2_a21oi_1 _08952_ (.A1(net1573),
    .A2(_02052_),
    .Y(_00146_),
    .B1(_02053_));
 sg13g2_and2_1 _08953_ (.A(\am_sdr0.am0.sum[10] ),
    .B(net1619),
    .X(_02054_));
 sg13g2_a21oi_1 _08954_ (.A1(\am_sdr0.am0.a[7] ),
    .A2(net1601),
    .Y(_02055_),
    .B1(_02054_));
 sg13g2_nor2_1 _08955_ (.A(net1448),
    .B(net1575),
    .Y(_02056_));
 sg13g2_a21oi_1 _08956_ (.A1(net1575),
    .A2(_02055_),
    .Y(_00147_),
    .B1(_02056_));
 sg13g2_and2_1 _08957_ (.A(\am_sdr0.am0.sum[11] ),
    .B(net1619),
    .X(_02057_));
 sg13g2_a21oi_1 _08958_ (.A1(\am_sdr0.am0.a[8] ),
    .A2(net1601),
    .Y(_02058_),
    .B1(_02057_));
 sg13g2_nor2_1 _08959_ (.A(net1317),
    .B(net1576),
    .Y(_02059_));
 sg13g2_a21oi_1 _08960_ (.A1(net1576),
    .A2(_02058_),
    .Y(_00148_),
    .B1(_02059_));
 sg13g2_and2_1 _08961_ (.A(net1480),
    .B(net1619),
    .X(_02060_));
 sg13g2_a21oi_1 _08962_ (.A1(net1448),
    .A2(net1601),
    .Y(_02061_),
    .B1(_02060_));
 sg13g2_nor2_1 _08963_ (.A(net1468),
    .B(net1574),
    .Y(_02062_));
 sg13g2_a21oi_1 _08964_ (.A1(net1574),
    .A2(_02061_),
    .Y(_00149_),
    .B1(_02062_));
 sg13g2_and2_1 _08965_ (.A(\am_sdr0.am0.sum[13] ),
    .B(net1619),
    .X(_02063_));
 sg13g2_a21oi_1 _08966_ (.A1(net1317),
    .A2(net1601),
    .Y(_02064_),
    .B1(_02063_));
 sg13g2_nor2_1 _08967_ (.A(net1358),
    .B(net1575),
    .Y(_02065_));
 sg13g2_a21oi_1 _08968_ (.A1(net1574),
    .A2(_02064_),
    .Y(_00150_),
    .B1(_02065_));
 sg13g2_and2_1 _08969_ (.A(\am_sdr0.am0.sum[14] ),
    .B(_01919_),
    .X(_02066_));
 sg13g2_a21oi_1 _08970_ (.A1(net1468),
    .A2(net1601),
    .Y(_02067_),
    .B1(_02066_));
 sg13g2_nor2_1 _08971_ (.A(net1377),
    .B(net1575),
    .Y(_02068_));
 sg13g2_a21oi_1 _08972_ (.A1(net1574),
    .A2(net1469),
    .Y(_00151_),
    .B1(_02068_));
 sg13g2_and2_1 _08973_ (.A(net2032),
    .B(_01919_),
    .X(_02069_));
 sg13g2_a21oi_1 _08974_ (.A1(net1358),
    .A2(net1601),
    .Y(_02070_),
    .B1(_02069_));
 sg13g2_nor2_1 _08975_ (.A(net1308),
    .B(net1574),
    .Y(_02071_));
 sg13g2_a21oi_1 _08976_ (.A1(net1574),
    .A2(_02070_),
    .Y(_00152_),
    .B1(_02071_));
 sg13g2_and2_1 _08977_ (.A(\am_sdr0.am0.sum[16] ),
    .B(_01919_),
    .X(_02072_));
 sg13g2_a21oi_1 _08978_ (.A1(net1377),
    .A2(net1601),
    .Y(_02073_),
    .B1(_02072_));
 sg13g2_nor2_1 _08979_ (.A(net1304),
    .B(net1574),
    .Y(_02074_));
 sg13g2_a21oi_1 _08980_ (.A1(net1574),
    .A2(net1378),
    .Y(_00153_),
    .B1(_02074_));
 sg13g2_nor2_1 _08981_ (.A(_01579_),
    .B(_01666_),
    .Y(_00154_));
 sg13g2_and2_1 _08982_ (.A(net1951),
    .B(net1179),
    .X(_00155_));
 sg13g2_and2_1 _08983_ (.A(net2013),
    .B(net1165),
    .X(_00156_));
 sg13g2_o21ai_1 _08984_ (.B1(net2013),
    .Y(_02075_),
    .A1(\am_sdr0.count[1] ),
    .A2(net2433));
 sg13g2_a21oi_1 _08985_ (.A1(\am_sdr0.count[1] ),
    .A2(net2433),
    .Y(_00157_),
    .B1(_02075_));
 sg13g2_a21oi_1 _08986_ (.A1(\am_sdr0.count[1] ),
    .A2(net2433),
    .Y(_02076_),
    .B1(net2526));
 sg13g2_nand3_1 _08987_ (.B(\am_sdr0.count[1] ),
    .C(net3226),
    .A(net2526),
    .Y(_02077_));
 sg13g2_nand2_1 _08988_ (.Y(_02078_),
    .A(net2013),
    .B(_02077_));
 sg13g2_nor2_1 _08989_ (.A(net2527),
    .B(_02078_),
    .Y(_00158_));
 sg13g2_and2_1 _08990_ (.A(_01586_),
    .B(_02077_),
    .X(_02079_));
 sg13g2_nor2_1 _08991_ (.A(_01586_),
    .B(_02077_),
    .Y(_02080_));
 sg13g2_nor3_1 _08992_ (.A(net1894),
    .B(_02079_),
    .C(_02080_),
    .Y(_00159_));
 sg13g2_nor3_2 _08993_ (.A(_01585_),
    .B(_01586_),
    .C(_02077_),
    .Y(_02081_));
 sg13g2_o21ai_1 _08994_ (.B1(net2014),
    .Y(_02082_),
    .A1(net3092),
    .A2(_02080_));
 sg13g2_nor2_1 _08995_ (.A(_02081_),
    .B(_02082_),
    .Y(_00160_));
 sg13g2_xnor2_1 _08996_ (.Y(_02083_),
    .A(net3074),
    .B(_02081_));
 sg13g2_nor2_1 _08997_ (.A(net1894),
    .B(_02083_),
    .Y(_00161_));
 sg13g2_a21oi_1 _08998_ (.A1(net3074),
    .A2(_02081_),
    .Y(_02084_),
    .B1(net1870));
 sg13g2_nand3_1 _08999_ (.B(net3074),
    .C(_02081_),
    .A(net1870),
    .Y(_02085_));
 sg13g2_nand2_1 _09000_ (.Y(_02086_),
    .A(net2014),
    .B(_02085_));
 sg13g2_nor2_1 _09001_ (.A(net3075),
    .B(_02086_),
    .Y(_00162_));
 sg13g2_o21ai_1 _09002_ (.B1(net2014),
    .Y(_02087_),
    .A1(net1621),
    .A2(_02085_));
 sg13g2_a21oi_1 _09003_ (.A1(net1621),
    .A2(_02085_),
    .Y(_00163_),
    .B1(_02087_));
 sg13g2_nand3_1 _09004_ (.B(net1603),
    .C(net1583),
    .A(net1172),
    .Y(_02088_));
 sg13g2_o21ai_1 _09005_ (.B1(_02088_),
    .Y(_00164_),
    .A1(_01190_),
    .A2(net1583));
 sg13g2_nand3_1 _09006_ (.B(net1603),
    .C(net1581),
    .A(net2301),
    .Y(_02089_));
 sg13g2_o21ai_1 _09007_ (.B1(_02089_),
    .Y(_00165_),
    .A1(_01189_),
    .A2(net1581));
 sg13g2_nand3_1 _09008_ (.B(net1603),
    .C(net1581),
    .A(net2139),
    .Y(_02090_));
 sg13g2_o21ai_1 _09009_ (.B1(_02090_),
    .Y(_00166_),
    .A1(_01187_),
    .A2(net1581));
 sg13g2_nand3_1 _09010_ (.B(net1603),
    .C(net1581),
    .A(net2127),
    .Y(_02091_));
 sg13g2_o21ai_1 _09011_ (.B1(_02091_),
    .Y(_00167_),
    .A1(_01185_),
    .A2(net1581));
 sg13g2_nand3_1 _09012_ (.B(net1603),
    .C(net1582),
    .A(net1522),
    .Y(_02092_));
 sg13g2_o21ai_1 _09013_ (.B1(_02092_),
    .Y(_00168_),
    .A1(_01183_),
    .A2(net1582));
 sg13g2_nand3_1 _09014_ (.B(net1603),
    .C(net1582),
    .A(net2168),
    .Y(_02093_));
 sg13g2_o21ai_1 _09015_ (.B1(_02093_),
    .Y(_00169_),
    .A1(_01181_),
    .A2(net1582));
 sg13g2_nand3_1 _09016_ (.B(net1603),
    .C(net1582),
    .A(net1488),
    .Y(_02094_));
 sg13g2_o21ai_1 _09017_ (.B1(_02094_),
    .Y(_00170_),
    .A1(_01179_),
    .A2(net1581));
 sg13g2_nand3_1 _09018_ (.B(net1603),
    .C(net1582),
    .A(net1435),
    .Y(_02095_));
 sg13g2_o21ai_1 _09019_ (.B1(_02095_),
    .Y(_00171_),
    .A1(_01177_),
    .A2(net1581));
 sg13g2_o21ai_1 _09020_ (.B1(\am_sdr0.am0.sqrt_state[1] ),
    .Y(_02096_),
    .A1(net2097),
    .A2(_01931_));
 sg13g2_inv_1 _09021_ (.Y(_02097_),
    .A(_02096_));
 sg13g2_o21ai_1 _09022_ (.B1(_01917_),
    .Y(_02098_),
    .A1(\am_sdr0.am0.sqrt_state[1] ),
    .A2(net1260));
 sg13g2_nor3_1 _09023_ (.A(_01923_),
    .B(_02097_),
    .C(_02098_),
    .Y(_00172_));
 sg13g2_and3_2 _09024_ (.X(_02099_),
    .A(\am_sdr0.am0.sqrt_state[1] ),
    .B(\am_sdr0.am0.sqrt_state[0] ),
    .C(net2025));
 sg13g2_nor2_1 _09025_ (.A(net1471),
    .B(_02099_),
    .Y(_02100_));
 sg13g2_a21oi_1 _09026_ (.A1(_01562_),
    .A2(_01917_),
    .Y(_00174_),
    .B1(net1472));
 sg13g2_nor3_1 _09027_ (.A(net1893),
    .B(net1618),
    .C(_02028_),
    .Y(_02101_));
 sg13g2_a22oi_1 _09028_ (.Y(_02102_),
    .B1(net1571),
    .B2(net1308),
    .A2(net1579),
    .A1(net1233));
 sg13g2_inv_1 _09029_ (.Y(_00175_),
    .A(_02102_));
 sg13g2_a22oi_1 _09030_ (.Y(_02103_),
    .B1(net1570),
    .B2(net1304),
    .A2(net1579),
    .A1(\am_sdr0.am0.left[1] ));
 sg13g2_inv_1 _09031_ (.Y(_00176_),
    .A(net1305));
 sg13g2_a22oi_1 _09032_ (.Y(_02104_),
    .B1(net1570),
    .B2(net1212),
    .A2(_02029_),
    .A1(\am_sdr0.am0.left[2] ));
 sg13g2_inv_1 _09033_ (.Y(_00177_),
    .A(net1213));
 sg13g2_a22oi_1 _09034_ (.Y(_02105_),
    .B1(net1570),
    .B2(net1217),
    .A2(net1579),
    .A1(\am_sdr0.am0.left[3] ));
 sg13g2_inv_1 _09035_ (.Y(_00178_),
    .A(net1218));
 sg13g2_a22oi_1 _09036_ (.Y(_02106_),
    .B1(net1570),
    .B2(net1210),
    .A2(net1579),
    .A1(\am_sdr0.am0.left[4] ));
 sg13g2_inv_1 _09037_ (.Y(_00179_),
    .A(net1211));
 sg13g2_a22oi_1 _09038_ (.Y(_02107_),
    .B1(net1571),
    .B2(net1222),
    .A2(net1578),
    .A1(\am_sdr0.am0.left[5] ));
 sg13g2_inv_1 _09039_ (.Y(_00180_),
    .A(net1223));
 sg13g2_a22oi_1 _09040_ (.Y(_02108_),
    .B1(net1570),
    .B2(net1224),
    .A2(net1577),
    .A1(\am_sdr0.am0.left[6] ));
 sg13g2_inv_1 _09041_ (.Y(_00181_),
    .A(net1225));
 sg13g2_a22oi_1 _09042_ (.Y(_02109_),
    .B1(net1571),
    .B2(net1313),
    .A2(net1578),
    .A1(\am_sdr0.am0.left[7] ));
 sg13g2_inv_1 _09043_ (.Y(_00182_),
    .A(net1314));
 sg13g2_a22oi_1 _09044_ (.Y(_02110_),
    .B1(net1569),
    .B2(net1200),
    .A2(net1577),
    .A1(\am_sdr0.am0.left[8] ));
 sg13g2_inv_1 _09045_ (.Y(_00183_),
    .A(net1201));
 sg13g2_a22oi_1 _09046_ (.Y(_02111_),
    .B1(net1569),
    .B2(net1352),
    .A2(net1577),
    .A1(\am_sdr0.am0.left[9] ));
 sg13g2_inv_1 _09047_ (.Y(_00184_),
    .A(net1353));
 sg13g2_a21o_1 _09048_ (.A2(net1579),
    .A1(net3029),
    .B1(net1570),
    .X(_00185_));
 sg13g2_a22oi_1 _09049_ (.Y(_02112_),
    .B1(net1570),
    .B2(net1872),
    .A2(net1579),
    .A1(net2317));
 sg13g2_inv_1 _09050_ (.Y(_00186_),
    .A(net2318));
 sg13g2_a22oi_1 _09051_ (.Y(_02113_),
    .B1(net1570),
    .B2(\am_sdr0.am0.q[0] ),
    .A2(net1578),
    .A1(net1474));
 sg13g2_inv_1 _09052_ (.Y(_00187_),
    .A(net1475));
 sg13g2_a22oi_1 _09053_ (.Y(_02114_),
    .B1(net1571),
    .B2(net2139),
    .A2(net1578),
    .A1(\am_sdr0.am0.right[3] ));
 sg13g2_inv_1 _09054_ (.Y(_00188_),
    .A(net2140));
 sg13g2_a22oi_1 _09055_ (.Y(_02115_),
    .B1(net1569),
    .B2(\am_sdr0.am0.q[2] ),
    .A2(net1578),
    .A1(net1395));
 sg13g2_inv_1 _09056_ (.Y(_00189_),
    .A(net1396));
 sg13g2_a22oi_1 _09057_ (.Y(_02116_),
    .B1(net1569),
    .B2(net1522),
    .A2(net1577),
    .A1(net1524));
 sg13g2_inv_1 _09058_ (.Y(_00190_),
    .A(_02116_));
 sg13g2_a22oi_1 _09059_ (.Y(_02117_),
    .B1(net1569),
    .B2(\am_sdr0.am0.q[4] ),
    .A2(net1577),
    .A1(net1364));
 sg13g2_inv_1 _09060_ (.Y(_00191_),
    .A(net1365));
 sg13g2_a22oi_1 _09061_ (.Y(_02118_),
    .B1(net1569),
    .B2(net1488),
    .A2(net1577),
    .A1(\am_sdr0.am0.right[7] ));
 sg13g2_inv_1 _09062_ (.Y(_00192_),
    .A(net1489));
 sg13g2_a22oi_1 _09063_ (.Y(_02119_),
    .B1(net1569),
    .B2(net1435),
    .A2(net1577),
    .A1(\am_sdr0.am0.right[8] ));
 sg13g2_inv_1 _09064_ (.Y(_00193_),
    .A(net1436));
 sg13g2_a22oi_1 _09065_ (.Y(_02120_),
    .B1(net1569),
    .B2(net1323),
    .A2(net1577),
    .A1(\am_sdr0.am0.right[9] ));
 sg13g2_inv_1 _09066_ (.Y(_00194_),
    .A(net1324));
 sg13g2_nand3_1 _09067_ (.B(net1243),
    .C(net1490),
    .A(net1738),
    .Y(_02121_));
 sg13g2_nor2_1 _09068_ (.A(_01479_),
    .B(_02121_),
    .Y(_02122_));
 sg13g2_and2_1 _09069_ (.A(net2591),
    .B(_02122_),
    .X(_02123_));
 sg13g2_and2_1 _09070_ (.A(net2601),
    .B(_02123_),
    .X(_02124_));
 sg13g2_nand2_1 _09071_ (.Y(_02125_),
    .A(net2861),
    .B(_02124_));
 sg13g2_nor3_2 _09072_ (.A(net1375),
    .B(net2094),
    .C(_02125_),
    .Y(_02126_));
 sg13g2_nand2_1 _09073_ (.Y(_02127_),
    .A(net1983),
    .B(_02126_));
 sg13g2_inv_1 _09074_ (.Y(_00195_),
    .A(net1532));
 sg13g2_nand3_1 _09075_ (.B(net1228),
    .C(net1397),
    .A(net1670),
    .Y(_02128_));
 sg13g2_nor2_1 _09076_ (.A(_01393_),
    .B(_02128_),
    .Y(_02129_));
 sg13g2_and2_1 _09077_ (.A(net2548),
    .B(_02129_),
    .X(_02130_));
 sg13g2_and2_1 _09078_ (.A(net2619),
    .B(_02130_),
    .X(_02131_));
 sg13g2_nand2_1 _09079_ (.Y(_02132_),
    .A(net2851),
    .B(_02131_));
 sg13g2_nor4_1 _09080_ (.A(net1328),
    .B(net2063),
    .C(net1888),
    .D(_02132_),
    .Y(_00409_));
 sg13g2_nor3_1 _09081_ (.A(net1328),
    .B(net2063),
    .C(_02132_),
    .Y(_02133_));
 sg13g2_and2_2 _09082_ (.A(net1963),
    .B(_02133_),
    .X(_02134_));
 sg13g2_mux2_1 _09083_ (.A0(net2422),
    .A1(net1464),
    .S(net1538),
    .X(_00196_));
 sg13g2_mux2_1 _09084_ (.A0(net2453),
    .A1(net2629),
    .S(net1538),
    .X(_00197_));
 sg13g2_mux2_1 _09085_ (.A0(net2599),
    .A1(net2604),
    .S(net1539),
    .X(_00198_));
 sg13g2_nor2_1 _09086_ (.A(net2137),
    .B(net1539),
    .Y(_02135_));
 sg13g2_a21oi_1 _09087_ (.A1(_01386_),
    .A2(_02134_),
    .Y(_00199_),
    .B1(_02135_));
 sg13g2_mux2_1 _09088_ (.A0(net2447),
    .A1(\am_sdr0.cic2.integ3[4] ),
    .S(net1539),
    .X(_00200_));
 sg13g2_nor2_1 _09089_ (.A(\am_sdr0.cic2.integ_sample[5] ),
    .B(net1539),
    .Y(_02136_));
 sg13g2_a21oi_1 _09090_ (.A1(_01385_),
    .A2(_02134_),
    .Y(_00201_),
    .B1(_02136_));
 sg13g2_mux2_1 _09091_ (.A0(net2374),
    .A1(net2704),
    .S(net1537),
    .X(_00202_));
 sg13g2_mux2_1 _09092_ (.A0(net2396),
    .A1(net2620),
    .S(net1537),
    .X(_00203_));
 sg13g2_mux2_1 _09093_ (.A0(net2151),
    .A1(net2338),
    .S(net1537),
    .X(_00204_));
 sg13g2_mux2_1 _09094_ (.A0(net2361),
    .A1(net2658),
    .S(net1537),
    .X(_00205_));
 sg13g2_mux2_1 _09095_ (.A0(net2077),
    .A1(net2519),
    .S(net1537),
    .X(_00206_));
 sg13g2_mux2_1 _09096_ (.A0(net2066),
    .A1(net2274),
    .S(net1537),
    .X(_00207_));
 sg13g2_mux2_1 _09097_ (.A0(net2356),
    .A1(\am_sdr0.cic2.integ3[12] ),
    .S(net1537),
    .X(_00208_));
 sg13g2_mux2_1 _09098_ (.A0(net2849),
    .A1(\am_sdr0.cic2.integ3[13] ),
    .S(net1537),
    .X(_00209_));
 sg13g2_mux2_1 _09099_ (.A0(net1384),
    .A1(\am_sdr0.cic2.integ3[14] ),
    .S(net1538),
    .X(_00210_));
 sg13g2_mux2_1 _09100_ (.A0(net2226),
    .A1(\am_sdr0.cic2.integ3[15] ),
    .S(net1538),
    .X(_00211_));
 sg13g2_mux2_1 _09101_ (.A0(net2296),
    .A1(\am_sdr0.cic2.integ3[16] ),
    .S(net1538),
    .X(_00212_));
 sg13g2_mux2_1 _09102_ (.A0(net2234),
    .A1(\am_sdr0.cic2.integ3[17] ),
    .S(net1538),
    .X(_00213_));
 sg13g2_mux2_1 _09103_ (.A0(net2342),
    .A1(\am_sdr0.cic2.integ3[18] ),
    .S(net1538),
    .X(_00214_));
 sg13g2_mux2_1 _09104_ (.A0(net1486),
    .A1(net2305),
    .S(net1538),
    .X(_00215_));
 sg13g2_o21ai_1 _09105_ (.B1(net2022),
    .Y(_02137_),
    .A1(net1864),
    .A2(\am_sdr0.am0.Q_in[0] ));
 sg13g2_a21oi_1 _09106_ (.A1(net1864),
    .A2(_01514_),
    .Y(_00216_),
    .B1(_02137_));
 sg13g2_o21ai_1 _09107_ (.B1(net2023),
    .Y(_02138_),
    .A1(net1864),
    .A2(\am_sdr0.am0.Q_in[1] ));
 sg13g2_a21oi_1 _09108_ (.A1(net1864),
    .A2(_01513_),
    .Y(_00217_),
    .B1(_02138_));
 sg13g2_o21ai_1 _09109_ (.B1(net2023),
    .Y(_02139_),
    .A1(net1867),
    .A2(\am_sdr0.am0.Q_in[2] ));
 sg13g2_a21oi_1 _09110_ (.A1(net1866),
    .A2(_01512_),
    .Y(_00218_),
    .B1(_02139_));
 sg13g2_o21ai_1 _09111_ (.B1(net2023),
    .Y(_02140_),
    .A1(net1867),
    .A2(\am_sdr0.am0.Q_in[3] ));
 sg13g2_a21oi_1 _09112_ (.A1(net1867),
    .A2(_01511_),
    .Y(_00219_),
    .B1(_02140_));
 sg13g2_o21ai_1 _09113_ (.B1(net2022),
    .Y(_02141_),
    .A1(net1864),
    .A2(\am_sdr0.am0.Q_in[4] ));
 sg13g2_a21oi_1 _09114_ (.A1(net1864),
    .A2(_01510_),
    .Y(_00220_),
    .B1(_02141_));
 sg13g2_o21ai_1 _09115_ (.B1(net2022),
    .Y(_02142_),
    .A1(net1858),
    .A2(\am_sdr0.am0.Q_in[5] ));
 sg13g2_a21oi_1 _09116_ (.A1(net1858),
    .A2(_01509_),
    .Y(_00221_),
    .B1(_02142_));
 sg13g2_o21ai_1 _09117_ (.B1(net2022),
    .Y(_02143_),
    .A1(net1858),
    .A2(\am_sdr0.am0.Q_in[6] ));
 sg13g2_a21oi_1 _09118_ (.A1(net1858),
    .A2(_01508_),
    .Y(_00222_),
    .B1(_02143_));
 sg13g2_o21ai_1 _09119_ (.B1(net2017),
    .Y(_02144_),
    .A1(net1857),
    .A2(\am_sdr0.am0.Q_in[7] ));
 sg13g2_a21oi_1 _09120_ (.A1(net1857),
    .A2(_01507_),
    .Y(_00223_),
    .B1(_02144_));
 sg13g2_nand2b_1 _09121_ (.Y(_02145_),
    .B(net2413),
    .A_N(net2262));
 sg13g2_a21oi_1 _09122_ (.A1(_01560_),
    .A2(net2262),
    .Y(_02146_),
    .B1(net1622));
 sg13g2_a221oi_1 _09123_ (.B2(_02146_),
    .C1(net1890),
    .B1(_02145_),
    .A1(net1622),
    .Y(_00224_),
    .A2(_01537_));
 sg13g2_nor2b_1 _09124_ (.A(net2372),
    .B_N(\am_sdr0.cic3.integ_sample[1] ),
    .Y(_02147_));
 sg13g2_xnor2_1 _09125_ (.Y(_02148_),
    .A(net2372),
    .B(net2349));
 sg13g2_xnor2_1 _09126_ (.Y(_02149_),
    .A(_02145_),
    .B(_02148_));
 sg13g2_o21ai_1 _09127_ (.B1(net1985),
    .Y(_02150_),
    .A1(net1836),
    .A2(net2347));
 sg13g2_a21oi_1 _09128_ (.A1(net1836),
    .A2(_02149_),
    .Y(_00225_),
    .B1(_02150_));
 sg13g2_nand2b_1 _09129_ (.Y(_02151_),
    .B(\am_sdr0.cic3.integ_sample[2] ),
    .A_N(\am_sdr0.cic3.comb1_in_del[2] ));
 sg13g2_xor2_1 _09130_ (.B(net2483),
    .A(net2602),
    .X(_02152_));
 sg13g2_a21oi_1 _09131_ (.A1(_02145_),
    .A2(_02148_),
    .Y(_02153_),
    .B1(_02147_));
 sg13g2_xnor2_1 _09132_ (.Y(_02154_),
    .A(_02152_),
    .B(_02153_));
 sg13g2_o21ai_1 _09133_ (.B1(net1985),
    .Y(_02155_),
    .A1(net1836),
    .A2(net2238));
 sg13g2_a21oi_1 _09134_ (.A1(net1836),
    .A2(_02154_),
    .Y(_00226_),
    .B1(_02155_));
 sg13g2_nor2_1 _09135_ (.A(net2506),
    .B(_01557_),
    .Y(_02156_));
 sg13g2_nand2_1 _09136_ (.Y(_02157_),
    .A(net2833),
    .B(_01557_));
 sg13g2_nand2b_1 _09137_ (.Y(_02158_),
    .B(_02157_),
    .A_N(_02156_));
 sg13g2_o21ai_1 _09138_ (.B1(_02151_),
    .Y(_02159_),
    .A1(_02152_),
    .A2(_02153_));
 sg13g2_xnor2_1 _09139_ (.Y(_02160_),
    .A(_02158_),
    .B(_02159_));
 sg13g2_o21ai_1 _09140_ (.B1(net1985),
    .Y(_02161_),
    .A1(net1622),
    .A2(_02160_));
 sg13g2_a21oi_1 _09141_ (.A1(net1622),
    .A2(_01533_),
    .Y(_00227_),
    .B1(_02161_));
 sg13g2_nor2_1 _09142_ (.A(\am_sdr0.cic3.comb1_in_del[4] ),
    .B(_01556_),
    .Y(_02162_));
 sg13g2_xor2_1 _09143_ (.B(net2513),
    .A(net2735),
    .X(_02163_));
 sg13g2_a21oi_1 _09144_ (.A1(_02157_),
    .A2(_02159_),
    .Y(_02164_),
    .B1(_02156_));
 sg13g2_or2_1 _09145_ (.X(_02165_),
    .B(_02164_),
    .A(_02163_));
 sg13g2_xnor2_1 _09146_ (.Y(_02166_),
    .A(_02163_),
    .B(_02164_));
 sg13g2_o21ai_1 _09147_ (.B1(net1985),
    .Y(_02167_),
    .A1(net1842),
    .A2(net2595));
 sg13g2_a21oi_1 _09148_ (.A1(net1838),
    .A2(_02166_),
    .Y(_00228_),
    .B1(_02167_));
 sg13g2_xor2_1 _09149_ (.B(net2891),
    .A(\am_sdr0.cic3.comb1_in_del[5] ),
    .X(_02168_));
 sg13g2_nor2b_1 _09150_ (.A(_02162_),
    .B_N(_02165_),
    .Y(_02169_));
 sg13g2_xnor2_1 _09151_ (.Y(_02170_),
    .A(_02168_),
    .B(_02169_));
 sg13g2_o21ai_1 _09152_ (.B1(net1985),
    .Y(_02171_),
    .A1(net1838),
    .A2(net2449));
 sg13g2_a21oi_1 _09153_ (.A1(net1842),
    .A2(net2892),
    .Y(_00229_),
    .B1(_02171_));
 sg13g2_nor2_1 _09154_ (.A(\am_sdr0.cic3.comb1_in_del[6] ),
    .B(_01553_),
    .Y(_02172_));
 sg13g2_xor2_1 _09155_ (.B(net2587),
    .A(net2635),
    .X(_02173_));
 sg13g2_a21oi_1 _09156_ (.A1(_01554_),
    .A2(\am_sdr0.cic3.integ_sample[5] ),
    .Y(_02174_),
    .B1(_02162_));
 sg13g2_a22oi_1 _09157_ (.Y(_02175_),
    .B1(_02165_),
    .B2(_02174_),
    .A2(_01555_),
    .A1(\am_sdr0.cic3.comb1_in_del[5] ));
 sg13g2_a221oi_1 _09158_ (.B2(_02174_),
    .C1(_02173_),
    .B1(_02165_),
    .A1(\am_sdr0.cic3.comb1_in_del[5] ),
    .Y(_02176_),
    .A2(_01555_));
 sg13g2_xor2_1 _09159_ (.B(_02175_),
    .A(_02173_),
    .X(_02177_));
 sg13g2_o21ai_1 _09160_ (.B1(net1991),
    .Y(_02178_),
    .A1(net1838),
    .A2(net2724));
 sg13g2_a21oi_1 _09161_ (.A1(net1838),
    .A2(_02177_),
    .Y(_00230_),
    .B1(_02178_));
 sg13g2_nand2b_1 _09162_ (.Y(_02179_),
    .B(\am_sdr0.cic3.integ_sample[7] ),
    .A_N(\am_sdr0.cic3.comb1_in_del[7] ));
 sg13g2_xnor2_1 _09163_ (.Y(_02180_),
    .A(\am_sdr0.cic3.comb1_in_del[7] ),
    .B(\am_sdr0.cic3.integ_sample[7] ));
 sg13g2_o21ai_1 _09164_ (.B1(_02180_),
    .Y(_02181_),
    .A1(_02172_),
    .A2(_02176_));
 sg13g2_or3_1 _09165_ (.A(_02172_),
    .B(_02176_),
    .C(_02180_),
    .X(_02182_));
 sg13g2_and2_1 _09166_ (.A(_02181_),
    .B(_02182_),
    .X(_02183_));
 sg13g2_o21ai_1 _09167_ (.B1(net1991),
    .Y(_02184_),
    .A1(net1624),
    .A2(_02183_));
 sg13g2_a21oi_1 _09168_ (.A1(net1624),
    .A2(_01528_),
    .Y(_00231_),
    .B1(_02184_));
 sg13g2_nand2_1 _09169_ (.Y(_02185_),
    .A(_02179_),
    .B(_02181_));
 sg13g2_nor2_1 _09170_ (.A(\am_sdr0.cic3.comb1_in_del[8] ),
    .B(_01551_),
    .Y(_02186_));
 sg13g2_xnor2_1 _09171_ (.Y(_02187_),
    .A(\am_sdr0.cic3.comb1_in_del[8] ),
    .B(net2504));
 sg13g2_inv_1 _09172_ (.Y(_02188_),
    .A(_02187_));
 sg13g2_xnor2_1 _09173_ (.Y(_02189_),
    .A(_02185_),
    .B(_02187_));
 sg13g2_o21ai_1 _09174_ (.B1(net1991),
    .Y(_02190_),
    .A1(net1845),
    .A2(net2727));
 sg13g2_a21oi_1 _09175_ (.A1(net1845),
    .A2(_02189_),
    .Y(_00232_),
    .B1(_02190_));
 sg13g2_xor2_1 _09176_ (.B(\am_sdr0.cic3.integ_sample[9] ),
    .A(net2889),
    .X(_02191_));
 sg13g2_a21oi_1 _09177_ (.A1(_02185_),
    .A2(_02187_),
    .Y(_02192_),
    .B1(_02186_));
 sg13g2_xnor2_1 _09178_ (.Y(_02193_),
    .A(net2890),
    .B(_02192_));
 sg13g2_o21ai_1 _09179_ (.B1(net1991),
    .Y(_02194_),
    .A1(net1843),
    .A2(net2776));
 sg13g2_a21oi_1 _09180_ (.A1(net1843),
    .A2(_02193_),
    .Y(_00233_),
    .B1(_02194_));
 sg13g2_nand2b_1 _09181_ (.Y(_02195_),
    .B(\am_sdr0.cic3.integ_sample[10] ),
    .A_N(\am_sdr0.cic3.comb1_in_del[10] ));
 sg13g2_xor2_1 _09182_ (.B(\am_sdr0.cic3.integ_sample[10] ),
    .A(\am_sdr0.cic3.comb1_in_del[10] ),
    .X(_02196_));
 sg13g2_a21oi_1 _09183_ (.A1(_01549_),
    .A2(\am_sdr0.cic3.integ_sample[9] ),
    .Y(_02197_),
    .B1(_02186_));
 sg13g2_a21oi_1 _09184_ (.A1(\am_sdr0.cic3.comb1_in_del[9] ),
    .A2(_01550_),
    .Y(_02198_),
    .B1(_02197_));
 sg13g2_nor2_1 _09185_ (.A(_02188_),
    .B(_02191_),
    .Y(_02199_));
 sg13g2_a21oi_1 _09186_ (.A1(_02185_),
    .A2(_02199_),
    .Y(_02200_),
    .B1(_02198_));
 sg13g2_xnor2_1 _09187_ (.Y(_02201_),
    .A(_02196_),
    .B(_02200_));
 sg13g2_o21ai_1 _09188_ (.B1(net1997),
    .Y(_02202_),
    .A1(net1843),
    .A2(net2379));
 sg13g2_a21oi_1 _09189_ (.A1(net1843),
    .A2(_02201_),
    .Y(_00234_),
    .B1(_02202_));
 sg13g2_nor2b_1 _09190_ (.A(\am_sdr0.cic3.integ_sample[11] ),
    .B_N(\am_sdr0.cic3.comb1_in_del[11] ),
    .Y(_02203_));
 sg13g2_nand2b_1 _09191_ (.Y(_02204_),
    .B(\am_sdr0.cic3.integ_sample[11] ),
    .A_N(\am_sdr0.cic3.comb1_in_del[11] ));
 sg13g2_nand2b_1 _09192_ (.Y(_02205_),
    .B(_02204_),
    .A_N(_02203_));
 sg13g2_o21ai_1 _09193_ (.B1(_02195_),
    .Y(_02206_),
    .A1(_02196_),
    .A2(_02200_));
 sg13g2_xor2_1 _09194_ (.B(_02206_),
    .A(_02205_),
    .X(_02207_));
 sg13g2_o21ai_1 _09195_ (.B1(net1997),
    .Y(_02208_),
    .A1(net1843),
    .A2(net2236));
 sg13g2_a21oi_1 _09196_ (.A1(net1843),
    .A2(_02207_),
    .Y(_00235_),
    .B1(_02208_));
 sg13g2_nor2_1 _09197_ (.A(\am_sdr0.cic3.comb1_in_del[12] ),
    .B(_01546_),
    .Y(_02209_));
 sg13g2_xor2_1 _09198_ (.B(\am_sdr0.cic3.integ_sample[12] ),
    .A(\am_sdr0.cic3.comb1_in_del[12] ),
    .X(_02210_));
 sg13g2_inv_1 _09199_ (.Y(_02211_),
    .A(_02210_));
 sg13g2_nor2_1 _09200_ (.A(_02196_),
    .B(_02205_),
    .Y(_02212_));
 sg13g2_o21ai_1 _09201_ (.B1(_02204_),
    .Y(_02213_),
    .A1(_02195_),
    .A2(_02203_));
 sg13g2_a21o_1 _09202_ (.A2(_02212_),
    .A1(_02198_),
    .B1(_02213_),
    .X(_02214_));
 sg13g2_nand2_1 _09203_ (.Y(_02215_),
    .A(_02199_),
    .B(_02212_));
 sg13g2_a21oi_2 _09204_ (.B1(_02215_),
    .Y(_02216_),
    .A2(_02181_),
    .A1(_02179_));
 sg13g2_o21ai_1 _09205_ (.B1(_02211_),
    .Y(_02217_),
    .A1(_02214_),
    .A2(_02216_));
 sg13g2_or3_1 _09206_ (.A(_02211_),
    .B(_02214_),
    .C(_02216_),
    .X(_02218_));
 sg13g2_nand2_1 _09207_ (.Y(_02219_),
    .A(_02217_),
    .B(_02218_));
 sg13g2_o21ai_1 _09208_ (.B1(net1997),
    .Y(_02220_),
    .A1(net1860),
    .A2(net2522));
 sg13g2_a21oi_1 _09209_ (.A1(net1860),
    .A2(_02219_),
    .Y(_00236_),
    .B1(_02220_));
 sg13g2_nor2b_1 _09210_ (.A(\am_sdr0.cic3.integ_sample[13] ),
    .B_N(\am_sdr0.cic3.comb1_in_del[13] ),
    .Y(_02221_));
 sg13g2_nor2_1 _09211_ (.A(\am_sdr0.cic3.comb1_in_del[13] ),
    .B(_01545_),
    .Y(_02222_));
 sg13g2_nor2_1 _09212_ (.A(_02221_),
    .B(_02222_),
    .Y(_02223_));
 sg13g2_nand2b_1 _09213_ (.Y(_02224_),
    .B(_02217_),
    .A_N(_02209_));
 sg13g2_xnor2_1 _09214_ (.Y(_02225_),
    .A(_02223_),
    .B(_02224_));
 sg13g2_o21ai_1 _09215_ (.B1(net1997),
    .Y(_02226_),
    .A1(net1860),
    .A2(net3030));
 sg13g2_a21oi_1 _09216_ (.A1(net1860),
    .A2(_02225_),
    .Y(_00237_),
    .B1(_02226_));
 sg13g2_nor2_1 _09217_ (.A(\am_sdr0.cic3.comb1_in_del[14] ),
    .B(_01544_),
    .Y(_02227_));
 sg13g2_xnor2_1 _09218_ (.Y(_02228_),
    .A(\am_sdr0.cic3.comb1_in_del[14] ),
    .B(net2762));
 sg13g2_inv_1 _09219_ (.Y(_02229_),
    .A(_02228_));
 sg13g2_nor2_1 _09220_ (.A(_02209_),
    .B(_02222_),
    .Y(_02230_));
 sg13g2_a21oi_1 _09221_ (.A1(_02217_),
    .A2(_02230_),
    .Y(_02231_),
    .B1(_02221_));
 sg13g2_a221oi_1 _09222_ (.B2(_02230_),
    .C1(_02229_),
    .B1(_02217_),
    .A1(\am_sdr0.cic3.comb1_in_del[13] ),
    .Y(_02232_),
    .A2(_01545_));
 sg13g2_xnor2_1 _09223_ (.Y(_02233_),
    .A(_02228_),
    .B(_02231_));
 sg13g2_o21ai_1 _09224_ (.B1(net1999),
    .Y(_02234_),
    .A1(net1861),
    .A2(net2321));
 sg13g2_a21oi_1 _09225_ (.A1(net1851),
    .A2(_02233_),
    .Y(_00238_),
    .B1(_02234_));
 sg13g2_nand2_1 _09226_ (.Y(_02235_),
    .A(_01542_),
    .B(\am_sdr0.cic3.integ_sample[15] ));
 sg13g2_xor2_1 _09227_ (.B(net3017),
    .A(net2813),
    .X(_02236_));
 sg13g2_o21ai_1 _09228_ (.B1(_02236_),
    .Y(_02237_),
    .A1(_02227_),
    .A2(_02232_));
 sg13g2_nor3_1 _09229_ (.A(_02227_),
    .B(_02232_),
    .C(_02236_),
    .Y(_02238_));
 sg13g2_nor2_1 _09230_ (.A(net1625),
    .B(_02238_),
    .Y(_02239_));
 sg13g2_a221oi_1 _09231_ (.B2(_02239_),
    .C1(net1890),
    .B1(_02237_),
    .A1(net1625),
    .Y(_00239_),
    .A2(_01519_));
 sg13g2_or2_1 _09232_ (.X(_02240_),
    .B(_02236_),
    .A(_02229_));
 sg13g2_nor4_1 _09233_ (.A(_02210_),
    .B(_02221_),
    .C(_02222_),
    .D(_02240_),
    .Y(_02241_));
 sg13g2_o21ai_1 _09234_ (.B1(_02227_),
    .Y(_02242_),
    .A1(_01542_),
    .A2(\am_sdr0.cic3.integ_sample[15] ));
 sg13g2_nor3_1 _09235_ (.A(_02221_),
    .B(_02230_),
    .C(_02240_),
    .Y(_02243_));
 sg13g2_a21oi_1 _09236_ (.A1(_02214_),
    .A2(_02241_),
    .Y(_02244_),
    .B1(_02243_));
 sg13g2_nand3_1 _09237_ (.B(_02242_),
    .C(_02244_),
    .A(_02235_),
    .Y(_02245_));
 sg13g2_a21o_1 _09238_ (.A2(_02241_),
    .A1(_02216_),
    .B1(_02245_),
    .X(_02246_));
 sg13g2_nor2_1 _09239_ (.A(\am_sdr0.cic3.comb1_in_del[16] ),
    .B(_01541_),
    .Y(_02247_));
 sg13g2_xnor2_1 _09240_ (.Y(_02248_),
    .A(\am_sdr0.cic3.comb1_in_del[16] ),
    .B(net2796));
 sg13g2_inv_1 _09241_ (.Y(_02249_),
    .A(_02248_));
 sg13g2_xnor2_1 _09242_ (.Y(_02250_),
    .A(_02246_),
    .B(_02248_));
 sg13g2_o21ai_1 _09243_ (.B1(net1999),
    .Y(_02251_),
    .A1(net1851),
    .A2(net2365));
 sg13g2_a21oi_1 _09244_ (.A1(net1851),
    .A2(_02250_),
    .Y(_00240_),
    .B1(_02251_));
 sg13g2_nand2_1 _09245_ (.Y(_02252_),
    .A(\am_sdr0.cic3.comb1_in_del[17] ),
    .B(_01540_));
 sg13g2_nor2_1 _09246_ (.A(\am_sdr0.cic3.comb1_in_del[17] ),
    .B(_01540_),
    .Y(_02253_));
 sg13g2_xor2_1 _09247_ (.B(\am_sdr0.cic3.integ_sample[17] ),
    .A(\am_sdr0.cic3.comb1_in_del[17] ),
    .X(_02254_));
 sg13g2_a21oi_1 _09248_ (.A1(_02246_),
    .A2(_02248_),
    .Y(_02255_),
    .B1(_02247_));
 sg13g2_xnor2_1 _09249_ (.Y(_02256_),
    .A(_02254_),
    .B(_02255_));
 sg13g2_o21ai_1 _09250_ (.B1(net1995),
    .Y(_02257_),
    .A1(net1851),
    .A2(net2736));
 sg13g2_a21oi_1 _09251_ (.A1(net1851),
    .A2(_02256_),
    .Y(_00241_),
    .B1(_02257_));
 sg13g2_nand2b_1 _09252_ (.Y(_02258_),
    .B(net2476),
    .A_N(\am_sdr0.cic3.comb1_in_del[18] ));
 sg13g2_xor2_1 _09253_ (.B(net2476),
    .A(net2853),
    .X(_02259_));
 sg13g2_nor2_1 _09254_ (.A(_02249_),
    .B(_02254_),
    .Y(_02260_));
 sg13g2_a221oi_1 _09255_ (.B2(_02246_),
    .C1(_02253_),
    .B1(_02260_),
    .A1(_02247_),
    .Y(_02261_),
    .A2(_02252_));
 sg13g2_xnor2_1 _09256_ (.Y(_02262_),
    .A(_02259_),
    .B(_02261_));
 sg13g2_o21ai_1 _09257_ (.B1(net1995),
    .Y(_02263_),
    .A1(net1854),
    .A2(net2363));
 sg13g2_a21oi_1 _09258_ (.A1(net1854),
    .A2(net2854),
    .Y(_00242_),
    .B1(_02263_));
 sg13g2_o21ai_1 _09259_ (.B1(_02258_),
    .Y(_02264_),
    .A1(_02259_),
    .A2(_02261_));
 sg13g2_xnor2_1 _09260_ (.Y(_02265_),
    .A(net2198),
    .B(net2194));
 sg13g2_xnor2_1 _09261_ (.Y(_02266_),
    .A(_02264_),
    .B(_02265_));
 sg13g2_o21ai_1 _09262_ (.B1(net1994),
    .Y(_02267_),
    .A1(net1853),
    .A2(net2798));
 sg13g2_a21oi_1 _09263_ (.A1(net1853),
    .A2(_02266_),
    .Y(_00243_),
    .B1(_02267_));
 sg13g2_o21ai_1 _09264_ (.B1(net1985),
    .Y(_02268_),
    .A1(net1831),
    .A2(net2413));
 sg13g2_a21oi_1 _09265_ (.A1(net1831),
    .A2(_01561_),
    .Y(_00244_),
    .B1(_02268_));
 sg13g2_o21ai_1 _09266_ (.B1(net1982),
    .Y(_02269_),
    .A1(net1831),
    .A2(net2372));
 sg13g2_a21oi_1 _09267_ (.A1(net1835),
    .A2(_01559_),
    .Y(_00245_),
    .B1(_02269_));
 sg13g2_o21ai_1 _09268_ (.B1(net1982),
    .Y(_02270_),
    .A1(net1831),
    .A2(net2602));
 sg13g2_a21oi_1 _09269_ (.A1(net1831),
    .A2(_01558_),
    .Y(_00246_),
    .B1(_02270_));
 sg13g2_o21ai_1 _09270_ (.B1(net1985),
    .Y(_02271_),
    .A1(net1831),
    .A2(net2506));
 sg13g2_a21oi_1 _09271_ (.A1(net1831),
    .A2(_01557_),
    .Y(_00247_),
    .B1(_02271_));
 sg13g2_o21ai_1 _09272_ (.B1(net1988),
    .Y(_02272_),
    .A1(net1832),
    .A2(net2735));
 sg13g2_a21oi_1 _09273_ (.A1(net1832),
    .A2(_01556_),
    .Y(_00248_),
    .B1(_02272_));
 sg13g2_o21ai_1 _09274_ (.B1(net1988),
    .Y(_02273_),
    .A1(net1832),
    .A2(net2957));
 sg13g2_a21oi_1 _09275_ (.A1(net1831),
    .A2(_01555_),
    .Y(_00249_),
    .B1(_02273_));
 sg13g2_o21ai_1 _09276_ (.B1(net1982),
    .Y(_02274_),
    .A1(net1832),
    .A2(net2635));
 sg13g2_a21oi_1 _09277_ (.A1(net1832),
    .A2(_01553_),
    .Y(_00250_),
    .B1(_02274_));
 sg13g2_o21ai_1 _09278_ (.B1(net1984),
    .Y(_02275_),
    .A1(net1833),
    .A2(net2552));
 sg13g2_a21oi_1 _09279_ (.A1(net1833),
    .A2(_01552_),
    .Y(_00251_),
    .B1(_02275_));
 sg13g2_o21ai_1 _09280_ (.B1(net1991),
    .Y(_02276_),
    .A1(net1833),
    .A2(net2728));
 sg13g2_a21oi_1 _09281_ (.A1(net1833),
    .A2(_01551_),
    .Y(_00252_),
    .B1(_02276_));
 sg13g2_o21ai_1 _09282_ (.B1(net1991),
    .Y(_02277_),
    .A1(net1833),
    .A2(net2889));
 sg13g2_a21oi_1 _09283_ (.A1(net1833),
    .A2(_01550_),
    .Y(_00253_),
    .B1(_02277_));
 sg13g2_o21ai_1 _09284_ (.B1(net1984),
    .Y(_02278_),
    .A1(net1833),
    .A2(net2696));
 sg13g2_a21oi_1 _09285_ (.A1(net1833),
    .A2(_01548_),
    .Y(_00254_),
    .B1(_02278_));
 sg13g2_o21ai_1 _09286_ (.B1(net1984),
    .Y(_02279_),
    .A1(net1834),
    .A2(net2306));
 sg13g2_a21oi_1 _09287_ (.A1(net1834),
    .A2(_01547_),
    .Y(_00255_),
    .B1(_02279_));
 sg13g2_o21ai_1 _09288_ (.B1(net1996),
    .Y(_02280_),
    .A1(net1834),
    .A2(net2769));
 sg13g2_a21oi_1 _09289_ (.A1(net1834),
    .A2(_01546_),
    .Y(_00256_),
    .B1(_02280_));
 sg13g2_o21ai_1 _09290_ (.B1(net1997),
    .Y(_02281_),
    .A1(net1850),
    .A2(net2939));
 sg13g2_a21oi_1 _09291_ (.A1(net1850),
    .A2(_01545_),
    .Y(_00257_),
    .B1(_02281_));
 sg13g2_o21ai_1 _09292_ (.B1(net1993),
    .Y(_02282_),
    .A1(net1850),
    .A2(\am_sdr0.cic3.comb1_in_del[14] ));
 sg13g2_a21oi_1 _09293_ (.A1(net1850),
    .A2(_01544_),
    .Y(_00258_),
    .B1(_02282_));
 sg13g2_o21ai_1 _09294_ (.B1(net1993),
    .Y(_02283_),
    .A1(net1850),
    .A2(net2813));
 sg13g2_a21oi_1 _09295_ (.A1(net1850),
    .A2(_01543_),
    .Y(_00259_),
    .B1(_02283_));
 sg13g2_o21ai_1 _09296_ (.B1(net1995),
    .Y(_02284_),
    .A1(net1852),
    .A2(\am_sdr0.cic3.comb1_in_del[16] ));
 sg13g2_a21oi_1 _09297_ (.A1(net1852),
    .A2(_01541_),
    .Y(_00260_),
    .B1(_02284_));
 sg13g2_o21ai_1 _09298_ (.B1(net1995),
    .Y(_02285_),
    .A1(net1852),
    .A2(net2887));
 sg13g2_a21oi_1 _09299_ (.A1(net1852),
    .A2(_01540_),
    .Y(_00261_),
    .B1(_02285_));
 sg13g2_o21ai_1 _09300_ (.B1(net1995),
    .Y(_02286_),
    .A1(net1852),
    .A2(\am_sdr0.cic3.comb1_in_del[18] ));
 sg13g2_a21oi_1 _09301_ (.A1(net1852),
    .A2(_01539_),
    .Y(_00262_),
    .B1(_02286_));
 sg13g2_o21ai_1 _09302_ (.B1(net1994),
    .Y(_02287_),
    .A1(net1853),
    .A2(net2198));
 sg13g2_a21oi_1 _09303_ (.A1(net1853),
    .A2(_01538_),
    .Y(_00263_),
    .B1(_02287_));
 sg13g2_nand2b_1 _09304_ (.Y(_02288_),
    .B(net2358),
    .A_N(net2260));
 sg13g2_a21oi_1 _09305_ (.A1(_01536_),
    .A2(net2260),
    .Y(_02289_),
    .B1(net1622));
 sg13g2_a221oi_1 _09306_ (.B2(_02289_),
    .C1(net1890),
    .B1(_02288_),
    .A1(net1623),
    .Y(_00264_),
    .A2(_01506_));
 sg13g2_nor2b_1 _09307_ (.A(net2772),
    .B_N(\am_sdr0.cic3.comb1[1] ),
    .Y(_02290_));
 sg13g2_xnor2_1 _09308_ (.Y(_02291_),
    .A(net2772),
    .B(net2347));
 sg13g2_xnor2_1 _09309_ (.Y(_02292_),
    .A(_02288_),
    .B(_02291_));
 sg13g2_o21ai_1 _09310_ (.B1(net1986),
    .Y(_02293_),
    .A1(net1839),
    .A2(net2045));
 sg13g2_a21oi_1 _09311_ (.A1(net1839),
    .A2(_02292_),
    .Y(_00265_),
    .B1(_02293_));
 sg13g2_nand2b_1 _09312_ (.Y(_02294_),
    .B(\am_sdr0.cic3.comb1[2] ),
    .A_N(\am_sdr0.cic3.comb2_in_del[2] ));
 sg13g2_xor2_1 _09313_ (.B(\am_sdr0.cic3.comb1[2] ),
    .A(\am_sdr0.cic3.comb2_in_del[2] ),
    .X(_02295_));
 sg13g2_a21oi_1 _09314_ (.A1(_02288_),
    .A2(_02291_),
    .Y(_02296_),
    .B1(_02290_));
 sg13g2_xnor2_1 _09315_ (.Y(_02297_),
    .A(_02295_),
    .B(_02296_));
 sg13g2_o21ai_1 _09316_ (.B1(net1986),
    .Y(_02298_),
    .A1(net1839),
    .A2(net2859));
 sg13g2_a21oi_1 _09317_ (.A1(net1839),
    .A2(_02297_),
    .Y(_00266_),
    .B1(_02298_));
 sg13g2_nor2_1 _09318_ (.A(\am_sdr0.cic3.comb2_in_del[3] ),
    .B(_01533_),
    .Y(_02299_));
 sg13g2_nand2_1 _09319_ (.Y(_02300_),
    .A(\am_sdr0.cic3.comb2_in_del[3] ),
    .B(_01533_));
 sg13g2_nand2b_1 _09320_ (.Y(_02301_),
    .B(_02300_),
    .A_N(_02299_));
 sg13g2_o21ai_1 _09321_ (.B1(_02294_),
    .Y(_02302_),
    .A1(_02295_),
    .A2(_02296_));
 sg13g2_xnor2_1 _09322_ (.Y(_02303_),
    .A(_02301_),
    .B(_02302_));
 sg13g2_o21ai_1 _09323_ (.B1(net1987),
    .Y(_02304_),
    .A1(net1623),
    .A2(_02303_));
 sg13g2_a21oi_1 _09324_ (.A1(net1622),
    .A2(_01503_),
    .Y(_00267_),
    .B1(_02304_));
 sg13g2_nor2_1 _09325_ (.A(net3322),
    .B(_01532_),
    .Y(_02305_));
 sg13g2_xor2_1 _09326_ (.B(net2595),
    .A(\am_sdr0.cic3.comb2_in_del[4] ),
    .X(_02306_));
 sg13g2_a21oi_1 _09327_ (.A1(_02300_),
    .A2(_02302_),
    .Y(_02307_),
    .B1(_02299_));
 sg13g2_or2_1 _09328_ (.X(_02308_),
    .B(_02307_),
    .A(_02306_));
 sg13g2_xnor2_1 _09329_ (.Y(_02309_),
    .A(net2596),
    .B(_02307_));
 sg13g2_o21ai_1 _09330_ (.B1(net1987),
    .Y(_02310_),
    .A1(net1840),
    .A2(net2228));
 sg13g2_a21oi_1 _09331_ (.A1(net1840),
    .A2(_02309_),
    .Y(_00268_),
    .B1(_02310_));
 sg13g2_xor2_1 _09332_ (.B(net2449),
    .A(\am_sdr0.cic3.comb2_in_del[5] ),
    .X(_02311_));
 sg13g2_nor2b_1 _09333_ (.A(_02305_),
    .B_N(_02308_),
    .Y(_02312_));
 sg13g2_xnor2_1 _09334_ (.Y(_02313_),
    .A(net2450),
    .B(_02312_));
 sg13g2_o21ai_1 _09335_ (.B1(net1987),
    .Y(_02314_),
    .A1(net1841),
    .A2(net2232));
 sg13g2_a21oi_1 _09336_ (.A1(net1841),
    .A2(_02313_),
    .Y(_00269_),
    .B1(_02314_));
 sg13g2_nor2_1 _09337_ (.A(\am_sdr0.cic3.comb2_in_del[6] ),
    .B(_01529_),
    .Y(_02315_));
 sg13g2_xor2_1 _09338_ (.B(\am_sdr0.cic3.comb1[6] ),
    .A(net2719),
    .X(_02316_));
 sg13g2_a21oi_1 _09339_ (.A1(_01530_),
    .A2(\am_sdr0.cic3.comb1[5] ),
    .Y(_02317_),
    .B1(_02305_));
 sg13g2_a22oi_1 _09340_ (.Y(_02318_),
    .B1(_02308_),
    .B2(_02317_),
    .A2(_01531_),
    .A1(\am_sdr0.cic3.comb2_in_del[5] ));
 sg13g2_a221oi_1 _09341_ (.B2(_02317_),
    .C1(_02316_),
    .B1(_02308_),
    .A1(\am_sdr0.cic3.comb2_in_del[5] ),
    .Y(_02319_),
    .A2(_01531_));
 sg13g2_xor2_1 _09342_ (.B(_02318_),
    .A(_02316_),
    .X(_02320_));
 sg13g2_o21ai_1 _09343_ (.B1(net1989),
    .Y(_02321_),
    .A1(net1848),
    .A2(net2770));
 sg13g2_a21oi_1 _09344_ (.A1(net1848),
    .A2(_02320_),
    .Y(_00270_),
    .B1(_02321_));
 sg13g2_nand2b_1 _09345_ (.Y(_02322_),
    .B(\am_sdr0.cic3.comb1[7] ),
    .A_N(\am_sdr0.cic3.comb2_in_del[7] ));
 sg13g2_xnor2_1 _09346_ (.Y(_02323_),
    .A(\am_sdr0.cic3.comb2_in_del[7] ),
    .B(\am_sdr0.cic3.comb1[7] ));
 sg13g2_o21ai_1 _09347_ (.B1(_02323_),
    .Y(_02324_),
    .A1(_02315_),
    .A2(_02319_));
 sg13g2_or3_1 _09348_ (.A(_02315_),
    .B(_02319_),
    .C(_02323_),
    .X(_02325_));
 sg13g2_and2_1 _09349_ (.A(_02324_),
    .B(_02325_),
    .X(_02326_));
 sg13g2_o21ai_1 _09350_ (.B1(net1989),
    .Y(_02327_),
    .A1(net1624),
    .A2(_02326_));
 sg13g2_a21oi_1 _09351_ (.A1(net1623),
    .A2(_01496_),
    .Y(_00271_),
    .B1(_02327_));
 sg13g2_nand2_1 _09352_ (.Y(_02328_),
    .A(_02322_),
    .B(_02324_));
 sg13g2_nor2_1 _09353_ (.A(\am_sdr0.cic3.comb2_in_del[8] ),
    .B(_01527_),
    .Y(_02329_));
 sg13g2_xnor2_1 _09354_ (.Y(_02330_),
    .A(\am_sdr0.cic3.comb2_in_del[8] ),
    .B(\am_sdr0.cic3.comb1[8] ));
 sg13g2_inv_1 _09355_ (.Y(_02331_),
    .A(_02330_));
 sg13g2_xnor2_1 _09356_ (.Y(_02332_),
    .A(_02328_),
    .B(_02330_));
 sg13g2_o21ai_1 _09357_ (.B1(net1990),
    .Y(_02333_),
    .A1(net1846),
    .A2(net2784));
 sg13g2_a21oi_1 _09358_ (.A1(net1846),
    .A2(_02332_),
    .Y(_00272_),
    .B1(_02333_));
 sg13g2_xor2_1 _09359_ (.B(\am_sdr0.cic3.comb1[9] ),
    .A(\am_sdr0.cic3.comb2_in_del[9] ),
    .X(_02334_));
 sg13g2_a21oi_1 _09360_ (.A1(_02328_),
    .A2(_02330_),
    .Y(_02335_),
    .B1(_02329_));
 sg13g2_xnor2_1 _09361_ (.Y(_02336_),
    .A(_02334_),
    .B(_02335_));
 sg13g2_o21ai_1 _09362_ (.B1(net1990),
    .Y(_02337_),
    .A1(net1846),
    .A2(net2650));
 sg13g2_a21oi_1 _09363_ (.A1(net1847),
    .A2(_02336_),
    .Y(_00273_),
    .B1(_02337_));
 sg13g2_nand2b_1 _09364_ (.Y(_02338_),
    .B(\am_sdr0.cic3.comb1[10] ),
    .A_N(\am_sdr0.cic3.comb2_in_del[10] ));
 sg13g2_xor2_1 _09365_ (.B(net2558),
    .A(\am_sdr0.cic3.comb2_in_del[10] ),
    .X(_02339_));
 sg13g2_a21oi_1 _09366_ (.A1(_01525_),
    .A2(\am_sdr0.cic3.comb1[9] ),
    .Y(_02340_),
    .B1(_02329_));
 sg13g2_a21oi_1 _09367_ (.A1(\am_sdr0.cic3.comb2_in_del[9] ),
    .A2(_01526_),
    .Y(_02341_),
    .B1(_02340_));
 sg13g2_nor2_1 _09368_ (.A(_02331_),
    .B(_02334_),
    .Y(_02342_));
 sg13g2_a21oi_1 _09369_ (.A1(_02328_),
    .A2(_02342_),
    .Y(_02343_),
    .B1(_02341_));
 sg13g2_xnor2_1 _09370_ (.Y(_02344_),
    .A(_02339_),
    .B(_02343_));
 sg13g2_o21ai_1 _09371_ (.B1(net1998),
    .Y(_02345_),
    .A1(net1847),
    .A2(net2757));
 sg13g2_a21oi_1 _09372_ (.A1(net1847),
    .A2(_02344_),
    .Y(_00274_),
    .B1(_02345_));
 sg13g2_nor2b_1 _09373_ (.A(\am_sdr0.cic3.comb1[11] ),
    .B_N(\am_sdr0.cic3.comb2_in_del[11] ),
    .Y(_02346_));
 sg13g2_nand2b_1 _09374_ (.Y(_02347_),
    .B(\am_sdr0.cic3.comb1[11] ),
    .A_N(\am_sdr0.cic3.comb2_in_del[11] ));
 sg13g2_nand2b_1 _09375_ (.Y(_02348_),
    .B(_02347_),
    .A_N(_02346_));
 sg13g2_o21ai_1 _09376_ (.B1(net2559),
    .Y(_02349_),
    .A1(_02339_),
    .A2(_02343_));
 sg13g2_xor2_1 _09377_ (.B(_02349_),
    .A(_02348_),
    .X(_02350_));
 sg13g2_o21ai_1 _09378_ (.B1(net1998),
    .Y(_02351_),
    .A1(net1846),
    .A2(net2213));
 sg13g2_a21oi_1 _09379_ (.A1(net1847),
    .A2(_02350_),
    .Y(_00275_),
    .B1(_02351_));
 sg13g2_nor2_2 _09380_ (.A(net2742),
    .B(_01522_),
    .Y(_02352_));
 sg13g2_nor2b_1 _09381_ (.A(\am_sdr0.cic3.comb1[12] ),
    .B_N(\am_sdr0.cic3.comb2_in_del[12] ),
    .Y(_02353_));
 sg13g2_nor2_1 _09382_ (.A(_02352_),
    .B(_02353_),
    .Y(_02354_));
 sg13g2_nor2_1 _09383_ (.A(_02339_),
    .B(_02348_),
    .Y(_02355_));
 sg13g2_o21ai_1 _09384_ (.B1(_02347_),
    .Y(_02356_),
    .A1(_02338_),
    .A2(_02346_));
 sg13g2_a21o_1 _09385_ (.A2(_02355_),
    .A1(_02341_),
    .B1(_02356_),
    .X(_02357_));
 sg13g2_nand2_1 _09386_ (.Y(_02358_),
    .A(_02342_),
    .B(_02355_));
 sg13g2_a21oi_2 _09387_ (.B1(_02358_),
    .Y(_02359_),
    .A2(_02324_),
    .A1(_02322_));
 sg13g2_o21ai_1 _09388_ (.B1(_02354_),
    .Y(_02360_),
    .A1(_02357_),
    .A2(_02359_));
 sg13g2_or3_1 _09389_ (.A(_02354_),
    .B(_02357_),
    .C(_02359_),
    .X(_02361_));
 sg13g2_nand2_1 _09390_ (.Y(_02362_),
    .A(_02360_),
    .B(_02361_));
 sg13g2_o21ai_1 _09391_ (.B1(net2001),
    .Y(_02363_),
    .A1(net1862),
    .A2(net2270));
 sg13g2_a21oi_1 _09392_ (.A1(net1862),
    .A2(_02362_),
    .Y(_00276_),
    .B1(_02363_));
 sg13g2_nor2_1 _09393_ (.A(_01521_),
    .B(\am_sdr0.cic3.comb1[13] ),
    .Y(_02364_));
 sg13g2_xor2_1 _09394_ (.B(\am_sdr0.cic3.comb1[13] ),
    .A(net2540),
    .X(_02365_));
 sg13g2_nor2b_1 _09395_ (.A(_02352_),
    .B_N(_02360_),
    .Y(_02366_));
 sg13g2_xnor2_1 _09396_ (.Y(_02367_),
    .A(_02365_),
    .B(_02366_));
 sg13g2_o21ai_1 _09397_ (.B1(net2001),
    .Y(_02368_),
    .A1(net1862),
    .A2(net2542));
 sg13g2_a21oi_1 _09398_ (.A1(net1862),
    .A2(_02367_),
    .Y(_00277_),
    .B1(_02368_));
 sg13g2_nor2_1 _09399_ (.A(\am_sdr0.cic3.comb2_in_del[14] ),
    .B(_01520_),
    .Y(_02369_));
 sg13g2_xnor2_1 _09400_ (.Y(_02370_),
    .A(\am_sdr0.cic3.comb2_in_del[14] ),
    .B(\am_sdr0.cic3.comb1[14] ));
 sg13g2_a21oi_1 _09401_ (.A1(_01521_),
    .A2(\am_sdr0.cic3.comb1[13] ),
    .Y(_02371_),
    .B1(_02352_));
 sg13g2_a21oi_1 _09402_ (.A1(_02360_),
    .A2(_02371_),
    .Y(_02372_),
    .B1(_02364_));
 sg13g2_xnor2_1 _09403_ (.Y(_02373_),
    .A(_02370_),
    .B(_02372_));
 sg13g2_o21ai_1 _09404_ (.B1(net2000),
    .Y(_02374_),
    .A1(net1865),
    .A2(net2300));
 sg13g2_a21oi_1 _09405_ (.A1(net1861),
    .A2(_02373_),
    .Y(_00278_),
    .B1(_02374_));
 sg13g2_nand2_1 _09406_ (.Y(_02375_),
    .A(\am_sdr0.cic3.comb2_in_del[15] ),
    .B(_01519_));
 sg13g2_nor2_1 _09407_ (.A(\am_sdr0.cic3.comb2_in_del[15] ),
    .B(_01519_),
    .Y(_02376_));
 sg13g2_xor2_1 _09408_ (.B(net2758),
    .A(\am_sdr0.cic3.comb2_in_del[15] ),
    .X(_02377_));
 sg13g2_a21oi_1 _09409_ (.A1(_02370_),
    .A2(_02372_),
    .Y(_02378_),
    .B1(_02369_));
 sg13g2_xnor2_1 _09410_ (.Y(_02379_),
    .A(_02377_),
    .B(_02378_));
 sg13g2_o21ai_1 _09411_ (.B1(net2000),
    .Y(_02380_),
    .A1(net1860),
    .A2(net2885));
 sg13g2_a21oi_1 _09412_ (.A1(net1860),
    .A2(_02379_),
    .Y(_00279_),
    .B1(_02380_));
 sg13g2_nor2_1 _09413_ (.A(\am_sdr0.cic3.comb2_in_del[16] ),
    .B(_01518_),
    .Y(_02381_));
 sg13g2_xnor2_1 _09414_ (.Y(_02382_),
    .A(\am_sdr0.cic3.comb2_in_del[16] ),
    .B(net2764));
 sg13g2_inv_1 _09415_ (.Y(_02383_),
    .A(_02382_));
 sg13g2_nand3b_1 _09416_ (.B(_02370_),
    .C(_02375_),
    .Y(_02384_),
    .A_N(_02376_));
 sg13g2_nor4_1 _09417_ (.A(_02352_),
    .B(_02353_),
    .C(_02365_),
    .D(_02384_),
    .Y(_02385_));
 sg13g2_nor3_1 _09418_ (.A(_02364_),
    .B(_02371_),
    .C(_02384_),
    .Y(_02386_));
 sg13g2_a221oi_1 _09419_ (.B2(_02357_),
    .C1(_02376_),
    .B1(_02385_),
    .A1(_02369_),
    .Y(_02387_),
    .A2(_02375_));
 sg13g2_nand2b_1 _09420_ (.Y(_02388_),
    .B(_02387_),
    .A_N(_02386_));
 sg13g2_a21o_1 _09421_ (.A2(_02385_),
    .A1(_02359_),
    .B1(_02388_),
    .X(_02389_));
 sg13g2_xnor2_1 _09422_ (.Y(_02390_),
    .A(_02382_),
    .B(_02389_));
 sg13g2_o21ai_1 _09423_ (.B1(net2000),
    .Y(_02391_),
    .A1(net1865),
    .A2(net2490));
 sg13g2_a21oi_1 _09424_ (.A1(net1865),
    .A2(_02390_),
    .Y(_00280_),
    .B1(_02391_));
 sg13g2_nand2_1 _09425_ (.Y(_02392_),
    .A(\am_sdr0.cic3.comb2_in_del[17] ),
    .B(_01517_));
 sg13g2_nor2_1 _09426_ (.A(\am_sdr0.cic3.comb2_in_del[17] ),
    .B(_01517_),
    .Y(_02393_));
 sg13g2_xor2_1 _09427_ (.B(net2862),
    .A(\am_sdr0.cic3.comb2_in_del[17] ),
    .X(_02394_));
 sg13g2_a21oi_1 _09428_ (.A1(_02382_),
    .A2(_02389_),
    .Y(_02395_),
    .B1(_02381_));
 sg13g2_xnor2_1 _09429_ (.Y(_02396_),
    .A(_02394_),
    .B(_02395_));
 sg13g2_o21ai_1 _09430_ (.B1(net1999),
    .Y(_02397_),
    .A1(net1856),
    .A2(net2203));
 sg13g2_a21oi_1 _09431_ (.A1(net1856),
    .A2(_02396_),
    .Y(_00281_),
    .B1(_02397_));
 sg13g2_nand2b_1 _09432_ (.Y(_02398_),
    .B(net3315),
    .A_N(\am_sdr0.cic3.comb2_in_del[18] ));
 sg13g2_xor2_1 _09433_ (.B(net2826),
    .A(\am_sdr0.cic3.comb2_in_del[18] ),
    .X(_02399_));
 sg13g2_nor2_1 _09434_ (.A(_02383_),
    .B(_02394_),
    .Y(_02400_));
 sg13g2_a221oi_1 _09435_ (.B2(_02389_),
    .C1(_02393_),
    .B1(_02400_),
    .A1(_02381_),
    .Y(_02401_),
    .A2(_02392_));
 sg13g2_xnor2_1 _09436_ (.Y(_02402_),
    .A(_02399_),
    .B(_02401_));
 sg13g2_o21ai_1 _09437_ (.B1(net2017),
    .Y(_02403_),
    .A1(net1856),
    .A2(net2423));
 sg13g2_a21oi_1 _09438_ (.A1(net1856),
    .A2(_02402_),
    .Y(_00282_),
    .B1(_02403_));
 sg13g2_o21ai_1 _09439_ (.B1(_02398_),
    .Y(_02404_),
    .A1(_02399_),
    .A2(_02401_));
 sg13g2_xnor2_1 _09440_ (.Y(_02405_),
    .A(net2435),
    .B(net2798));
 sg13g2_xnor2_1 _09441_ (.Y(_02406_),
    .A(_02404_),
    .B(_02405_));
 sg13g2_o21ai_1 _09442_ (.B1(net2017),
    .Y(_02407_),
    .A1(net2191),
    .A2(net1853));
 sg13g2_a21oi_1 _09443_ (.A1(net1854),
    .A2(_02406_),
    .Y(_00283_),
    .B1(_02407_));
 sg13g2_o21ai_1 _09444_ (.B1(net1985),
    .Y(_02408_),
    .A1(net1836),
    .A2(\am_sdr0.cic3.comb2_in_del[0] ));
 sg13g2_a21oi_1 _09445_ (.A1(net1836),
    .A2(_01537_),
    .Y(_00284_),
    .B1(_02408_));
 sg13g2_o21ai_1 _09446_ (.B1(net1986),
    .Y(_02409_),
    .A1(net1837),
    .A2(\am_sdr0.cic3.comb2_in_del[1] ));
 sg13g2_a21oi_1 _09447_ (.A1(net1837),
    .A2(_01535_),
    .Y(_00285_),
    .B1(_02409_));
 sg13g2_o21ai_1 _09448_ (.B1(net1986),
    .Y(_02410_),
    .A1(net1837),
    .A2(\am_sdr0.cic3.comb2_in_del[2] ));
 sg13g2_a21oi_1 _09449_ (.A1(net1837),
    .A2(_01534_),
    .Y(_00286_),
    .B1(_02410_));
 sg13g2_o21ai_1 _09450_ (.B1(net1987),
    .Y(_02411_),
    .A1(net1836),
    .A2(net2533));
 sg13g2_a21oi_1 _09451_ (.A1(net1836),
    .A2(_01533_),
    .Y(_00287_),
    .B1(_02411_));
 sg13g2_o21ai_1 _09452_ (.B1(net1987),
    .Y(_02412_),
    .A1(net1838),
    .A2(net2708));
 sg13g2_a21oi_1 _09453_ (.A1(net1838),
    .A2(_01532_),
    .Y(_00288_),
    .B1(_02412_));
 sg13g2_o21ai_1 _09454_ (.B1(net1989),
    .Y(_02413_),
    .A1(net1840),
    .A2(net2945));
 sg13g2_a21oi_1 _09455_ (.A1(net1840),
    .A2(_01531_),
    .Y(_00289_),
    .B1(_02413_));
 sg13g2_o21ai_1 _09456_ (.B1(net1989),
    .Y(_02414_),
    .A1(net1845),
    .A2(net2719));
 sg13g2_a21oi_1 _09457_ (.A1(net1845),
    .A2(_01529_),
    .Y(_00290_),
    .B1(_02414_));
 sg13g2_o21ai_1 _09458_ (.B1(net1989),
    .Y(_02415_),
    .A1(net1845),
    .A2(\am_sdr0.cic3.comb2_in_del[7] ));
 sg13g2_a21oi_1 _09459_ (.A1(net1845),
    .A2(_01528_),
    .Y(_00291_),
    .B1(_02415_));
 sg13g2_o21ai_1 _09460_ (.B1(net1990),
    .Y(_02416_),
    .A1(net1845),
    .A2(net2665));
 sg13g2_a21oi_1 _09461_ (.A1(net1845),
    .A2(_01527_),
    .Y(_00292_),
    .B1(_02416_));
 sg13g2_o21ai_1 _09462_ (.B1(net1990),
    .Y(_02417_),
    .A1(net1843),
    .A2(\am_sdr0.cic3.comb2_in_del[9] ));
 sg13g2_a21oi_1 _09463_ (.A1(net1843),
    .A2(_01526_),
    .Y(_00293_),
    .B1(_02417_));
 sg13g2_o21ai_1 _09464_ (.B1(net1997),
    .Y(_02418_),
    .A1(net1844),
    .A2(\am_sdr0.cic3.comb2_in_del[10] ));
 sg13g2_a21oi_1 _09465_ (.A1(net1844),
    .A2(_01524_),
    .Y(_00294_),
    .B1(_02418_));
 sg13g2_o21ai_1 _09466_ (.B1(net1998),
    .Y(_02419_),
    .A1(net1844),
    .A2(\am_sdr0.cic3.comb2_in_del[11] ));
 sg13g2_a21oi_1 _09467_ (.A1(net1844),
    .A2(_01523_),
    .Y(_00295_),
    .B1(_02419_));
 sg13g2_o21ai_1 _09468_ (.B1(net1997),
    .Y(_02420_),
    .A1(net1860),
    .A2(net2742));
 sg13g2_a21oi_1 _09469_ (.A1(net1860),
    .A2(_01522_),
    .Y(_00296_),
    .B1(_02420_));
 sg13g2_o21ai_1 _09470_ (.B1(net1997),
    .Y(_02421_),
    .A1(net1625),
    .A2(\am_sdr0.cic3.comb1[13] ));
 sg13g2_a21oi_1 _09471_ (.A1(net1625),
    .A2(_01521_),
    .Y(_00297_),
    .B1(_02421_));
 sg13g2_o21ai_1 _09472_ (.B1(net1999),
    .Y(_02422_),
    .A1(net1861),
    .A2(\am_sdr0.cic3.comb2_in_del[14] ));
 sg13g2_a21oi_1 _09473_ (.A1(net1861),
    .A2(_01520_),
    .Y(_00298_),
    .B1(_02422_));
 sg13g2_o21ai_1 _09474_ (.B1(net1999),
    .Y(_02423_),
    .A1(net1861),
    .A2(\am_sdr0.cic3.comb2_in_del[15] ));
 sg13g2_a21oi_1 _09475_ (.A1(net1861),
    .A2(_01519_),
    .Y(_00299_),
    .B1(_02423_));
 sg13g2_o21ai_1 _09476_ (.B1(net1999),
    .Y(_02424_),
    .A1(net1850),
    .A2(\am_sdr0.cic3.comb2_in_del[16] ));
 sg13g2_a21oi_1 _09477_ (.A1(net1850),
    .A2(_01518_),
    .Y(_00300_),
    .B1(_02424_));
 sg13g2_o21ai_1 _09478_ (.B1(net1999),
    .Y(_02425_),
    .A1(net1859),
    .A2(net2933));
 sg13g2_a21oi_1 _09479_ (.A1(net1859),
    .A2(_01517_),
    .Y(_00301_),
    .B1(_02425_));
 sg13g2_o21ai_1 _09480_ (.B1(net1995),
    .Y(_02426_),
    .A1(net1854),
    .A2(\am_sdr0.cic3.comb2_in_del[18] ));
 sg13g2_a21oi_1 _09481_ (.A1(net1853),
    .A2(_01516_),
    .Y(_00302_),
    .B1(_02426_));
 sg13g2_o21ai_1 _09482_ (.B1(net2017),
    .Y(_02427_),
    .A1(net1853),
    .A2(net2435));
 sg13g2_a21oi_1 _09483_ (.A1(net1853),
    .A2(_01515_),
    .Y(_00303_),
    .B1(_02427_));
 sg13g2_nor2_1 _09484_ (.A(\am_sdr0.cic3.comb3_in_del[12] ),
    .B(_01488_),
    .Y(_02428_));
 sg13g2_xor2_1 _09485_ (.B(\am_sdr0.cic3.comb2[12] ),
    .A(\am_sdr0.cic3.comb3_in_del[12] ),
    .X(_02429_));
 sg13g2_nand2b_1 _09486_ (.Y(_02430_),
    .B(\am_sdr0.cic3.comb3_in_del[1] ),
    .A_N(\am_sdr0.cic3.comb2[1] ));
 sg13g2_nand2b_1 _09487_ (.Y(_02431_),
    .B(\am_sdr0.cic3.comb3_in_del[0] ),
    .A_N(\am_sdr0.cic3.comb2[0] ));
 sg13g2_nor2b_1 _09488_ (.A(\am_sdr0.cic3.comb3_in_del[1] ),
    .B_N(\am_sdr0.cic3.comb2[1] ),
    .Y(_02432_));
 sg13g2_a221oi_1 _09489_ (.B2(_02431_),
    .C1(_02432_),
    .B1(_02430_),
    .A1(_01504_),
    .Y(_02433_),
    .A2(\am_sdr0.cic3.comb2[2] ));
 sg13g2_nand2b_1 _09490_ (.Y(_02434_),
    .B(\am_sdr0.cic3.comb3_in_del[3] ),
    .A_N(\am_sdr0.cic3.comb2[3] ));
 sg13g2_o21ai_1 _09491_ (.B1(_02434_),
    .Y(_02435_),
    .A1(_01504_),
    .A2(\am_sdr0.cic3.comb2[2] ));
 sg13g2_a22oi_1 _09492_ (.Y(_02436_),
    .B1(_01502_),
    .B2(\am_sdr0.cic3.comb2[3] ),
    .A2(\am_sdr0.cic3.comb2[4] ),
    .A1(_01500_));
 sg13g2_o21ai_1 _09493_ (.B1(_02436_),
    .Y(_02437_),
    .A1(_02433_),
    .A2(_02435_));
 sg13g2_a22oi_1 _09494_ (.Y(_02438_),
    .B1(\am_sdr0.cic3.comb3_in_del[4] ),
    .B2(_01501_),
    .A2(_01499_),
    .A1(\am_sdr0.cic3.comb3_in_del[5] ));
 sg13g2_a22oi_1 _09495_ (.Y(_02439_),
    .B1(_02437_),
    .B2(_02438_),
    .A2(\am_sdr0.cic3.comb2[5] ),
    .A1(_01498_));
 sg13g2_nor2_1 _09496_ (.A(_01497_),
    .B(\am_sdr0.cic3.comb2[6] ),
    .Y(_02440_));
 sg13g2_a22oi_1 _09497_ (.Y(_02441_),
    .B1(_01497_),
    .B2(\am_sdr0.cic3.comb2[6] ),
    .A2(\am_sdr0.cic3.comb2[7] ),
    .A1(_01495_));
 sg13g2_o21ai_1 _09498_ (.B1(_02441_),
    .Y(_02442_),
    .A1(_02439_),
    .A2(_02440_));
 sg13g2_a22oi_1 _09499_ (.Y(_02443_),
    .B1(_01491_),
    .B2(\am_sdr0.cic3.comb2[10] ),
    .A2(\am_sdr0.cic3.comb2[11] ),
    .A1(_01489_));
 sg13g2_a22oi_1 _09500_ (.Y(_02444_),
    .B1(_01494_),
    .B2(\am_sdr0.cic3.comb2[8] ),
    .A2(\am_sdr0.cic3.comb2[9] ),
    .A1(_01493_));
 sg13g2_nand2_1 _09501_ (.Y(_02445_),
    .A(_02443_),
    .B(_02444_));
 sg13g2_nor2_1 _09502_ (.A(_01495_),
    .B(\am_sdr0.cic3.comb2[7] ),
    .Y(_02446_));
 sg13g2_nand2_1 _09503_ (.Y(_02447_),
    .A(\am_sdr0.cic3.comb3_in_del[11] ),
    .B(_01490_));
 sg13g2_o21ai_1 _09504_ (.B1(_02447_),
    .Y(_02448_),
    .A1(_01494_),
    .A2(\am_sdr0.cic3.comb2[8] ));
 sg13g2_nand2b_1 _09505_ (.Y(_02449_),
    .B(\am_sdr0.cic3.comb3_in_del[9] ),
    .A_N(\am_sdr0.cic3.comb2[9] ));
 sg13g2_o21ai_1 _09506_ (.B1(_02449_),
    .Y(_02450_),
    .A1(_01491_),
    .A2(\am_sdr0.cic3.comb2[10] ));
 sg13g2_nor4_1 _09507_ (.A(_02445_),
    .B(_02446_),
    .C(_02448_),
    .D(_02450_),
    .Y(_02451_));
 sg13g2_o21ai_1 _09508_ (.B1(_02443_),
    .Y(_02452_),
    .A1(_02444_),
    .A2(_02450_));
 sg13g2_a22oi_1 _09509_ (.Y(_02453_),
    .B1(_02452_),
    .B2(_02447_),
    .A2(_02451_),
    .A1(_02442_));
 sg13g2_nor2_1 _09510_ (.A(_02429_),
    .B(_02453_),
    .Y(_02454_));
 sg13g2_xnor2_1 _09511_ (.Y(_02455_),
    .A(_02429_),
    .B(_02453_));
 sg13g2_o21ai_1 _09512_ (.B1(net2023),
    .Y(_02456_),
    .A1(net1867),
    .A2(net1516));
 sg13g2_a21oi_1 _09513_ (.A1(net1866),
    .A2(_02455_),
    .Y(_00304_),
    .B1(_02456_));
 sg13g2_or2_1 _09514_ (.X(_02457_),
    .B(_02454_),
    .A(_02428_));
 sg13g2_nand2_1 _09515_ (.Y(_02458_),
    .A(\am_sdr0.cic3.comb3_in_del[13] ),
    .B(_01487_));
 sg13g2_nor2_1 _09516_ (.A(\am_sdr0.cic3.comb3_in_del[13] ),
    .B(_01487_),
    .Y(_02459_));
 sg13g2_xor2_1 _09517_ (.B(\am_sdr0.cic3.comb2[13] ),
    .A(\am_sdr0.cic3.comb3_in_del[13] ),
    .X(_02460_));
 sg13g2_or2_1 _09518_ (.X(_02461_),
    .B(net2543),
    .A(_02457_));
 sg13g2_a21oi_1 _09519_ (.A1(_02457_),
    .A2(net2543),
    .Y(_02462_),
    .B1(net1624));
 sg13g2_a221oi_1 _09520_ (.B2(_02462_),
    .C1(net1890),
    .B1(_02461_),
    .A1(net1624),
    .Y(_00305_),
    .A2(_01513_));
 sg13g2_nand2b_1 _09521_ (.Y(_02463_),
    .B(\am_sdr0.cic3.comb2[14] ),
    .A_N(\am_sdr0.cic3.comb3_in_del[14] ));
 sg13g2_xor2_1 _09522_ (.B(\am_sdr0.cic3.comb2[14] ),
    .A(\am_sdr0.cic3.comb3_in_del[14] ),
    .X(_02464_));
 sg13g2_or2_1 _09523_ (.X(_02465_),
    .B(_02460_),
    .A(_02429_));
 sg13g2_o21ai_1 _09524_ (.B1(_02458_),
    .Y(_02466_),
    .A1(_02428_),
    .A2(_02459_));
 sg13g2_o21ai_1 _09525_ (.B1(_02466_),
    .Y(_02467_),
    .A1(_02453_),
    .A2(_02465_));
 sg13g2_o21ai_1 _09526_ (.B1(_02458_),
    .Y(_02468_),
    .A1(_02457_),
    .A2(_02459_));
 sg13g2_xor2_1 _09527_ (.B(_02467_),
    .A(_02464_),
    .X(_02469_));
 sg13g2_o21ai_1 _09528_ (.B1(net2023),
    .Y(_02470_),
    .A1(net1866),
    .A2(net1452));
 sg13g2_a21oi_1 _09529_ (.A1(net1866),
    .A2(_02469_),
    .Y(_00306_),
    .B1(_02470_));
 sg13g2_nor2b_1 _09530_ (.A(\am_sdr0.cic3.comb2[15] ),
    .B_N(\am_sdr0.cic3.comb3_in_del[15] ),
    .Y(_02471_));
 sg13g2_nand2b_1 _09531_ (.Y(_02472_),
    .B(\am_sdr0.cic3.comb2[15] ),
    .A_N(\am_sdr0.cic3.comb3_in_del[15] ));
 sg13g2_nand2b_1 _09532_ (.Y(_02473_),
    .B(_02472_),
    .A_N(_02471_));
 sg13g2_o21ai_1 _09533_ (.B1(_02463_),
    .Y(_02474_),
    .A1(_02464_),
    .A2(_02468_));
 sg13g2_xor2_1 _09534_ (.B(_02474_),
    .A(_02473_),
    .X(_02475_));
 sg13g2_o21ai_1 _09535_ (.B1(net2023),
    .Y(_02476_),
    .A1(net1866),
    .A2(net1462));
 sg13g2_a21oi_1 _09536_ (.A1(net1866),
    .A2(_02475_),
    .Y(_00307_),
    .B1(_02476_));
 sg13g2_nor2_1 _09537_ (.A(\am_sdr0.cic3.comb3_in_del[16] ),
    .B(_01484_),
    .Y(_02477_));
 sg13g2_xnor2_1 _09538_ (.Y(_02478_),
    .A(\am_sdr0.cic3.comb3_in_del[16] ),
    .B(net2536));
 sg13g2_a21oi_1 _09539_ (.A1(_02463_),
    .A2(_02472_),
    .Y(_02479_),
    .B1(_02471_));
 sg13g2_nor2_1 _09540_ (.A(_02464_),
    .B(_02473_),
    .Y(_02480_));
 sg13g2_a21o_1 _09541_ (.A2(_02480_),
    .A1(_02467_),
    .B1(_02479_),
    .X(_02481_));
 sg13g2_xnor2_1 _09542_ (.Y(_02482_),
    .A(_02478_),
    .B(_02481_));
 sg13g2_o21ai_1 _09543_ (.B1(net2022),
    .Y(_02483_),
    .A1(net1864),
    .A2(net1319));
 sg13g2_a21oi_1 _09544_ (.A1(net1864),
    .A2(_02482_),
    .Y(_00308_),
    .B1(_02483_));
 sg13g2_a21oi_1 _09545_ (.A1(_02478_),
    .A2(_02481_),
    .Y(_02484_),
    .B1(_02477_));
 sg13g2_nor2b_1 _09546_ (.A(\am_sdr0.cic3.comb2[17] ),
    .B_N(\am_sdr0.cic3.comb3_in_del[17] ),
    .Y(_02485_));
 sg13g2_nand2b_1 _09547_ (.Y(_02486_),
    .B(net2353),
    .A_N(\am_sdr0.cic3.comb3_in_del[17] ));
 sg13g2_nand2b_1 _09548_ (.Y(_02487_),
    .B(_02486_),
    .A_N(_02485_));
 sg13g2_xnor2_1 _09549_ (.Y(_02488_),
    .A(_02484_),
    .B(_02487_));
 sg13g2_o21ai_1 _09550_ (.B1(net2022),
    .Y(_02489_),
    .A1(net1857),
    .A2(net1349));
 sg13g2_a21oi_1 _09551_ (.A1(net1857),
    .A2(_02488_),
    .Y(_00309_),
    .B1(_02489_));
 sg13g2_nor2_1 _09552_ (.A(\am_sdr0.cic3.comb3_in_del[18] ),
    .B(_01482_),
    .Y(_02490_));
 sg13g2_xnor2_1 _09553_ (.Y(_02491_),
    .A(\am_sdr0.cic3.comb3_in_del[18] ),
    .B(net2423));
 sg13g2_a21oi_1 _09554_ (.A1(_02484_),
    .A2(_02486_),
    .Y(_02492_),
    .B1(_02485_));
 sg13g2_xnor2_1 _09555_ (.Y(_02493_),
    .A(_02491_),
    .B(_02492_));
 sg13g2_o21ai_1 _09556_ (.B1(net2022),
    .Y(_02494_),
    .A1(net1857),
    .A2(net1355));
 sg13g2_a21oi_1 _09557_ (.A1(net1857),
    .A2(net2424),
    .Y(_00310_),
    .B1(_02494_));
 sg13g2_a21oi_1 _09558_ (.A1(_02491_),
    .A2(_02492_),
    .Y(_02495_),
    .B1(_02490_));
 sg13g2_xor2_1 _09559_ (.B(net2191),
    .A(net2474),
    .X(_02496_));
 sg13g2_xnor2_1 _09560_ (.Y(_02497_),
    .A(_02495_),
    .B(_02496_));
 sg13g2_o21ai_1 _09561_ (.B1(net2017),
    .Y(_02498_),
    .A1(net1857),
    .A2(net1332));
 sg13g2_a21oi_1 _09562_ (.A1(net1857),
    .A2(net2475),
    .Y(_00311_),
    .B1(_02498_));
 sg13g2_o21ai_1 _09563_ (.B1(net1986),
    .Y(_02499_),
    .A1(net1839),
    .A2(\am_sdr0.cic3.comb3_in_del[0] ));
 sg13g2_a21oi_1 _09564_ (.A1(net1839),
    .A2(_01506_),
    .Y(_00312_),
    .B1(_02499_));
 sg13g2_o21ai_1 _09565_ (.B1(net1986),
    .Y(_02500_),
    .A1(net1839),
    .A2(\am_sdr0.cic3.comb3_in_del[1] ));
 sg13g2_a21oi_1 _09566_ (.A1(net1841),
    .A2(_01505_),
    .Y(_00313_),
    .B1(_02500_));
 sg13g2_o21ai_1 _09567_ (.B1(net1986),
    .Y(_02501_),
    .A1(net1622),
    .A2(\am_sdr0.cic3.comb2[2] ));
 sg13g2_a21oi_1 _09568_ (.A1(net1622),
    .A2(_01504_),
    .Y(_00314_),
    .B1(_02501_));
 sg13g2_o21ai_1 _09569_ (.B1(net1987),
    .Y(_02502_),
    .A1(net1839),
    .A2(net2215));
 sg13g2_a21oi_1 _09570_ (.A1(net1841),
    .A2(_01503_),
    .Y(_00315_),
    .B1(_02502_));
 sg13g2_o21ai_1 _09571_ (.B1(net1987),
    .Y(_02503_),
    .A1(net1840),
    .A2(\am_sdr0.cic3.comb3_in_del[4] ));
 sg13g2_a21oi_1 _09572_ (.A1(net1840),
    .A2(_01501_),
    .Y(_00316_),
    .B1(_02503_));
 sg13g2_o21ai_1 _09573_ (.B1(net1986),
    .Y(_02504_),
    .A1(net1840),
    .A2(\am_sdr0.cic3.comb3_in_del[5] ));
 sg13g2_a21oi_1 _09574_ (.A1(net1840),
    .A2(_01499_),
    .Y(_00317_),
    .B1(_02504_));
 sg13g2_o21ai_1 _09575_ (.B1(net1989),
    .Y(_02505_),
    .A1(net1623),
    .A2(\am_sdr0.cic3.comb2[6] ));
 sg13g2_a21oi_1 _09576_ (.A1(net1623),
    .A2(_01497_),
    .Y(_00318_),
    .B1(_02505_));
 sg13g2_o21ai_1 _09577_ (.B1(net1990),
    .Y(_02506_),
    .A1(net1848),
    .A2(net2155));
 sg13g2_a21oi_1 _09578_ (.A1(net1848),
    .A2(_01496_),
    .Y(_00319_),
    .B1(_02506_));
 sg13g2_o21ai_1 _09579_ (.B1(net1989),
    .Y(_02507_),
    .A1(net1623),
    .A2(\am_sdr0.cic3.comb2[8] ));
 sg13g2_a21oi_1 _09580_ (.A1(net1623),
    .A2(_01494_),
    .Y(_00320_),
    .B1(_02507_));
 sg13g2_o21ai_1 _09581_ (.B1(net1989),
    .Y(_02508_),
    .A1(net1624),
    .A2(\am_sdr0.cic3.comb2[9] ));
 sg13g2_a21oi_1 _09582_ (.A1(net1624),
    .A2(_01493_),
    .Y(_00321_),
    .B1(_02508_));
 sg13g2_o21ai_1 _09583_ (.B1(net1998),
    .Y(_02509_),
    .A1(net1846),
    .A2(net2294));
 sg13g2_a21oi_1 _09584_ (.A1(net1846),
    .A2(_01492_),
    .Y(_00322_),
    .B1(_02509_));
 sg13g2_o21ai_1 _09585_ (.B1(net1998),
    .Y(_02510_),
    .A1(net1846),
    .A2(\am_sdr0.cic3.comb3_in_del[11] ));
 sg13g2_a21oi_1 _09586_ (.A1(net1846),
    .A2(_01490_),
    .Y(_00323_),
    .B1(_02510_));
 sg13g2_o21ai_1 _09587_ (.B1(net2000),
    .Y(_02511_),
    .A1(net1862),
    .A2(\am_sdr0.cic3.comb3_in_del[12] ));
 sg13g2_a21oi_1 _09588_ (.A1(net1862),
    .A2(_01488_),
    .Y(_00324_),
    .B1(_02511_));
 sg13g2_o21ai_1 _09589_ (.B1(net2000),
    .Y(_02512_),
    .A1(net1862),
    .A2(net2837));
 sg13g2_a21oi_1 _09590_ (.A1(net1862),
    .A2(_01487_),
    .Y(_00325_),
    .B1(_02512_));
 sg13g2_o21ai_1 _09591_ (.B1(net2000),
    .Y(_02513_),
    .A1(net1865),
    .A2(net2438));
 sg13g2_a21oi_1 _09592_ (.A1(net1865),
    .A2(_01486_),
    .Y(_00326_),
    .B1(_02513_));
 sg13g2_o21ai_1 _09593_ (.B1(net2000),
    .Y(_02514_),
    .A1(net1866),
    .A2(net2285));
 sg13g2_a21oi_1 _09594_ (.A1(net1866),
    .A2(_01485_),
    .Y(_00327_),
    .B1(_02514_));
 sg13g2_o21ai_1 _09595_ (.B1(net1999),
    .Y(_02515_),
    .A1(net1865),
    .A2(\am_sdr0.cic3.comb3_in_del[16] ));
 sg13g2_a21oi_1 _09596_ (.A1(net1865),
    .A2(_01484_),
    .Y(_00328_),
    .B1(_02515_));
 sg13g2_o21ai_1 _09597_ (.B1(net2022),
    .Y(_02516_),
    .A1(net1856),
    .A2(\am_sdr0.cic3.comb3_in_del[17] ));
 sg13g2_a21oi_1 _09598_ (.A1(net1856),
    .A2(_01483_),
    .Y(_00329_),
    .B1(_02516_));
 sg13g2_o21ai_1 _09599_ (.B1(net2017),
    .Y(_02517_),
    .A1(net1856),
    .A2(net2623));
 sg13g2_a21oi_1 _09600_ (.A1(net1856),
    .A2(_01482_),
    .Y(_00330_),
    .B1(_02517_));
 sg13g2_o21ai_1 _09601_ (.B1(net2017),
    .Y(_02518_),
    .A1(\am_sdr0.cic3.comb3_in_del[19] ),
    .A2(net1855));
 sg13g2_a21oi_1 _09602_ (.A1(_01480_),
    .A2(net1855),
    .Y(_00331_),
    .B1(_02518_));
 sg13g2_o21ai_1 _09603_ (.B1(net1968),
    .Y(_02519_),
    .A1(net1737),
    .A2(net1490));
 sg13g2_a21oi_1 _09604_ (.A1(net1737),
    .A2(net1490),
    .Y(_00332_),
    .B1(_02519_));
 sg13g2_a21oi_1 _09605_ (.A1(net1739),
    .A2(\am_sdr0.cic3.count[0] ),
    .Y(_02520_),
    .B1(net1243));
 sg13g2_nand2_1 _09606_ (.Y(_02521_),
    .A(net1966),
    .B(_02121_));
 sg13g2_nor2_1 _09607_ (.A(net1244),
    .B(_02521_),
    .Y(_00333_));
 sg13g2_a21oi_1 _09608_ (.A1(_01479_),
    .A2(_02121_),
    .Y(_02522_),
    .B1(net1889));
 sg13g2_nor2b_1 _09609_ (.A(_02122_),
    .B_N(_02522_),
    .Y(_00334_));
 sg13g2_o21ai_1 _09610_ (.B1(net1967),
    .Y(_02523_),
    .A1(net2591),
    .A2(_02122_));
 sg13g2_nor2_1 _09611_ (.A(_02123_),
    .B(net2592),
    .Y(_00335_));
 sg13g2_o21ai_1 _09612_ (.B1(net1967),
    .Y(_02524_),
    .A1(net2601),
    .A2(_02123_));
 sg13g2_nor2_1 _09613_ (.A(_02124_),
    .B(_02524_),
    .Y(_00336_));
 sg13g2_o21ai_1 _09614_ (.B1(net1968),
    .Y(_02525_),
    .A1(net2861),
    .A2(_02124_));
 sg13g2_nor2b_1 _09615_ (.A(_02525_),
    .B_N(_02125_),
    .Y(_00337_));
 sg13g2_a21oi_1 _09616_ (.A1(\am_sdr0.cic3.count[5] ),
    .A2(_02124_),
    .Y(_02526_),
    .B1(net2094));
 sg13g2_and3_1 _09617_ (.X(_02527_),
    .A(net2094),
    .B(\am_sdr0.cic3.count[5] ),
    .C(_02124_));
 sg13g2_nor4_1 _09618_ (.A(net1889),
    .B(_02126_),
    .C(net2095),
    .D(_02527_),
    .Y(_00338_));
 sg13g2_o21ai_1 _09619_ (.B1(net1968),
    .Y(_02528_),
    .A1(net1375),
    .A2(_02527_));
 sg13g2_a21oi_1 _09620_ (.A1(net1375),
    .A2(_02527_),
    .Y(_00339_),
    .B1(_02528_));
 sg13g2_a21oi_1 _09621_ (.A1(\am_sdr0.cic1.x_out[8] ),
    .A2(net1737),
    .Y(_02529_),
    .B1(net1277));
 sg13g2_nand2_1 _09622_ (.Y(_02530_),
    .A(\am_sdr0.cic1.x_out[8] ),
    .B(net1277));
 sg13g2_nor2_1 _09623_ (.A(net1627),
    .B(_02530_),
    .Y(_02531_));
 sg13g2_nor3_1 _09624_ (.A(net1888),
    .B(net1278),
    .C(_02531_),
    .Y(_00340_));
 sg13g2_nand2_1 _09625_ (.Y(_02532_),
    .A(\am_sdr0.cic1.x_out[9] ),
    .B(net3299));
 sg13g2_xnor2_1 _09626_ (.Y(_02533_),
    .A(\am_sdr0.cic1.x_out[9] ),
    .B(net2805));
 sg13g2_xnor2_1 _09627_ (.Y(_02534_),
    .A(_02530_),
    .B(_02533_));
 sg13g2_o21ai_1 _09628_ (.B1(net1965),
    .Y(_02535_),
    .A1(net1737),
    .A2(net2805));
 sg13g2_a21oi_1 _09629_ (.A1(net1737),
    .A2(_02534_),
    .Y(_00341_),
    .B1(_02535_));
 sg13g2_and2_1 _09630_ (.A(\am_sdr0.cic1.x_out[10] ),
    .B(\am_sdr0.cic3.integ1[2] ),
    .X(_02536_));
 sg13g2_xor2_1 _09631_ (.B(net2699),
    .A(\am_sdr0.cic1.x_out[10] ),
    .X(_02537_));
 sg13g2_o21ai_1 _09632_ (.B1(_02532_),
    .Y(_02538_),
    .A1(_02530_),
    .A2(_02533_));
 sg13g2_xnor2_1 _09633_ (.Y(_02539_),
    .A(_02537_),
    .B(_02538_));
 sg13g2_o21ai_1 _09634_ (.B1(net1965),
    .Y(_02540_),
    .A1(net1735),
    .A2(net2699));
 sg13g2_a21oi_1 _09635_ (.A1(net1735),
    .A2(_02539_),
    .Y(_00342_),
    .B1(_02540_));
 sg13g2_nand2_1 _09636_ (.Y(_02541_),
    .A(\am_sdr0.cic1.x_out[11] ),
    .B(\am_sdr0.cic3.integ1[3] ));
 sg13g2_xnor2_1 _09637_ (.Y(_02542_),
    .A(\am_sdr0.cic1.x_out[11] ),
    .B(\am_sdr0.cic3.integ1[3] ));
 sg13g2_a21oi_1 _09638_ (.A1(_02537_),
    .A2(_02538_),
    .Y(_02543_),
    .B1(_02536_));
 sg13g2_xnor2_1 _09639_ (.Y(_02544_),
    .A(_02542_),
    .B(_02543_));
 sg13g2_o21ai_1 _09640_ (.B1(net1962),
    .Y(_02545_),
    .A1(net1735),
    .A2(net3035));
 sg13g2_a21oi_1 _09641_ (.A1(net1735),
    .A2(_02544_),
    .Y(_00343_),
    .B1(_02545_));
 sg13g2_o21ai_1 _09642_ (.B1(_02541_),
    .Y(_02546_),
    .A1(_02542_),
    .A2(_02543_));
 sg13g2_nand2_1 _09643_ (.Y(_02547_),
    .A(\am_sdr0.cic1.x_out[12] ),
    .B(\am_sdr0.cic3.integ1[4] ));
 sg13g2_xor2_1 _09644_ (.B(\am_sdr0.cic3.integ1[4] ),
    .A(\am_sdr0.cic1.x_out[12] ),
    .X(_02548_));
 sg13g2_nand2_1 _09645_ (.Y(_02549_),
    .A(_02546_),
    .B(_02548_));
 sg13g2_xnor2_1 _09646_ (.Y(_02550_),
    .A(_02546_),
    .B(_02548_));
 sg13g2_o21ai_1 _09647_ (.B1(net1962),
    .Y(_02551_),
    .A1(net1736),
    .A2(net3132));
 sg13g2_a21oi_1 _09648_ (.A1(net1736),
    .A2(_02550_),
    .Y(_00344_),
    .B1(_02551_));
 sg13g2_nor2_1 _09649_ (.A(\am_sdr0.cic1.x_out[13] ),
    .B(\am_sdr0.cic3.integ1[5] ),
    .Y(_02552_));
 sg13g2_and2_1 _09650_ (.A(\am_sdr0.cic1.x_out[13] ),
    .B(\am_sdr0.cic3.integ1[5] ),
    .X(_02553_));
 sg13g2_nor2_1 _09651_ (.A(_02552_),
    .B(_02553_),
    .Y(_02554_));
 sg13g2_nand2_1 _09652_ (.Y(_02555_),
    .A(_02547_),
    .B(_02549_));
 sg13g2_xnor2_1 _09653_ (.Y(_02556_),
    .A(_02554_),
    .B(_02555_));
 sg13g2_o21ai_1 _09654_ (.B1(net1962),
    .Y(_02557_),
    .A1(net1736),
    .A2(net2966));
 sg13g2_a21oi_1 _09655_ (.A1(net1736),
    .A2(_02556_),
    .Y(_00345_),
    .B1(_02557_));
 sg13g2_nand2_1 _09656_ (.Y(_02558_),
    .A(\am_sdr0.cic1.x_out[14] ),
    .B(\am_sdr0.cic3.integ1[6] ));
 sg13g2_or2_1 _09657_ (.X(_02559_),
    .B(\am_sdr0.cic3.integ1[6] ),
    .A(\am_sdr0.cic1.x_out[14] ));
 sg13g2_nand2_1 _09658_ (.Y(_02560_),
    .A(_02558_),
    .B(_02559_));
 sg13g2_a21oi_1 _09659_ (.A1(\am_sdr0.cic1.x_out[12] ),
    .A2(\am_sdr0.cic3.integ1[4] ),
    .Y(_02561_),
    .B1(_02553_));
 sg13g2_and2_1 _09660_ (.A(_02548_),
    .B(_02554_),
    .X(_02562_));
 sg13g2_nor2_1 _09661_ (.A(_02547_),
    .B(_02552_),
    .Y(_02563_));
 sg13g2_a21oi_1 _09662_ (.A1(_02549_),
    .A2(_02561_),
    .Y(_02564_),
    .B1(_02552_));
 sg13g2_nand2b_1 _09663_ (.Y(_02565_),
    .B(_02564_),
    .A_N(_02560_));
 sg13g2_xor2_1 _09664_ (.B(_02564_),
    .A(_02560_),
    .X(_02566_));
 sg13g2_o21ai_1 _09665_ (.B1(net1966),
    .Y(_02567_),
    .A1(net1736),
    .A2(net2935));
 sg13g2_a21oi_1 _09666_ (.A1(net1736),
    .A2(_02566_),
    .Y(_00346_),
    .B1(_02567_));
 sg13g2_and2_1 _09667_ (.A(net1758),
    .B(\am_sdr0.cic3.integ1[7] ),
    .X(_02568_));
 sg13g2_nor2_1 _09668_ (.A(net1758),
    .B(\am_sdr0.cic3.integ1[7] ),
    .Y(_02569_));
 sg13g2_inv_1 _09669_ (.Y(_02570_),
    .A(_02569_));
 sg13g2_nand2_1 _09670_ (.Y(_02571_),
    .A(_02558_),
    .B(_02565_));
 sg13g2_o21ai_1 _09671_ (.B1(_02571_),
    .Y(_02572_),
    .A1(_02568_),
    .A2(_02569_));
 sg13g2_nor3_1 _09672_ (.A(_02568_),
    .B(_02569_),
    .C(_02571_),
    .Y(_02573_));
 sg13g2_nor2_1 _09673_ (.A(net1627),
    .B(_02573_),
    .Y(_02574_));
 sg13g2_o21ai_1 _09674_ (.B1(net1966),
    .Y(_02575_),
    .A1(net1738),
    .A2(net3111));
 sg13g2_a21oi_1 _09675_ (.A1(_02572_),
    .A2(_02574_),
    .Y(_00347_),
    .B1(_02575_));
 sg13g2_nor2_1 _09676_ (.A(_02558_),
    .B(_02569_),
    .Y(_02576_));
 sg13g2_or4_1 _09677_ (.A(_02553_),
    .B(_02563_),
    .C(_02568_),
    .D(_02576_),
    .X(_02577_));
 sg13g2_a21oi_1 _09678_ (.A1(_02546_),
    .A2(_02562_),
    .Y(_02578_),
    .B1(_02577_));
 sg13g2_o21ai_1 _09679_ (.B1(_02570_),
    .Y(_02579_),
    .A1(_02559_),
    .A2(_02568_));
 sg13g2_or2_1 _09680_ (.X(_02580_),
    .B(_02579_),
    .A(_02578_));
 sg13g2_xor2_1 _09681_ (.B(\am_sdr0.cic3.integ1[8] ),
    .A(net1756),
    .X(_02581_));
 sg13g2_nand2b_1 _09682_ (.Y(_02582_),
    .B(_02581_),
    .A_N(_02580_));
 sg13g2_xor2_1 _09683_ (.B(_02581_),
    .A(_02580_),
    .X(_02583_));
 sg13g2_o21ai_1 _09684_ (.B1(net1966),
    .Y(_02584_),
    .A1(net1738),
    .A2(net3089));
 sg13g2_a21oi_1 _09685_ (.A1(net1738),
    .A2(_02583_),
    .Y(_00348_),
    .B1(_02584_));
 sg13g2_xor2_1 _09686_ (.B(\am_sdr0.cic3.integ1[9] ),
    .A(net1756),
    .X(_02585_));
 sg13g2_inv_1 _09687_ (.Y(_02586_),
    .A(_02585_));
 sg13g2_o21ai_1 _09688_ (.B1(_02582_),
    .Y(_02587_),
    .A1(_01383_),
    .A2(_01478_));
 sg13g2_xnor2_1 _09689_ (.Y(_02588_),
    .A(_02585_),
    .B(_02587_));
 sg13g2_o21ai_1 _09690_ (.B1(net1967),
    .Y(_02589_),
    .A1(net1740),
    .A2(net3054));
 sg13g2_a21oi_1 _09691_ (.A1(net1740),
    .A2(_02588_),
    .Y(_00349_),
    .B1(_02589_));
 sg13g2_and2_1 _09692_ (.A(net1756),
    .B(\am_sdr0.cic3.integ1[10] ),
    .X(_02590_));
 sg13g2_xor2_1 _09693_ (.B(\am_sdr0.cic3.integ1[10] ),
    .A(net1756),
    .X(_02591_));
 sg13g2_o21ai_1 _09694_ (.B1(net1756),
    .Y(_02592_),
    .A1(\am_sdr0.cic3.integ1[9] ),
    .A2(\am_sdr0.cic3.integ1[8] ));
 sg13g2_o21ai_1 _09695_ (.B1(_02592_),
    .Y(_02593_),
    .A1(_02582_),
    .A2(_02586_));
 sg13g2_xnor2_1 _09696_ (.Y(_02594_),
    .A(_02591_),
    .B(_02593_));
 sg13g2_o21ai_1 _09697_ (.B1(net1969),
    .Y(_02595_),
    .A1(net1740),
    .A2(net3062));
 sg13g2_a21oi_1 _09698_ (.A1(net1740),
    .A2(_02594_),
    .Y(_00350_),
    .B1(_02595_));
 sg13g2_a21oi_1 _09699_ (.A1(_02591_),
    .A2(_02593_),
    .Y(_02596_),
    .B1(_02590_));
 sg13g2_xor2_1 _09700_ (.B(\am_sdr0.cic3.integ1[11] ),
    .A(net1756),
    .X(_02597_));
 sg13g2_xor2_1 _09701_ (.B(_02597_),
    .A(_02596_),
    .X(_02598_));
 sg13g2_o21ai_1 _09702_ (.B1(net1969),
    .Y(_02599_),
    .A1(net1741),
    .A2(net3078));
 sg13g2_a21oi_1 _09703_ (.A1(net1741),
    .A2(_02598_),
    .Y(_00351_),
    .B1(_02599_));
 sg13g2_xor2_1 _09704_ (.B(\am_sdr0.cic3.integ1[12] ),
    .A(net1757),
    .X(_02600_));
 sg13g2_nand4_1 _09705_ (.B(_02585_),
    .C(_02591_),
    .A(_02581_),
    .Y(_02601_),
    .D(_02597_));
 sg13g2_nor3_1 _09706_ (.A(_02578_),
    .B(_02579_),
    .C(_02601_),
    .Y(_02602_));
 sg13g2_o21ai_1 _09707_ (.B1(net1756),
    .Y(_02603_),
    .A1(\am_sdr0.cic3.integ1[11] ),
    .A2(\am_sdr0.cic3.integ1[10] ));
 sg13g2_and2_1 _09708_ (.A(_02592_),
    .B(_02603_),
    .X(_02604_));
 sg13g2_nand2b_1 _09709_ (.Y(_02605_),
    .B(_02604_),
    .A_N(_02602_));
 sg13g2_and2_1 _09710_ (.A(_02600_),
    .B(_02605_),
    .X(_02606_));
 sg13g2_xnor2_1 _09711_ (.Y(_02607_),
    .A(_02600_),
    .B(_02605_));
 sg13g2_o21ai_1 _09712_ (.B1(net1969),
    .Y(_02608_),
    .A1(net1740),
    .A2(net3053));
 sg13g2_a21oi_1 _09713_ (.A1(net1740),
    .A2(_02607_),
    .Y(_00352_),
    .B1(_02608_));
 sg13g2_xor2_1 _09714_ (.B(\am_sdr0.cic3.integ1[13] ),
    .A(net1757),
    .X(_02609_));
 sg13g2_a21oi_1 _09715_ (.A1(net1757),
    .A2(\am_sdr0.cic3.integ1[12] ),
    .Y(_02610_),
    .B1(_02606_));
 sg13g2_xor2_1 _09716_ (.B(_02610_),
    .A(_02609_),
    .X(_02611_));
 sg13g2_o21ai_1 _09717_ (.B1(net1967),
    .Y(_02612_),
    .A1(net1742),
    .A2(net3091));
 sg13g2_a21oi_1 _09718_ (.A1(net1743),
    .A2(_02611_),
    .Y(_00353_),
    .B1(_02612_));
 sg13g2_nand2_1 _09719_ (.Y(_02613_),
    .A(net1757),
    .B(\am_sdr0.cic3.integ1[14] ));
 sg13g2_xnor2_1 _09720_ (.Y(_02614_),
    .A(net1757),
    .B(\am_sdr0.cic3.integ1[14] ));
 sg13g2_o21ai_1 _09721_ (.B1(net1757),
    .Y(_02615_),
    .A1(\am_sdr0.cic3.integ1[13] ),
    .A2(\am_sdr0.cic3.integ1[12] ));
 sg13g2_inv_1 _09722_ (.Y(_02616_),
    .A(_02615_));
 sg13g2_a21oi_1 _09723_ (.A1(_02606_),
    .A2(_02609_),
    .Y(_02617_),
    .B1(_02616_));
 sg13g2_xnor2_1 _09724_ (.Y(_02618_),
    .A(_02614_),
    .B(_02617_));
 sg13g2_o21ai_1 _09725_ (.B1(net1967),
    .Y(_02619_),
    .A1(net1742),
    .A2(net3152));
 sg13g2_a21oi_1 _09726_ (.A1(net1742),
    .A2(_02618_),
    .Y(_00354_),
    .B1(_02619_));
 sg13g2_xnor2_1 _09727_ (.Y(_02620_),
    .A(net1757),
    .B(\am_sdr0.cic3.integ1[15] ));
 sg13g2_o21ai_1 _09728_ (.B1(_02613_),
    .Y(_02621_),
    .A1(_02614_),
    .A2(_02617_));
 sg13g2_or2_1 _09729_ (.X(_02622_),
    .B(_02621_),
    .A(_02620_));
 sg13g2_a21oi_1 _09730_ (.A1(_02620_),
    .A2(_02621_),
    .Y(_02623_),
    .B1(net1626));
 sg13g2_o21ai_1 _09731_ (.B1(net1969),
    .Y(_02624_),
    .A1(net1742),
    .A2(net3127));
 sg13g2_a21oi_1 _09732_ (.A1(_02622_),
    .A2(_02623_),
    .Y(_00355_),
    .B1(_02624_));
 sg13g2_nand2_1 _09733_ (.Y(_02625_),
    .A(_02600_),
    .B(_02609_));
 sg13g2_nor3_1 _09734_ (.A(_02614_),
    .B(_02620_),
    .C(_02625_),
    .Y(_02626_));
 sg13g2_o21ai_1 _09735_ (.B1(net1757),
    .Y(_02627_),
    .A1(\am_sdr0.cic3.integ1[15] ),
    .A2(\am_sdr0.cic3.integ1[14] ));
 sg13g2_nand3_1 _09736_ (.B(_02615_),
    .C(_02627_),
    .A(_02604_),
    .Y(_02628_));
 sg13g2_a21oi_2 _09737_ (.B1(_02628_),
    .Y(_02629_),
    .A2(_02626_),
    .A1(_02602_));
 sg13g2_xnor2_1 _09738_ (.Y(_02630_),
    .A(net1759),
    .B(\am_sdr0.cic3.integ1[16] ));
 sg13g2_nor2_1 _09739_ (.A(_02629_),
    .B(_02630_),
    .Y(_02631_));
 sg13g2_inv_1 _09740_ (.Y(_02632_),
    .A(_02631_));
 sg13g2_xnor2_1 _09741_ (.Y(_02633_),
    .A(_02629_),
    .B(_02630_));
 sg13g2_o21ai_1 _09742_ (.B1(net1968),
    .Y(_02634_),
    .A1(net1743),
    .A2(net3055));
 sg13g2_a21oi_1 _09743_ (.A1(net1743),
    .A2(_02633_),
    .Y(_00356_),
    .B1(_02634_));
 sg13g2_xnor2_1 _09744_ (.Y(_02635_),
    .A(net1761),
    .B(\am_sdr0.cic3.integ1[17] ));
 sg13g2_a21oi_1 _09745_ (.A1(net1759),
    .A2(\am_sdr0.cic3.integ1[16] ),
    .Y(_02636_),
    .B1(_02631_));
 sg13g2_xnor2_1 _09746_ (.Y(_02637_),
    .A(_02635_),
    .B(_02636_));
 sg13g2_o21ai_1 _09747_ (.B1(net1969),
    .Y(_02638_),
    .A1(net1742),
    .A2(net3050));
 sg13g2_a21oi_1 _09748_ (.A1(net1742),
    .A2(_02637_),
    .Y(_00357_),
    .B1(_02638_));
 sg13g2_or2_1 _09749_ (.X(_02639_),
    .B(\am_sdr0.cic3.integ1[18] ),
    .A(net1759));
 sg13g2_and2_1 _09750_ (.A(net1759),
    .B(\am_sdr0.cic3.integ1[18] ),
    .X(_02640_));
 sg13g2_xnor2_1 _09751_ (.Y(_02641_),
    .A(net1759),
    .B(\am_sdr0.cic3.integ1[18] ));
 sg13g2_o21ai_1 _09752_ (.B1(net1759),
    .Y(_02642_),
    .A1(\am_sdr0.cic3.integ1[17] ),
    .A2(\am_sdr0.cic3.integ1[16] ));
 sg13g2_o21ai_1 _09753_ (.B1(_02642_),
    .Y(_02643_),
    .A1(_02632_),
    .A2(_02635_));
 sg13g2_xor2_1 _09754_ (.B(_02643_),
    .A(_02641_),
    .X(_02644_));
 sg13g2_o21ai_1 _09755_ (.B1(net1969),
    .Y(_02645_),
    .A1(net1742),
    .A2(net3154));
 sg13g2_a21oi_1 _09756_ (.A1(net1742),
    .A2(_02644_),
    .Y(_00358_),
    .B1(_02645_));
 sg13g2_xnor2_1 _09757_ (.Y(_02646_),
    .A(net1759),
    .B(\am_sdr0.cic3.integ1[19] ));
 sg13g2_a21oi_1 _09758_ (.A1(_02639_),
    .A2(_02643_),
    .Y(_02647_),
    .B1(_02640_));
 sg13g2_xnor2_1 _09759_ (.Y(_02648_),
    .A(_02646_),
    .B(_02647_));
 sg13g2_o21ai_1 _09760_ (.B1(net1968),
    .Y(_02649_),
    .A1(net1749),
    .A2(net3039));
 sg13g2_a21oi_1 _09761_ (.A1(net1749),
    .A2(_02648_),
    .Y(_00359_),
    .B1(_02649_));
 sg13g2_xor2_1 _09762_ (.B(\am_sdr0.cic3.integ1[20] ),
    .A(net1760),
    .X(_02650_));
 sg13g2_nor4_1 _09763_ (.A(_02630_),
    .B(_02635_),
    .C(_02641_),
    .D(_02646_),
    .Y(_02651_));
 sg13g2_nor2b_2 _09764_ (.A(_02629_),
    .B_N(_02651_),
    .Y(_02652_));
 sg13g2_o21ai_1 _09765_ (.B1(net1759),
    .Y(_02653_),
    .A1(\am_sdr0.cic3.integ1[19] ),
    .A2(\am_sdr0.cic3.integ1[18] ));
 sg13g2_and2_1 _09766_ (.A(_02642_),
    .B(_02653_),
    .X(_02654_));
 sg13g2_inv_1 _09767_ (.Y(_02655_),
    .A(_02654_));
 sg13g2_nor3_1 _09768_ (.A(_02650_),
    .B(_02652_),
    .C(_02655_),
    .Y(_02656_));
 sg13g2_o21ai_1 _09769_ (.B1(_02650_),
    .Y(_02657_),
    .A1(_02652_),
    .A2(_02655_));
 sg13g2_nor2b_1 _09770_ (.A(_02656_),
    .B_N(_02657_),
    .Y(_02658_));
 sg13g2_o21ai_1 _09771_ (.B1(net1976),
    .Y(_02659_),
    .A1(net1627),
    .A2(_02658_));
 sg13g2_a21oi_1 _09772_ (.A1(net1627),
    .A2(_01477_),
    .Y(_00360_),
    .B1(_02659_));
 sg13g2_xor2_1 _09773_ (.B(\am_sdr0.cic3.integ1[21] ),
    .A(net1760),
    .X(_02660_));
 sg13g2_inv_1 _09774_ (.Y(_02661_),
    .A(_02660_));
 sg13g2_o21ai_1 _09775_ (.B1(_02657_),
    .Y(_02662_),
    .A1(_01383_),
    .A2(_01477_));
 sg13g2_xnor2_1 _09776_ (.Y(_02663_),
    .A(_02660_),
    .B(_02662_));
 sg13g2_o21ai_1 _09777_ (.B1(net1979),
    .Y(_02664_),
    .A1(net1750),
    .A2(net3052));
 sg13g2_a21oi_1 _09778_ (.A1(net1749),
    .A2(_02663_),
    .Y(_00361_),
    .B1(_02664_));
 sg13g2_or2_1 _09779_ (.X(_02665_),
    .B(\am_sdr0.cic3.integ1[22] ),
    .A(net1760));
 sg13g2_and2_1 _09780_ (.A(net1760),
    .B(\am_sdr0.cic3.integ1[22] ),
    .X(_02666_));
 sg13g2_xnor2_1 _09781_ (.Y(_02667_),
    .A(net1760),
    .B(\am_sdr0.cic3.integ1[22] ));
 sg13g2_o21ai_1 _09782_ (.B1(net1760),
    .Y(_02668_),
    .A1(\am_sdr0.cic3.integ1[21] ),
    .A2(\am_sdr0.cic3.integ1[20] ));
 sg13g2_o21ai_1 _09783_ (.B1(_02668_),
    .Y(_02669_),
    .A1(_02657_),
    .A2(_02661_));
 sg13g2_xor2_1 _09784_ (.B(_02669_),
    .A(_02667_),
    .X(_02670_));
 sg13g2_o21ai_1 _09785_ (.B1(net1976),
    .Y(_02671_),
    .A1(net1749),
    .A2(net3195));
 sg13g2_a21oi_1 _09786_ (.A1(net1749),
    .A2(_02670_),
    .Y(_00362_),
    .B1(_02671_));
 sg13g2_xnor2_1 _09787_ (.Y(_02672_),
    .A(net1760),
    .B(\am_sdr0.cic3.integ1[23] ));
 sg13g2_a21oi_1 _09788_ (.A1(_02665_),
    .A2(_02669_),
    .Y(_02673_),
    .B1(_02666_));
 sg13g2_xnor2_1 _09789_ (.Y(_02674_),
    .A(_02672_),
    .B(_02673_));
 sg13g2_o21ai_1 _09790_ (.B1(net1976),
    .Y(_02675_),
    .A1(net1749),
    .A2(net3000));
 sg13g2_a21oi_1 _09791_ (.A1(net1749),
    .A2(_02674_),
    .Y(_00363_),
    .B1(_02675_));
 sg13g2_nand2_1 _09792_ (.Y(_02676_),
    .A(_02650_),
    .B(_02660_));
 sg13g2_nor3_1 _09793_ (.A(_02667_),
    .B(_02672_),
    .C(_02676_),
    .Y(_02677_));
 sg13g2_o21ai_1 _09794_ (.B1(net1760),
    .Y(_02678_),
    .A1(\am_sdr0.cic3.integ1[23] ),
    .A2(\am_sdr0.cic3.integ1[22] ));
 sg13g2_nand3_1 _09795_ (.B(_02668_),
    .C(_02678_),
    .A(_02654_),
    .Y(_02679_));
 sg13g2_a21oi_2 _09796_ (.B1(_02679_),
    .Y(_02680_),
    .A2(_02677_),
    .A1(_02652_));
 sg13g2_xnor2_1 _09797_ (.Y(_02681_),
    .A(net1761),
    .B(\am_sdr0.cic3.integ1[24] ));
 sg13g2_xnor2_1 _09798_ (.Y(_02682_),
    .A(_02680_),
    .B(_02681_));
 sg13g2_o21ai_1 _09799_ (.B1(net1976),
    .Y(_02683_),
    .A1(net1750),
    .A2(net3138));
 sg13g2_a21oi_1 _09800_ (.A1(net1750),
    .A2(_02682_),
    .Y(_00364_),
    .B1(_02683_));
 sg13g2_a21o_1 _09801_ (.A2(\am_sdr0.cic3.integ1[24] ),
    .A1(_01383_),
    .B1(_02680_),
    .X(_02684_));
 sg13g2_o21ai_1 _09802_ (.B1(_02680_),
    .Y(_02685_),
    .A1(_01383_),
    .A2(\am_sdr0.cic3.integ1[24] ));
 sg13g2_and3_1 _09803_ (.X(_02686_),
    .A(net1750),
    .B(_02684_),
    .C(_02685_));
 sg13g2_o21ai_1 _09804_ (.B1(net1979),
    .Y(_02687_),
    .A1(net1297),
    .A2(_02686_));
 sg13g2_a21oi_1 _09805_ (.A1(net1297),
    .A2(_02686_),
    .Y(_00365_),
    .B1(_02687_));
 sg13g2_a21oi_1 _09806_ (.A1(net1735),
    .A2(\am_sdr0.cic3.integ1[3] ),
    .Y(_02688_),
    .B1(net1321));
 sg13g2_nand2_1 _09807_ (.Y(_02689_),
    .A(net1321),
    .B(\am_sdr0.cic3.integ1[3] ));
 sg13g2_nor2_1 _09808_ (.A(net1627),
    .B(_02689_),
    .Y(_02690_));
 sg13g2_nor3_1 _09809_ (.A(net1888),
    .B(net1322),
    .C(_02690_),
    .Y(_00366_));
 sg13g2_nand2_1 _09810_ (.Y(_02691_),
    .A(\am_sdr0.cic3.integ2[1] ),
    .B(\am_sdr0.cic3.integ1[4] ));
 sg13g2_xnor2_1 _09811_ (.Y(_02692_),
    .A(net2741),
    .B(\am_sdr0.cic3.integ1[4] ));
 sg13g2_xnor2_1 _09812_ (.Y(_02693_),
    .A(_02689_),
    .B(_02692_));
 sg13g2_o21ai_1 _09813_ (.B1(net1962),
    .Y(_02694_),
    .A1(net1735),
    .A2(net2741));
 sg13g2_a21oi_1 _09814_ (.A1(net1735),
    .A2(_02693_),
    .Y(_00367_),
    .B1(_02694_));
 sg13g2_and2_1 _09815_ (.A(\am_sdr0.cic3.integ2[2] ),
    .B(\am_sdr0.cic3.integ1[5] ),
    .X(_02695_));
 sg13g2_xor2_1 _09816_ (.B(\am_sdr0.cic3.integ1[5] ),
    .A(net2652),
    .X(_02696_));
 sg13g2_o21ai_1 _09817_ (.B1(_02691_),
    .Y(_02697_),
    .A1(_02689_),
    .A2(_02692_));
 sg13g2_and2_1 _09818_ (.A(_02696_),
    .B(_02697_),
    .X(_02698_));
 sg13g2_xnor2_1 _09819_ (.Y(_02699_),
    .A(_02696_),
    .B(_02697_));
 sg13g2_o21ai_1 _09820_ (.B1(net1962),
    .Y(_02700_),
    .A1(net1736),
    .A2(net2652));
 sg13g2_a21oi_1 _09821_ (.A1(net1735),
    .A2(_02699_),
    .Y(_00368_),
    .B1(_02700_));
 sg13g2_nand2_1 _09822_ (.Y(_02701_),
    .A(\am_sdr0.cic3.integ2[3] ),
    .B(net2935));
 sg13g2_xor2_1 _09823_ (.B(\am_sdr0.cic3.integ1[6] ),
    .A(\am_sdr0.cic3.integ2[3] ),
    .X(_02702_));
 sg13g2_nor2_1 _09824_ (.A(_02695_),
    .B(_02698_),
    .Y(_02703_));
 sg13g2_o21ai_1 _09825_ (.B1(_02702_),
    .Y(_02704_),
    .A1(_02695_),
    .A2(_02698_));
 sg13g2_xnor2_1 _09826_ (.Y(_02705_),
    .A(_02702_),
    .B(_02703_));
 sg13g2_o21ai_1 _09827_ (.B1(net1966),
    .Y(_02706_),
    .A1(net1627),
    .A2(_02705_));
 sg13g2_a21oi_1 _09828_ (.A1(net1627),
    .A2(_01476_),
    .Y(_00369_),
    .B1(_02706_));
 sg13g2_nand2_1 _09829_ (.Y(_02707_),
    .A(\am_sdr0.cic3.integ2[4] ),
    .B(\am_sdr0.cic3.integ1[7] ));
 sg13g2_xnor2_1 _09830_ (.Y(_02708_),
    .A(\am_sdr0.cic3.integ2[4] ),
    .B(\am_sdr0.cic3.integ1[7] ));
 sg13g2_nand3_1 _09831_ (.B(_02704_),
    .C(_02708_),
    .A(_02701_),
    .Y(_02709_));
 sg13g2_a21o_1 _09832_ (.A2(_02704_),
    .A1(_02701_),
    .B1(_02708_),
    .X(_02710_));
 sg13g2_nand2_1 _09833_ (.Y(_02711_),
    .A(_02709_),
    .B(_02710_));
 sg13g2_o21ai_1 _09834_ (.B1(net1966),
    .Y(_02712_),
    .A1(net1738),
    .A2(net3129));
 sg13g2_a21oi_1 _09835_ (.A1(net1738),
    .A2(_02711_),
    .Y(_00370_),
    .B1(_02712_));
 sg13g2_xor2_1 _09836_ (.B(\am_sdr0.cic3.integ1[8] ),
    .A(\am_sdr0.cic3.integ2[5] ),
    .X(_02713_));
 sg13g2_nand2_1 _09837_ (.Y(_02714_),
    .A(_02707_),
    .B(_02710_));
 sg13g2_xnor2_1 _09838_ (.Y(_02715_),
    .A(_02713_),
    .B(_02714_));
 sg13g2_o21ai_1 _09839_ (.B1(net1966),
    .Y(_02716_),
    .A1(net1738),
    .A2(net3140));
 sg13g2_a21oi_1 _09840_ (.A1(net1738),
    .A2(_02715_),
    .Y(_00371_),
    .B1(_02716_));
 sg13g2_and2_1 _09841_ (.A(\am_sdr0.cic3.integ2[6] ),
    .B(\am_sdr0.cic3.integ1[9] ),
    .X(_02717_));
 sg13g2_xor2_1 _09842_ (.B(\am_sdr0.cic3.integ1[9] ),
    .A(\am_sdr0.cic3.integ2[6] ),
    .X(_02718_));
 sg13g2_inv_1 _09843_ (.Y(_02719_),
    .A(_02718_));
 sg13g2_a22oi_1 _09844_ (.Y(_02720_),
    .B1(\am_sdr0.cic3.integ1[7] ),
    .B2(\am_sdr0.cic3.integ2[4] ),
    .A2(\am_sdr0.cic3.integ1[8] ),
    .A1(\am_sdr0.cic3.integ2[5] ));
 sg13g2_a22oi_1 _09845_ (.Y(_02721_),
    .B1(_02710_),
    .B2(_02720_),
    .A2(_01478_),
    .A1(_01475_));
 sg13g2_a221oi_1 _09846_ (.B2(_02720_),
    .C1(_02719_),
    .B1(_02710_),
    .A1(_01475_),
    .Y(_02722_),
    .A2(_01478_));
 sg13g2_xnor2_1 _09847_ (.Y(_02723_),
    .A(_02718_),
    .B(_02721_));
 sg13g2_o21ai_1 _09848_ (.B1(net1967),
    .Y(_02724_),
    .A1(net1740),
    .A2(net3076));
 sg13g2_a21oi_1 _09849_ (.A1(net1740),
    .A2(_02723_),
    .Y(_00372_),
    .B1(_02724_));
 sg13g2_nand2_1 _09850_ (.Y(_02725_),
    .A(\am_sdr0.cic3.integ2[7] ),
    .B(\am_sdr0.cic3.integ1[10] ));
 sg13g2_xnor2_1 _09851_ (.Y(_02726_),
    .A(\am_sdr0.cic3.integ2[7] ),
    .B(\am_sdr0.cic3.integ1[10] ));
 sg13g2_inv_1 _09852_ (.Y(_02727_),
    .A(_02726_));
 sg13g2_o21ai_1 _09853_ (.B1(_02727_),
    .Y(_02728_),
    .A1(_02717_),
    .A2(_02722_));
 sg13g2_or3_1 _09854_ (.A(_02717_),
    .B(_02722_),
    .C(_02727_),
    .X(_02729_));
 sg13g2_nand2_1 _09855_ (.Y(_02730_),
    .A(_02728_),
    .B(_02729_));
 sg13g2_o21ai_1 _09856_ (.B1(net1967),
    .Y(_02731_),
    .A1(net1741),
    .A2(net3049));
 sg13g2_a21oi_1 _09857_ (.A1(net1741),
    .A2(_02730_),
    .Y(_00373_),
    .B1(_02731_));
 sg13g2_xor2_1 _09858_ (.B(\am_sdr0.cic3.integ1[11] ),
    .A(\am_sdr0.cic3.integ2[8] ),
    .X(_02732_));
 sg13g2_inv_1 _09859_ (.Y(_02733_),
    .A(_02732_));
 sg13g2_and3_1 _09860_ (.X(_02734_),
    .A(_02725_),
    .B(_02728_),
    .C(_02733_));
 sg13g2_a21oi_1 _09861_ (.A1(_02725_),
    .A2(_02728_),
    .Y(_02735_),
    .B1(_02733_));
 sg13g2_or2_1 _09862_ (.X(_02736_),
    .B(_02735_),
    .A(_02734_));
 sg13g2_o21ai_1 _09863_ (.B1(net1981),
    .Y(_02737_),
    .A1(net1741),
    .A2(net3145));
 sg13g2_a21oi_1 _09864_ (.A1(net1741),
    .A2(_02736_),
    .Y(_00374_),
    .B1(_02737_));
 sg13g2_nor2_1 _09865_ (.A(\am_sdr0.cic3.integ2[9] ),
    .B(\am_sdr0.cic3.integ1[12] ),
    .Y(_02738_));
 sg13g2_or2_1 _09866_ (.X(_02739_),
    .B(\am_sdr0.cic3.integ1[12] ),
    .A(\am_sdr0.cic3.integ2[9] ));
 sg13g2_a21oi_1 _09867_ (.A1(\am_sdr0.cic3.integ2[8] ),
    .A2(\am_sdr0.cic3.integ1[11] ),
    .Y(_02740_),
    .B1(_02735_));
 sg13g2_and2_1 _09868_ (.A(\am_sdr0.cic3.integ2[9] ),
    .B(\am_sdr0.cic3.integ1[12] ),
    .X(_02741_));
 sg13g2_nor2_1 _09869_ (.A(_02738_),
    .B(_02741_),
    .Y(_02742_));
 sg13g2_xor2_1 _09870_ (.B(_02742_),
    .A(_02740_),
    .X(_02743_));
 sg13g2_o21ai_1 _09871_ (.B1(net1982),
    .Y(_02744_),
    .A1(net1744),
    .A2(net3016));
 sg13g2_a21oi_1 _09872_ (.A1(net1744),
    .A2(_02743_),
    .Y(_00375_),
    .B1(_02744_));
 sg13g2_nand2_1 _09873_ (.Y(_02745_),
    .A(\am_sdr0.cic3.integ2[10] ),
    .B(\am_sdr0.cic3.integ1[13] ));
 sg13g2_xnor2_1 _09874_ (.Y(_02746_),
    .A(\am_sdr0.cic3.integ2[10] ),
    .B(\am_sdr0.cic3.integ1[13] ));
 sg13g2_a21oi_1 _09875_ (.A1(\am_sdr0.cic3.integ2[8] ),
    .A2(\am_sdr0.cic3.integ1[11] ),
    .Y(_02747_),
    .B1(_02741_));
 sg13g2_nor2_1 _09876_ (.A(_02738_),
    .B(_02747_),
    .Y(_02748_));
 sg13g2_a21oi_1 _09877_ (.A1(_02735_),
    .A2(_02739_),
    .Y(_02749_),
    .B1(_02748_));
 sg13g2_xnor2_1 _09878_ (.Y(_02750_),
    .A(_02746_),
    .B(_02749_));
 sg13g2_o21ai_1 _09879_ (.B1(net1982),
    .Y(_02751_),
    .A1(net1744),
    .A2(net3097));
 sg13g2_a21oi_1 _09880_ (.A1(net1744),
    .A2(_02750_),
    .Y(_00376_),
    .B1(_02751_));
 sg13g2_nor2_1 _09881_ (.A(\am_sdr0.cic3.integ2[11] ),
    .B(\am_sdr0.cic3.integ1[14] ),
    .Y(_02752_));
 sg13g2_xnor2_1 _09882_ (.Y(_02753_),
    .A(\am_sdr0.cic3.integ2[11] ),
    .B(\am_sdr0.cic3.integ1[14] ));
 sg13g2_o21ai_1 _09883_ (.B1(_02745_),
    .Y(_02754_),
    .A1(_02746_),
    .A2(_02749_));
 sg13g2_xor2_1 _09884_ (.B(_02754_),
    .A(_02753_),
    .X(_02755_));
 sg13g2_o21ai_1 _09885_ (.B1(net1981),
    .Y(_02756_),
    .A1(net1747),
    .A2(net3038));
 sg13g2_a21oi_1 _09886_ (.A1(net1747),
    .A2(_02755_),
    .Y(_00377_),
    .B1(_02756_));
 sg13g2_nand2_1 _09887_ (.Y(_02757_),
    .A(\am_sdr0.cic3.integ2[12] ),
    .B(\am_sdr0.cic3.integ1[15] ));
 sg13g2_xor2_1 _09888_ (.B(\am_sdr0.cic3.integ1[15] ),
    .A(\am_sdr0.cic3.integ2[12] ),
    .X(_02758_));
 sg13g2_xnor2_1 _09889_ (.Y(_02759_),
    .A(\am_sdr0.cic3.integ2[12] ),
    .B(\am_sdr0.cic3.integ1[15] ));
 sg13g2_nor2_1 _09890_ (.A(_02746_),
    .B(_02753_),
    .Y(_02760_));
 sg13g2_a22oi_1 _09891_ (.Y(_02761_),
    .B1(\am_sdr0.cic3.integ1[13] ),
    .B2(\am_sdr0.cic3.integ2[10] ),
    .A2(\am_sdr0.cic3.integ1[14] ),
    .A1(\am_sdr0.cic3.integ2[11] ));
 sg13g2_nor2_1 _09892_ (.A(_02752_),
    .B(_02761_),
    .Y(_02762_));
 sg13g2_a21oi_1 _09893_ (.A1(_02748_),
    .A2(_02760_),
    .Y(_02763_),
    .B1(_02762_));
 sg13g2_inv_1 _09894_ (.Y(_02764_),
    .A(_02763_));
 sg13g2_and3_1 _09895_ (.X(_02765_),
    .A(_02732_),
    .B(_02742_),
    .C(_02760_));
 sg13g2_inv_1 _09896_ (.Y(_02766_),
    .A(_02765_));
 sg13g2_a21oi_2 _09897_ (.B1(_02766_),
    .Y(_02767_),
    .A2(_02728_),
    .A1(_02725_));
 sg13g2_nor3_1 _09898_ (.A(_02758_),
    .B(_02764_),
    .C(_02767_),
    .Y(_02768_));
 sg13g2_o21ai_1 _09899_ (.B1(_02758_),
    .Y(_02769_),
    .A1(_02764_),
    .A2(_02767_));
 sg13g2_nand2b_1 _09900_ (.Y(_02770_),
    .B(_02769_),
    .A_N(_02768_));
 sg13g2_o21ai_1 _09901_ (.B1(net1983),
    .Y(_02771_),
    .A1(net1743),
    .A2(net3077));
 sg13g2_a21oi_1 _09902_ (.A1(net1743),
    .A2(_02770_),
    .Y(_00378_),
    .B1(_02771_));
 sg13g2_nor2_1 _09903_ (.A(\am_sdr0.cic3.integ2[13] ),
    .B(\am_sdr0.cic3.integ1[16] ),
    .Y(_02772_));
 sg13g2_nand2_1 _09904_ (.Y(_02773_),
    .A(\am_sdr0.cic3.integ2[13] ),
    .B(\am_sdr0.cic3.integ1[16] ));
 sg13g2_nand2b_1 _09905_ (.Y(_02774_),
    .B(_02773_),
    .A_N(_02772_));
 sg13g2_nand2_1 _09906_ (.Y(_02775_),
    .A(_02757_),
    .B(_02769_));
 sg13g2_xor2_1 _09907_ (.B(_02775_),
    .A(_02774_),
    .X(_02776_));
 sg13g2_o21ai_1 _09908_ (.B1(net1983),
    .Y(_02777_),
    .A1(net1747),
    .A2(net3061));
 sg13g2_a21oi_1 _09909_ (.A1(net1747),
    .A2(_02776_),
    .Y(_00379_),
    .B1(_02777_));
 sg13g2_and2_1 _09910_ (.A(\am_sdr0.cic3.integ2[14] ),
    .B(\am_sdr0.cic3.integ1[17] ),
    .X(_02778_));
 sg13g2_xnor2_1 _09911_ (.Y(_02779_),
    .A(\am_sdr0.cic3.integ2[14] ),
    .B(\am_sdr0.cic3.integ1[17] ));
 sg13g2_o21ai_1 _09912_ (.B1(_02773_),
    .Y(_02780_),
    .A1(_02757_),
    .A2(_02772_));
 sg13g2_inv_1 _09913_ (.Y(_02781_),
    .A(_02780_));
 sg13g2_nor2_1 _09914_ (.A(_02759_),
    .B(_02774_),
    .Y(_02782_));
 sg13g2_o21ai_1 _09915_ (.B1(_02782_),
    .Y(_02783_),
    .A1(_02764_),
    .A2(_02767_));
 sg13g2_a21oi_1 _09916_ (.A1(_02781_),
    .A2(_02783_),
    .Y(_02784_),
    .B1(_02779_));
 sg13g2_nand3_1 _09917_ (.B(_02781_),
    .C(_02783_),
    .A(_02779_),
    .Y(_02785_));
 sg13g2_nand2b_1 _09918_ (.Y(_02786_),
    .B(_02785_),
    .A_N(_02784_));
 sg13g2_o21ai_1 _09919_ (.B1(net1983),
    .Y(_02787_),
    .A1(net1747),
    .A2(net3069));
 sg13g2_a21oi_1 _09920_ (.A1(net1747),
    .A2(_02786_),
    .Y(_00380_),
    .B1(_02787_));
 sg13g2_or2_1 _09921_ (.X(_02788_),
    .B(\am_sdr0.cic3.integ1[18] ),
    .A(\am_sdr0.cic3.integ2[15] ));
 sg13g2_and2_1 _09922_ (.A(\am_sdr0.cic3.integ2[15] ),
    .B(\am_sdr0.cic3.integ1[18] ),
    .X(_02789_));
 sg13g2_xnor2_1 _09923_ (.Y(_02790_),
    .A(\am_sdr0.cic3.integ2[15] ),
    .B(\am_sdr0.cic3.integ1[18] ));
 sg13g2_nor3_1 _09924_ (.A(_02778_),
    .B(_02784_),
    .C(_02790_),
    .Y(_02791_));
 sg13g2_o21ai_1 _09925_ (.B1(_02790_),
    .Y(_02792_),
    .A1(_02778_),
    .A2(_02784_));
 sg13g2_nor2_1 _09926_ (.A(net1626),
    .B(_02791_),
    .Y(_02793_));
 sg13g2_o21ai_1 _09927_ (.B1(net1983),
    .Y(_02794_),
    .A1(net1749),
    .A2(net3147));
 sg13g2_a21oi_1 _09928_ (.A1(_02792_),
    .A2(_02793_),
    .Y(_00381_),
    .B1(_02794_));
 sg13g2_nand2_1 _09929_ (.Y(_02795_),
    .A(\am_sdr0.cic3.integ2[16] ),
    .B(\am_sdr0.cic3.integ1[19] ));
 sg13g2_xnor2_1 _09930_ (.Y(_02796_),
    .A(\am_sdr0.cic3.integ2[16] ),
    .B(\am_sdr0.cic3.integ1[19] ));
 sg13g2_or2_1 _09931_ (.X(_02797_),
    .B(_02790_),
    .A(_02779_));
 sg13g2_nor3_1 _09932_ (.A(_02759_),
    .B(_02774_),
    .C(_02797_),
    .Y(_02798_));
 sg13g2_a221oi_1 _09933_ (.B2(_02764_),
    .C1(_02789_),
    .B1(_02798_),
    .A1(_02778_),
    .Y(_02799_),
    .A2(_02788_));
 sg13g2_o21ai_1 _09934_ (.B1(_02799_),
    .Y(_02800_),
    .A1(_02781_),
    .A2(_02797_));
 sg13g2_a21oi_2 _09935_ (.B1(_02800_),
    .Y(_02801_),
    .A2(_02798_),
    .A1(_02767_));
 sg13g2_xnor2_1 _09936_ (.Y(_02802_),
    .A(_02796_),
    .B(_02801_));
 sg13g2_o21ai_1 _09937_ (.B1(net1983),
    .Y(_02803_),
    .A1(net1751),
    .A2(net3128));
 sg13g2_a21oi_1 _09938_ (.A1(net1751),
    .A2(_02802_),
    .Y(_00382_),
    .B1(_02803_));
 sg13g2_or2_1 _09939_ (.X(_02804_),
    .B(\am_sdr0.cic3.integ1[20] ),
    .A(\am_sdr0.cic3.integ2[17] ));
 sg13g2_nand2_1 _09940_ (.Y(_02805_),
    .A(\am_sdr0.cic3.integ2[17] ),
    .B(\am_sdr0.cic3.integ1[20] ));
 sg13g2_nand2_1 _09941_ (.Y(_02806_),
    .A(_02804_),
    .B(_02805_));
 sg13g2_o21ai_1 _09942_ (.B1(_02795_),
    .Y(_02807_),
    .A1(_02796_),
    .A2(_02801_));
 sg13g2_xor2_1 _09943_ (.B(_02807_),
    .A(_02806_),
    .X(_02808_));
 sg13g2_o21ai_1 _09944_ (.B1(net1993),
    .Y(_02809_),
    .A1(net1751),
    .A2(net2989));
 sg13g2_a21oi_1 _09945_ (.A1(net1751),
    .A2(_02808_),
    .Y(_00383_),
    .B1(_02809_));
 sg13g2_and2_1 _09946_ (.A(\am_sdr0.cic3.integ2[18] ),
    .B(\am_sdr0.cic3.integ1[21] ),
    .X(_02810_));
 sg13g2_xor2_1 _09947_ (.B(\am_sdr0.cic3.integ1[21] ),
    .A(\am_sdr0.cic3.integ2[18] ),
    .X(_02811_));
 sg13g2_or2_1 _09948_ (.X(_02812_),
    .B(_02806_),
    .A(_02796_));
 sg13g2_nand3_1 _09949_ (.B(\am_sdr0.cic3.integ1[19] ),
    .C(_02804_),
    .A(\am_sdr0.cic3.integ2[16] ),
    .Y(_02813_));
 sg13g2_and2_1 _09950_ (.A(_02805_),
    .B(_02813_),
    .X(_02814_));
 sg13g2_o21ai_1 _09951_ (.B1(_02814_),
    .Y(_02815_),
    .A1(_02801_),
    .A2(_02812_));
 sg13g2_xnor2_1 _09952_ (.Y(_02816_),
    .A(_02811_),
    .B(_02815_));
 sg13g2_o21ai_1 _09953_ (.B1(net1993),
    .Y(_02817_),
    .A1(net1751),
    .A2(net3137));
 sg13g2_a21oi_1 _09954_ (.A1(net1751),
    .A2(_02816_),
    .Y(_00384_),
    .B1(_02817_));
 sg13g2_nand2_1 _09955_ (.Y(_02818_),
    .A(\am_sdr0.cic3.integ2[19] ),
    .B(\am_sdr0.cic3.integ1[22] ));
 sg13g2_xor2_1 _09956_ (.B(\am_sdr0.cic3.integ1[22] ),
    .A(\am_sdr0.cic3.integ2[19] ),
    .X(_02819_));
 sg13g2_a21oi_1 _09957_ (.A1(_02811_),
    .A2(_02815_),
    .Y(_02820_),
    .B1(_02810_));
 sg13g2_xor2_1 _09958_ (.B(_02820_),
    .A(_02819_),
    .X(_02821_));
 sg13g2_o21ai_1 _09959_ (.B1(net1993),
    .Y(_02822_),
    .A1(net1753),
    .A2(net3098));
 sg13g2_a21oi_1 _09960_ (.A1(net1753),
    .A2(_02821_),
    .Y(_00385_),
    .B1(_02822_));
 sg13g2_nand2_1 _09961_ (.Y(_02823_),
    .A(_02811_),
    .B(_02819_));
 sg13g2_or2_1 _09962_ (.X(_02824_),
    .B(_02823_),
    .A(_02812_));
 sg13g2_o21ai_1 _09963_ (.B1(_02810_),
    .Y(_02825_),
    .A1(\am_sdr0.cic3.integ2[19] ),
    .A2(\am_sdr0.cic3.integ1[22] ));
 sg13g2_o21ai_1 _09964_ (.B1(_02818_),
    .Y(_02826_),
    .A1(_02814_),
    .A2(_02823_));
 sg13g2_nor2b_1 _09965_ (.A(_02826_),
    .B_N(_02825_),
    .Y(_02827_));
 sg13g2_o21ai_1 _09966_ (.B1(_02827_),
    .Y(_02828_),
    .A1(_02801_),
    .A2(_02824_));
 sg13g2_nor2_1 _09967_ (.A(\am_sdr0.cic3.integ2[20] ),
    .B(\am_sdr0.cic3.integ1[23] ),
    .Y(_02829_));
 sg13g2_and2_1 _09968_ (.A(\am_sdr0.cic3.integ2[20] ),
    .B(\am_sdr0.cic3.integ1[23] ),
    .X(_02830_));
 sg13g2_nor2_1 _09969_ (.A(_02829_),
    .B(_02830_),
    .Y(_02831_));
 sg13g2_xnor2_1 _09970_ (.Y(_02832_),
    .A(_02828_),
    .B(_02831_));
 sg13g2_o21ai_1 _09971_ (.B1(net1993),
    .Y(_02833_),
    .A1(net1753),
    .A2(net3041));
 sg13g2_a21oi_1 _09972_ (.A1(net1753),
    .A2(_02832_),
    .Y(_00386_),
    .B1(_02833_));
 sg13g2_or2_1 _09973_ (.X(_02834_),
    .B(\am_sdr0.cic3.integ1[24] ),
    .A(\am_sdr0.cic3.integ2[21] ));
 sg13g2_and2_1 _09974_ (.A(\am_sdr0.cic3.integ2[21] ),
    .B(\am_sdr0.cic3.integ1[24] ),
    .X(_02835_));
 sg13g2_xnor2_1 _09975_ (.Y(_02836_),
    .A(\am_sdr0.cic3.integ2[21] ),
    .B(\am_sdr0.cic3.integ1[24] ));
 sg13g2_a21oi_1 _09976_ (.A1(_02828_),
    .A2(_02831_),
    .Y(_02837_),
    .B1(_02830_));
 sg13g2_xnor2_1 _09977_ (.Y(_02838_),
    .A(_02836_),
    .B(_02837_));
 sg13g2_o21ai_1 _09978_ (.B1(net1994),
    .Y(_02839_),
    .A1(net1754),
    .A2(net3024));
 sg13g2_a21oi_1 _09979_ (.A1(net1754),
    .A2(_02838_),
    .Y(_00387_),
    .B1(_02839_));
 sg13g2_nor3_1 _09980_ (.A(_02829_),
    .B(_02830_),
    .C(_02836_),
    .Y(_02840_));
 sg13g2_a221oi_1 _09981_ (.B2(_02828_),
    .C1(_02835_),
    .B1(_02840_),
    .A1(_02830_),
    .Y(_02841_),
    .A2(_02834_));
 sg13g2_xor2_1 _09982_ (.B(net1297),
    .A(net2896),
    .X(_02842_));
 sg13g2_or2_1 _09983_ (.X(_02843_),
    .B(_02842_),
    .A(_02841_));
 sg13g2_a21oi_1 _09984_ (.A1(_02841_),
    .A2(_02842_),
    .Y(_02844_),
    .B1(_01470_));
 sg13g2_o21ai_1 _09985_ (.B1(net1994),
    .Y(_02845_),
    .A1(net1750),
    .A2(net2896));
 sg13g2_a21oi_1 _09986_ (.A1(_02843_),
    .A2(_02844_),
    .Y(_00388_),
    .B1(_02845_));
 sg13g2_a21oi_1 _09987_ (.A1(net1741),
    .A2(\am_sdr0.cic3.integ2[3] ),
    .Y(_02846_),
    .B1(net2116));
 sg13g2_nand2_1 _09988_ (.Y(_02847_),
    .A(net2116),
    .B(\am_sdr0.cic3.integ2[3] ));
 sg13g2_nor2_1 _09989_ (.A(net1626),
    .B(_02847_),
    .Y(_02848_));
 sg13g2_nor3_1 _09990_ (.A(net1890),
    .B(net2117),
    .C(_02848_),
    .Y(_00389_));
 sg13g2_nand2_1 _09991_ (.Y(_02849_),
    .A(\am_sdr0.cic3.integ3[1] ),
    .B(\am_sdr0.cic3.integ2[4] ));
 sg13g2_xnor2_1 _09992_ (.Y(_02850_),
    .A(\am_sdr0.cic3.integ3[1] ),
    .B(\am_sdr0.cic3.integ2[4] ));
 sg13g2_xnor2_1 _09993_ (.Y(_02851_),
    .A(_02847_),
    .B(_02850_));
 sg13g2_o21ai_1 _09994_ (.B1(net1981),
    .Y(_02852_),
    .A1(net1744),
    .A2(net3015));
 sg13g2_a21oi_1 _09995_ (.A1(net1744),
    .A2(_02851_),
    .Y(_00390_),
    .B1(_02852_));
 sg13g2_and2_1 _09996_ (.A(\am_sdr0.cic3.integ3[2] ),
    .B(\am_sdr0.cic3.integ2[5] ),
    .X(_02853_));
 sg13g2_xor2_1 _09997_ (.B(\am_sdr0.cic3.integ2[5] ),
    .A(\am_sdr0.cic3.integ3[2] ),
    .X(_02854_));
 sg13g2_o21ai_1 _09998_ (.B1(_02849_),
    .Y(_02855_),
    .A1(_02847_),
    .A2(_02850_));
 sg13g2_and2_1 _09999_ (.A(_02854_),
    .B(_02855_),
    .X(_02856_));
 sg13g2_xnor2_1 _10000_ (.Y(_02857_),
    .A(_02854_),
    .B(_02855_));
 sg13g2_o21ai_1 _10001_ (.B1(net1981),
    .Y(_02858_),
    .A1(net1744),
    .A2(net2974));
 sg13g2_a21oi_1 _10002_ (.A1(net1744),
    .A2(_02857_),
    .Y(_00391_),
    .B1(_02858_));
 sg13g2_nand2_1 _10003_ (.Y(_02859_),
    .A(net2467),
    .B(\am_sdr0.cic3.integ2[6] ));
 sg13g2_xor2_1 _10004_ (.B(\am_sdr0.cic3.integ2[6] ),
    .A(\am_sdr0.cic3.integ3[3] ),
    .X(_02860_));
 sg13g2_nor2_1 _10005_ (.A(_02853_),
    .B(_02856_),
    .Y(_02861_));
 sg13g2_o21ai_1 _10006_ (.B1(_02860_),
    .Y(_02862_),
    .A1(_02853_),
    .A2(_02856_));
 sg13g2_xnor2_1 _10007_ (.Y(_02863_),
    .A(_02860_),
    .B(_02861_));
 sg13g2_o21ai_1 _10008_ (.B1(net1981),
    .Y(_02864_),
    .A1(net1626),
    .A2(_02863_));
 sg13g2_a21oi_1 _10009_ (.A1(net1626),
    .A2(_01473_),
    .Y(_00392_),
    .B1(_02864_));
 sg13g2_nand2_1 _10010_ (.Y(_02865_),
    .A(\am_sdr0.cic3.integ3[4] ),
    .B(\am_sdr0.cic3.integ2[7] ));
 sg13g2_xnor2_1 _10011_ (.Y(_02866_),
    .A(\am_sdr0.cic3.integ3[4] ),
    .B(\am_sdr0.cic3.integ2[7] ));
 sg13g2_nand3_1 _10012_ (.B(_02862_),
    .C(_02866_),
    .A(_02859_),
    .Y(_02867_));
 sg13g2_a21o_1 _10013_ (.A2(_02862_),
    .A1(_02859_),
    .B1(_02866_),
    .X(_02868_));
 sg13g2_nand2_1 _10014_ (.Y(_02869_),
    .A(_02867_),
    .B(_02868_));
 sg13g2_o21ai_1 _10015_ (.B1(net1981),
    .Y(_02870_),
    .A1(net1745),
    .A2(net3007));
 sg13g2_a21oi_1 _10016_ (.A1(net1745),
    .A2(_02869_),
    .Y(_00393_),
    .B1(_02870_));
 sg13g2_xor2_1 _10017_ (.B(\am_sdr0.cic3.integ2[8] ),
    .A(net2980),
    .X(_02871_));
 sg13g2_nand2_1 _10018_ (.Y(_02872_),
    .A(_02865_),
    .B(_02868_));
 sg13g2_xnor2_1 _10019_ (.Y(_02873_),
    .A(_02871_),
    .B(_02872_));
 sg13g2_o21ai_1 _10020_ (.B1(net1982),
    .Y(_02874_),
    .A1(net1745),
    .A2(net2765));
 sg13g2_a21oi_1 _10021_ (.A1(net1745),
    .A2(net2981),
    .Y(_00394_),
    .B1(_02874_));
 sg13g2_and2_1 _10022_ (.A(\am_sdr0.cic3.integ3[6] ),
    .B(\am_sdr0.cic3.integ2[9] ),
    .X(_02875_));
 sg13g2_xnor2_1 _10023_ (.Y(_02876_),
    .A(\am_sdr0.cic3.integ3[6] ),
    .B(\am_sdr0.cic3.integ2[9] ));
 sg13g2_a22oi_1 _10024_ (.Y(_02877_),
    .B1(\am_sdr0.cic3.integ2[7] ),
    .B2(\am_sdr0.cic3.integ3[4] ),
    .A2(\am_sdr0.cic3.integ2[8] ),
    .A1(\am_sdr0.cic3.integ3[5] ));
 sg13g2_a22oi_1 _10025_ (.Y(_02878_),
    .B1(_02868_),
    .B2(_02877_),
    .A2(_01474_),
    .A1(_01472_));
 sg13g2_a221oi_1 _10026_ (.B2(_02877_),
    .C1(_02876_),
    .B1(_02868_),
    .A1(_01472_),
    .Y(_02879_),
    .A2(_01474_));
 sg13g2_xnor2_1 _10027_ (.Y(_02880_),
    .A(_02876_),
    .B(_02878_));
 sg13g2_o21ai_1 _10028_ (.B1(net1981),
    .Y(_02881_),
    .A1(net1626),
    .A2(_02880_));
 sg13g2_a21oi_1 _10029_ (.A1(net1626),
    .A2(_01471_),
    .Y(_00395_),
    .B1(_02881_));
 sg13g2_nand2_1 _10030_ (.Y(_02882_),
    .A(\am_sdr0.cic3.integ3[7] ),
    .B(\am_sdr0.cic3.integ2[10] ));
 sg13g2_xor2_1 _10031_ (.B(\am_sdr0.cic3.integ2[10] ),
    .A(\am_sdr0.cic3.integ3[7] ),
    .X(_02883_));
 sg13g2_o21ai_1 _10032_ (.B1(_02883_),
    .Y(_02884_),
    .A1(_02875_),
    .A2(_02879_));
 sg13g2_or3_1 _10033_ (.A(_02875_),
    .B(_02879_),
    .C(_02883_),
    .X(_02885_));
 sg13g2_a21oi_1 _10034_ (.A1(_02884_),
    .A2(_02885_),
    .Y(_02886_),
    .B1(net1626));
 sg13g2_o21ai_1 _10035_ (.B1(net1981),
    .Y(_02887_),
    .A1(net1746),
    .A2(net2977));
 sg13g2_nor2_1 _10036_ (.A(_02886_),
    .B(_02887_),
    .Y(_00396_));
 sg13g2_nand2_1 _10037_ (.Y(_02888_),
    .A(_02882_),
    .B(_02884_));
 sg13g2_and2_1 _10038_ (.A(\am_sdr0.cic3.integ3[8] ),
    .B(\am_sdr0.cic3.integ2[11] ),
    .X(_02889_));
 sg13g2_xor2_1 _10039_ (.B(\am_sdr0.cic3.integ2[11] ),
    .A(\am_sdr0.cic3.integ3[8] ),
    .X(_02890_));
 sg13g2_xnor2_1 _10040_ (.Y(_02891_),
    .A(_02888_),
    .B(_02890_));
 sg13g2_o21ai_1 _10041_ (.B1(net1984),
    .Y(_02892_),
    .A1(net1746),
    .A2(net2967));
 sg13g2_a21oi_1 _10042_ (.A1(net1746),
    .A2(_02891_),
    .Y(_00397_),
    .B1(_02892_));
 sg13g2_or2_1 _10043_ (.X(_02893_),
    .B(\am_sdr0.cic3.integ2[12] ),
    .A(\am_sdr0.cic3.integ3[9] ));
 sg13g2_nand2_1 _10044_ (.Y(_02894_),
    .A(net2755),
    .B(\am_sdr0.cic3.integ2[12] ));
 sg13g2_nand2_1 _10045_ (.Y(_02895_),
    .A(_02893_),
    .B(_02894_));
 sg13g2_a21oi_1 _10046_ (.A1(_02888_),
    .A2(_02890_),
    .Y(_02896_),
    .B1(_02889_));
 sg13g2_xnor2_1 _10047_ (.Y(_02897_),
    .A(_02895_),
    .B(_02896_));
 sg13g2_o21ai_1 _10048_ (.B1(net1984),
    .Y(_02898_),
    .A1(net1746),
    .A2(net2405));
 sg13g2_a21oi_1 _10049_ (.A1(net1746),
    .A2(_02897_),
    .Y(_00398_),
    .B1(_02898_));
 sg13g2_nand2_1 _10050_ (.Y(_02899_),
    .A(\am_sdr0.cic3.integ3[10] ),
    .B(\am_sdr0.cic3.integ2[13] ));
 sg13g2_xnor2_1 _10051_ (.Y(_02900_),
    .A(\am_sdr0.cic3.integ3[10] ),
    .B(\am_sdr0.cic3.integ2[13] ));
 sg13g2_nand2_1 _10052_ (.Y(_02901_),
    .A(_02889_),
    .B(_02893_));
 sg13g2_nand2_1 _10053_ (.Y(_02902_),
    .A(_02894_),
    .B(_02901_));
 sg13g2_and3_1 _10054_ (.X(_02903_),
    .A(_02890_),
    .B(_02893_),
    .C(_02894_));
 sg13g2_a21oi_1 _10055_ (.A1(_02888_),
    .A2(_02903_),
    .Y(_02904_),
    .B1(_02902_));
 sg13g2_xnor2_1 _10056_ (.Y(_02905_),
    .A(_02900_),
    .B(_02904_));
 sg13g2_o21ai_1 _10057_ (.B1(net1983),
    .Y(_02906_),
    .A1(net1747),
    .A2(net2995));
 sg13g2_a21oi_1 _10058_ (.A1(net1746),
    .A2(_02905_),
    .Y(_00399_),
    .B1(_02906_));
 sg13g2_or2_1 _10059_ (.X(_02907_),
    .B(\am_sdr0.cic3.integ2[14] ),
    .A(\am_sdr0.cic3.integ3[11] ));
 sg13g2_xnor2_1 _10060_ (.Y(_02908_),
    .A(\am_sdr0.cic3.integ3[11] ),
    .B(\am_sdr0.cic3.integ2[14] ));
 sg13g2_o21ai_1 _10061_ (.B1(_02899_),
    .Y(_02909_),
    .A1(_02900_),
    .A2(_02904_));
 sg13g2_xor2_1 _10062_ (.B(_02909_),
    .A(_02908_),
    .X(_02910_));
 sg13g2_o21ai_1 _10063_ (.B1(net1983),
    .Y(_02911_),
    .A1(net1746),
    .A2(net2959));
 sg13g2_a21oi_1 _10064_ (.A1(net1746),
    .A2(_02910_),
    .Y(_00400_),
    .B1(_02911_));
 sg13g2_nand2_1 _10065_ (.Y(_02912_),
    .A(net3040),
    .B(\am_sdr0.cic3.integ2[15] ));
 sg13g2_xor2_1 _10066_ (.B(\am_sdr0.cic3.integ2[15] ),
    .A(\am_sdr0.cic3.integ3[12] ),
    .X(_02913_));
 sg13g2_inv_1 _10067_ (.Y(_02914_),
    .A(_02913_));
 sg13g2_nor2_1 _10068_ (.A(_02900_),
    .B(_02908_),
    .Y(_02915_));
 sg13g2_and3_1 _10069_ (.X(_02916_),
    .A(\am_sdr0.cic3.integ3[10] ),
    .B(\am_sdr0.cic3.integ2[13] ),
    .C(_02907_));
 sg13g2_a221oi_1 _10070_ (.B2(_02915_),
    .C1(_02916_),
    .B1(_02902_),
    .A1(\am_sdr0.cic3.integ3[11] ),
    .Y(_02917_),
    .A2(\am_sdr0.cic3.integ2[14] ));
 sg13g2_inv_1 _10071_ (.Y(_02918_),
    .A(_02917_));
 sg13g2_and2_1 _10072_ (.A(_02903_),
    .B(_02915_),
    .X(_02919_));
 sg13g2_inv_1 _10073_ (.Y(_02920_),
    .A(_02919_));
 sg13g2_a21oi_2 _10074_ (.B1(_02920_),
    .Y(_02921_),
    .A2(_02884_),
    .A1(_02882_));
 sg13g2_nor3_1 _10075_ (.A(_02913_),
    .B(_02918_),
    .C(_02921_),
    .Y(_02922_));
 sg13g2_o21ai_1 _10076_ (.B1(_02913_),
    .Y(_02923_),
    .A1(_02918_),
    .A2(_02921_));
 sg13g2_nand2b_1 _10077_ (.Y(_02924_),
    .B(_02923_),
    .A_N(_02922_));
 sg13g2_o21ai_1 _10078_ (.B1(net1984),
    .Y(_02925_),
    .A1(net1752),
    .A2(net2984));
 sg13g2_a21oi_1 _10079_ (.A1(net1752),
    .A2(_02924_),
    .Y(_00401_),
    .B1(_02925_));
 sg13g2_nor2_1 _10080_ (.A(\am_sdr0.cic3.integ3[13] ),
    .B(\am_sdr0.cic3.integ2[16] ),
    .Y(_02926_));
 sg13g2_xnor2_1 _10081_ (.Y(_02927_),
    .A(\am_sdr0.cic3.integ3[13] ),
    .B(\am_sdr0.cic3.integ2[16] ));
 sg13g2_nand2_1 _10082_ (.Y(_02928_),
    .A(_02912_),
    .B(_02923_));
 sg13g2_xor2_1 _10083_ (.B(_02928_),
    .A(_02927_),
    .X(_02929_));
 sg13g2_o21ai_1 _10084_ (.B1(net1996),
    .Y(_02930_),
    .A1(net1751),
    .A2(net2787));
 sg13g2_a21oi_1 _10085_ (.A1(net1751),
    .A2(_02929_),
    .Y(_00402_),
    .B1(_02930_));
 sg13g2_and2_1 _10086_ (.A(net2899),
    .B(\am_sdr0.cic3.integ2[17] ),
    .X(_02931_));
 sg13g2_xor2_1 _10087_ (.B(\am_sdr0.cic3.integ2[17] ),
    .A(\am_sdr0.cic3.integ3[14] ),
    .X(_02932_));
 sg13g2_inv_1 _10088_ (.Y(_02933_),
    .A(_02932_));
 sg13g2_a22oi_1 _10089_ (.Y(_02934_),
    .B1(\am_sdr0.cic3.integ2[15] ),
    .B2(\am_sdr0.cic3.integ3[12] ),
    .A2(\am_sdr0.cic3.integ2[16] ),
    .A1(\am_sdr0.cic3.integ3[13] ));
 sg13g2_a21oi_1 _10090_ (.A1(_02923_),
    .A2(_02934_),
    .Y(_02935_),
    .B1(_02926_));
 sg13g2_xnor2_1 _10091_ (.Y(_02936_),
    .A(net2900),
    .B(_02935_));
 sg13g2_o21ai_1 _10092_ (.B1(net1996),
    .Y(_02937_),
    .A1(net1752),
    .A2(net2279));
 sg13g2_a21oi_1 _10093_ (.A1(net1752),
    .A2(_02936_),
    .Y(_00403_),
    .B1(_02937_));
 sg13g2_nand2_1 _10094_ (.Y(_02938_),
    .A(\am_sdr0.cic3.integ3[15] ),
    .B(\am_sdr0.cic3.integ2[18] ));
 sg13g2_xnor2_1 _10095_ (.Y(_02939_),
    .A(\am_sdr0.cic3.integ3[15] ),
    .B(\am_sdr0.cic3.integ2[18] ));
 sg13g2_a21oi_1 _10096_ (.A1(_02932_),
    .A2(_02935_),
    .Y(_02940_),
    .B1(_02931_));
 sg13g2_xnor2_1 _10097_ (.Y(_02941_),
    .A(_02939_),
    .B(_02940_));
 sg13g2_o21ai_1 _10098_ (.B1(net1993),
    .Y(_02942_),
    .A1(net1752),
    .A2(net2733));
 sg13g2_a21oi_1 _10099_ (.A1(net1752),
    .A2(_02941_),
    .Y(_00404_),
    .B1(_02942_));
 sg13g2_nand2_1 _10100_ (.Y(_02943_),
    .A(net2954),
    .B(\am_sdr0.cic3.integ2[19] ));
 sg13g2_xnor2_1 _10101_ (.Y(_02944_),
    .A(\am_sdr0.cic3.integ3[16] ),
    .B(\am_sdr0.cic3.integ2[19] ));
 sg13g2_nor4_2 _10102_ (.A(_02914_),
    .B(_02927_),
    .C(_02933_),
    .Y(_02945_),
    .D(_02939_));
 sg13g2_o21ai_1 _10103_ (.B1(_02931_),
    .Y(_02946_),
    .A1(\am_sdr0.cic3.integ3[15] ),
    .A2(\am_sdr0.cic3.integ2[18] ));
 sg13g2_nor4_1 _10104_ (.A(_02926_),
    .B(_02933_),
    .C(_02934_),
    .D(_02939_),
    .Y(_02947_));
 sg13g2_a21oi_1 _10105_ (.A1(_02918_),
    .A2(_02945_),
    .Y(_02948_),
    .B1(_02947_));
 sg13g2_nand3_1 _10106_ (.B(_02946_),
    .C(_02948_),
    .A(_02938_),
    .Y(_02949_));
 sg13g2_a21oi_2 _10107_ (.B1(_02949_),
    .Y(_02950_),
    .A2(_02945_),
    .A1(_02921_));
 sg13g2_xnor2_1 _10108_ (.Y(_02951_),
    .A(_02944_),
    .B(_02950_));
 sg13g2_o21ai_1 _10109_ (.B1(net1993),
    .Y(_02952_),
    .A1(net1754),
    .A2(net2517));
 sg13g2_a21oi_1 _10110_ (.A1(net1754),
    .A2(_02951_),
    .Y(_00405_),
    .B1(_02952_));
 sg13g2_nor2_1 _10111_ (.A(\am_sdr0.cic3.integ3[17] ),
    .B(\am_sdr0.cic3.integ2[20] ),
    .Y(_02953_));
 sg13g2_xnor2_1 _10112_ (.Y(_02954_),
    .A(\am_sdr0.cic3.integ3[17] ),
    .B(\am_sdr0.cic3.integ2[20] ));
 sg13g2_o21ai_1 _10113_ (.B1(_02943_),
    .Y(_02955_),
    .A1(_02944_),
    .A2(_02950_));
 sg13g2_xor2_1 _10114_ (.B(_02955_),
    .A(_02954_),
    .X(_02956_));
 sg13g2_o21ai_1 _10115_ (.B1(net1994),
    .Y(_02957_),
    .A1(net1754),
    .A2(net2791));
 sg13g2_a21oi_1 _10116_ (.A1(net1754),
    .A2(_02956_),
    .Y(_00406_),
    .B1(_02957_));
 sg13g2_and2_1 _10117_ (.A(\am_sdr0.cic3.integ3[18] ),
    .B(\am_sdr0.cic3.integ2[21] ),
    .X(_02958_));
 sg13g2_or2_1 _10118_ (.X(_02959_),
    .B(\am_sdr0.cic3.integ2[21] ),
    .A(\am_sdr0.cic3.integ3[18] ));
 sg13g2_nor2b_1 _10119_ (.A(_02958_),
    .B_N(_02959_),
    .Y(_02960_));
 sg13g2_or2_1 _10120_ (.X(_02961_),
    .B(_02954_),
    .A(_02944_));
 sg13g2_nor2_1 _10121_ (.A(_02943_),
    .B(_02953_),
    .Y(_02962_));
 sg13g2_a21oi_1 _10122_ (.A1(\am_sdr0.cic3.integ3[17] ),
    .A2(\am_sdr0.cic3.integ2[20] ),
    .Y(_02963_),
    .B1(_02962_));
 sg13g2_o21ai_1 _10123_ (.B1(_02963_),
    .Y(_02964_),
    .A1(_02950_),
    .A2(_02961_));
 sg13g2_xnor2_1 _10124_ (.Y(_02965_),
    .A(_02960_),
    .B(_02964_));
 sg13g2_o21ai_1 _10125_ (.B1(net1994),
    .Y(_02966_),
    .A1(net1753),
    .A2(net2230));
 sg13g2_a21oi_1 _10126_ (.A1(net1753),
    .A2(_02965_),
    .Y(_00407_),
    .B1(_02966_));
 sg13g2_a21oi_1 _10127_ (.A1(_02959_),
    .A2(_02964_),
    .Y(_02967_),
    .B1(_02958_));
 sg13g2_xnor2_1 _10128_ (.Y(_02968_),
    .A(net2874),
    .B(\am_sdr0.cic3.integ2[22] ));
 sg13g2_xnor2_1 _10129_ (.Y(_02969_),
    .A(_02967_),
    .B(_02968_));
 sg13g2_o21ai_1 _10130_ (.B1(net1994),
    .Y(_02970_),
    .A1(net2874),
    .A2(net1753));
 sg13g2_a21oi_1 _10131_ (.A1(net1753),
    .A2(_02969_),
    .Y(_00408_),
    .B1(_02970_));
 sg13g2_nor2_1 _10132_ (.A(net1634),
    .B(net1892),
    .Y(_00410_));
 sg13g2_and3_1 _10133_ (.X(_02971_),
    .A(\am_sdr0.cic1.count[0] ),
    .B(\am_sdr0.cic1.count[1] ),
    .C(net1202));
 sg13g2_and2_1 _10134_ (.A(net1439),
    .B(_02971_),
    .X(_02972_));
 sg13g2_and2_1 _10135_ (.A(net1429),
    .B(_02972_),
    .X(_02973_));
 sg13g2_nand2_1 _10136_ (.Y(_02974_),
    .A(net2857),
    .B(_02973_));
 sg13g2_or2_1 _10137_ (.X(_02975_),
    .B(\am_sdr0.cic1.count[6] ),
    .A(\am_sdr0.cic1.count[7] ));
 sg13g2_nor3_1 _10138_ (.A(net1877),
    .B(_02974_),
    .C(_02975_),
    .Y(_00624_));
 sg13g2_mux2_1 _10139_ (.A0(\am_sdr0.cic1.integ_sample[0] ),
    .A1(net2407),
    .S(net1552),
    .X(_00411_));
 sg13g2_nand2_1 _10140_ (.Y(_02976_),
    .A(net1389),
    .B(net1550));
 sg13g2_o21ai_1 _10141_ (.B1(_02976_),
    .Y(_00412_),
    .A1(_01381_),
    .A2(net1550));
 sg13g2_nand2_1 _10142_ (.Y(_02977_),
    .A(net2081),
    .B(net1550));
 sg13g2_o21ai_1 _10143_ (.B1(_02977_),
    .Y(_00413_),
    .A1(_01380_),
    .A2(net1550));
 sg13g2_nand2_1 _10144_ (.Y(_02978_),
    .A(net2070),
    .B(net1550));
 sg13g2_o21ai_1 _10145_ (.B1(_02978_),
    .Y(_00414_),
    .A1(_01379_),
    .A2(net1550));
 sg13g2_nand2_1 _10146_ (.Y(_02979_),
    .A(net2159),
    .B(net1550));
 sg13g2_o21ai_1 _10147_ (.B1(_02979_),
    .Y(_00415_),
    .A1(_01378_),
    .A2(net1550));
 sg13g2_nand2_1 _10148_ (.Y(_02980_),
    .A(net2085),
    .B(net1551));
 sg13g2_o21ai_1 _10149_ (.B1(_02980_),
    .Y(_00416_),
    .A1(_01377_),
    .A2(net1551));
 sg13g2_nand2_1 _10150_ (.Y(_02981_),
    .A(net1334),
    .B(net1551));
 sg13g2_o21ai_1 _10151_ (.B1(_02981_),
    .Y(_00417_),
    .A1(_01375_),
    .A2(net1551));
 sg13g2_nand2_1 _10152_ (.Y(_02982_),
    .A(net1441),
    .B(net1551));
 sg13g2_o21ai_1 _10153_ (.B1(_02982_),
    .Y(_00418_),
    .A1(_01374_),
    .A2(net1551));
 sg13g2_nand2_1 _10154_ (.Y(_02983_),
    .A(net1476),
    .B(net1551));
 sg13g2_o21ai_1 _10155_ (.B1(_02983_),
    .Y(_00419_),
    .A1(_01373_),
    .A2(net1551));
 sg13g2_nand2_1 _10156_ (.Y(_02984_),
    .A(net1423),
    .B(net1548));
 sg13g2_o21ai_1 _10157_ (.B1(_02984_),
    .Y(_00420_),
    .A1(_01372_),
    .A2(net1548));
 sg13g2_nand2_1 _10158_ (.Y(_02985_),
    .A(net1497),
    .B(net1548));
 sg13g2_o21ai_1 _10159_ (.B1(_02985_),
    .Y(_00421_),
    .A1(_01370_),
    .A2(net1548));
 sg13g2_nand2_1 _10160_ (.Y(_02986_),
    .A(net2114),
    .B(net1548));
 sg13g2_o21ai_1 _10161_ (.B1(_02986_),
    .Y(_00422_),
    .A1(_01369_),
    .A2(net1548));
 sg13g2_mux2_1 _10162_ (.A0(\am_sdr0.cic1.integ_sample[12] ),
    .A1(net2645),
    .S(net1548),
    .X(_00423_));
 sg13g2_nand2_1 _10163_ (.Y(_02987_),
    .A(net1398),
    .B(net1549));
 sg13g2_o21ai_1 _10164_ (.B1(_02987_),
    .Y(_00424_),
    .A1(_01367_),
    .A2(net1548));
 sg13g2_nand2_1 _10165_ (.Y(_02988_),
    .A(net2354),
    .B(net1547));
 sg13g2_o21ai_1 _10166_ (.B1(_02988_),
    .Y(_00425_),
    .A1(_01366_),
    .A2(net1546));
 sg13g2_nand2_1 _10167_ (.Y(_02989_),
    .A(net2176),
    .B(net1546));
 sg13g2_o21ai_1 _10168_ (.B1(_02989_),
    .Y(_00426_),
    .A1(_01365_),
    .A2(net1546));
 sg13g2_nand2_1 _10169_ (.Y(_02990_),
    .A(net2157),
    .B(net1547));
 sg13g2_o21ai_1 _10170_ (.B1(_02990_),
    .Y(_00427_),
    .A1(_01364_),
    .A2(net1547));
 sg13g2_nor2_1 _10171_ (.A(net2351),
    .B(net1546),
    .Y(_02991_));
 sg13g2_a21oi_1 _10172_ (.A1(_01591_),
    .A2(net1546),
    .Y(_00428_),
    .B1(_02991_));
 sg13g2_nand2_1 _10173_ (.Y(_02992_),
    .A(net1406),
    .B(net1547));
 sg13g2_o21ai_1 _10174_ (.B1(_02992_),
    .Y(_00429_),
    .A1(_01362_),
    .A2(net1547));
 sg13g2_nand2_1 _10175_ (.Y(_02993_),
    .A(net1379),
    .B(net1546));
 sg13g2_o21ai_1 _10176_ (.B1(_02993_),
    .Y(_00430_),
    .A1(_01361_),
    .A2(net1546));
 sg13g2_o21ai_1 _10177_ (.B1(net2018),
    .Y(_02994_),
    .A1(net1823),
    .A2(\am_sdr0.am0.I_in[0] ));
 sg13g2_a21oi_1 _10178_ (.A1(net1822),
    .A2(_01425_),
    .Y(_00431_),
    .B1(_02994_));
 sg13g2_o21ai_1 _10179_ (.B1(net2018),
    .Y(_02995_),
    .A1(net1824),
    .A2(\am_sdr0.am0.I_in[1] ));
 sg13g2_a21oi_1 _10180_ (.A1(net1823),
    .A2(_01424_),
    .Y(_00432_),
    .B1(_02995_));
 sg13g2_o21ai_1 _10181_ (.B1(net2018),
    .Y(_02996_),
    .A1(net1823),
    .A2(\am_sdr0.am0.I_in[2] ));
 sg13g2_a21oi_1 _10182_ (.A1(net1823),
    .A2(_01423_),
    .Y(_00433_),
    .B1(_02996_));
 sg13g2_o21ai_1 _10183_ (.B1(net2018),
    .Y(_02997_),
    .A1(net1823),
    .A2(\am_sdr0.am0.I_in[3] ));
 sg13g2_a21oi_1 _10184_ (.A1(net1823),
    .A2(_01422_),
    .Y(_00434_),
    .B1(_02997_));
 sg13g2_o21ai_1 _10185_ (.B1(net2021),
    .Y(_02998_),
    .A1(net1824),
    .A2(\am_sdr0.am0.I_in[4] ));
 sg13g2_a21oi_1 _10186_ (.A1(net1824),
    .A2(_01421_),
    .Y(_00435_),
    .B1(_02998_));
 sg13g2_o21ai_1 _10187_ (.B1(net2020),
    .Y(_02999_),
    .A1(net1825),
    .A2(\am_sdr0.am0.I_in[5] ));
 sg13g2_a21oi_1 _10188_ (.A1(net1825),
    .A2(_01420_),
    .Y(_00436_),
    .B1(_02999_));
 sg13g2_o21ai_1 _10189_ (.B1(net2020),
    .Y(_03000_),
    .A1(net1829),
    .A2(\am_sdr0.am0.I_in[6] ));
 sg13g2_a21oi_1 _10190_ (.A1(net1829),
    .A2(_01419_),
    .Y(_00437_),
    .B1(_03000_));
 sg13g2_o21ai_1 _10191_ (.B1(net2020),
    .Y(_03001_),
    .A1(net1829),
    .A2(\am_sdr0.am0.I_in[7] ));
 sg13g2_a21oi_1 _10192_ (.A1(net1829),
    .A2(_01418_),
    .Y(_00438_),
    .B1(_03001_));
 sg13g2_nand2b_1 _10193_ (.Y(_03002_),
    .B(net2068),
    .A_N(net2422));
 sg13g2_a21oi_1 _10194_ (.A1(_01469_),
    .A2(net2422),
    .Y(_03003_),
    .B1(net1630));
 sg13g2_a221oi_1 _10195_ (.B2(_03003_),
    .C1(net1891),
    .B1(_03002_),
    .A1(net1630),
    .Y(_00439_),
    .A2(_01448_));
 sg13g2_nor2b_1 _10196_ (.A(net2870),
    .B_N(\am_sdr0.cic2.integ_sample[1] ),
    .Y(_03004_));
 sg13g2_xnor2_1 _10197_ (.Y(_03005_),
    .A(net2870),
    .B(net2453));
 sg13g2_xnor2_1 _10198_ (.Y(_03006_),
    .A(_03002_),
    .B(_03005_));
 sg13g2_o21ai_1 _10199_ (.B1(net2014),
    .Y(_03007_),
    .A1(net1814),
    .A2(net2312));
 sg13g2_a21oi_1 _10200_ (.A1(net1813),
    .A2(_03006_),
    .Y(_00440_),
    .B1(_03007_));
 sg13g2_nand2b_1 _10201_ (.Y(_03008_),
    .B(\am_sdr0.cic2.integ_sample[2] ),
    .A_N(\am_sdr0.cic2.comb1_in_del[2] ));
 sg13g2_xor2_1 _10202_ (.B(net2599),
    .A(net2992),
    .X(_03009_));
 sg13g2_a21oi_1 _10203_ (.A1(_03002_),
    .A2(_03005_),
    .Y(_03010_),
    .B1(_03004_));
 sg13g2_xnor2_1 _10204_ (.Y(_03011_),
    .A(_03009_),
    .B(_03010_));
 sg13g2_o21ai_1 _10205_ (.B1(net2006),
    .Y(_03012_),
    .A1(net1814),
    .A2(net2420));
 sg13g2_a21oi_1 _10206_ (.A1(net1813),
    .A2(_03011_),
    .Y(_00441_),
    .B1(_03012_));
 sg13g2_nor2_1 _10207_ (.A(\am_sdr0.cic2.comb1_in_del[3] ),
    .B(_01466_),
    .Y(_03013_));
 sg13g2_nand2_1 _10208_ (.Y(_03014_),
    .A(\am_sdr0.cic2.comb1_in_del[3] ),
    .B(_01466_));
 sg13g2_nor2b_1 _10209_ (.A(_03013_),
    .B_N(_03014_),
    .Y(_03015_));
 sg13g2_o21ai_1 _10210_ (.B1(_03008_),
    .Y(_03016_),
    .A1(_03009_),
    .A2(_03010_));
 sg13g2_xnor2_1 _10211_ (.Y(_03017_),
    .A(_03015_),
    .B(_03016_));
 sg13g2_o21ai_1 _10212_ (.B1(net2005),
    .Y(_03018_),
    .A1(net1812),
    .A2(net2581));
 sg13g2_a21oi_1 _10213_ (.A1(net1812),
    .A2(_03017_),
    .Y(_00442_),
    .B1(_03018_));
 sg13g2_nor2_1 _10214_ (.A(\am_sdr0.cic2.comb1_in_del[4] ),
    .B(_01465_),
    .Y(_03019_));
 sg13g2_xor2_1 _10215_ (.B(\am_sdr0.cic2.integ_sample[4] ),
    .A(\am_sdr0.cic2.comb1_in_del[4] ),
    .X(_03020_));
 sg13g2_a21oi_2 _10216_ (.B1(_03013_),
    .Y(_03021_),
    .A2(_03016_),
    .A1(_03014_));
 sg13g2_nor2_1 _10217_ (.A(_03020_),
    .B(_03021_),
    .Y(_03022_));
 sg13g2_xnor2_1 _10218_ (.Y(_03023_),
    .A(_03020_),
    .B(_03021_));
 sg13g2_o21ai_1 _10219_ (.B1(net2009),
    .Y(_03024_),
    .A1(net1812),
    .A2(net2222));
 sg13g2_a21oi_1 _10220_ (.A1(net1812),
    .A2(_03023_),
    .Y(_00443_),
    .B1(_03024_));
 sg13g2_nor2_1 _10221_ (.A(_01464_),
    .B(\am_sdr0.cic2.integ_sample[5] ),
    .Y(_03025_));
 sg13g2_xor2_1 _10222_ (.B(\am_sdr0.cic2.integ_sample[5] ),
    .A(\am_sdr0.cic2.comb1_in_del[5] ),
    .X(_03026_));
 sg13g2_nor2_1 _10223_ (.A(_03019_),
    .B(_03022_),
    .Y(_03027_));
 sg13g2_xnor2_1 _10224_ (.Y(_03028_),
    .A(_03026_),
    .B(_03027_));
 sg13g2_o21ai_1 _10225_ (.B1(net2009),
    .Y(_03029_),
    .A1(net1807),
    .A2(net2386));
 sg13g2_a21oi_1 _10226_ (.A1(net1812),
    .A2(_03028_),
    .Y(_00444_),
    .B1(_03029_));
 sg13g2_nand2b_1 _10227_ (.Y(_03030_),
    .B(net2374),
    .A_N(\am_sdr0.cic2.comb1_in_del[6] ));
 sg13g2_xnor2_1 _10228_ (.Y(_03031_),
    .A(\am_sdr0.cic2.comb1_in_del[6] ),
    .B(net2869));
 sg13g2_a21oi_1 _10229_ (.A1(_01464_),
    .A2(\am_sdr0.cic2.integ_sample[5] ),
    .Y(_03032_),
    .B1(_03019_));
 sg13g2_o21ai_1 _10230_ (.B1(_03032_),
    .Y(_03033_),
    .A1(_03020_),
    .A2(_03021_));
 sg13g2_nor2b_1 _10231_ (.A(_03025_),
    .B_N(_03033_),
    .Y(_03034_));
 sg13g2_nand3b_1 _10232_ (.B(_03031_),
    .C(_03033_),
    .Y(_03035_),
    .A_N(_03025_));
 sg13g2_xnor2_1 _10233_ (.Y(_03036_),
    .A(_03031_),
    .B(_03034_));
 sg13g2_o21ai_1 _10234_ (.B1(net1978),
    .Y(_03037_),
    .A1(net1801),
    .A2(net2394));
 sg13g2_a21oi_1 _10235_ (.A1(net1801),
    .A2(_03036_),
    .Y(_00445_),
    .B1(_03037_));
 sg13g2_nand2b_1 _10236_ (.Y(_03038_),
    .B(\am_sdr0.cic2.integ_sample[7] ),
    .A_N(\am_sdr0.cic2.comb1_in_del[7] ));
 sg13g2_xor2_1 _10237_ (.B(\am_sdr0.cic2.integ_sample[7] ),
    .A(\am_sdr0.cic2.comb1_in_del[7] ),
    .X(_03039_));
 sg13g2_a21o_1 _10238_ (.A2(_03035_),
    .A1(_03030_),
    .B1(_03039_),
    .X(_03040_));
 sg13g2_nand3_1 _10239_ (.B(_03035_),
    .C(_03039_),
    .A(_03030_),
    .Y(_03041_));
 sg13g2_a21oi_1 _10240_ (.A1(_03040_),
    .A2(_03041_),
    .Y(_03042_),
    .B1(net1628));
 sg13g2_o21ai_1 _10241_ (.B1(net1978),
    .Y(_03043_),
    .A1(net1801),
    .A2(net2520));
 sg13g2_nor2_1 _10242_ (.A(_03042_),
    .B(_03043_),
    .Y(_00446_));
 sg13g2_nand2_2 _10243_ (.Y(_03044_),
    .A(_03038_),
    .B(_03040_));
 sg13g2_nor2_1 _10244_ (.A(\am_sdr0.cic2.comb1_in_del[8] ),
    .B(_01461_),
    .Y(_03045_));
 sg13g2_xnor2_1 _10245_ (.Y(_03046_),
    .A(\am_sdr0.cic2.comb1_in_del[8] ),
    .B(net2934));
 sg13g2_inv_1 _10246_ (.Y(_03047_),
    .A(_03046_));
 sg13g2_xnor2_1 _10247_ (.Y(_03048_),
    .A(_03044_),
    .B(_03046_));
 sg13g2_o21ai_1 _10248_ (.B1(net1975),
    .Y(_03049_),
    .A1(net1799),
    .A2(net2479));
 sg13g2_a21oi_1 _10249_ (.A1(net1799),
    .A2(_03048_),
    .Y(_00447_),
    .B1(_03049_));
 sg13g2_xor2_1 _10250_ (.B(net2361),
    .A(\am_sdr0.cic2.comb1_in_del[9] ),
    .X(_03050_));
 sg13g2_a21oi_1 _10251_ (.A1(_03044_),
    .A2(_03046_),
    .Y(_03051_),
    .B1(_03045_));
 sg13g2_xnor2_1 _10252_ (.Y(_03052_),
    .A(_03050_),
    .B(_03051_));
 sg13g2_o21ai_1 _10253_ (.B1(net1975),
    .Y(_03053_),
    .A1(net1799),
    .A2(net2281));
 sg13g2_a21oi_1 _10254_ (.A1(net1797),
    .A2(_03052_),
    .Y(_00448_),
    .B1(_03053_));
 sg13g2_nand2b_1 _10255_ (.Y(_03054_),
    .B(\am_sdr0.cic2.integ_sample[10] ),
    .A_N(\am_sdr0.cic2.comb1_in_del[10] ));
 sg13g2_xor2_1 _10256_ (.B(net2768),
    .A(\am_sdr0.cic2.comb1_in_del[10] ),
    .X(_03055_));
 sg13g2_a21oi_1 _10257_ (.A1(_01459_),
    .A2(\am_sdr0.cic2.integ_sample[9] ),
    .Y(_03056_),
    .B1(_03045_));
 sg13g2_a21oi_1 _10258_ (.A1(\am_sdr0.cic2.comb1_in_del[9] ),
    .A2(_01460_),
    .Y(_03057_),
    .B1(_03056_));
 sg13g2_nor2_1 _10259_ (.A(_03047_),
    .B(_03050_),
    .Y(_03058_));
 sg13g2_a21oi_1 _10260_ (.A1(_03044_),
    .A2(_03058_),
    .Y(_03059_),
    .B1(_03057_));
 sg13g2_xnor2_1 _10261_ (.Y(_03060_),
    .A(_03055_),
    .B(_03059_));
 sg13g2_o21ai_1 _10262_ (.B1(net1975),
    .Y(_03061_),
    .A1(net1799),
    .A2(net2496));
 sg13g2_a21oi_1 _10263_ (.A1(net1797),
    .A2(_03060_),
    .Y(_00449_),
    .B1(_03061_));
 sg13g2_nor2b_1 _10264_ (.A(\am_sdr0.cic2.integ_sample[11] ),
    .B_N(\am_sdr0.cic2.comb1_in_del[11] ),
    .Y(_03062_));
 sg13g2_nand2b_1 _10265_ (.Y(_03063_),
    .B(\am_sdr0.cic2.integ_sample[11] ),
    .A_N(\am_sdr0.cic2.comb1_in_del[11] ));
 sg13g2_nand2b_1 _10266_ (.Y(_03064_),
    .B(_03063_),
    .A_N(_03062_));
 sg13g2_o21ai_1 _10267_ (.B1(_03054_),
    .Y(_03065_),
    .A1(_03055_),
    .A2(_03059_));
 sg13g2_xor2_1 _10268_ (.B(_03065_),
    .A(_03064_),
    .X(_03066_));
 sg13g2_o21ai_1 _10269_ (.B1(net1975),
    .Y(_03067_),
    .A1(net1798),
    .A2(net2251));
 sg13g2_a21oi_1 _10270_ (.A1(net1798),
    .A2(_03066_),
    .Y(_00450_),
    .B1(_03067_));
 sg13g2_nor2_1 _10271_ (.A(\am_sdr0.cic2.comb1_in_del[12] ),
    .B(_01456_),
    .Y(_03068_));
 sg13g2_xor2_1 _10272_ (.B(\am_sdr0.cic2.integ_sample[12] ),
    .A(\am_sdr0.cic2.comb1_in_del[12] ),
    .X(_03069_));
 sg13g2_inv_1 _10273_ (.Y(_03070_),
    .A(_03069_));
 sg13g2_nor2_1 _10274_ (.A(_03055_),
    .B(_03064_),
    .Y(_03071_));
 sg13g2_o21ai_1 _10275_ (.B1(_03063_),
    .Y(_03072_),
    .A1(_03054_),
    .A2(_03062_));
 sg13g2_a21o_2 _10276_ (.A2(_03071_),
    .A1(_03057_),
    .B1(_03072_),
    .X(_03073_));
 sg13g2_nand2_1 _10277_ (.Y(_03074_),
    .A(_03058_),
    .B(_03071_));
 sg13g2_a21oi_2 _10278_ (.B1(_03074_),
    .Y(_03075_),
    .A2(_03040_),
    .A1(_03038_));
 sg13g2_nor3_1 _10279_ (.A(_03070_),
    .B(_03073_),
    .C(_03075_),
    .Y(_03076_));
 sg13g2_o21ai_1 _10280_ (.B1(_03070_),
    .Y(_03077_),
    .A1(_03073_),
    .A2(_03075_));
 sg13g2_nand2b_1 _10281_ (.Y(_03078_),
    .B(_03077_),
    .A_N(_03076_));
 sg13g2_o21ai_1 _10282_ (.B1(net2008),
    .Y(_03079_),
    .A1(net1802),
    .A2(net2794));
 sg13g2_a21oi_1 _10283_ (.A1(net1802),
    .A2(_03078_),
    .Y(_00451_),
    .B1(_03079_));
 sg13g2_nor2_1 _10284_ (.A(_01455_),
    .B(\am_sdr0.cic2.integ_sample[13] ),
    .Y(_03080_));
 sg13g2_xor2_1 _10285_ (.B(\am_sdr0.cic2.integ_sample[13] ),
    .A(\am_sdr0.cic2.comb1_in_del[13] ),
    .X(_03081_));
 sg13g2_nor2b_1 _10286_ (.A(_03068_),
    .B_N(_03077_),
    .Y(_03082_));
 sg13g2_xnor2_1 _10287_ (.Y(_03083_),
    .A(_03081_),
    .B(_03082_));
 sg13g2_o21ai_1 _10288_ (.B1(net2008),
    .Y(_03084_),
    .A1(net1819),
    .A2(net2538));
 sg13g2_a21oi_1 _10289_ (.A1(net1804),
    .A2(_03083_),
    .Y(_00452_),
    .B1(_03084_));
 sg13g2_nor2_1 _10290_ (.A(net2884),
    .B(_01454_),
    .Y(_03085_));
 sg13g2_nand2_1 _10291_ (.Y(_03086_),
    .A(net2304),
    .B(_01454_));
 sg13g2_nand2b_2 _10292_ (.Y(_03087_),
    .B(_03086_),
    .A_N(_03085_));
 sg13g2_a21oi_1 _10293_ (.A1(_01455_),
    .A2(\am_sdr0.cic2.integ_sample[13] ),
    .Y(_03088_),
    .B1(_03068_));
 sg13g2_a21oi_1 _10294_ (.A1(_03077_),
    .A2(_03088_),
    .Y(_03089_),
    .B1(_03080_));
 sg13g2_xor2_1 _10295_ (.B(_03089_),
    .A(_03087_),
    .X(_03090_));
 sg13g2_o21ai_1 _10296_ (.B1(net2008),
    .Y(_03091_),
    .A1(net1819),
    .A2(net2567));
 sg13g2_a21oi_1 _10297_ (.A1(net1808),
    .A2(_03090_),
    .Y(_00453_),
    .B1(_03091_));
 sg13g2_nand2_1 _10298_ (.Y(_03092_),
    .A(\am_sdr0.cic2.comb1_in_del[15] ),
    .B(_01453_));
 sg13g2_nor2_1 _10299_ (.A(\am_sdr0.cic2.comb1_in_del[15] ),
    .B(_01453_),
    .Y(_03093_));
 sg13g2_xor2_1 _10300_ (.B(\am_sdr0.cic2.integ_sample[15] ),
    .A(\am_sdr0.cic2.comb1_in_del[15] ),
    .X(_03094_));
 sg13g2_a21oi_1 _10301_ (.A1(_03086_),
    .A2(_03089_),
    .Y(_03095_),
    .B1(_03085_));
 sg13g2_xnor2_1 _10302_ (.Y(_03096_),
    .A(_03094_),
    .B(_03095_));
 sg13g2_o21ai_1 _10303_ (.B1(net2008),
    .Y(_03097_),
    .A1(net1808),
    .A2(net2855));
 sg13g2_a21oi_1 _10304_ (.A1(net1807),
    .A2(_03096_),
    .Y(_00454_),
    .B1(_03097_));
 sg13g2_nor2_1 _10305_ (.A(\am_sdr0.cic2.comb1_in_del[16] ),
    .B(_01452_),
    .Y(_03098_));
 sg13g2_xor2_1 _10306_ (.B(\am_sdr0.cic2.integ_sample[16] ),
    .A(\am_sdr0.cic2.comb1_in_del[16] ),
    .X(_03099_));
 sg13g2_nor4_2 _10307_ (.A(_03069_),
    .B(_03081_),
    .C(_03087_),
    .Y(_03100_),
    .D(_03094_));
 sg13g2_nor4_1 _10308_ (.A(_03080_),
    .B(_03087_),
    .C(_03088_),
    .D(_03094_),
    .Y(_03101_));
 sg13g2_a221oi_1 _10309_ (.B2(_03073_),
    .C1(_03093_),
    .B1(_03100_),
    .A1(_03085_),
    .Y(_03102_),
    .A2(_03092_));
 sg13g2_nand2b_1 _10310_ (.Y(_03103_),
    .B(_03102_),
    .A_N(_03101_));
 sg13g2_a21oi_2 _10311_ (.B1(_03103_),
    .Y(_03104_),
    .A2(_03100_),
    .A1(_03075_));
 sg13g2_nor2_1 _10312_ (.A(_03099_),
    .B(_03104_),
    .Y(_03105_));
 sg13g2_xnor2_1 _10313_ (.Y(_03106_),
    .A(_03099_),
    .B(_03104_));
 sg13g2_o21ai_1 _10314_ (.B1(net2010),
    .Y(_03107_),
    .A1(net1809),
    .A2(net2631));
 sg13g2_a21oi_1 _10315_ (.A1(net1809),
    .A2(_03106_),
    .Y(_00455_),
    .B1(_03107_));
 sg13g2_nand2_1 _10316_ (.Y(_03108_),
    .A(\am_sdr0.cic2.comb1_in_del[17] ),
    .B(_01451_));
 sg13g2_nor2_1 _10317_ (.A(\am_sdr0.cic2.comb1_in_del[17] ),
    .B(_01451_),
    .Y(_03109_));
 sg13g2_xnor2_1 _10318_ (.Y(_03110_),
    .A(\am_sdr0.cic2.comb1_in_del[17] ),
    .B(\am_sdr0.cic2.integ_sample[17] ));
 sg13g2_nor2_1 _10319_ (.A(_03098_),
    .B(_03105_),
    .Y(_03111_));
 sg13g2_xor2_1 _10320_ (.B(_03111_),
    .A(_03110_),
    .X(_03112_));
 sg13g2_o21ai_1 _10321_ (.B1(net2010),
    .Y(_03113_),
    .A1(net1818),
    .A2(net2659));
 sg13g2_a21oi_1 _10322_ (.A1(net1818),
    .A2(_03112_),
    .Y(_00456_),
    .B1(_03113_));
 sg13g2_nor2_1 _10323_ (.A(net2499),
    .B(_01450_),
    .Y(_03114_));
 sg13g2_xnor2_1 _10324_ (.Y(_03115_),
    .A(net2499),
    .B(net2342));
 sg13g2_nand2b_1 _10325_ (.Y(_03116_),
    .B(_03110_),
    .A_N(_03099_));
 sg13g2_a21oi_1 _10326_ (.A1(_03098_),
    .A2(_03108_),
    .Y(_03117_),
    .B1(_03109_));
 sg13g2_o21ai_1 _10327_ (.B1(_03117_),
    .Y(_03118_),
    .A1(_03104_),
    .A2(_03116_));
 sg13g2_xnor2_1 _10328_ (.Y(_03119_),
    .A(_03115_),
    .B(_03118_));
 sg13g2_o21ai_1 _10329_ (.B1(net2012),
    .Y(_03120_),
    .A1(net1816),
    .A2(net2245));
 sg13g2_a21oi_1 _10330_ (.A1(net1816),
    .A2(_03119_),
    .Y(_00457_),
    .B1(_03120_));
 sg13g2_a21oi_1 _10331_ (.A1(_03115_),
    .A2(_03118_),
    .Y(_03121_),
    .B1(_03114_));
 sg13g2_xor2_1 _10332_ (.B(net1486),
    .A(net2669),
    .X(_03122_));
 sg13g2_inv_1 _10333_ (.Y(_03123_),
    .A(_03122_));
 sg13g2_nand2b_1 _10334_ (.Y(_03124_),
    .B(_03122_),
    .A_N(_03121_));
 sg13g2_a21oi_1 _10335_ (.A1(_03121_),
    .A2(_03123_),
    .Y(_03125_),
    .B1(net1630));
 sg13g2_a221oi_1 _10336_ (.B2(_03125_),
    .C1(net1891),
    .B1(_03124_),
    .A1(net1630),
    .Y(_00458_),
    .A2(_01426_));
 sg13g2_o21ai_1 _10337_ (.B1(net2013),
    .Y(_03126_),
    .A1(net1630),
    .A2(\am_sdr0.cic2.integ_sample[0] ));
 sg13g2_a21oi_1 _10338_ (.A1(net1630),
    .A2(_01469_),
    .Y(_00459_),
    .B1(_03126_));
 sg13g2_o21ai_1 _10339_ (.B1(net2013),
    .Y(_03127_),
    .A1(net1813),
    .A2(\am_sdr0.cic2.comb1_in_del[1] ));
 sg13g2_a21oi_1 _10340_ (.A1(net1813),
    .A2(_01468_),
    .Y(_00460_),
    .B1(_03127_));
 sg13g2_o21ai_1 _10341_ (.B1(net2014),
    .Y(_03128_),
    .A1(net1813),
    .A2(\am_sdr0.cic2.comb1_in_del[2] ));
 sg13g2_a21oi_1 _10342_ (.A1(net1813),
    .A2(_01467_),
    .Y(_00461_),
    .B1(_03128_));
 sg13g2_o21ai_1 _10343_ (.B1(net2004),
    .Y(_03129_),
    .A1(net1812),
    .A2(net2535));
 sg13g2_a21oi_1 _10344_ (.A1(net1812),
    .A2(_01466_),
    .Y(_00462_),
    .B1(_03129_));
 sg13g2_o21ai_1 _10345_ (.B1(net1973),
    .Y(_03130_),
    .A1(net1803),
    .A2(net2564));
 sg13g2_a21oi_1 _10346_ (.A1(net1803),
    .A2(_01465_),
    .Y(_00463_),
    .B1(_03130_));
 sg13g2_o21ai_1 _10347_ (.B1(net1973),
    .Y(_03131_),
    .A1(net1628),
    .A2(\am_sdr0.cic2.integ_sample[5] ));
 sg13g2_a21oi_1 _10348_ (.A1(net1628),
    .A2(_01464_),
    .Y(_00464_),
    .B1(_03131_));
 sg13g2_o21ai_1 _10349_ (.B1(net1975),
    .Y(_03132_),
    .A1(net1800),
    .A2(\am_sdr0.cic2.comb1_in_del[6] ));
 sg13g2_a21oi_1 _10350_ (.A1(net1800),
    .A2(_01463_),
    .Y(_00465_),
    .B1(_03132_));
 sg13g2_o21ai_1 _10351_ (.B1(net1975),
    .Y(_03133_),
    .A1(net1800),
    .A2(\am_sdr0.cic2.comb1_in_del[7] ));
 sg13g2_a21oi_1 _10352_ (.A1(net1800),
    .A2(_01462_),
    .Y(_00466_),
    .B1(_03133_));
 sg13g2_o21ai_1 _10353_ (.B1(net1968),
    .Y(_03134_),
    .A1(net1797),
    .A2(\am_sdr0.cic2.comb1_in_del[8] ));
 sg13g2_a21oi_1 _10354_ (.A1(net1797),
    .A2(_01461_),
    .Y(_00467_),
    .B1(_03134_));
 sg13g2_o21ai_1 _10355_ (.B1(net1968),
    .Y(_03135_),
    .A1(net1797),
    .A2(\am_sdr0.cic2.comb1_in_del[9] ));
 sg13g2_a21oi_1 _10356_ (.A1(net1797),
    .A2(_01460_),
    .Y(_00468_),
    .B1(_03135_));
 sg13g2_o21ai_1 _10357_ (.B1(net1968),
    .Y(_03136_),
    .A1(net1797),
    .A2(\am_sdr0.cic2.comb1_in_del[10] ));
 sg13g2_a21oi_1 _10358_ (.A1(net1797),
    .A2(_01458_),
    .Y(_00469_),
    .B1(_03136_));
 sg13g2_o21ai_1 _10359_ (.B1(net1975),
    .Y(_03137_),
    .A1(net1800),
    .A2(\am_sdr0.cic2.comb1_in_del[11] ));
 sg13g2_a21oi_1 _10360_ (.A1(net1800),
    .A2(_01457_),
    .Y(_00470_),
    .B1(_03137_));
 sg13g2_o21ai_1 _10361_ (.B1(net1978),
    .Y(_03138_),
    .A1(net1802),
    .A2(net2466));
 sg13g2_a21oi_1 _10362_ (.A1(net1802),
    .A2(_01456_),
    .Y(_00471_),
    .B1(_03138_));
 sg13g2_o21ai_1 _10363_ (.B1(net1978),
    .Y(_03139_),
    .A1(net1628),
    .A2(\am_sdr0.cic2.integ_sample[13] ));
 sg13g2_a21oi_1 _10364_ (.A1(net1628),
    .A2(_01455_),
    .Y(_00472_),
    .B1(_03139_));
 sg13g2_o21ai_1 _10365_ (.B1(net2009),
    .Y(_03140_),
    .A1(net1807),
    .A2(net2304));
 sg13g2_a21oi_1 _10366_ (.A1(net1807),
    .A2(_01454_),
    .Y(_00473_),
    .B1(_03140_));
 sg13g2_o21ai_1 _10367_ (.B1(net2009),
    .Y(_03141_),
    .A1(net1807),
    .A2(net2761));
 sg13g2_a21oi_1 _10368_ (.A1(net1807),
    .A2(_01453_),
    .Y(_00474_),
    .B1(_03141_));
 sg13g2_o21ai_1 _10369_ (.B1(net2011),
    .Y(_03142_),
    .A1(net1809),
    .A2(net2525));
 sg13g2_a21oi_1 _10370_ (.A1(net1809),
    .A2(_01452_),
    .Y(_00475_),
    .B1(_03142_));
 sg13g2_o21ai_1 _10371_ (.B1(net2011),
    .Y(_03143_),
    .A1(net1816),
    .A2(net2795));
 sg13g2_a21oi_1 _10372_ (.A1(net1816),
    .A2(_01451_),
    .Y(_00476_),
    .B1(_03143_));
 sg13g2_o21ai_1 _10373_ (.B1(net2011),
    .Y(_03144_),
    .A1(net1816),
    .A2(net2499));
 sg13g2_a21oi_1 _10374_ (.A1(net1816),
    .A2(_01450_),
    .Y(_00477_),
    .B1(_03144_));
 sg13g2_o21ai_1 _10375_ (.B1(net2013),
    .Y(_03145_),
    .A1(net1814),
    .A2(\am_sdr0.cic2.comb1_in_del[19] ));
 sg13g2_a21oi_1 _10376_ (.A1(net1813),
    .A2(_01449_),
    .Y(_00478_),
    .B1(_03145_));
 sg13g2_nand2b_1 _10377_ (.Y(_03146_),
    .B(net2416),
    .A_N(net2383));
 sg13g2_a21oi_1 _10378_ (.A1(_01447_),
    .A2(net2383),
    .Y(_03147_),
    .B1(net1630));
 sg13g2_a221oi_1 _10379_ (.B2(net2384),
    .C1(net1891),
    .B1(_03146_),
    .A1(net1630),
    .Y(_00479_),
    .A2(_01417_));
 sg13g2_nor2b_1 _10380_ (.A(net2639),
    .B_N(\am_sdr0.cic2.comb1[1] ),
    .Y(_03148_));
 sg13g2_xnor2_1 _10381_ (.Y(_03149_),
    .A(net2639),
    .B(net2312));
 sg13g2_xnor2_1 _10382_ (.Y(_03150_),
    .A(_03146_),
    .B(_03149_));
 sg13g2_o21ai_1 _10383_ (.B1(net2015),
    .Y(_03151_),
    .A1(net1817),
    .A2(net2083));
 sg13g2_a21oi_1 _10384_ (.A1(net1817),
    .A2(_03150_),
    .Y(_00480_),
    .B1(_03151_));
 sg13g2_nand2b_1 _10385_ (.Y(_03152_),
    .B(\am_sdr0.cic2.comb1[2] ),
    .A_N(\am_sdr0.cic2.comb2_in_del[2] ));
 sg13g2_xor2_1 _10386_ (.B(\am_sdr0.cic2.comb1[2] ),
    .A(\am_sdr0.cic2.comb2_in_del[2] ),
    .X(_03153_));
 sg13g2_a21oi_1 _10387_ (.A1(_03146_),
    .A2(_03149_),
    .Y(_03154_),
    .B1(_03148_));
 sg13g2_xnor2_1 _10388_ (.Y(_03155_),
    .A(_03153_),
    .B(_03154_));
 sg13g2_o21ai_1 _10389_ (.B1(net2015),
    .Y(_03156_),
    .A1(net1817),
    .A2(net2871));
 sg13g2_a21oi_1 _10390_ (.A1(net1817),
    .A2(_03155_),
    .Y(_00481_),
    .B1(_03156_));
 sg13g2_nor2_1 _10391_ (.A(\am_sdr0.cic2.comb2_in_del[3] ),
    .B(_01444_),
    .Y(_03157_));
 sg13g2_nand2_1 _10392_ (.Y(_03158_),
    .A(\am_sdr0.cic2.comb2_in_del[3] ),
    .B(_01444_));
 sg13g2_nor2b_1 _10393_ (.A(_03157_),
    .B_N(_03158_),
    .Y(_03159_));
 sg13g2_o21ai_1 _10394_ (.B1(_03152_),
    .Y(_03160_),
    .A1(_03153_),
    .A2(_03154_));
 sg13g2_xnor2_1 _10395_ (.Y(_03161_),
    .A(_03159_),
    .B(_03160_));
 sg13g2_o21ai_1 _10396_ (.B1(net2011),
    .Y(_03162_),
    .A1(net1816),
    .A2(net2839));
 sg13g2_a21oi_1 _10397_ (.A1(net1816),
    .A2(_03161_),
    .Y(_00482_),
    .B1(_03162_));
 sg13g2_nor2_1 _10398_ (.A(\am_sdr0.cic2.comb2_in_del[4] ),
    .B(_01443_),
    .Y(_03163_));
 sg13g2_xor2_1 _10399_ (.B(net2222),
    .A(\am_sdr0.cic2.comb2_in_del[4] ),
    .X(_03164_));
 sg13g2_a21oi_2 _10400_ (.B1(_03157_),
    .Y(_03165_),
    .A2(_03160_),
    .A1(_03158_));
 sg13g2_nor2_1 _10401_ (.A(_03164_),
    .B(_03165_),
    .Y(_03166_));
 sg13g2_xnor2_1 _10402_ (.Y(_03167_),
    .A(_03164_),
    .B(_03165_));
 sg13g2_o21ai_1 _10403_ (.B1(net2011),
    .Y(_03168_),
    .A1(net1810),
    .A2(net2529));
 sg13g2_a21oi_1 _10404_ (.A1(net1809),
    .A2(_03167_),
    .Y(_00483_),
    .B1(_03168_));
 sg13g2_nand2b_1 _10405_ (.Y(_03169_),
    .B(net2386),
    .A_N(net2750));
 sg13g2_nand2_1 _10406_ (.Y(_03170_),
    .A(net2750),
    .B(_01442_));
 sg13g2_nor2_1 _10407_ (.A(_03163_),
    .B(_03166_),
    .Y(_03171_));
 sg13g2_a21oi_1 _10408_ (.A1(_03169_),
    .A2(_03170_),
    .Y(_03172_),
    .B1(_03171_));
 sg13g2_nand3_1 _10409_ (.B(_03170_),
    .C(_03171_),
    .A(_03169_),
    .Y(_03173_));
 sg13g2_nor2_1 _10410_ (.A(net1632),
    .B(_03172_),
    .Y(_03174_));
 sg13g2_a221oi_1 _10411_ (.B2(_03174_),
    .C1(net1891),
    .B1(_03173_),
    .A1(net1632),
    .Y(_00484_),
    .A2(_01411_));
 sg13g2_nand2b_1 _10412_ (.Y(_03175_),
    .B(\am_sdr0.cic2.comb1[6] ),
    .A_N(\am_sdr0.cic2.comb2_in_del[6] ));
 sg13g2_xnor2_1 _10413_ (.Y(_03176_),
    .A(\am_sdr0.cic2.comb2_in_del[6] ),
    .B(\am_sdr0.cic2.comb1[6] ));
 sg13g2_nor2b_1 _10414_ (.A(_03163_),
    .B_N(_03169_),
    .Y(_03177_));
 sg13g2_o21ai_1 _10415_ (.B1(_03177_),
    .Y(_03178_),
    .A1(_03164_),
    .A2(_03165_));
 sg13g2_nand3_1 _10416_ (.B(_03176_),
    .C(_03178_),
    .A(_03170_),
    .Y(_03179_));
 sg13g2_a21o_1 _10417_ (.A2(_03178_),
    .A1(_03170_),
    .B1(_03176_),
    .X(_03180_));
 sg13g2_nand2_1 _10418_ (.Y(_03181_),
    .A(_03179_),
    .B(_03180_));
 sg13g2_o21ai_1 _10419_ (.B1(net2009),
    .Y(_03182_),
    .A1(net1808),
    .A2(net2876));
 sg13g2_a21oi_1 _10420_ (.A1(net1808),
    .A2(_03181_),
    .Y(_00485_),
    .B1(_03182_));
 sg13g2_nand2b_1 _10421_ (.Y(_03183_),
    .B(\am_sdr0.cic2.comb1[7] ),
    .A_N(\am_sdr0.cic2.comb2_in_del[7] ));
 sg13g2_xor2_1 _10422_ (.B(\am_sdr0.cic2.comb1[7] ),
    .A(\am_sdr0.cic2.comb2_in_del[7] ),
    .X(_03184_));
 sg13g2_a21o_1 _10423_ (.A2(_03179_),
    .A1(_03175_),
    .B1(_03184_),
    .X(_03185_));
 sg13g2_nand3_1 _10424_ (.B(_03179_),
    .C(_03184_),
    .A(_03175_),
    .Y(_03186_));
 sg13g2_a21oi_1 _10425_ (.A1(_03185_),
    .A2(_03186_),
    .Y(_03187_),
    .B1(net1628));
 sg13g2_o21ai_1 _10426_ (.B1(net1978),
    .Y(_03188_),
    .A1(net1802),
    .A2(net2785));
 sg13g2_nor2_1 _10427_ (.A(_03187_),
    .B(_03188_),
    .Y(_00486_));
 sg13g2_nand2_1 _10428_ (.Y(_03189_),
    .A(_03183_),
    .B(_03185_));
 sg13g2_nand2b_1 _10429_ (.Y(_03190_),
    .B(net3310),
    .A_N(\am_sdr0.cic2.comb2_in_del[8] ));
 sg13g2_xnor2_1 _10430_ (.Y(_03191_),
    .A(\am_sdr0.cic2.comb2_in_del[8] ),
    .B(\am_sdr0.cic2.comb1[8] ));
 sg13g2_inv_1 _10431_ (.Y(_03192_),
    .A(_03191_));
 sg13g2_nand2_1 _10432_ (.Y(_03193_),
    .A(_03189_),
    .B(_03191_));
 sg13g2_xnor2_1 _10433_ (.Y(_03194_),
    .A(_03189_),
    .B(_03191_));
 sg13g2_o21ai_1 _10434_ (.B1(net1977),
    .Y(_03195_),
    .A1(net1802),
    .A2(net2325));
 sg13g2_a21oi_1 _10435_ (.A1(net1801),
    .A2(_03194_),
    .Y(_00487_),
    .B1(_03195_));
 sg13g2_nor2b_1 _10436_ (.A(\am_sdr0.cic2.comb1[9] ),
    .B_N(\am_sdr0.cic2.comb2_in_del[9] ),
    .Y(_03196_));
 sg13g2_nand2b_1 _10437_ (.Y(_03197_),
    .B(\am_sdr0.cic2.comb1[9] ),
    .A_N(\am_sdr0.cic2.comb2_in_del[9] ));
 sg13g2_nand2b_1 _10438_ (.Y(_03198_),
    .B(_03197_),
    .A_N(_03196_));
 sg13g2_nand2_1 _10439_ (.Y(_03199_),
    .A(_03190_),
    .B(_03193_));
 sg13g2_o21ai_1 _10440_ (.B1(net1805),
    .Y(_03200_),
    .A1(_03198_),
    .A2(_03199_));
 sg13g2_a21oi_1 _10441_ (.A1(_03198_),
    .A2(_03199_),
    .Y(_03201_),
    .B1(_03200_));
 sg13g2_o21ai_1 _10442_ (.B1(net1977),
    .Y(_03202_),
    .A1(net1805),
    .A2(net2172));
 sg13g2_nor2_1 _10443_ (.A(_03201_),
    .B(_03202_),
    .Y(_00488_));
 sg13g2_nand2b_1 _10444_ (.Y(_03203_),
    .B(\am_sdr0.cic2.comb1[10] ),
    .A_N(\am_sdr0.cic2.comb2_in_del[10] ));
 sg13g2_xor2_1 _10445_ (.B(\am_sdr0.cic2.comb1[10] ),
    .A(\am_sdr0.cic2.comb2_in_del[10] ),
    .X(_03204_));
 sg13g2_o21ai_1 _10446_ (.B1(_03197_),
    .Y(_03205_),
    .A1(_03190_),
    .A2(_03196_));
 sg13g2_nor2_1 _10447_ (.A(_03192_),
    .B(_03198_),
    .Y(_03206_));
 sg13g2_a21oi_1 _10448_ (.A1(_03189_),
    .A2(_03206_),
    .Y(_03207_),
    .B1(_03205_));
 sg13g2_xnor2_1 _10449_ (.Y(_03208_),
    .A(_03204_),
    .B(_03207_));
 sg13g2_o21ai_1 _10450_ (.B1(net1977),
    .Y(_03209_),
    .A1(net1805),
    .A2(net2333));
 sg13g2_a21oi_1 _10451_ (.A1(net1805),
    .A2(_03208_),
    .Y(_00489_),
    .B1(_03209_));
 sg13g2_nor2b_1 _10452_ (.A(\am_sdr0.cic2.comb1[11] ),
    .B_N(\am_sdr0.cic2.comb2_in_del[11] ),
    .Y(_03210_));
 sg13g2_nand2b_1 _10453_ (.Y(_03211_),
    .B(\am_sdr0.cic2.comb1[11] ),
    .A_N(\am_sdr0.cic2.comb2_in_del[11] ));
 sg13g2_nand2b_1 _10454_ (.Y(_03212_),
    .B(_03211_),
    .A_N(_03210_));
 sg13g2_o21ai_1 _10455_ (.B1(_03203_),
    .Y(_03213_),
    .A1(_03204_),
    .A2(_03207_));
 sg13g2_or2_1 _10456_ (.X(_03214_),
    .B(_03213_),
    .A(_03212_));
 sg13g2_a21oi_1 _10457_ (.A1(_03212_),
    .A2(_03213_),
    .Y(_03215_),
    .B1(net1629));
 sg13g2_a221oi_1 _10458_ (.B2(_03215_),
    .C1(net1889),
    .B1(_03214_),
    .A1(net1629),
    .Y(_00490_),
    .A2(_01403_));
 sg13g2_xor2_1 _10459_ (.B(\am_sdr0.cic2.comb1[12] ),
    .A(\am_sdr0.cic2.comb2_in_del[12] ),
    .X(_03216_));
 sg13g2_inv_1 _10460_ (.Y(_03217_),
    .A(_03216_));
 sg13g2_nor2_1 _10461_ (.A(_03204_),
    .B(_03212_),
    .Y(_03218_));
 sg13g2_o21ai_1 _10462_ (.B1(_03211_),
    .Y(_03219_),
    .A1(_03203_),
    .A2(_03210_));
 sg13g2_a21o_2 _10463_ (.A2(_03218_),
    .A1(_03205_),
    .B1(_03219_),
    .X(_03220_));
 sg13g2_nand2_1 _10464_ (.Y(_03221_),
    .A(_03206_),
    .B(_03218_));
 sg13g2_a21oi_2 _10465_ (.B1(_03221_),
    .Y(_03222_),
    .A2(_03185_),
    .A1(_03183_));
 sg13g2_o21ai_1 _10466_ (.B1(_03217_),
    .Y(_03223_),
    .A1(_03220_),
    .A2(_03222_));
 sg13g2_or3_1 _10467_ (.A(_03217_),
    .B(_03220_),
    .C(_03222_),
    .X(_03224_));
 sg13g2_nand2_1 _10468_ (.Y(_03225_),
    .A(_03223_),
    .B(_03224_));
 sg13g2_o21ai_1 _10469_ (.B1(net1994),
    .Y(_03226_),
    .A1(net1806),
    .A2(net2674));
 sg13g2_a21oi_1 _10470_ (.A1(net1806),
    .A2(_03225_),
    .Y(_00491_),
    .B1(_03226_));
 sg13g2_nor2_1 _10471_ (.A(_01432_),
    .B(\am_sdr0.cic2.comb1[13] ),
    .Y(_03227_));
 sg13g2_xor2_1 _10472_ (.B(net2538),
    .A(\am_sdr0.cic2.comb2_in_del[13] ),
    .X(_03228_));
 sg13g2_o21ai_1 _10473_ (.B1(_03223_),
    .Y(_03229_),
    .A1(net2675),
    .A2(_01435_));
 sg13g2_o21ai_1 _10474_ (.B1(net1820),
    .Y(_03230_),
    .A1(_03228_),
    .A2(_03229_));
 sg13g2_a21oi_1 _10475_ (.A1(_03228_),
    .A2(net2676),
    .Y(_03231_),
    .B1(_03230_));
 sg13g2_o21ai_1 _10476_ (.B1(net2019),
    .Y(_03232_),
    .A1(net1819),
    .A2(net2509));
 sg13g2_nor2_1 _10477_ (.A(net2677),
    .B(_03232_),
    .Y(_00492_));
 sg13g2_nor2_1 _10478_ (.A(net2952),
    .B(_01431_),
    .Y(_03233_));
 sg13g2_xor2_1 _10479_ (.B(net3320),
    .A(\am_sdr0.cic2.comb2_in_del[14] ),
    .X(_03234_));
 sg13g2_a22oi_1 _10480_ (.Y(_03235_),
    .B1(_01434_),
    .B2(\am_sdr0.cic2.comb1[12] ),
    .A2(\am_sdr0.cic2.comb1[13] ),
    .A1(_01432_));
 sg13g2_a21oi_1 _10481_ (.A1(_03223_),
    .A2(_03235_),
    .Y(_03236_),
    .B1(net2539));
 sg13g2_a221oi_1 _10482_ (.B2(_03235_),
    .C1(_03234_),
    .B1(_03223_),
    .A1(\am_sdr0.cic2.comb2_in_del[13] ),
    .Y(_03237_),
    .A2(_01433_));
 sg13g2_xor2_1 _10483_ (.B(_03236_),
    .A(_03234_),
    .X(_03238_));
 sg13g2_o21ai_1 _10484_ (.B1(net2019),
    .Y(_03239_),
    .A1(net1819),
    .A2(net2314));
 sg13g2_a21oi_1 _10485_ (.A1(net1820),
    .A2(_03238_),
    .Y(_00493_),
    .B1(_03239_));
 sg13g2_nand2_1 _10486_ (.Y(_03240_),
    .A(\am_sdr0.cic2.comb2_in_del[15] ),
    .B(_01430_));
 sg13g2_nor2_1 _10487_ (.A(\am_sdr0.cic2.comb2_in_del[15] ),
    .B(_01430_),
    .Y(_03241_));
 sg13g2_xor2_1 _10488_ (.B(net2855),
    .A(\am_sdr0.cic2.comb2_in_del[15] ),
    .X(_03242_));
 sg13g2_o21ai_1 _10489_ (.B1(_03242_),
    .Y(_03243_),
    .A1(_03233_),
    .A2(_03237_));
 sg13g2_nor3_1 _10490_ (.A(_03233_),
    .B(_03237_),
    .C(_03242_),
    .Y(_03244_));
 sg13g2_nor2_1 _10491_ (.A(net1629),
    .B(_03244_),
    .Y(_03245_));
 sg13g2_a221oi_1 _10492_ (.B2(_03245_),
    .C1(net1892),
    .B1(net2953),
    .A1(net1629),
    .Y(_00494_),
    .A2(_01399_));
 sg13g2_nor2_1 _10493_ (.A(\am_sdr0.cic2.comb2_in_del[16] ),
    .B(_01429_),
    .Y(_03246_));
 sg13g2_xnor2_1 _10494_ (.Y(_03247_),
    .A(\am_sdr0.cic2.comb2_in_del[16] ),
    .B(net2866));
 sg13g2_or4_1 _10495_ (.A(_03216_),
    .B(_03228_),
    .C(_03234_),
    .D(_03242_),
    .X(_03248_));
 sg13g2_inv_1 _10496_ (.Y(_03249_),
    .A(_03248_));
 sg13g2_nor4_1 _10497_ (.A(_03227_),
    .B(_03234_),
    .C(_03235_),
    .D(_03242_),
    .Y(_03250_));
 sg13g2_a221oi_1 _10498_ (.B2(_03220_),
    .C1(_03241_),
    .B1(_03249_),
    .A1(_03233_),
    .Y(_03251_),
    .A2(_03240_));
 sg13g2_nand2b_1 _10499_ (.Y(_03252_),
    .B(_03251_),
    .A_N(_03250_));
 sg13g2_a21o_1 _10500_ (.A2(_03249_),
    .A1(_03222_),
    .B1(_03252_),
    .X(_03253_));
 sg13g2_xnor2_1 _10501_ (.Y(_03254_),
    .A(_03247_),
    .B(_03253_));
 sg13g2_o21ai_1 _10502_ (.B1(net2010),
    .Y(_03255_),
    .A1(net1821),
    .A2(net2344));
 sg13g2_a21oi_1 _10503_ (.A1(net1826),
    .A2(_03254_),
    .Y(_00495_),
    .B1(_03255_));
 sg13g2_nand2_1 _10504_ (.Y(_03256_),
    .A(\am_sdr0.cic2.comb2_in_del[17] ),
    .B(_01428_));
 sg13g2_nor2_1 _10505_ (.A(\am_sdr0.cic2.comb2_in_del[17] ),
    .B(_01428_),
    .Y(_03257_));
 sg13g2_xnor2_1 _10506_ (.Y(_03258_),
    .A(\am_sdr0.cic2.comb2_in_del[17] ),
    .B(net2659));
 sg13g2_a21oi_1 _10507_ (.A1(_03247_),
    .A2(_03253_),
    .Y(_03259_),
    .B1(_03246_));
 sg13g2_or2_1 _10508_ (.X(_03260_),
    .B(_03259_),
    .A(_03258_));
 sg13g2_a21oi_1 _10509_ (.A1(_03258_),
    .A2(_03259_),
    .Y(_03261_),
    .B1(net1633));
 sg13g2_a221oi_1 _10510_ (.B2(_03261_),
    .C1(net1892),
    .B1(_03260_),
    .A1(net1633),
    .Y(_00496_),
    .A2(_01397_));
 sg13g2_nand2b_1 _10511_ (.Y(_03262_),
    .B(net2245),
    .A_N(\am_sdr0.cic2.comb2_in_del[18] ));
 sg13g2_xor2_1 _10512_ (.B(net2789),
    .A(\am_sdr0.cic2.comb2_in_del[18] ),
    .X(_03263_));
 sg13g2_and2_1 _10513_ (.A(_03247_),
    .B(_03258_),
    .X(_03264_));
 sg13g2_a221oi_1 _10514_ (.B2(_03253_),
    .C1(_03257_),
    .B1(_03264_),
    .A1(_03246_),
    .Y(_03265_),
    .A2(_03256_));
 sg13g2_xnor2_1 _10515_ (.Y(_03266_),
    .A(net2790),
    .B(_03265_));
 sg13g2_o21ai_1 _10516_ (.B1(net2010),
    .Y(_03267_),
    .A1(net1828),
    .A2(net2339));
 sg13g2_a21oi_1 _10517_ (.A1(net1827),
    .A2(_03266_),
    .Y(_00497_),
    .B1(_03267_));
 sg13g2_o21ai_1 _10518_ (.B1(_03262_),
    .Y(_03268_),
    .A1(_03263_),
    .A2(_03265_));
 sg13g2_xor2_1 _10519_ (.B(net2315),
    .A(net2615),
    .X(_03269_));
 sg13g2_or2_1 _10520_ (.X(_03270_),
    .B(_03269_),
    .A(_03268_));
 sg13g2_a21oi_1 _10521_ (.A1(_03268_),
    .A2(_03269_),
    .Y(_03271_),
    .B1(net1634));
 sg13g2_a221oi_1 _10522_ (.B2(_03271_),
    .C1(net1893),
    .B1(_03270_),
    .A1(_01394_),
    .Y(_00498_),
    .A2(net1634));
 sg13g2_o21ai_1 _10523_ (.B1(net2014),
    .Y(_03272_),
    .A1(net1813),
    .A2(net2416));
 sg13g2_a21oi_1 _10524_ (.A1(net1814),
    .A2(_01448_),
    .Y(_00499_),
    .B1(_03272_));
 sg13g2_o21ai_1 _10525_ (.B1(net2013),
    .Y(_03273_),
    .A1(net1814),
    .A2(\am_sdr0.cic2.comb2_in_del[1] ));
 sg13g2_a21oi_1 _10526_ (.A1(net1814),
    .A2(_01446_),
    .Y(_00500_),
    .B1(_03273_));
 sg13g2_o21ai_1 _10527_ (.B1(net2011),
    .Y(_03274_),
    .A1(net1815),
    .A2(\am_sdr0.cic2.comb2_in_del[2] ));
 sg13g2_a21oi_1 _10528_ (.A1(net1815),
    .A2(_01445_),
    .Y(_00501_),
    .B1(_03274_));
 sg13g2_o21ai_1 _10529_ (.B1(net2011),
    .Y(_03275_),
    .A1(net1815),
    .A2(net2515));
 sg13g2_a21oi_1 _10530_ (.A1(net1815),
    .A2(_01444_),
    .Y(_00502_),
    .B1(_03275_));
 sg13g2_o21ai_1 _10531_ (.B1(net2009),
    .Y(_03276_),
    .A1(net1809),
    .A2(\am_sdr0.cic2.comb2_in_del[4] ));
 sg13g2_a21oi_1 _10532_ (.A1(net1809),
    .A2(_01443_),
    .Y(_00503_),
    .B1(_03276_));
 sg13g2_o21ai_1 _10533_ (.B1(net2009),
    .Y(_03277_),
    .A1(net1807),
    .A2(\am_sdr0.cic2.comb2_in_del[5] ));
 sg13g2_a21oi_1 _10534_ (.A1(net1807),
    .A2(_01442_),
    .Y(_00504_),
    .B1(_03277_));
 sg13g2_o21ai_1 _10535_ (.B1(net1978),
    .Y(_03278_),
    .A1(net1801),
    .A2(\am_sdr0.cic2.comb2_in_del[6] ));
 sg13g2_a21oi_1 _10536_ (.A1(net1801),
    .A2(_01441_),
    .Y(_00505_),
    .B1(_03278_));
 sg13g2_o21ai_1 _10537_ (.B1(net1978),
    .Y(_03279_),
    .A1(net1801),
    .A2(\am_sdr0.cic2.comb2_in_del[7] ));
 sg13g2_a21oi_1 _10538_ (.A1(net1801),
    .A2(_01440_),
    .Y(_00506_),
    .B1(_03279_));
 sg13g2_o21ai_1 _10539_ (.B1(net1976),
    .Y(_03280_),
    .A1(net1798),
    .A2(net2369));
 sg13g2_a21oi_1 _10540_ (.A1(net1798),
    .A2(_01439_),
    .Y(_00507_),
    .B1(_03280_));
 sg13g2_o21ai_1 _10541_ (.B1(net1976),
    .Y(_03281_),
    .A1(net1799),
    .A2(\am_sdr0.cic2.comb2_in_del[9] ));
 sg13g2_a21oi_1 _10542_ (.A1(net1799),
    .A2(_01438_),
    .Y(_00508_),
    .B1(_03281_));
 sg13g2_o21ai_1 _10543_ (.B1(net1976),
    .Y(_03282_),
    .A1(net1798),
    .A2(\am_sdr0.cic2.comb2_in_del[10] ));
 sg13g2_a21oi_1 _10544_ (.A1(net1798),
    .A2(_01437_),
    .Y(_00509_),
    .B1(_03282_));
 sg13g2_o21ai_1 _10545_ (.B1(net1975),
    .Y(_03283_),
    .A1(net1798),
    .A2(\am_sdr0.cic2.comb2_in_del[11] ));
 sg13g2_a21oi_1 _10546_ (.A1(net1798),
    .A2(_01436_),
    .Y(_00510_),
    .B1(_03283_));
 sg13g2_o21ai_1 _10547_ (.B1(net2008),
    .Y(_03284_),
    .A1(net1804),
    .A2(net2675));
 sg13g2_a21oi_1 _10548_ (.A1(net1804),
    .A2(_01435_),
    .Y(_00511_),
    .B1(_03284_));
 sg13g2_o21ai_1 _10549_ (.B1(net2008),
    .Y(_03285_),
    .A1(net1820),
    .A2(net2783));
 sg13g2_a21oi_1 _10550_ (.A1(net1820),
    .A2(_01433_),
    .Y(_00512_),
    .B1(_03285_));
 sg13g2_o21ai_1 _10551_ (.B1(net2012),
    .Y(_03286_),
    .A1(net1819),
    .A2(\am_sdr0.cic2.comb2_in_del[14] ));
 sg13g2_a21oi_1 _10552_ (.A1(net1819),
    .A2(_01431_),
    .Y(_00513_),
    .B1(_03286_));
 sg13g2_o21ai_1 _10553_ (.B1(net2008),
    .Y(_03287_),
    .A1(net1819),
    .A2(\am_sdr0.cic2.comb2_in_del[15] ));
 sg13g2_a21oi_1 _10554_ (.A1(net1819),
    .A2(_01430_),
    .Y(_00514_),
    .B1(_03287_));
 sg13g2_o21ai_1 _10555_ (.B1(net2010),
    .Y(_03288_),
    .A1(net1821),
    .A2(\am_sdr0.cic2.comb2_in_del[16] ));
 sg13g2_a21oi_1 _10556_ (.A1(net1826),
    .A2(_01429_),
    .Y(_00515_),
    .B1(_03288_));
 sg13g2_o21ai_1 _10557_ (.B1(net2010),
    .Y(_03289_),
    .A1(net1827),
    .A2(net2907));
 sg13g2_a21oi_1 _10558_ (.A1(net1827),
    .A2(_01428_),
    .Y(_00516_),
    .B1(_03289_));
 sg13g2_o21ai_1 _10559_ (.B1(net2010),
    .Y(_03290_),
    .A1(net1828),
    .A2(\am_sdr0.cic2.comb2_in_del[18] ));
 sg13g2_a21oi_1 _10560_ (.A1(net1828),
    .A2(_01427_),
    .Y(_00517_),
    .B1(_03290_));
 sg13g2_o21ai_1 _10561_ (.B1(net2016),
    .Y(_03291_),
    .A1(net1818),
    .A2(\am_sdr0.cic2.comb2_in_del[19] ));
 sg13g2_a21oi_1 _10562_ (.A1(net1818),
    .A2(_01426_),
    .Y(_00518_),
    .B1(_03291_));
 sg13g2_nand2_1 _10563_ (.Y(_03292_),
    .A(\am_sdr0.cic2.comb3_in_del[4] ),
    .B(_01413_));
 sg13g2_nand2b_1 _10564_ (.Y(_03293_),
    .B(\am_sdr0.cic2.comb3_in_del[1] ),
    .A_N(\am_sdr0.cic2.comb2[1] ));
 sg13g2_nand2b_1 _10565_ (.Y(_03294_),
    .B(\am_sdr0.cic2.comb3_in_del[0] ),
    .A_N(\am_sdr0.cic2.comb2[0] ));
 sg13g2_nor2b_1 _10566_ (.A(\am_sdr0.cic2.comb3_in_del[1] ),
    .B_N(\am_sdr0.cic2.comb2[1] ),
    .Y(_03295_));
 sg13g2_a221oi_1 _10567_ (.B2(_03294_),
    .C1(_03295_),
    .B1(_03293_),
    .A1(_01415_),
    .Y(_03296_),
    .A2(\am_sdr0.cic2.comb2[2] ));
 sg13g2_nand2b_1 _10568_ (.Y(_03297_),
    .B(\am_sdr0.cic2.comb3_in_del[3] ),
    .A_N(\am_sdr0.cic2.comb2[3] ));
 sg13g2_o21ai_1 _10569_ (.B1(_03297_),
    .Y(_03298_),
    .A1(_01415_),
    .A2(\am_sdr0.cic2.comb2[2] ));
 sg13g2_a22oi_1 _10570_ (.Y(_03299_),
    .B1(_01414_),
    .B2(\am_sdr0.cic2.comb2[3] ),
    .A2(\am_sdr0.cic2.comb2[4] ),
    .A1(_01412_));
 sg13g2_o21ai_1 _10571_ (.B1(_03299_),
    .Y(_03300_),
    .A1(_03296_),
    .A2(_03298_));
 sg13g2_a22oi_1 _10572_ (.Y(_03301_),
    .B1(_03292_),
    .B2(_03300_),
    .A2(\am_sdr0.cic2.comb2[5] ),
    .A1(_01410_));
 sg13g2_nand2_1 _10573_ (.Y(_03302_),
    .A(\am_sdr0.cic2.comb3_in_del[5] ),
    .B(_01411_));
 sg13g2_o21ai_1 _10574_ (.B1(_03302_),
    .Y(_03303_),
    .A1(_01409_),
    .A2(\am_sdr0.cic2.comb2[6] ));
 sg13g2_a22oi_1 _10575_ (.Y(_03304_),
    .B1(_01409_),
    .B2(\am_sdr0.cic2.comb2[6] ),
    .A2(\am_sdr0.cic2.comb2[7] ),
    .A1(_01407_));
 sg13g2_o21ai_1 _10576_ (.B1(_03304_),
    .Y(_03305_),
    .A1(_03301_),
    .A2(_03303_));
 sg13g2_nand2b_1 _10577_ (.Y(_03306_),
    .B(\am_sdr0.cic2.comb2[11] ),
    .A_N(\am_sdr0.cic2.comb3_in_del[11] ));
 sg13g2_nand2_1 _10578_ (.Y(_03307_),
    .A(\am_sdr0.cic2.comb3_in_del[11] ),
    .B(_01403_));
 sg13g2_nand2b_1 _10579_ (.Y(_03308_),
    .B(\am_sdr0.cic2.comb2[10] ),
    .A_N(\am_sdr0.cic2.comb3_in_del[10] ));
 sg13g2_a22oi_1 _10580_ (.Y(_03309_),
    .B1(\am_sdr0.cic2.comb3_in_del[9] ),
    .B2(_01405_),
    .A2(_01404_),
    .A1(\am_sdr0.cic2.comb3_in_del[10] ));
 sg13g2_nand4_1 _10581_ (.B(_03307_),
    .C(_03308_),
    .A(_03306_),
    .Y(_03310_),
    .D(_03309_));
 sg13g2_nand2b_1 _10582_ (.Y(_03311_),
    .B(\am_sdr0.cic2.comb2[9] ),
    .A_N(\am_sdr0.cic2.comb3_in_del[9] ));
 sg13g2_o21ai_1 _10583_ (.B1(_03311_),
    .Y(_03312_),
    .A1(\am_sdr0.cic2.comb3_in_del[8] ),
    .A2(_01406_));
 sg13g2_a221oi_1 _10584_ (.B2(_01408_),
    .C1(_03312_),
    .B1(\am_sdr0.cic2.comb3_in_del[7] ),
    .A1(\am_sdr0.cic2.comb3_in_del[8] ),
    .Y(_03313_),
    .A2(_01406_));
 sg13g2_nor2b_1 _10585_ (.A(_03310_),
    .B_N(_03313_),
    .Y(_03314_));
 sg13g2_nand2b_1 _10586_ (.Y(_03315_),
    .B(_03312_),
    .A_N(_03310_));
 sg13g2_nand3b_1 _10587_ (.B(\am_sdr0.cic2.comb2[10] ),
    .C(_03307_),
    .Y(_03316_),
    .A_N(\am_sdr0.cic2.comb3_in_del[10] ));
 sg13g2_nand3_1 _10588_ (.B(_03315_),
    .C(_03316_),
    .A(_03306_),
    .Y(_03317_));
 sg13g2_a21oi_2 _10589_ (.B1(_03317_),
    .Y(_03318_),
    .A2(_03314_),
    .A1(_03305_));
 sg13g2_xnor2_1 _10590_ (.Y(_03319_),
    .A(\am_sdr0.cic2.comb3_in_del[12] ),
    .B(\am_sdr0.cic2.comb2[12] ));
 sg13g2_nor2b_1 _10591_ (.A(_03318_),
    .B_N(_03319_),
    .Y(_03320_));
 sg13g2_xor2_1 _10592_ (.B(_03319_),
    .A(_03318_),
    .X(_03321_));
 sg13g2_o21ai_1 _10593_ (.B1(net2017),
    .Y(_03322_),
    .A1(net1826),
    .A2(net1231));
 sg13g2_a21oi_1 _10594_ (.A1(net1822),
    .A2(_03321_),
    .Y(_00519_),
    .B1(_03322_));
 sg13g2_nand2_1 _10595_ (.Y(_03323_),
    .A(\am_sdr0.cic2.comb3_in_del[13] ),
    .B(_01401_));
 sg13g2_xnor2_1 _10596_ (.Y(_03324_),
    .A(\am_sdr0.cic2.comb3_in_del[13] ),
    .B(net2509));
 sg13g2_a21oi_1 _10597_ (.A1(_01402_),
    .A2(net3296),
    .Y(_03325_),
    .B1(_03320_));
 sg13g2_o21ai_1 _10598_ (.B1(net1822),
    .Y(_03326_),
    .A1(_03324_),
    .A2(_03325_));
 sg13g2_a21oi_1 _10599_ (.A1(net2510),
    .A2(_03325_),
    .Y(_03327_),
    .B1(_03326_));
 sg13g2_o21ai_1 _10600_ (.B1(net2019),
    .Y(_03328_),
    .A1(net1822),
    .A2(net1369));
 sg13g2_nor2_1 _10601_ (.A(_03327_),
    .B(_03328_),
    .Y(_00520_));
 sg13g2_nand2b_1 _10602_ (.Y(_03329_),
    .B(net2314),
    .A_N(\am_sdr0.cic2.comb3_in_del[14] ));
 sg13g2_inv_1 _10603_ (.Y(_03330_),
    .A(_03329_));
 sg13g2_nand2_1 _10604_ (.Y(_03331_),
    .A(net3318),
    .B(_01400_));
 sg13g2_nand2_1 _10605_ (.Y(_03332_),
    .A(_03329_),
    .B(_03331_));
 sg13g2_nand3_1 _10606_ (.B(\am_sdr0.cic2.comb2[12] ),
    .C(_03323_),
    .A(_01402_),
    .Y(_03333_));
 sg13g2_o21ai_1 _10607_ (.B1(_03333_),
    .Y(_03334_),
    .A1(\am_sdr0.cic2.comb3_in_del[13] ),
    .A2(_01401_));
 sg13g2_nand3b_1 _10608_ (.B(_03319_),
    .C(_03324_),
    .Y(_03335_),
    .A_N(_03318_));
 sg13g2_nand2b_1 _10609_ (.Y(_03336_),
    .B(_03335_),
    .A_N(_03334_));
 sg13g2_xor2_1 _10610_ (.B(_03336_),
    .A(_03332_),
    .X(_03337_));
 sg13g2_o21ai_1 _10611_ (.B1(net2018),
    .Y(_03338_),
    .A1(net1823),
    .A2(net1295));
 sg13g2_a21oi_1 _10612_ (.A1(net1823),
    .A2(_03337_),
    .Y(_00521_),
    .B1(_03338_));
 sg13g2_nand2b_1 _10613_ (.Y(_03339_),
    .B(net2104),
    .A_N(\am_sdr0.cic2.comb3_in_del[15] ));
 sg13g2_nand2_1 _10614_ (.Y(_03340_),
    .A(net3319),
    .B(_01399_));
 sg13g2_a21oi_1 _10615_ (.A1(_03331_),
    .A2(_03336_),
    .Y(_03341_),
    .B1(_03330_));
 sg13g2_a21oi_1 _10616_ (.A1(_03339_),
    .A2(_03340_),
    .Y(_03342_),
    .B1(_03341_));
 sg13g2_nand3_1 _10617_ (.B(_03340_),
    .C(_03341_),
    .A(net2105),
    .Y(_03343_));
 sg13g2_nor2_1 _10618_ (.A(net1633),
    .B(_03342_),
    .Y(_03344_));
 sg13g2_a221oi_1 _10619_ (.B2(_03344_),
    .C1(net1892),
    .B1(net2106),
    .A1(net1633),
    .Y(_00522_),
    .A2(_01422_));
 sg13g2_nor2_1 _10620_ (.A(\am_sdr0.cic2.comb3_in_del[16] ),
    .B(_01398_),
    .Y(_03345_));
 sg13g2_xnor2_1 _10621_ (.Y(_03346_),
    .A(\am_sdr0.cic2.comb3_in_del[16] ),
    .B(net2344));
 sg13g2_nor2b_1 _10622_ (.A(_03331_),
    .B_N(_03339_),
    .Y(_03347_));
 sg13g2_nand2_1 _10623_ (.Y(_03348_),
    .A(_03330_),
    .B(_03340_));
 sg13g2_nand2_1 _10624_ (.Y(_03349_),
    .A(_03339_),
    .B(_03348_));
 sg13g2_nor2_1 _10625_ (.A(_03334_),
    .B(_03349_),
    .Y(_03350_));
 sg13g2_a221oi_1 _10626_ (.B2(_03350_),
    .C1(_03347_),
    .B1(_03335_),
    .A1(\am_sdr0.cic2.comb3_in_del[15] ),
    .Y(_03351_),
    .A2(_01399_));
 sg13g2_xnor2_1 _10627_ (.Y(_03352_),
    .A(net2345),
    .B(_03351_));
 sg13g2_o21ai_1 _10628_ (.B1(net2020),
    .Y(_03353_),
    .A1(net1825),
    .A2(net1262));
 sg13g2_a21oi_1 _10629_ (.A1(net1825),
    .A2(net2346),
    .Y(_00523_),
    .B1(_03353_));
 sg13g2_a21oi_1 _10630_ (.A1(_03346_),
    .A2(_03351_),
    .Y(_03354_),
    .B1(_03345_));
 sg13g2_nand2b_1 _10631_ (.Y(_03355_),
    .B(\am_sdr0.cic2.comb2[17] ),
    .A_N(\am_sdr0.cic2.comb3_in_del[17] ));
 sg13g2_nor2b_1 _10632_ (.A(net2039),
    .B_N(\am_sdr0.cic2.comb3_in_del[17] ),
    .Y(_03356_));
 sg13g2_xnor2_1 _10633_ (.Y(_03357_),
    .A(\am_sdr0.cic2.comb3_in_del[17] ),
    .B(net2039));
 sg13g2_nor2_1 _10634_ (.A(_03354_),
    .B(_03357_),
    .Y(_03358_));
 sg13g2_nand2_1 _10635_ (.Y(_03359_),
    .A(_03354_),
    .B(net2040));
 sg13g2_nor2_1 _10636_ (.A(net1633),
    .B(_03358_),
    .Y(_03360_));
 sg13g2_a221oi_1 _10637_ (.B2(_03360_),
    .C1(net1892),
    .B1(net2041),
    .A1(net1633),
    .Y(_00524_),
    .A2(_01420_));
 sg13g2_nor2_1 _10638_ (.A(\am_sdr0.cic2.comb3_in_del[18] ),
    .B(_01396_),
    .Y(_03361_));
 sg13g2_xnor2_1 _10639_ (.Y(_03362_),
    .A(\am_sdr0.cic2.comb3_in_del[18] ),
    .B(net2339));
 sg13g2_a21oi_1 _10640_ (.A1(_03354_),
    .A2(_03355_),
    .Y(_03363_),
    .B1(_03356_));
 sg13g2_xnor2_1 _10641_ (.Y(_03364_),
    .A(net2340),
    .B(_03363_));
 sg13g2_o21ai_1 _10642_ (.B1(net2020),
    .Y(_03365_),
    .A1(net1829),
    .A2(net1246));
 sg13g2_a21oi_1 _10643_ (.A1(net1829),
    .A2(net2341),
    .Y(_00525_),
    .B1(_03365_));
 sg13g2_a21oi_1 _10644_ (.A1(_03362_),
    .A2(_03363_),
    .Y(_03366_),
    .B1(_03361_));
 sg13g2_xnor2_1 _10645_ (.Y(_03367_),
    .A(\am_sdr0.cic2.comb3_in_del[19] ),
    .B(net2057));
 sg13g2_or2_1 _10646_ (.X(_03368_),
    .B(net2058),
    .A(_03366_));
 sg13g2_a21oi_1 _10647_ (.A1(_03366_),
    .A2(net2058),
    .Y(_03369_),
    .B1(net1633));
 sg13g2_a221oi_1 _10648_ (.B2(_03369_),
    .C1(net1892),
    .B1(net2059),
    .A1(net1633),
    .Y(_00526_),
    .A2(_01418_));
 sg13g2_o21ai_1 _10649_ (.B1(net2015),
    .Y(_03370_),
    .A1(net1817),
    .A2(\am_sdr0.cic2.comb3_in_del[0] ));
 sg13g2_a21oi_1 _10650_ (.A1(net1817),
    .A2(_01417_),
    .Y(_00527_),
    .B1(_03370_));
 sg13g2_o21ai_1 _10651_ (.B1(net2015),
    .Y(_03371_),
    .A1(net1817),
    .A2(\am_sdr0.cic2.comb3_in_del[1] ));
 sg13g2_a21oi_1 _10652_ (.A1(net1817),
    .A2(_01416_),
    .Y(_00528_),
    .B1(_03371_));
 sg13g2_o21ai_1 _10653_ (.B1(net2015),
    .Y(_03372_),
    .A1(net1631),
    .A2(\am_sdr0.cic2.comb2[2] ));
 sg13g2_a21oi_1 _10654_ (.A1(net1631),
    .A2(_01415_),
    .Y(_00529_),
    .B1(_03372_));
 sg13g2_o21ai_1 _10655_ (.B1(net2011),
    .Y(_03373_),
    .A1(net1631),
    .A2(\am_sdr0.cic2.comb2[3] ));
 sg13g2_a21oi_1 _10656_ (.A1(net1631),
    .A2(_01414_),
    .Y(_00530_),
    .B1(_03373_));
 sg13g2_o21ai_1 _10657_ (.B1(net2010),
    .Y(_03374_),
    .A1(net1810),
    .A2(\am_sdr0.cic2.comb3_in_del[4] ));
 sg13g2_a21oi_1 _10658_ (.A1(net1810),
    .A2(_01413_),
    .Y(_00531_),
    .B1(_03374_));
 sg13g2_o21ai_1 _10659_ (.B1(net2008),
    .Y(_03375_),
    .A1(net1810),
    .A2(\am_sdr0.cic2.comb3_in_del[5] ));
 sg13g2_a21oi_1 _10660_ (.A1(net1809),
    .A2(_01411_),
    .Y(_00532_),
    .B1(_03375_));
 sg13g2_o21ai_1 _10661_ (.B1(net2012),
    .Y(_03376_),
    .A1(net1628),
    .A2(\am_sdr0.cic2.comb2[6] ));
 sg13g2_a21oi_1 _10662_ (.A1(net1629),
    .A2(_01409_),
    .Y(_00533_),
    .B1(_03376_));
 sg13g2_o21ai_1 _10663_ (.B1(net1977),
    .Y(_03377_),
    .A1(net1802),
    .A2(net2585));
 sg13g2_a21oi_1 _10664_ (.A1(net1804),
    .A2(_01408_),
    .Y(_00534_),
    .B1(_03377_));
 sg13g2_o21ai_1 _10665_ (.B1(net1977),
    .Y(_03378_),
    .A1(net1804),
    .A2(\am_sdr0.cic2.comb3_in_del[8] ));
 sg13g2_a21oi_1 _10666_ (.A1(net1804),
    .A2(_01406_),
    .Y(_00535_),
    .B1(_03378_));
 sg13g2_o21ai_1 _10667_ (.B1(net1977),
    .Y(_03379_),
    .A1(net1804),
    .A2(\am_sdr0.cic2.comb3_in_del[9] ));
 sg13g2_a21oi_1 _10668_ (.A1(net1804),
    .A2(_01405_),
    .Y(_00536_),
    .B1(_03379_));
 sg13g2_o21ai_1 _10669_ (.B1(net1977),
    .Y(_03380_),
    .A1(net1805),
    .A2(\am_sdr0.cic2.comb3_in_del[10] ));
 sg13g2_a21oi_1 _10670_ (.A1(net1805),
    .A2(_01404_),
    .Y(_00537_),
    .B1(_03380_));
 sg13g2_o21ai_1 _10671_ (.B1(net1977),
    .Y(_03381_),
    .A1(net1805),
    .A2(net2511));
 sg13g2_a21oi_1 _10672_ (.A1(net1805),
    .A2(_01403_),
    .Y(_00538_),
    .B1(_03381_));
 sg13g2_o21ai_1 _10673_ (.B1(net2019),
    .Y(_03382_),
    .A1(net1628),
    .A2(net2674));
 sg13g2_a21oi_1 _10674_ (.A1(net1629),
    .A2(_01402_),
    .Y(_00539_),
    .B1(_03382_));
 sg13g2_o21ai_1 _10675_ (.B1(net2019),
    .Y(_03383_),
    .A1(net1822),
    .A2(net2797));
 sg13g2_a21oi_1 _10676_ (.A1(net1822),
    .A2(_01401_),
    .Y(_00540_),
    .B1(_03383_));
 sg13g2_o21ai_1 _10677_ (.B1(net2019),
    .Y(_03384_),
    .A1(net1822),
    .A2(net2437));
 sg13g2_a21oi_1 _10678_ (.A1(net1822),
    .A2(_01400_),
    .Y(_00541_),
    .B1(_03384_));
 sg13g2_o21ai_1 _10679_ (.B1(net2019),
    .Y(_03385_),
    .A1(net1821),
    .A2(net2707));
 sg13g2_a21oi_1 _10680_ (.A1(net1821),
    .A2(_01399_),
    .Y(_00542_),
    .B1(_03385_));
 sg13g2_o21ai_1 _10681_ (.B1(net2020),
    .Y(_03386_),
    .A1(net1821),
    .A2(net2531));
 sg13g2_a21oi_1 _10682_ (.A1(net1821),
    .A2(_01398_),
    .Y(_00543_),
    .B1(_03386_));
 sg13g2_o21ai_1 _10683_ (.B1(net2020),
    .Y(_03387_),
    .A1(net1827),
    .A2(net2647));
 sg13g2_a21oi_1 _10684_ (.A1(net1827),
    .A2(_01397_),
    .Y(_00544_),
    .B1(_03387_));
 sg13g2_o21ai_1 _10685_ (.B1(net2020),
    .Y(_03388_),
    .A1(net1827),
    .A2(net2532));
 sg13g2_a21oi_1 _10686_ (.A1(net1827),
    .A2(_01396_),
    .Y(_00545_),
    .B1(_03388_));
 sg13g2_o21ai_1 _10687_ (.B1(net2015),
    .Y(_03389_),
    .A1(net2391),
    .A2(net1828));
 sg13g2_a21oi_1 _10688_ (.A1(_01394_),
    .A2(net1828),
    .Y(_00546_),
    .B1(_03389_));
 sg13g2_o21ai_1 _10689_ (.B1(net1914),
    .Y(_03390_),
    .A1(net1670),
    .A2(net1397));
 sg13g2_a21oi_1 _10690_ (.A1(net1670),
    .A2(net1397),
    .Y(_00547_),
    .B1(_03390_));
 sg13g2_a21oi_1 _10691_ (.A1(net1670),
    .A2(\am_sdr0.cic2.count[0] ),
    .Y(_03391_),
    .B1(net1228));
 sg13g2_nand2_1 _10692_ (.Y(_03392_),
    .A(net1914),
    .B(_02128_));
 sg13g2_nor2_1 _10693_ (.A(net1229),
    .B(_03392_),
    .Y(_00548_));
 sg13g2_a21oi_1 _10694_ (.A1(_01393_),
    .A2(_02128_),
    .Y(_03393_),
    .B1(net1888));
 sg13g2_nor2b_1 _10695_ (.A(_02129_),
    .B_N(_03393_),
    .Y(_00549_));
 sg13g2_o21ai_1 _10696_ (.B1(net1964),
    .Y(_03394_),
    .A1(net2548),
    .A2(_02129_));
 sg13g2_nor2_1 _10697_ (.A(_02130_),
    .B(net2549),
    .Y(_00550_));
 sg13g2_o21ai_1 _10698_ (.B1(net1963),
    .Y(_03395_),
    .A1(net2619),
    .A2(_02130_));
 sg13g2_nor2_1 _10699_ (.A(_02131_),
    .B(_03395_),
    .Y(_00551_));
 sg13g2_o21ai_1 _10700_ (.B1(net1963),
    .Y(_03396_),
    .A1(net2851),
    .A2(_02131_));
 sg13g2_nor2b_1 _10701_ (.A(_03396_),
    .B_N(_02132_),
    .Y(_00552_));
 sg13g2_a21oi_1 _10702_ (.A1(\am_sdr0.cic2.count[5] ),
    .A2(_02131_),
    .Y(_03397_),
    .B1(net2063));
 sg13g2_and3_1 _10703_ (.X(_03398_),
    .A(net2063),
    .B(\am_sdr0.cic2.count[5] ),
    .C(_02131_));
 sg13g2_nor4_1 _10704_ (.A(net1888),
    .B(_02133_),
    .C(net2064),
    .D(_03398_),
    .Y(_00553_));
 sg13g2_o21ai_1 _10705_ (.B1(net1963),
    .Y(_03399_),
    .A1(net1328),
    .A2(_03398_));
 sg13g2_a21oi_1 _10706_ (.A1(net1328),
    .A2(_03398_),
    .Y(_00554_),
    .B1(_03399_));
 sg13g2_a21oi_1 _10707_ (.A1(\am_sdr0.cic0.x_out[8] ),
    .A2(net1692),
    .Y(_03400_),
    .B1(net1280));
 sg13g2_nand2_1 _10708_ (.Y(_03401_),
    .A(\am_sdr0.cic0.x_out[8] ),
    .B(net1280));
 sg13g2_nor2_1 _10709_ (.A(net1636),
    .B(_03401_),
    .Y(_03402_));
 sg13g2_nor3_1 _10710_ (.A(net1891),
    .B(net1281),
    .C(_03402_),
    .Y(_00555_));
 sg13g2_nand2_1 _10711_ (.Y(_03403_),
    .A(\am_sdr0.cic0.x_out[9] ),
    .B(\am_sdr0.cic2.integ1[1] ));
 sg13g2_xnor2_1 _10712_ (.Y(_03404_),
    .A(\am_sdr0.cic0.x_out[9] ),
    .B(net2840));
 sg13g2_xnor2_1 _10713_ (.Y(_03405_),
    .A(_03401_),
    .B(_03404_));
 sg13g2_o21ai_1 _10714_ (.B1(net2005),
    .Y(_03406_),
    .A1(net1692),
    .A2(net2840));
 sg13g2_a21oi_1 _10715_ (.A1(net1689),
    .A2(_03405_),
    .Y(_00556_),
    .B1(_03406_));
 sg13g2_and2_1 _10716_ (.A(\am_sdr0.cic0.x_out[10] ),
    .B(\am_sdr0.cic2.integ1[2] ),
    .X(_03407_));
 sg13g2_xor2_1 _10717_ (.B(net2802),
    .A(\am_sdr0.cic0.x_out[10] ),
    .X(_03408_));
 sg13g2_o21ai_1 _10718_ (.B1(_03403_),
    .Y(_03409_),
    .A1(_03401_),
    .A2(_03404_));
 sg13g2_xnor2_1 _10719_ (.Y(_03410_),
    .A(_03408_),
    .B(_03409_));
 sg13g2_o21ai_1 _10720_ (.B1(net2005),
    .Y(_03411_),
    .A1(net1689),
    .A2(net2802));
 sg13g2_a21oi_1 _10721_ (.A1(net1689),
    .A2(_03410_),
    .Y(_00557_),
    .B1(_03411_));
 sg13g2_nand2_1 _10722_ (.Y(_03412_),
    .A(\am_sdr0.cic0.x_out[11] ),
    .B(\am_sdr0.cic2.integ1[3] ));
 sg13g2_xnor2_1 _10723_ (.Y(_03413_),
    .A(\am_sdr0.cic0.x_out[11] ),
    .B(\am_sdr0.cic2.integ1[3] ));
 sg13g2_a21oi_1 _10724_ (.A1(_03408_),
    .A2(_03409_),
    .Y(_03414_),
    .B1(_03407_));
 sg13g2_xnor2_1 _10725_ (.Y(_03415_),
    .A(_03413_),
    .B(_03414_));
 sg13g2_o21ai_1 _10726_ (.B1(net2005),
    .Y(_03416_),
    .A1(net1689),
    .A2(net2961));
 sg13g2_a21oi_1 _10727_ (.A1(net1689),
    .A2(_03415_),
    .Y(_00558_),
    .B1(_03416_));
 sg13g2_o21ai_1 _10728_ (.B1(_03412_),
    .Y(_03417_),
    .A1(_03413_),
    .A2(_03414_));
 sg13g2_nand2_1 _10729_ (.Y(_03418_),
    .A(\am_sdr0.cic0.x_out[12] ),
    .B(\am_sdr0.cic2.integ1[4] ));
 sg13g2_xor2_1 _10730_ (.B(\am_sdr0.cic2.integ1[4] ),
    .A(\am_sdr0.cic0.x_out[12] ),
    .X(_03419_));
 sg13g2_inv_1 _10731_ (.Y(_03420_),
    .A(_03419_));
 sg13g2_nand2_1 _10732_ (.Y(_03421_),
    .A(_03417_),
    .B(_03419_));
 sg13g2_xnor2_1 _10733_ (.Y(_03422_),
    .A(_03417_),
    .B(_03419_));
 sg13g2_o21ai_1 _10734_ (.B1(net1946),
    .Y(_03423_),
    .A1(net1684),
    .A2(net3063));
 sg13g2_a21oi_1 _10735_ (.A1(net1684),
    .A2(_03422_),
    .Y(_00559_),
    .B1(_03423_));
 sg13g2_nor2_1 _10736_ (.A(\am_sdr0.cic0.x_out[13] ),
    .B(\am_sdr0.cic2.integ1[5] ),
    .Y(_03424_));
 sg13g2_nand2_1 _10737_ (.Y(_03425_),
    .A(\am_sdr0.cic0.x_out[13] ),
    .B(\am_sdr0.cic2.integ1[5] ));
 sg13g2_nand2b_1 _10738_ (.Y(_03426_),
    .B(_03425_),
    .A_N(_03424_));
 sg13g2_nand2_1 _10739_ (.Y(_03427_),
    .A(_03418_),
    .B(_03421_));
 sg13g2_o21ai_1 _10740_ (.B1(net1683),
    .Y(_03428_),
    .A1(_03426_),
    .A2(_03427_));
 sg13g2_a21oi_1 _10741_ (.A1(_03426_),
    .A2(_03427_),
    .Y(_03429_),
    .B1(_03428_));
 sg13g2_o21ai_1 _10742_ (.B1(net1945),
    .Y(_03430_),
    .A1(net1683),
    .A2(net2978));
 sg13g2_nor2_1 _10743_ (.A(_03429_),
    .B(_03430_),
    .Y(_00560_));
 sg13g2_nand2_1 _10744_ (.Y(_03431_),
    .A(\am_sdr0.cic0.x_out[14] ),
    .B(\am_sdr0.cic2.integ1[6] ));
 sg13g2_or2_1 _10745_ (.X(_03432_),
    .B(\am_sdr0.cic2.integ1[6] ),
    .A(\am_sdr0.cic0.x_out[14] ));
 sg13g2_nand2_1 _10746_ (.Y(_03433_),
    .A(_03431_),
    .B(_03432_));
 sg13g2_nor2_1 _10747_ (.A(_03420_),
    .B(_03426_),
    .Y(_03434_));
 sg13g2_o21ai_1 _10748_ (.B1(_03425_),
    .Y(_03435_),
    .A1(_03418_),
    .A2(_03424_));
 sg13g2_a21o_1 _10749_ (.A2(_03434_),
    .A1(_03417_),
    .B1(_03435_),
    .X(_03436_));
 sg13g2_nand2b_1 _10750_ (.Y(_03437_),
    .B(_03436_),
    .A_N(_03433_));
 sg13g2_xor2_1 _10751_ (.B(_03436_),
    .A(_03433_),
    .X(_03438_));
 sg13g2_o21ai_1 _10752_ (.B1(net1946),
    .Y(_03439_),
    .A1(net1683),
    .A2(net2993));
 sg13g2_a21oi_1 _10753_ (.A1(net1683),
    .A2(_03438_),
    .Y(_00561_),
    .B1(_03439_));
 sg13g2_nor2_1 _10754_ (.A(net1698),
    .B(\am_sdr0.cic2.integ1[7] ),
    .Y(_03440_));
 sg13g2_inv_1 _10755_ (.Y(_03441_),
    .A(_03440_));
 sg13g2_and2_1 _10756_ (.A(net1698),
    .B(\am_sdr0.cic2.integ1[7] ),
    .X(_03442_));
 sg13g2_nand2_1 _10757_ (.Y(_03443_),
    .A(_03431_),
    .B(_03437_));
 sg13g2_nor3_1 _10758_ (.A(_03440_),
    .B(_03442_),
    .C(_03443_),
    .Y(_03444_));
 sg13g2_o21ai_1 _10759_ (.B1(_03443_),
    .Y(_03445_),
    .A1(_03440_),
    .A2(_03442_));
 sg13g2_nor2_1 _10760_ (.A(net1635),
    .B(_03444_),
    .Y(_03446_));
 sg13g2_o21ai_1 _10761_ (.B1(net1924),
    .Y(_03447_),
    .A1(net1683),
    .A2(net3002));
 sg13g2_a21oi_1 _10762_ (.A1(_03445_),
    .A2(_03446_),
    .Y(_00562_),
    .B1(_03447_));
 sg13g2_nor2_1 _10763_ (.A(_03431_),
    .B(_03440_),
    .Y(_03448_));
 sg13g2_or3_1 _10764_ (.A(_03435_),
    .B(_03442_),
    .C(_03448_),
    .X(_03449_));
 sg13g2_a21oi_2 _10765_ (.B1(_03449_),
    .Y(_03450_),
    .A2(_03434_),
    .A1(_03417_));
 sg13g2_o21ai_1 _10766_ (.B1(_03441_),
    .Y(_03451_),
    .A1(_03432_),
    .A2(_03442_));
 sg13g2_or2_1 _10767_ (.X(_03452_),
    .B(_03451_),
    .A(_03450_));
 sg13g2_xor2_1 _10768_ (.B(\am_sdr0.cic2.integ1[8] ),
    .A(net1694),
    .X(_03453_));
 sg13g2_nand2b_1 _10769_ (.Y(_03454_),
    .B(_03453_),
    .A_N(_03452_));
 sg13g2_xor2_1 _10770_ (.B(_03453_),
    .A(_03452_),
    .X(_03455_));
 sg13g2_o21ai_1 _10771_ (.B1(net1924),
    .Y(_03456_),
    .A1(net1681),
    .A2(net3065));
 sg13g2_a21oi_1 _10772_ (.A1(net1678),
    .A2(_03455_),
    .Y(_00563_),
    .B1(_03456_));
 sg13g2_xor2_1 _10773_ (.B(\am_sdr0.cic2.integ1[9] ),
    .A(net1694),
    .X(_03457_));
 sg13g2_inv_1 _10774_ (.Y(_03458_),
    .A(_03457_));
 sg13g2_o21ai_1 _10775_ (.B1(_03454_),
    .Y(_03459_),
    .A1(_01304_),
    .A2(_01392_));
 sg13g2_xnor2_1 _10776_ (.Y(_03460_),
    .A(_03457_),
    .B(_03459_));
 sg13g2_o21ai_1 _10777_ (.B1(net1924),
    .Y(_03461_),
    .A1(net1677),
    .A2(net3010));
 sg13g2_a21oi_1 _10778_ (.A1(net1677),
    .A2(_03460_),
    .Y(_00564_),
    .B1(_03461_));
 sg13g2_and2_1 _10779_ (.A(net1694),
    .B(\am_sdr0.cic2.integ1[10] ),
    .X(_03462_));
 sg13g2_xor2_1 _10780_ (.B(\am_sdr0.cic2.integ1[10] ),
    .A(net1694),
    .X(_03463_));
 sg13g2_o21ai_1 _10781_ (.B1(net1694),
    .Y(_03464_),
    .A1(\am_sdr0.cic2.integ1[9] ),
    .A2(\am_sdr0.cic2.integ1[8] ));
 sg13g2_o21ai_1 _10782_ (.B1(_03464_),
    .Y(_03465_),
    .A1(_03454_),
    .A2(_03458_));
 sg13g2_xnor2_1 _10783_ (.Y(_03466_),
    .A(_03463_),
    .B(_03465_));
 sg13g2_o21ai_1 _10784_ (.B1(net1924),
    .Y(_03467_),
    .A1(net1677),
    .A2(net3125));
 sg13g2_a21oi_1 _10785_ (.A1(net1677),
    .A2(_03466_),
    .Y(_00565_),
    .B1(_03467_));
 sg13g2_xor2_1 _10786_ (.B(\am_sdr0.cic2.integ1[11] ),
    .A(net1694),
    .X(_03468_));
 sg13g2_a21oi_1 _10787_ (.A1(_03463_),
    .A2(_03465_),
    .Y(_03469_),
    .B1(_03462_));
 sg13g2_xor2_1 _10788_ (.B(_03469_),
    .A(_03468_),
    .X(_03470_));
 sg13g2_o21ai_1 _10789_ (.B1(net1925),
    .Y(_03471_),
    .A1(net1677),
    .A2(net3023));
 sg13g2_a21oi_1 _10790_ (.A1(net1677),
    .A2(_03470_),
    .Y(_00566_),
    .B1(_03471_));
 sg13g2_xor2_1 _10791_ (.B(\am_sdr0.cic2.integ1[12] ),
    .A(net1693),
    .X(_03472_));
 sg13g2_nand4_1 _10792_ (.B(_03457_),
    .C(_03463_),
    .A(_03453_),
    .Y(_03473_),
    .D(_03468_));
 sg13g2_nor3_2 _10793_ (.A(_03450_),
    .B(_03451_),
    .C(_03473_),
    .Y(_03474_));
 sg13g2_o21ai_1 _10794_ (.B1(net1694),
    .Y(_03475_),
    .A1(\am_sdr0.cic2.integ1[11] ),
    .A2(\am_sdr0.cic2.integ1[10] ));
 sg13g2_and2_1 _10795_ (.A(_03464_),
    .B(_03475_),
    .X(_03476_));
 sg13g2_nand2b_1 _10796_ (.Y(_03477_),
    .B(_03476_),
    .A_N(_03474_));
 sg13g2_and2_1 _10797_ (.A(_03472_),
    .B(_03477_),
    .X(_03478_));
 sg13g2_xnor2_1 _10798_ (.Y(_03479_),
    .A(_03472_),
    .B(_03477_));
 sg13g2_o21ai_1 _10799_ (.B1(net1922),
    .Y(_03480_),
    .A1(net1672),
    .A2(net3014));
 sg13g2_a21oi_1 _10800_ (.A1(net1672),
    .A2(_03479_),
    .Y(_00567_),
    .B1(_03480_));
 sg13g2_xnor2_1 _10801_ (.Y(_03481_),
    .A(net1693),
    .B(\am_sdr0.cic2.integ1[13] ));
 sg13g2_inv_1 _10802_ (.Y(_03482_),
    .A(_03481_));
 sg13g2_a21oi_1 _10803_ (.A1(net1693),
    .A2(net3317),
    .Y(_03483_),
    .B1(_03478_));
 sg13g2_xnor2_1 _10804_ (.Y(_03484_),
    .A(_03481_),
    .B(_03483_));
 sg13g2_o21ai_1 _10805_ (.B1(net1922),
    .Y(_03485_),
    .A1(net1672),
    .A2(net3001));
 sg13g2_a21oi_1 _10806_ (.A1(net1672),
    .A2(_03484_),
    .Y(_00568_),
    .B1(_03485_));
 sg13g2_xnor2_1 _10807_ (.Y(_03486_),
    .A(net1693),
    .B(\am_sdr0.cic2.integ1[14] ));
 sg13g2_o21ai_1 _10808_ (.B1(net1693),
    .Y(_03487_),
    .A1(\am_sdr0.cic2.integ1[13] ),
    .A2(\am_sdr0.cic2.integ1[12] ));
 sg13g2_nand2_1 _10809_ (.Y(_03488_),
    .A(_03478_),
    .B(_03482_));
 sg13g2_a21oi_1 _10810_ (.A1(_03487_),
    .A2(_03488_),
    .Y(_03489_),
    .B1(_03486_));
 sg13g2_nand3_1 _10811_ (.B(_03487_),
    .C(_03488_),
    .A(_03486_),
    .Y(_03490_));
 sg13g2_nand2b_1 _10812_ (.Y(_03491_),
    .B(_03490_),
    .A_N(_03489_));
 sg13g2_o21ai_1 _10813_ (.B1(net1922),
    .Y(_03492_),
    .A1(net1670),
    .A2(net3121));
 sg13g2_a21oi_1 _10814_ (.A1(net1670),
    .A2(_03491_),
    .Y(_00569_),
    .B1(_03492_));
 sg13g2_xnor2_1 _10815_ (.Y(_03493_),
    .A(net1693),
    .B(\am_sdr0.cic2.integ1[15] ));
 sg13g2_a21oi_1 _10816_ (.A1(net1693),
    .A2(\am_sdr0.cic2.integ1[14] ),
    .Y(_03494_),
    .B1(_03489_));
 sg13g2_xnor2_1 _10817_ (.Y(_03495_),
    .A(_03493_),
    .B(_03494_));
 sg13g2_o21ai_1 _10818_ (.B1(net1922),
    .Y(_03496_),
    .A1(net1670),
    .A2(net3146));
 sg13g2_a21oi_1 _10819_ (.A1(net1670),
    .A2(_03495_),
    .Y(_00570_),
    .B1(_03496_));
 sg13g2_nor2_1 _10820_ (.A(_03486_),
    .B(_03493_),
    .Y(_03497_));
 sg13g2_and3_1 _10821_ (.X(_03498_),
    .A(_03472_),
    .B(_03482_),
    .C(_03497_));
 sg13g2_o21ai_1 _10822_ (.B1(net1693),
    .Y(_03499_),
    .A1(\am_sdr0.cic2.integ1[15] ),
    .A2(\am_sdr0.cic2.integ1[14] ));
 sg13g2_nand3_1 _10823_ (.B(_03487_),
    .C(_03499_),
    .A(_03476_),
    .Y(_03500_));
 sg13g2_a21oi_2 _10824_ (.B1(_03500_),
    .Y(_03501_),
    .A2(_03498_),
    .A1(_03474_));
 sg13g2_xnor2_1 _10825_ (.Y(_03502_),
    .A(net1695),
    .B(\am_sdr0.cic2.integ1[16] ));
 sg13g2_nor2_1 _10826_ (.A(_03501_),
    .B(_03502_),
    .Y(_03503_));
 sg13g2_inv_1 _10827_ (.Y(_03504_),
    .A(_03503_));
 sg13g2_xnor2_1 _10828_ (.Y(_03505_),
    .A(_03501_),
    .B(_03502_));
 sg13g2_o21ai_1 _10829_ (.B1(net1970),
    .Y(_03506_),
    .A1(net1675),
    .A2(net3156));
 sg13g2_a21oi_1 _10830_ (.A1(net1675),
    .A2(_03505_),
    .Y(_00571_),
    .B1(_03506_));
 sg13g2_xnor2_1 _10831_ (.Y(_03507_),
    .A(net1695),
    .B(\am_sdr0.cic2.integ1[17] ));
 sg13g2_a21oi_1 _10832_ (.A1(net1696),
    .A2(\am_sdr0.cic2.integ1[16] ),
    .Y(_03508_),
    .B1(_03503_));
 sg13g2_xnor2_1 _10833_ (.Y(_03509_),
    .A(_03507_),
    .B(_03508_));
 sg13g2_o21ai_1 _10834_ (.B1(net1971),
    .Y(_03510_),
    .A1(net1675),
    .A2(net3064));
 sg13g2_a21oi_1 _10835_ (.A1(net1675),
    .A2(_03509_),
    .Y(_00572_),
    .B1(_03510_));
 sg13g2_or2_1 _10836_ (.X(_03511_),
    .B(\am_sdr0.cic2.integ1[18] ),
    .A(net1695));
 sg13g2_and2_1 _10837_ (.A(net1695),
    .B(\am_sdr0.cic2.integ1[18] ),
    .X(_03512_));
 sg13g2_xnor2_1 _10838_ (.Y(_03513_),
    .A(net1695),
    .B(\am_sdr0.cic2.integ1[18] ));
 sg13g2_o21ai_1 _10839_ (.B1(net1695),
    .Y(_03514_),
    .A1(\am_sdr0.cic2.integ1[17] ),
    .A2(\am_sdr0.cic2.integ1[16] ));
 sg13g2_o21ai_1 _10840_ (.B1(_03514_),
    .Y(_03515_),
    .A1(_03504_),
    .A2(_03507_));
 sg13g2_xor2_1 _10841_ (.B(_03515_),
    .A(_03513_),
    .X(_03516_));
 sg13g2_o21ai_1 _10842_ (.B1(net1971),
    .Y(_03517_),
    .A1(net1676),
    .A2(net3187));
 sg13g2_a21oi_1 _10843_ (.A1(net1676),
    .A2(_03516_),
    .Y(_00573_),
    .B1(_03517_));
 sg13g2_xnor2_1 _10844_ (.Y(_03518_),
    .A(net1695),
    .B(\am_sdr0.cic2.integ1[19] ));
 sg13g2_a21oi_1 _10845_ (.A1(_03511_),
    .A2(_03515_),
    .Y(_03519_),
    .B1(_03512_));
 sg13g2_xnor2_1 _10846_ (.Y(_03520_),
    .A(_03518_),
    .B(_03519_));
 sg13g2_o21ai_1 _10847_ (.B1(net1970),
    .Y(_03521_),
    .A1(net1679),
    .A2(net3037));
 sg13g2_a21oi_1 _10848_ (.A1(net1679),
    .A2(_03520_),
    .Y(_00574_),
    .B1(_03521_));
 sg13g2_xor2_1 _10849_ (.B(\am_sdr0.cic2.integ1[20] ),
    .A(net1697),
    .X(_03522_));
 sg13g2_nor4_1 _10850_ (.A(_03502_),
    .B(_03507_),
    .C(_03513_),
    .D(_03518_),
    .Y(_03523_));
 sg13g2_nor2b_2 _10851_ (.A(_03501_),
    .B_N(_03523_),
    .Y(_03524_));
 sg13g2_o21ai_1 _10852_ (.B1(net1695),
    .Y(_03525_),
    .A1(\am_sdr0.cic2.integ1[19] ),
    .A2(\am_sdr0.cic2.integ1[18] ));
 sg13g2_and2_1 _10853_ (.A(_03514_),
    .B(_03525_),
    .X(_03526_));
 sg13g2_inv_1 _10854_ (.Y(_03527_),
    .A(_03526_));
 sg13g2_nor3_1 _10855_ (.A(_03522_),
    .B(_03524_),
    .C(_03527_),
    .Y(_03528_));
 sg13g2_o21ai_1 _10856_ (.B1(_03522_),
    .Y(_03529_),
    .A1(_03524_),
    .A2(_03527_));
 sg13g2_nor2b_1 _10857_ (.A(_03528_),
    .B_N(_03529_),
    .Y(_03530_));
 sg13g2_o21ai_1 _10858_ (.B1(net2003),
    .Y(_03531_),
    .A1(net1636),
    .A2(_03530_));
 sg13g2_a21oi_1 _10859_ (.A1(net1636),
    .A2(_01391_),
    .Y(_00575_),
    .B1(_03531_));
 sg13g2_xor2_1 _10860_ (.B(\am_sdr0.cic2.integ1[21] ),
    .A(net1697),
    .X(_03532_));
 sg13g2_inv_1 _10861_ (.Y(_03533_),
    .A(_03532_));
 sg13g2_o21ai_1 _10862_ (.B1(_03529_),
    .Y(_03534_),
    .A1(_01304_),
    .A2(_01391_));
 sg13g2_xnor2_1 _10863_ (.Y(_03535_),
    .A(_03532_),
    .B(_03534_));
 sg13g2_o21ai_1 _10864_ (.B1(net2003),
    .Y(_03536_),
    .A1(net1686),
    .A2(net2919));
 sg13g2_a21oi_1 _10865_ (.A1(net1686),
    .A2(_03535_),
    .Y(_00576_),
    .B1(_03536_));
 sg13g2_or2_1 _10866_ (.X(_03537_),
    .B(\am_sdr0.cic2.integ1[22] ),
    .A(net1698));
 sg13g2_and2_1 _10867_ (.A(net1697),
    .B(\am_sdr0.cic2.integ1[22] ),
    .X(_03538_));
 sg13g2_xnor2_1 _10868_ (.Y(_03539_),
    .A(net1697),
    .B(\am_sdr0.cic2.integ1[22] ));
 sg13g2_o21ai_1 _10869_ (.B1(net1697),
    .Y(_03540_),
    .A1(\am_sdr0.cic2.integ1[21] ),
    .A2(\am_sdr0.cic2.integ1[20] ));
 sg13g2_o21ai_1 _10870_ (.B1(_03540_),
    .Y(_03541_),
    .A1(_03529_),
    .A2(_03533_));
 sg13g2_xor2_1 _10871_ (.B(_03541_),
    .A(_03539_),
    .X(_03542_));
 sg13g2_o21ai_1 _10872_ (.B1(net2004),
    .Y(_03543_),
    .A1(net1685),
    .A2(net3161));
 sg13g2_a21oi_1 _10873_ (.A1(net1685),
    .A2(_03542_),
    .Y(_00577_),
    .B1(_03543_));
 sg13g2_xnor2_1 _10874_ (.Y(_03544_),
    .A(net1697),
    .B(\am_sdr0.cic2.integ1[23] ));
 sg13g2_a21oi_1 _10875_ (.A1(_03537_),
    .A2(_03541_),
    .Y(_03545_),
    .B1(_03538_));
 sg13g2_xnor2_1 _10876_ (.Y(_03546_),
    .A(_03544_),
    .B(_03545_));
 sg13g2_o21ai_1 _10877_ (.B1(net2003),
    .Y(_03547_),
    .A1(net1685),
    .A2(net3056));
 sg13g2_a21oi_1 _10878_ (.A1(net1685),
    .A2(_03546_),
    .Y(_00578_),
    .B1(_03547_));
 sg13g2_nand2_1 _10879_ (.Y(_03548_),
    .A(_03522_),
    .B(_03532_));
 sg13g2_nor3_1 _10880_ (.A(_03539_),
    .B(_03544_),
    .C(_03548_),
    .Y(_03549_));
 sg13g2_o21ai_1 _10881_ (.B1(net1697),
    .Y(_03550_),
    .A1(\am_sdr0.cic2.integ1[23] ),
    .A2(\am_sdr0.cic2.integ1[22] ));
 sg13g2_nand3_1 _10882_ (.B(_03540_),
    .C(_03550_),
    .A(_03526_),
    .Y(_03551_));
 sg13g2_a21oi_2 _10883_ (.B1(_03551_),
    .Y(_03552_),
    .A2(_03549_),
    .A1(_03524_));
 sg13g2_xnor2_1 _10884_ (.Y(_03553_),
    .A(net1697),
    .B(\am_sdr0.cic2.integ1[24] ));
 sg13g2_xnor2_1 _10885_ (.Y(_03554_),
    .A(_03552_),
    .B(_03553_));
 sg13g2_o21ai_1 _10886_ (.B1(net2003),
    .Y(_03555_),
    .A1(net1685),
    .A2(net3158));
 sg13g2_a21oi_1 _10887_ (.A1(net1685),
    .A2(_03554_),
    .Y(_00579_),
    .B1(_03555_));
 sg13g2_a21o_1 _10888_ (.A2(\am_sdr0.cic2.integ1[24] ),
    .A1(_01304_),
    .B1(_03552_),
    .X(_03556_));
 sg13g2_o21ai_1 _10889_ (.B1(_03552_),
    .Y(_03557_),
    .A1(_01304_),
    .A2(\am_sdr0.cic2.integ1[24] ));
 sg13g2_and3_1 _10890_ (.X(_03558_),
    .A(net1685),
    .B(_03556_),
    .C(_03557_));
 sg13g2_o21ai_1 _10891_ (.B1(net2005),
    .Y(_03559_),
    .A1(net1351),
    .A2(_03558_));
 sg13g2_a21oi_1 _10892_ (.A1(net1351),
    .A2(_03558_),
    .Y(_00580_),
    .B1(_03559_));
 sg13g2_a21oi_1 _10893_ (.A1(net1689),
    .A2(\am_sdr0.cic2.integ1[3] ),
    .Y(_03560_),
    .B1(net1300));
 sg13g2_nand2_1 _10894_ (.Y(_03561_),
    .A(net1300),
    .B(\am_sdr0.cic2.integ1[3] ));
 sg13g2_nor2_1 _10895_ (.A(net1636),
    .B(_03561_),
    .Y(_03562_));
 sg13g2_nor3_1 _10896_ (.A(net1891),
    .B(net1301),
    .C(_03562_),
    .Y(_00581_));
 sg13g2_nand2_1 _10897_ (.Y(_03563_),
    .A(\am_sdr0.cic2.integ2[1] ),
    .B(\am_sdr0.cic2.integ1[4] ));
 sg13g2_xnor2_1 _10898_ (.Y(_03564_),
    .A(net2815),
    .B(\am_sdr0.cic2.integ1[4] ));
 sg13g2_xnor2_1 _10899_ (.Y(_03565_),
    .A(_03561_),
    .B(_03564_));
 sg13g2_o21ai_1 _10900_ (.B1(net2003),
    .Y(_03566_),
    .A1(net1684),
    .A2(net2815));
 sg13g2_a21oi_1 _10901_ (.A1(net1683),
    .A2(_03565_),
    .Y(_00582_),
    .B1(_03566_));
 sg13g2_and2_1 _10902_ (.A(\am_sdr0.cic2.integ2[2] ),
    .B(\am_sdr0.cic2.integ1[5] ),
    .X(_03567_));
 sg13g2_xor2_1 _10903_ (.B(\am_sdr0.cic2.integ1[5] ),
    .A(net2715),
    .X(_03568_));
 sg13g2_o21ai_1 _10904_ (.B1(_03563_),
    .Y(_03569_),
    .A1(_03561_),
    .A2(_03564_));
 sg13g2_and2_1 _10905_ (.A(_03568_),
    .B(_03569_),
    .X(_03570_));
 sg13g2_xnor2_1 _10906_ (.Y(_03571_),
    .A(_03568_),
    .B(_03569_));
 sg13g2_o21ai_1 _10907_ (.B1(net2003),
    .Y(_03572_),
    .A1(net1684),
    .A2(net2715));
 sg13g2_a21oi_1 _10908_ (.A1(net1684),
    .A2(_03571_),
    .Y(_00583_),
    .B1(_03572_));
 sg13g2_nand2_1 _10909_ (.Y(_03573_),
    .A(\am_sdr0.cic2.integ2[3] ),
    .B(\am_sdr0.cic2.integ1[6] ));
 sg13g2_xor2_1 _10910_ (.B(\am_sdr0.cic2.integ1[6] ),
    .A(\am_sdr0.cic2.integ2[3] ),
    .X(_03574_));
 sg13g2_nor2_1 _10911_ (.A(_03567_),
    .B(_03570_),
    .Y(_03575_));
 sg13g2_o21ai_1 _10912_ (.B1(_03574_),
    .Y(_03576_),
    .A1(_03567_),
    .A2(_03570_));
 sg13g2_xnor2_1 _10913_ (.Y(_03577_),
    .A(_03574_),
    .B(_03575_));
 sg13g2_o21ai_1 _10914_ (.B1(net2003),
    .Y(_03578_),
    .A1(net1636),
    .A2(_03577_));
 sg13g2_a21oi_1 _10915_ (.A1(net1636),
    .A2(_01390_),
    .Y(_00584_),
    .B1(_03578_));
 sg13g2_nand2_1 _10916_ (.Y(_03579_),
    .A(\am_sdr0.cic2.integ2[4] ),
    .B(\am_sdr0.cic2.integ1[7] ));
 sg13g2_xnor2_1 _10917_ (.Y(_03580_),
    .A(\am_sdr0.cic2.integ2[4] ),
    .B(\am_sdr0.cic2.integ1[7] ));
 sg13g2_nand3_1 _10918_ (.B(_03576_),
    .C(_03580_),
    .A(_03573_),
    .Y(_03581_));
 sg13g2_a21o_1 _10919_ (.A2(_03576_),
    .A1(_03573_),
    .B1(_03580_),
    .X(_03582_));
 sg13g2_nand2_1 _10920_ (.Y(_03583_),
    .A(_03581_),
    .B(_03582_));
 sg13g2_o21ai_1 _10921_ (.B1(net2003),
    .Y(_03584_),
    .A1(net1683),
    .A2(net3172));
 sg13g2_a21oi_1 _10922_ (.A1(net1683),
    .A2(_03583_),
    .Y(_00585_),
    .B1(_03584_));
 sg13g2_xor2_1 _10923_ (.B(\am_sdr0.cic2.integ1[8] ),
    .A(\am_sdr0.cic2.integ2[5] ),
    .X(_03585_));
 sg13g2_nand2_1 _10924_ (.Y(_03586_),
    .A(_03579_),
    .B(_03582_));
 sg13g2_xnor2_1 _10925_ (.Y(_03587_),
    .A(_03585_),
    .B(_03586_));
 sg13g2_o21ai_1 _10926_ (.B1(net1972),
    .Y(_03588_),
    .A1(net1678),
    .A2(net3107));
 sg13g2_a21oi_1 _10927_ (.A1(net1678),
    .A2(_03587_),
    .Y(_00586_),
    .B1(_03588_));
 sg13g2_and2_1 _10928_ (.A(\am_sdr0.cic2.integ2[6] ),
    .B(\am_sdr0.cic2.integ1[9] ),
    .X(_03589_));
 sg13g2_xnor2_1 _10929_ (.Y(_03590_),
    .A(\am_sdr0.cic2.integ2[6] ),
    .B(\am_sdr0.cic2.integ1[9] ));
 sg13g2_a22oi_1 _10930_ (.Y(_03591_),
    .B1(\am_sdr0.cic2.integ1[7] ),
    .B2(\am_sdr0.cic2.integ2[4] ),
    .A2(\am_sdr0.cic2.integ1[8] ),
    .A1(\am_sdr0.cic2.integ2[5] ));
 sg13g2_a22oi_1 _10931_ (.Y(_03592_),
    .B1(_03582_),
    .B2(_03591_),
    .A2(_01392_),
    .A1(_01389_));
 sg13g2_a221oi_1 _10932_ (.B2(_03591_),
    .C1(_03590_),
    .B1(_03582_),
    .A1(_01389_),
    .Y(_03593_),
    .A2(_01392_));
 sg13g2_xnor2_1 _10933_ (.Y(_03594_),
    .A(_03590_),
    .B(_03592_));
 sg13g2_o21ai_1 _10934_ (.B1(net1972),
    .Y(_03595_),
    .A1(net1635),
    .A2(_03594_));
 sg13g2_a21oi_1 _10935_ (.A1(net1635),
    .A2(_01388_),
    .Y(_00587_),
    .B1(_03595_));
 sg13g2_nand2_2 _10936_ (.Y(_03596_),
    .A(\am_sdr0.cic2.integ2[7] ),
    .B(\am_sdr0.cic2.integ1[10] ));
 sg13g2_xor2_1 _10937_ (.B(\am_sdr0.cic2.integ1[10] ),
    .A(\am_sdr0.cic2.integ2[7] ),
    .X(_03597_));
 sg13g2_o21ai_1 _10938_ (.B1(_03597_),
    .Y(_03598_),
    .A1(_03589_),
    .A2(_03593_));
 sg13g2_or3_1 _10939_ (.A(_03589_),
    .B(_03593_),
    .C(_03597_),
    .X(_03599_));
 sg13g2_a21oi_1 _10940_ (.A1(_03598_),
    .A2(_03599_),
    .Y(_03600_),
    .B1(net1635));
 sg13g2_o21ai_1 _10941_ (.B1(net1972),
    .Y(_03601_),
    .A1(net1678),
    .A2(net3155));
 sg13g2_nor2_1 _10942_ (.A(_03600_),
    .B(_03601_),
    .Y(_00588_));
 sg13g2_and2_1 _10943_ (.A(\am_sdr0.cic2.integ2[8] ),
    .B(\am_sdr0.cic2.integ1[11] ),
    .X(_03602_));
 sg13g2_xnor2_1 _10944_ (.Y(_03603_),
    .A(\am_sdr0.cic2.integ2[8] ),
    .B(\am_sdr0.cic2.integ1[11] ));
 sg13g2_a21oi_2 _10945_ (.B1(_03603_),
    .Y(_03604_),
    .A2(_03598_),
    .A1(_03596_));
 sg13g2_and3_1 _10946_ (.X(_03605_),
    .A(_03596_),
    .B(_03598_),
    .C(_03603_));
 sg13g2_o21ai_1 _10947_ (.B1(net1671),
    .Y(_03606_),
    .A1(_03604_),
    .A2(_03605_));
 sg13g2_o21ai_1 _10948_ (.B1(_03606_),
    .Y(_03607_),
    .A1(net1677),
    .A2(net3120));
 sg13g2_nor2_1 _10949_ (.A(net1889),
    .B(_03607_),
    .Y(_00589_));
 sg13g2_or2_1 _10950_ (.X(_03608_),
    .B(\am_sdr0.cic2.integ1[12] ),
    .A(\am_sdr0.cic2.integ2[9] ));
 sg13g2_nand2_1 _10951_ (.Y(_03609_),
    .A(\am_sdr0.cic2.integ2[9] ),
    .B(\am_sdr0.cic2.integ1[12] ));
 sg13g2_and2_1 _10952_ (.A(_03608_),
    .B(_03609_),
    .X(_03610_));
 sg13g2_nor2_1 _10953_ (.A(_03602_),
    .B(_03604_),
    .Y(_03611_));
 sg13g2_xnor2_1 _10954_ (.Y(_03612_),
    .A(_03610_),
    .B(_03611_));
 sg13g2_nor2_1 _10955_ (.A(net1635),
    .B(_03612_),
    .Y(_03613_));
 sg13g2_o21ai_1 _10956_ (.B1(net1970),
    .Y(_03614_),
    .A1(net1671),
    .A2(net2968));
 sg13g2_nor2_1 _10957_ (.A(_03613_),
    .B(_03614_),
    .Y(_00590_));
 sg13g2_and2_1 _10958_ (.A(\am_sdr0.cic2.integ2[10] ),
    .B(\am_sdr0.cic2.integ1[13] ),
    .X(_03615_));
 sg13g2_xnor2_1 _10959_ (.Y(_03616_),
    .A(\am_sdr0.cic2.integ2[10] ),
    .B(\am_sdr0.cic2.integ1[13] ));
 sg13g2_o21ai_1 _10960_ (.B1(_03608_),
    .Y(_03617_),
    .A1(_03602_),
    .A2(_03604_));
 sg13g2_nand2_1 _10961_ (.Y(_03618_),
    .A(_03609_),
    .B(_03617_));
 sg13g2_a21oi_1 _10962_ (.A1(_03609_),
    .A2(_03617_),
    .Y(_03619_),
    .B1(_03616_));
 sg13g2_xor2_1 _10963_ (.B(_03618_),
    .A(_03616_),
    .X(_03620_));
 sg13g2_o21ai_1 _10964_ (.B1(net1970),
    .Y(_03621_),
    .A1(net1671),
    .A2(net3060));
 sg13g2_a21oi_1 _10965_ (.A1(net1671),
    .A2(_03620_),
    .Y(_00591_),
    .B1(_03621_));
 sg13g2_xnor2_1 _10966_ (.Y(_03622_),
    .A(\am_sdr0.cic2.integ2[11] ),
    .B(\am_sdr0.cic2.integ1[14] ));
 sg13g2_nor3_1 _10967_ (.A(_03615_),
    .B(_03619_),
    .C(_03622_),
    .Y(_03623_));
 sg13g2_o21ai_1 _10968_ (.B1(_03622_),
    .Y(_03624_),
    .A1(_03615_),
    .A2(_03619_));
 sg13g2_nor2_1 _10969_ (.A(net1635),
    .B(_03623_),
    .Y(_03625_));
 sg13g2_o21ai_1 _10970_ (.B1(net1970),
    .Y(_03626_),
    .A1(net1671),
    .A2(net3186));
 sg13g2_a21oi_1 _10971_ (.A1(_03624_),
    .A2(_03625_),
    .Y(_00592_),
    .B1(_03626_));
 sg13g2_nand2_1 _10972_ (.Y(_03627_),
    .A(\am_sdr0.cic2.integ2[12] ),
    .B(\am_sdr0.cic2.integ1[15] ));
 sg13g2_xor2_1 _10973_ (.B(\am_sdr0.cic2.integ1[15] ),
    .A(\am_sdr0.cic2.integ2[12] ),
    .X(_03628_));
 sg13g2_nor2_1 _10974_ (.A(_03616_),
    .B(_03622_),
    .Y(_03629_));
 sg13g2_nand2_1 _10975_ (.Y(_03630_),
    .A(_03602_),
    .B(_03608_));
 sg13g2_nand2_1 _10976_ (.Y(_03631_),
    .A(_03609_),
    .B(_03630_));
 sg13g2_o21ai_1 _10977_ (.B1(_03615_),
    .Y(_03632_),
    .A1(\am_sdr0.cic2.integ2[11] ),
    .A2(\am_sdr0.cic2.integ1[14] ));
 sg13g2_a22oi_1 _10978_ (.Y(_03633_),
    .B1(_03629_),
    .B2(_03631_),
    .A2(\am_sdr0.cic2.integ1[14] ),
    .A1(\am_sdr0.cic2.integ2[11] ));
 sg13g2_nand2_1 _10979_ (.Y(_03634_),
    .A(_03632_),
    .B(_03633_));
 sg13g2_nand3b_1 _10980_ (.B(_03610_),
    .C(_03629_),
    .Y(_03635_),
    .A_N(_03603_));
 sg13g2_a21oi_2 _10981_ (.B1(_03635_),
    .Y(_03636_),
    .A2(_03598_),
    .A1(_03596_));
 sg13g2_o21ai_1 _10982_ (.B1(_03628_),
    .Y(_03637_),
    .A1(_03634_),
    .A2(_03636_));
 sg13g2_or3_1 _10983_ (.A(_03628_),
    .B(_03634_),
    .C(_03636_),
    .X(_03638_));
 sg13g2_nand2_1 _10984_ (.Y(_03639_),
    .A(_03637_),
    .B(_03638_));
 sg13g2_o21ai_1 _10985_ (.B1(net1964),
    .Y(_03640_),
    .A1(net1674),
    .A2(net3139));
 sg13g2_a21oi_1 _10986_ (.A1(net1674),
    .A2(_03639_),
    .Y(_00593_),
    .B1(_03640_));
 sg13g2_nor2_1 _10987_ (.A(\am_sdr0.cic2.integ2[13] ),
    .B(\am_sdr0.cic2.integ1[16] ),
    .Y(_03641_));
 sg13g2_xor2_1 _10988_ (.B(\am_sdr0.cic2.integ1[16] ),
    .A(\am_sdr0.cic2.integ2[13] ),
    .X(_03642_));
 sg13g2_nand2_1 _10989_ (.Y(_03643_),
    .A(_03627_),
    .B(_03637_));
 sg13g2_xnor2_1 _10990_ (.Y(_03644_),
    .A(_03642_),
    .B(_03643_));
 sg13g2_o21ai_1 _10991_ (.B1(net1964),
    .Y(_03645_),
    .A1(net1674),
    .A2(net3141));
 sg13g2_a21oi_1 _10992_ (.A1(net1674),
    .A2(_03644_),
    .Y(_00594_),
    .B1(_03645_));
 sg13g2_and2_1 _10993_ (.A(\am_sdr0.cic2.integ2[14] ),
    .B(\am_sdr0.cic2.integ1[17] ),
    .X(_03646_));
 sg13g2_xor2_1 _10994_ (.B(\am_sdr0.cic2.integ1[17] ),
    .A(\am_sdr0.cic2.integ2[14] ),
    .X(_03647_));
 sg13g2_a22oi_1 _10995_ (.Y(_03648_),
    .B1(\am_sdr0.cic2.integ1[15] ),
    .B2(\am_sdr0.cic2.integ2[12] ),
    .A2(\am_sdr0.cic2.integ1[16] ),
    .A1(\am_sdr0.cic2.integ2[13] ));
 sg13g2_nor2_1 _10996_ (.A(_03641_),
    .B(_03648_),
    .Y(_03649_));
 sg13g2_a21oi_1 _10997_ (.A1(_03637_),
    .A2(_03648_),
    .Y(_03650_),
    .B1(_03641_));
 sg13g2_xnor2_1 _10998_ (.Y(_03651_),
    .A(_03647_),
    .B(_03650_));
 sg13g2_o21ai_1 _10999_ (.B1(net1971),
    .Y(_03652_),
    .A1(net1674),
    .A2(net3080));
 sg13g2_a21oi_1 _11000_ (.A1(net1676),
    .A2(_03651_),
    .Y(_00595_),
    .B1(_03652_));
 sg13g2_nand2_1 _11001_ (.Y(_03653_),
    .A(\am_sdr0.cic2.integ2[15] ),
    .B(\am_sdr0.cic2.integ1[18] ));
 sg13g2_xor2_1 _11002_ (.B(\am_sdr0.cic2.integ1[18] ),
    .A(\am_sdr0.cic2.integ2[15] ),
    .X(_03654_));
 sg13g2_a21oi_1 _11003_ (.A1(_03647_),
    .A2(_03650_),
    .Y(_03655_),
    .B1(_03646_));
 sg13g2_xor2_1 _11004_ (.B(_03655_),
    .A(_03654_),
    .X(_03656_));
 sg13g2_o21ai_1 _11005_ (.B1(net1971),
    .Y(_03657_),
    .A1(net1675),
    .A2(net3185));
 sg13g2_a21oi_1 _11006_ (.A1(net1675),
    .A2(_03656_),
    .Y(_00596_),
    .B1(_03657_));
 sg13g2_nand2_1 _11007_ (.Y(_03658_),
    .A(\am_sdr0.cic2.integ2[16] ),
    .B(\am_sdr0.cic2.integ1[19] ));
 sg13g2_xnor2_1 _11008_ (.Y(_03659_),
    .A(\am_sdr0.cic2.integ2[16] ),
    .B(\am_sdr0.cic2.integ1[19] ));
 sg13g2_and2_1 _11009_ (.A(_03647_),
    .B(_03654_),
    .X(_03660_));
 sg13g2_and3_1 _11010_ (.X(_03661_),
    .A(_03628_),
    .B(_03642_),
    .C(_03660_));
 sg13g2_o21ai_1 _11011_ (.B1(_03646_),
    .Y(_03662_),
    .A1(\am_sdr0.cic2.integ2[15] ),
    .A2(\am_sdr0.cic2.integ1[18] ));
 sg13g2_nand2_1 _11012_ (.Y(_03663_),
    .A(_03634_),
    .B(_03661_));
 sg13g2_nand3_1 _11013_ (.B(_03662_),
    .C(_03663_),
    .A(_03653_),
    .Y(_03664_));
 sg13g2_a221oi_1 _11014_ (.B2(_03636_),
    .C1(_03664_),
    .B1(_03661_),
    .A1(_03649_),
    .Y(_03665_),
    .A2(_03660_));
 sg13g2_xnor2_1 _11015_ (.Y(_03666_),
    .A(_03659_),
    .B(_03665_));
 sg13g2_o21ai_1 _11016_ (.B1(net1973),
    .Y(_03667_),
    .A1(net1679),
    .A2(net3070));
 sg13g2_a21oi_1 _11017_ (.A1(net1679),
    .A2(_03666_),
    .Y(_00597_),
    .B1(_03667_));
 sg13g2_or2_1 _11018_ (.X(_03668_),
    .B(\am_sdr0.cic2.integ1[20] ),
    .A(\am_sdr0.cic2.integ2[17] ));
 sg13g2_nand2_1 _11019_ (.Y(_03669_),
    .A(\am_sdr0.cic2.integ2[17] ),
    .B(\am_sdr0.cic2.integ1[20] ));
 sg13g2_nand2_1 _11020_ (.Y(_03670_),
    .A(_03668_),
    .B(_03669_));
 sg13g2_o21ai_1 _11021_ (.B1(_03658_),
    .Y(_03671_),
    .A1(_03659_),
    .A2(_03665_));
 sg13g2_xor2_1 _11022_ (.B(_03671_),
    .A(_03670_),
    .X(_03672_));
 sg13g2_o21ai_1 _11023_ (.B1(net1973),
    .Y(_03673_),
    .A1(net1686),
    .A2(net3028));
 sg13g2_a21oi_1 _11024_ (.A1(net1686),
    .A2(_03672_),
    .Y(_00598_),
    .B1(_03673_));
 sg13g2_and2_1 _11025_ (.A(\am_sdr0.cic2.integ2[18] ),
    .B(\am_sdr0.cic2.integ1[21] ),
    .X(_03674_));
 sg13g2_or2_1 _11026_ (.X(_03675_),
    .B(\am_sdr0.cic2.integ1[21] ),
    .A(\am_sdr0.cic2.integ2[18] ));
 sg13g2_nand2b_1 _11027_ (.Y(_03676_),
    .B(_03675_),
    .A_N(_03674_));
 sg13g2_or2_1 _11028_ (.X(_03677_),
    .B(_03670_),
    .A(_03659_));
 sg13g2_nand2_1 _11029_ (.Y(_03678_),
    .A(_03658_),
    .B(_03669_));
 sg13g2_nand2_1 _11030_ (.Y(_03679_),
    .A(_03668_),
    .B(_03678_));
 sg13g2_o21ai_1 _11031_ (.B1(_03679_),
    .Y(_03680_),
    .A1(_03665_),
    .A2(_03677_));
 sg13g2_xor2_1 _11032_ (.B(_03680_),
    .A(_03676_),
    .X(_03681_));
 sg13g2_o21ai_1 _11033_ (.B1(net2004),
    .Y(_03682_),
    .A1(net1686),
    .A2(net3079));
 sg13g2_a21oi_1 _11034_ (.A1(net1686),
    .A2(_03681_),
    .Y(_00599_),
    .B1(_03682_));
 sg13g2_nand2_1 _11035_ (.Y(_03683_),
    .A(\am_sdr0.cic2.integ2[19] ),
    .B(\am_sdr0.cic2.integ1[22] ));
 sg13g2_xnor2_1 _11036_ (.Y(_03684_),
    .A(\am_sdr0.cic2.integ2[19] ),
    .B(\am_sdr0.cic2.integ1[22] ));
 sg13g2_a21oi_1 _11037_ (.A1(_03675_),
    .A2(_03680_),
    .Y(_03685_),
    .B1(_03674_));
 sg13g2_xnor2_1 _11038_ (.Y(_03686_),
    .A(_03684_),
    .B(_03685_));
 sg13g2_o21ai_1 _11039_ (.B1(net2004),
    .Y(_03687_),
    .A1(net1687),
    .A2(net3068));
 sg13g2_a21oi_1 _11040_ (.A1(net1687),
    .A2(_03686_),
    .Y(_00600_),
    .B1(_03687_));
 sg13g2_or3_1 _11041_ (.A(_03676_),
    .B(_03677_),
    .C(_03684_),
    .X(_03688_));
 sg13g2_nor3_1 _11042_ (.A(_03676_),
    .B(_03679_),
    .C(_03684_),
    .Y(_03689_));
 sg13g2_o21ai_1 _11043_ (.B1(_03674_),
    .Y(_03690_),
    .A1(\am_sdr0.cic2.integ2[19] ),
    .A2(\am_sdr0.cic2.integ1[22] ));
 sg13g2_nand2_1 _11044_ (.Y(_03691_),
    .A(_03683_),
    .B(_03690_));
 sg13g2_nor2_1 _11045_ (.A(_03689_),
    .B(_03691_),
    .Y(_03692_));
 sg13g2_o21ai_1 _11046_ (.B1(_03692_),
    .Y(_03693_),
    .A1(_03665_),
    .A2(_03688_));
 sg13g2_or2_1 _11047_ (.X(_03694_),
    .B(\am_sdr0.cic2.integ1[23] ),
    .A(\am_sdr0.cic2.integ2[20] ));
 sg13g2_and2_1 _11048_ (.A(\am_sdr0.cic2.integ2[20] ),
    .B(\am_sdr0.cic2.integ1[23] ),
    .X(_03695_));
 sg13g2_xnor2_1 _11049_ (.Y(_03696_),
    .A(\am_sdr0.cic2.integ2[20] ),
    .B(\am_sdr0.cic2.integ1[23] ));
 sg13g2_xor2_1 _11050_ (.B(_03696_),
    .A(_03693_),
    .X(_03697_));
 sg13g2_o21ai_1 _11051_ (.B1(net2006),
    .Y(_03698_),
    .A1(net1690),
    .A2(net3101));
 sg13g2_a21oi_1 _11052_ (.A1(net1691),
    .A2(_03697_),
    .Y(_00601_),
    .B1(_03698_));
 sg13g2_xnor2_1 _11053_ (.Y(_03699_),
    .A(\am_sdr0.cic2.integ2[21] ),
    .B(\am_sdr0.cic2.integ1[24] ));
 sg13g2_a21oi_1 _11054_ (.A1(_03693_),
    .A2(_03694_),
    .Y(_03700_),
    .B1(_03695_));
 sg13g2_xnor2_1 _11055_ (.Y(_03701_),
    .A(_03699_),
    .B(_03700_));
 sg13g2_o21ai_1 _11056_ (.B1(net2006),
    .Y(_03702_),
    .A1(net1690),
    .A2(net2923));
 sg13g2_a21oi_1 _11057_ (.A1(net1690),
    .A2(_03701_),
    .Y(_00602_),
    .B1(_03702_));
 sg13g2_nor2_1 _11058_ (.A(_03696_),
    .B(_03699_),
    .Y(_03703_));
 sg13g2_o21ai_1 _11059_ (.B1(_03695_),
    .Y(_03704_),
    .A1(\am_sdr0.cic2.integ2[21] ),
    .A2(\am_sdr0.cic2.integ1[24] ));
 sg13g2_inv_1 _11060_ (.Y(_03705_),
    .A(_03704_));
 sg13g2_a221oi_1 _11061_ (.B2(_03703_),
    .C1(_03705_),
    .B1(_03693_),
    .A1(\am_sdr0.cic2.integ2[21] ),
    .Y(_03706_),
    .A2(\am_sdr0.cic2.integ1[24] ));
 sg13g2_xor2_1 _11062_ (.B(net1351),
    .A(net2809),
    .X(_03707_));
 sg13g2_or2_1 _11063_ (.X(_03708_),
    .B(_03707_),
    .A(_03706_));
 sg13g2_a21oi_1 _11064_ (.A1(_03706_),
    .A2(_03707_),
    .Y(_03709_),
    .B1(net1636));
 sg13g2_o21ai_1 _11065_ (.B1(net2005),
    .Y(_03710_),
    .A1(net1690),
    .A2(net2809));
 sg13g2_a21oi_1 _11066_ (.A1(_03708_),
    .A2(_03709_),
    .Y(_00603_),
    .B1(_03710_));
 sg13g2_a21oi_1 _11067_ (.A1(net1692),
    .A2(\am_sdr0.cic2.integ2[3] ),
    .Y(_03711_),
    .B1(net1464));
 sg13g2_nand2_1 _11068_ (.Y(_03712_),
    .A(net1464),
    .B(\am_sdr0.cic2.integ2[3] ));
 sg13g2_nor2_1 _11069_ (.A(net1636),
    .B(_03712_),
    .Y(_03713_));
 sg13g2_nor3_1 _11070_ (.A(net1891),
    .B(net1465),
    .C(_03713_),
    .Y(_00604_));
 sg13g2_nand2_1 _11071_ (.Y(_03714_),
    .A(\am_sdr0.cic2.integ3[1] ),
    .B(\am_sdr0.cic2.integ2[4] ));
 sg13g2_xnor2_1 _11072_ (.Y(_03715_),
    .A(net2629),
    .B(\am_sdr0.cic2.integ2[4] ));
 sg13g2_xnor2_1 _11073_ (.Y(_03716_),
    .A(_03712_),
    .B(_03715_));
 sg13g2_o21ai_1 _11074_ (.B1(net2005),
    .Y(_03717_),
    .A1(net1689),
    .A2(net2629));
 sg13g2_a21oi_1 _11075_ (.A1(net1689),
    .A2(_03716_),
    .Y(_00605_),
    .B1(_03717_));
 sg13g2_and2_1 _11076_ (.A(\am_sdr0.cic2.integ3[2] ),
    .B(\am_sdr0.cic2.integ2[5] ),
    .X(_03718_));
 sg13g2_xor2_1 _11077_ (.B(\am_sdr0.cic2.integ2[5] ),
    .A(\am_sdr0.cic2.integ3[2] ),
    .X(_03719_));
 sg13g2_o21ai_1 _11078_ (.B1(_03714_),
    .Y(_03720_),
    .A1(_03712_),
    .A2(_03715_));
 sg13g2_and2_1 _11079_ (.A(_03719_),
    .B(_03720_),
    .X(_03721_));
 sg13g2_xnor2_1 _11080_ (.Y(_03722_),
    .A(_03719_),
    .B(_03720_));
 sg13g2_o21ai_1 _11081_ (.B1(net1972),
    .Y(_03723_),
    .A1(net1678),
    .A2(net2604));
 sg13g2_a21oi_1 _11082_ (.A1(net1678),
    .A2(_03722_),
    .Y(_00606_),
    .B1(_03723_));
 sg13g2_nand2_1 _11083_ (.Y(_03724_),
    .A(net2634),
    .B(net2834));
 sg13g2_xor2_1 _11084_ (.B(\am_sdr0.cic2.integ2[6] ),
    .A(\am_sdr0.cic2.integ3[3] ),
    .X(_03725_));
 sg13g2_nor2_1 _11085_ (.A(_03718_),
    .B(_03721_),
    .Y(_03726_));
 sg13g2_o21ai_1 _11086_ (.B1(_03725_),
    .Y(_03727_),
    .A1(_03718_),
    .A2(_03721_));
 sg13g2_xnor2_1 _11087_ (.Y(_03728_),
    .A(_03725_),
    .B(_03726_));
 sg13g2_o21ai_1 _11088_ (.B1(net1972),
    .Y(_03729_),
    .A1(net1635),
    .A2(_03728_));
 sg13g2_a21oi_1 _11089_ (.A1(net1635),
    .A2(_01386_),
    .Y(_00607_),
    .B1(_03729_));
 sg13g2_nand2_1 _11090_ (.Y(_03730_),
    .A(\am_sdr0.cic2.integ3[4] ),
    .B(\am_sdr0.cic2.integ2[7] ));
 sg13g2_xnor2_1 _11091_ (.Y(_03731_),
    .A(\am_sdr0.cic2.integ3[4] ),
    .B(\am_sdr0.cic2.integ2[7] ));
 sg13g2_nand3_1 _11092_ (.B(_03727_),
    .C(_03731_),
    .A(_03724_),
    .Y(_03732_));
 sg13g2_a21o_1 _11093_ (.A2(_03727_),
    .A1(_03724_),
    .B1(_03731_),
    .X(_03733_));
 sg13g2_nand2_1 _11094_ (.Y(_03734_),
    .A(_03732_),
    .B(_03733_));
 sg13g2_o21ai_1 _11095_ (.B1(net1972),
    .Y(_03735_),
    .A1(net1679),
    .A2(net2818));
 sg13g2_a21oi_1 _11096_ (.A1(net1679),
    .A2(_03734_),
    .Y(_00608_),
    .B1(_03735_));
 sg13g2_xor2_1 _11097_ (.B(\am_sdr0.cic2.integ2[8] ),
    .A(net2811),
    .X(_03736_));
 sg13g2_nand2_1 _11098_ (.Y(_03737_),
    .A(_03730_),
    .B(_03733_));
 sg13g2_xnor2_1 _11099_ (.Y(_03738_),
    .A(_03736_),
    .B(_03737_));
 sg13g2_o21ai_1 _11100_ (.B1(net1970),
    .Y(_03739_),
    .A1(net1678),
    .A2(net2811));
 sg13g2_a21oi_1 _11101_ (.A1(net1677),
    .A2(_03738_),
    .Y(_00609_),
    .B1(_03739_));
 sg13g2_and2_1 _11102_ (.A(\am_sdr0.cic2.integ3[6] ),
    .B(\am_sdr0.cic2.integ2[9] ),
    .X(_03740_));
 sg13g2_xor2_1 _11103_ (.B(\am_sdr0.cic2.integ2[9] ),
    .A(net2991),
    .X(_03741_));
 sg13g2_inv_1 _11104_ (.Y(_03742_),
    .A(_03741_));
 sg13g2_a22oi_1 _11105_ (.Y(_03743_),
    .B1(\am_sdr0.cic2.integ2[7] ),
    .B2(\am_sdr0.cic2.integ3[4] ),
    .A2(\am_sdr0.cic2.integ2[8] ),
    .A1(\am_sdr0.cic2.integ3[5] ));
 sg13g2_a22oi_1 _11106_ (.Y(_03744_),
    .B1(_03733_),
    .B2(_03743_),
    .A2(_01387_),
    .A1(_01385_));
 sg13g2_a221oi_1 _11107_ (.B2(_03743_),
    .C1(_03742_),
    .B1(_03733_),
    .A1(_01385_),
    .Y(_03745_),
    .A2(_01387_));
 sg13g2_xnor2_1 _11108_ (.Y(_03746_),
    .A(_03741_),
    .B(_03744_));
 sg13g2_o21ai_1 _11109_ (.B1(net1970),
    .Y(_03747_),
    .A1(net1671),
    .A2(net2704));
 sg13g2_a21oi_1 _11110_ (.A1(net1671),
    .A2(_03746_),
    .Y(_00610_),
    .B1(_03747_));
 sg13g2_nand2_1 _11111_ (.Y(_03748_),
    .A(\am_sdr0.cic2.integ3[7] ),
    .B(\am_sdr0.cic2.integ2[10] ));
 sg13g2_xnor2_1 _11112_ (.Y(_03749_),
    .A(\am_sdr0.cic2.integ3[7] ),
    .B(\am_sdr0.cic2.integ2[10] ));
 sg13g2_inv_1 _11113_ (.Y(_03750_),
    .A(_03749_));
 sg13g2_o21ai_1 _11114_ (.B1(_03750_),
    .Y(_03751_),
    .A1(_03740_),
    .A2(_03745_));
 sg13g2_or3_1 _11115_ (.A(_03740_),
    .B(_03745_),
    .C(_03750_),
    .X(_03752_));
 sg13g2_nand2_1 _11116_ (.Y(_03753_),
    .A(_03751_),
    .B(_03752_));
 sg13g2_o21ai_1 _11117_ (.B1(net1970),
    .Y(_03754_),
    .A1(net1675),
    .A2(net2620));
 sg13g2_a21oi_1 _11118_ (.A1(net1675),
    .A2(_03753_),
    .Y(_00611_),
    .B1(_03754_));
 sg13g2_xor2_1 _11119_ (.B(\am_sdr0.cic2.integ2[11] ),
    .A(\am_sdr0.cic2.integ3[8] ),
    .X(_03755_));
 sg13g2_inv_1 _11120_ (.Y(_03756_),
    .A(_03755_));
 sg13g2_and3_1 _11121_ (.X(_03757_),
    .A(_03748_),
    .B(_03751_),
    .C(_03756_));
 sg13g2_a21oi_1 _11122_ (.A1(_03748_),
    .A2(_03751_),
    .Y(_03758_),
    .B1(_03756_));
 sg13g2_or2_1 _11123_ (.X(_03759_),
    .B(_03758_),
    .A(_03757_));
 sg13g2_o21ai_1 _11124_ (.B1(net1964),
    .Y(_03760_),
    .A1(net1673),
    .A2(net2338));
 sg13g2_a21oi_1 _11125_ (.A1(net1673),
    .A2(_03759_),
    .Y(_00612_),
    .B1(_03760_));
 sg13g2_nor2_1 _11126_ (.A(\am_sdr0.cic2.integ3[9] ),
    .B(\am_sdr0.cic2.integ2[12] ),
    .Y(_03761_));
 sg13g2_or2_1 _11127_ (.X(_03762_),
    .B(\am_sdr0.cic2.integ2[12] ),
    .A(\am_sdr0.cic2.integ3[9] ));
 sg13g2_a21oi_1 _11128_ (.A1(net2949),
    .A2(\am_sdr0.cic2.integ2[11] ),
    .Y(_03763_),
    .B1(_03758_));
 sg13g2_and2_1 _11129_ (.A(\am_sdr0.cic2.integ3[9] ),
    .B(\am_sdr0.cic2.integ2[12] ),
    .X(_03764_));
 sg13g2_nor2_1 _11130_ (.A(_03761_),
    .B(_03764_),
    .Y(_03765_));
 sg13g2_xor2_1 _11131_ (.B(_03765_),
    .A(_03763_),
    .X(_03766_));
 sg13g2_o21ai_1 _11132_ (.B1(net1964),
    .Y(_03767_),
    .A1(net1673),
    .A2(net2658));
 sg13g2_a21oi_1 _11133_ (.A1(net1673),
    .A2(_03766_),
    .Y(_00613_),
    .B1(_03767_));
 sg13g2_nand2_1 _11134_ (.Y(_03768_),
    .A(net3008),
    .B(\am_sdr0.cic2.integ2[13] ));
 sg13g2_xnor2_1 _11135_ (.Y(_03769_),
    .A(\am_sdr0.cic2.integ3[10] ),
    .B(\am_sdr0.cic2.integ2[13] ));
 sg13g2_a21oi_1 _11136_ (.A1(\am_sdr0.cic2.integ3[8] ),
    .A2(\am_sdr0.cic2.integ2[11] ),
    .Y(_03770_),
    .B1(_03764_));
 sg13g2_nor2_1 _11137_ (.A(_03761_),
    .B(_03770_),
    .Y(_03771_));
 sg13g2_a21oi_1 _11138_ (.A1(_03758_),
    .A2(_03762_),
    .Y(_03772_),
    .B1(_03771_));
 sg13g2_xnor2_1 _11139_ (.Y(_03773_),
    .A(_03769_),
    .B(_03772_));
 sg13g2_o21ai_1 _11140_ (.B1(net1964),
    .Y(_03774_),
    .A1(net1673),
    .A2(net2519));
 sg13g2_a21oi_1 _11141_ (.A1(net1673),
    .A2(_03773_),
    .Y(_00614_),
    .B1(_03774_));
 sg13g2_nor2_1 _11142_ (.A(\am_sdr0.cic2.integ3[11] ),
    .B(\am_sdr0.cic2.integ2[14] ),
    .Y(_03775_));
 sg13g2_xnor2_1 _11143_ (.Y(_03776_),
    .A(\am_sdr0.cic2.integ3[11] ),
    .B(\am_sdr0.cic2.integ2[14] ));
 sg13g2_o21ai_1 _11144_ (.B1(_03768_),
    .Y(_03777_),
    .A1(_03769_),
    .A2(_03772_));
 sg13g2_xor2_1 _11145_ (.B(_03777_),
    .A(_03776_),
    .X(_03778_));
 sg13g2_o21ai_1 _11146_ (.B1(net1964),
    .Y(_03779_),
    .A1(net1673),
    .A2(net2274));
 sg13g2_a21oi_1 _11147_ (.A1(net1673),
    .A2(_03778_),
    .Y(_00615_),
    .B1(_03779_));
 sg13g2_xor2_1 _11148_ (.B(\am_sdr0.cic2.integ2[15] ),
    .A(\am_sdr0.cic2.integ3[12] ),
    .X(_03780_));
 sg13g2_inv_1 _11149_ (.Y(_03781_),
    .A(_03780_));
 sg13g2_nor2_1 _11150_ (.A(_03769_),
    .B(_03776_),
    .Y(_03782_));
 sg13g2_a22oi_1 _11151_ (.Y(_03783_),
    .B1(\am_sdr0.cic2.integ2[13] ),
    .B2(\am_sdr0.cic2.integ3[10] ),
    .A2(\am_sdr0.cic2.integ2[14] ),
    .A1(\am_sdr0.cic2.integ3[11] ));
 sg13g2_nor2_1 _11152_ (.A(_03775_),
    .B(_03783_),
    .Y(_03784_));
 sg13g2_a21oi_2 _11153_ (.B1(_03784_),
    .Y(_03785_),
    .A2(_03782_),
    .A1(_03771_));
 sg13g2_nand3_1 _11154_ (.B(_03765_),
    .C(_03782_),
    .A(_03755_),
    .Y(_03786_));
 sg13g2_a21o_2 _11155_ (.A2(_03751_),
    .A1(_03748_),
    .B1(_03786_),
    .X(_03787_));
 sg13g2_nand2_1 _11156_ (.Y(_03788_),
    .A(_03785_),
    .B(_03787_));
 sg13g2_a21oi_1 _11157_ (.A1(_03785_),
    .A2(_03787_),
    .Y(_03789_),
    .B1(_03781_));
 sg13g2_xnor2_1 _11158_ (.Y(_03790_),
    .A(_03780_),
    .B(_03788_));
 sg13g2_o21ai_1 _11159_ (.B1(net1973),
    .Y(_03791_),
    .A1(net1680),
    .A2(net2996));
 sg13g2_a21oi_1 _11160_ (.A1(net1680),
    .A2(_03790_),
    .Y(_00616_),
    .B1(_03791_));
 sg13g2_nor2_1 _11161_ (.A(\am_sdr0.cic2.integ3[13] ),
    .B(\am_sdr0.cic2.integ2[16] ),
    .Y(_03792_));
 sg13g2_xor2_1 _11162_ (.B(\am_sdr0.cic2.integ2[16] ),
    .A(\am_sdr0.cic2.integ3[13] ),
    .X(_03793_));
 sg13g2_a21oi_1 _11163_ (.A1(\am_sdr0.cic2.integ3[12] ),
    .A2(\am_sdr0.cic2.integ2[15] ),
    .Y(_03794_),
    .B1(_03789_));
 sg13g2_xor2_1 _11164_ (.B(_03794_),
    .A(_03793_),
    .X(_03795_));
 sg13g2_o21ai_1 _11165_ (.B1(net1972),
    .Y(_03796_),
    .A1(net1680),
    .A2(net2987));
 sg13g2_a21oi_1 _11166_ (.A1(net1680),
    .A2(_03795_),
    .Y(_00617_),
    .B1(_03796_));
 sg13g2_nand2_1 _11167_ (.Y(_03797_),
    .A(net2912),
    .B(\am_sdr0.cic2.integ2[17] ));
 sg13g2_xnor2_1 _11168_ (.Y(_03798_),
    .A(\am_sdr0.cic2.integ3[14] ),
    .B(\am_sdr0.cic2.integ2[17] ));
 sg13g2_a22oi_1 _11169_ (.Y(_03799_),
    .B1(\am_sdr0.cic2.integ2[15] ),
    .B2(\am_sdr0.cic2.integ3[12] ),
    .A2(\am_sdr0.cic2.integ2[16] ),
    .A1(\am_sdr0.cic2.integ3[13] ));
 sg13g2_nor2_1 _11170_ (.A(_03792_),
    .B(_03799_),
    .Y(_03800_));
 sg13g2_a21oi_1 _11171_ (.A1(_03789_),
    .A2(_03793_),
    .Y(_03801_),
    .B1(_03800_));
 sg13g2_xnor2_1 _11172_ (.Y(_03802_),
    .A(_03798_),
    .B(_03801_));
 sg13g2_o21ai_1 _11173_ (.B1(net1972),
    .Y(_03803_),
    .A1(net1686),
    .A2(net2912));
 sg13g2_a21oi_1 _11174_ (.A1(net1686),
    .A2(_03802_),
    .Y(_00618_),
    .B1(_03803_));
 sg13g2_nor2_1 _11175_ (.A(\am_sdr0.cic2.integ3[15] ),
    .B(\am_sdr0.cic2.integ2[18] ),
    .Y(_03804_));
 sg13g2_xor2_1 _11176_ (.B(\am_sdr0.cic2.integ2[18] ),
    .A(\am_sdr0.cic2.integ3[15] ),
    .X(_03805_));
 sg13g2_o21ai_1 _11177_ (.B1(_03797_),
    .Y(_03806_),
    .A1(_03798_),
    .A2(_03801_));
 sg13g2_xnor2_1 _11178_ (.Y(_03807_),
    .A(_03805_),
    .B(_03806_));
 sg13g2_o21ai_1 _11179_ (.B1(net1973),
    .Y(_03808_),
    .A1(net1679),
    .A2(net3021));
 sg13g2_a21oi_1 _11180_ (.A1(net1679),
    .A2(_03807_),
    .Y(_00619_),
    .B1(_03808_));
 sg13g2_nand2_1 _11181_ (.Y(_03809_),
    .A(\am_sdr0.cic2.integ3[16] ),
    .B(\am_sdr0.cic2.integ2[19] ));
 sg13g2_xnor2_1 _11182_ (.Y(_03810_),
    .A(\am_sdr0.cic2.integ3[16] ),
    .B(\am_sdr0.cic2.integ2[19] ));
 sg13g2_nor2b_1 _11183_ (.A(_03798_),
    .B_N(_03805_),
    .Y(_03811_));
 sg13g2_and3_1 _11184_ (.X(_03812_),
    .A(_03780_),
    .B(_03793_),
    .C(_03811_));
 sg13g2_nor2_1 _11185_ (.A(_03797_),
    .B(_03804_),
    .Y(_03813_));
 sg13g2_a221oi_1 _11186_ (.B2(_03811_),
    .C1(_03813_),
    .B1(_03800_),
    .A1(\am_sdr0.cic2.integ3[15] ),
    .Y(_03814_),
    .A2(\am_sdr0.cic2.integ2[18] ));
 sg13g2_nor2b_1 _11187_ (.A(_03812_),
    .B_N(_03814_),
    .Y(_03815_));
 sg13g2_and2_1 _11188_ (.A(_03785_),
    .B(_03814_),
    .X(_03816_));
 sg13g2_a21o_2 _11189_ (.A2(_03816_),
    .A1(_03787_),
    .B1(_03815_),
    .X(_03817_));
 sg13g2_xnor2_1 _11190_ (.Y(_03818_),
    .A(_03810_),
    .B(_03817_));
 sg13g2_o21ai_1 _11191_ (.B1(net2004),
    .Y(_03819_),
    .A1(net1685),
    .A2(net2908));
 sg13g2_a21oi_1 _11192_ (.A1(net1687),
    .A2(_03818_),
    .Y(_00620_),
    .B1(_03819_));
 sg13g2_nor2_1 _11193_ (.A(\am_sdr0.cic2.integ3[17] ),
    .B(\am_sdr0.cic2.integ2[20] ),
    .Y(_03820_));
 sg13g2_xor2_1 _11194_ (.B(\am_sdr0.cic2.integ2[20] ),
    .A(\am_sdr0.cic2.integ3[17] ),
    .X(_03821_));
 sg13g2_o21ai_1 _11195_ (.B1(_03809_),
    .Y(_03822_),
    .A1(_03810_),
    .A2(_03817_));
 sg13g2_xnor2_1 _11196_ (.Y(_03823_),
    .A(_03821_),
    .B(_03822_));
 sg13g2_o21ai_1 _11197_ (.B1(net2006),
    .Y(_03824_),
    .A1(net1690),
    .A2(net2969));
 sg13g2_a21oi_1 _11198_ (.A1(net1690),
    .A2(_03823_),
    .Y(_00621_),
    .B1(_03824_));
 sg13g2_and2_1 _11199_ (.A(net3302),
    .B(\am_sdr0.cic2.integ2[21] ),
    .X(_03825_));
 sg13g2_xor2_1 _11200_ (.B(\am_sdr0.cic2.integ2[21] ),
    .A(net2958),
    .X(_03826_));
 sg13g2_nand2b_1 _11201_ (.Y(_03827_),
    .B(_03821_),
    .A_N(_03810_));
 sg13g2_nor2_1 _11202_ (.A(_03809_),
    .B(_03820_),
    .Y(_03828_));
 sg13g2_a21oi_1 _11203_ (.A1(\am_sdr0.cic2.integ3[17] ),
    .A2(\am_sdr0.cic2.integ2[20] ),
    .Y(_03829_),
    .B1(_03828_));
 sg13g2_o21ai_1 _11204_ (.B1(_03829_),
    .Y(_03830_),
    .A1(_03817_),
    .A2(_03827_));
 sg13g2_xnor2_1 _11205_ (.Y(_03831_),
    .A(_03826_),
    .B(_03830_));
 sg13g2_o21ai_1 _11206_ (.B1(net2006),
    .Y(_03832_),
    .A1(net1690),
    .A2(net2958));
 sg13g2_a21oi_1 _11207_ (.A1(net1690),
    .A2(_03831_),
    .Y(_00622_),
    .B1(_03832_));
 sg13g2_a21oi_1 _11208_ (.A1(_03826_),
    .A2(_03830_),
    .Y(_03833_),
    .B1(_03825_));
 sg13g2_xnor2_1 _11209_ (.Y(_03834_),
    .A(net2305),
    .B(net2809));
 sg13g2_xnor2_1 _11210_ (.Y(_03835_),
    .A(_03833_),
    .B(_03834_));
 sg13g2_o21ai_1 _11211_ (.B1(net2006),
    .Y(_03836_),
    .A1(net2305),
    .A2(net1691));
 sg13g2_a21oi_1 _11212_ (.A1(net1691),
    .A2(_03835_),
    .Y(_00623_),
    .B1(_03836_));
 sg13g2_nand2_1 _11213_ (.Y(_03837_),
    .A(net2588),
    .B(net2407));
 sg13g2_o21ai_1 _11214_ (.B1(net1904),
    .Y(_03838_),
    .A1(net2588),
    .A2(net2407));
 sg13g2_nor2b_1 _11215_ (.A(_03838_),
    .B_N(_03837_),
    .Y(_00625_));
 sg13g2_nand2_1 _11216_ (.Y(_03839_),
    .A(net2976),
    .B(net1389));
 sg13g2_xnor2_1 _11217_ (.Y(_03840_),
    .A(net2976),
    .B(net1389));
 sg13g2_o21ai_1 _11218_ (.B1(net1905),
    .Y(_03841_),
    .A1(_03837_),
    .A2(_03840_));
 sg13g2_a21oi_1 _11219_ (.A1(_03837_),
    .A2(_03840_),
    .Y(_00626_),
    .B1(_03841_));
 sg13g2_and2_1 _11220_ (.A(\am_sdr0.cic1.integ2[5] ),
    .B(net2081),
    .X(_03842_));
 sg13g2_xor2_1 _11221_ (.B(net2081),
    .A(net3169),
    .X(_03843_));
 sg13g2_o21ai_1 _11222_ (.B1(_03839_),
    .Y(_03844_),
    .A1(_03837_),
    .A2(_03840_));
 sg13g2_nor2_1 _11223_ (.A(_03843_),
    .B(_03844_),
    .Y(_03845_));
 sg13g2_a21oi_1 _11224_ (.A1(_03843_),
    .A2(_03844_),
    .Y(_03846_),
    .B1(net1876));
 sg13g2_nor2b_1 _11225_ (.A(_03845_),
    .B_N(_03846_),
    .Y(_00627_));
 sg13g2_nand2_1 _11226_ (.Y(_03847_),
    .A(net3313),
    .B(\am_sdr0.cic1.integ3[3] ));
 sg13g2_xnor2_1 _11227_ (.Y(_03848_),
    .A(net3130),
    .B(net2070));
 sg13g2_a21oi_1 _11228_ (.A1(_03843_),
    .A2(_03844_),
    .Y(_03849_),
    .B1(_03842_));
 sg13g2_o21ai_1 _11229_ (.B1(net1903),
    .Y(_03850_),
    .A1(_03848_),
    .A2(_03849_));
 sg13g2_a21oi_1 _11230_ (.A1(_03848_),
    .A2(_03849_),
    .Y(_00628_),
    .B1(_03850_));
 sg13g2_and2_1 _11231_ (.A(\am_sdr0.cic1.integ2[7] ),
    .B(net2159),
    .X(_03851_));
 sg13g2_xor2_1 _11232_ (.B(\am_sdr0.cic1.integ3[4] ),
    .A(\am_sdr0.cic1.integ2[7] ),
    .X(_03852_));
 sg13g2_o21ai_1 _11233_ (.B1(net3314),
    .Y(_03853_),
    .A1(_03848_),
    .A2(_03849_));
 sg13g2_or2_1 _11234_ (.X(_03854_),
    .B(_03853_),
    .A(_03852_));
 sg13g2_a21oi_1 _11235_ (.A1(_03852_),
    .A2(_03853_),
    .Y(_03855_),
    .B1(net1876));
 sg13g2_and2_1 _11236_ (.A(_03854_),
    .B(_03855_),
    .X(_00629_));
 sg13g2_a21oi_1 _11237_ (.A1(_03852_),
    .A2(_03853_),
    .Y(_03856_),
    .B1(_03851_));
 sg13g2_nor2_1 _11238_ (.A(\am_sdr0.cic1.integ2[8] ),
    .B(net3252),
    .Y(_03857_));
 sg13g2_xnor2_1 _11239_ (.Y(_03858_),
    .A(net3105),
    .B(net2085));
 sg13g2_o21ai_1 _11240_ (.B1(net1903),
    .Y(_03859_),
    .A1(_03856_),
    .A2(_03858_));
 sg13g2_a21oi_1 _11241_ (.A1(_03856_),
    .A2(_03858_),
    .Y(_00630_),
    .B1(_03859_));
 sg13g2_and2_1 _11242_ (.A(net3243),
    .B(net1334),
    .X(_03860_));
 sg13g2_xnor2_1 _11243_ (.Y(_03861_),
    .A(\am_sdr0.cic1.integ2[9] ),
    .B(net1334));
 sg13g2_a221oi_1 _11244_ (.B2(_03853_),
    .C1(_03851_),
    .B1(_03852_),
    .A1(\am_sdr0.cic1.integ2[8] ),
    .Y(_03862_),
    .A2(\am_sdr0.cic1.integ3[5] ));
 sg13g2_o21ai_1 _11245_ (.B1(_03861_),
    .Y(_03863_),
    .A1(_03857_),
    .A2(_03862_));
 sg13g2_nor3_2 _11246_ (.A(_03857_),
    .B(_03861_),
    .C(_03862_),
    .Y(_03864_));
 sg13g2_nand2_1 _11247_ (.Y(_03865_),
    .A(net1903),
    .B(_03863_));
 sg13g2_nor2_1 _11248_ (.A(net3253),
    .B(_03865_),
    .Y(_00631_));
 sg13g2_nand2_1 _11249_ (.Y(_03866_),
    .A(\am_sdr0.cic1.integ2[10] ),
    .B(\am_sdr0.cic1.integ3[7] ));
 sg13g2_xnor2_1 _11250_ (.Y(_03867_),
    .A(\am_sdr0.cic1.integ2[10] ),
    .B(net1441));
 sg13g2_inv_1 _11251_ (.Y(_03868_),
    .A(_03867_));
 sg13g2_nor3_1 _11252_ (.A(_03860_),
    .B(_03864_),
    .C(_03868_),
    .Y(_03869_));
 sg13g2_o21ai_1 _11253_ (.B1(_03868_),
    .Y(_03870_),
    .A1(_03860_),
    .A2(_03864_));
 sg13g2_nand2_1 _11254_ (.Y(_03871_),
    .A(net1898),
    .B(_03870_));
 sg13g2_nor2_1 _11255_ (.A(_03869_),
    .B(_03871_),
    .Y(_00632_));
 sg13g2_nand2_1 _11256_ (.Y(_03872_),
    .A(_03866_),
    .B(_03870_));
 sg13g2_nand2_1 _11257_ (.Y(_03873_),
    .A(net3227),
    .B(net1476));
 sg13g2_xor2_1 _11258_ (.B(net1476),
    .A(net3251),
    .X(_03874_));
 sg13g2_inv_1 _11259_ (.Y(_03875_),
    .A(_03874_));
 sg13g2_nand2_1 _11260_ (.Y(_03876_),
    .A(_03872_),
    .B(_03874_));
 sg13g2_o21ai_1 _11261_ (.B1(net1899),
    .Y(_03877_),
    .A1(_03872_),
    .A2(_03874_));
 sg13g2_nor2b_1 _11262_ (.A(_03877_),
    .B_N(_03876_),
    .Y(_00633_));
 sg13g2_nor2_1 _11263_ (.A(\am_sdr0.cic1.integ2[12] ),
    .B(net1423),
    .Y(_03878_));
 sg13g2_nand2_1 _11264_ (.Y(_03879_),
    .A(\am_sdr0.cic1.integ2[12] ),
    .B(net1423));
 sg13g2_nand2b_1 _11265_ (.Y(_03880_),
    .B(_03879_),
    .A_N(_03878_));
 sg13g2_and2_1 _11266_ (.A(_03873_),
    .B(_03876_),
    .X(_03881_));
 sg13g2_o21ai_1 _11267_ (.B1(net1898),
    .Y(_03882_),
    .A1(_03880_),
    .A2(_03881_));
 sg13g2_a21oi_1 _11268_ (.A1(_03880_),
    .A2(_03881_),
    .Y(_00634_),
    .B1(_03882_));
 sg13g2_nand2_1 _11269_ (.Y(_03883_),
    .A(net3133),
    .B(net1497));
 sg13g2_xnor2_1 _11270_ (.Y(_03884_),
    .A(net3133),
    .B(net1497));
 sg13g2_o21ai_1 _11271_ (.B1(_03879_),
    .Y(_03885_),
    .A1(_03873_),
    .A2(_03878_));
 sg13g2_nor2_1 _11272_ (.A(_03875_),
    .B(_03880_),
    .Y(_03886_));
 sg13g2_a21oi_1 _11273_ (.A1(_03872_),
    .A2(_03886_),
    .Y(_03887_),
    .B1(_03885_));
 sg13g2_or2_1 _11274_ (.X(_03888_),
    .B(_03887_),
    .A(_03884_));
 sg13g2_nand2_1 _11275_ (.Y(_03889_),
    .A(net1899),
    .B(_03888_));
 sg13g2_a21oi_1 _11276_ (.A1(_03884_),
    .A2(_03887_),
    .Y(_00635_),
    .B1(_03889_));
 sg13g2_nor2_1 _11277_ (.A(\am_sdr0.cic1.integ2[14] ),
    .B(\am_sdr0.cic1.integ3[11] ),
    .Y(_03890_));
 sg13g2_xnor2_1 _11278_ (.Y(_03891_),
    .A(net3212),
    .B(net2114));
 sg13g2_nand3_1 _11279_ (.B(_03888_),
    .C(_03891_),
    .A(_03883_),
    .Y(_03892_));
 sg13g2_a21oi_1 _11280_ (.A1(_03883_),
    .A2(_03888_),
    .Y(_03893_),
    .B1(_03891_));
 sg13g2_nand2_1 _11281_ (.Y(_03894_),
    .A(net1899),
    .B(_03892_));
 sg13g2_nor2_1 _11282_ (.A(_03893_),
    .B(_03894_),
    .Y(_00636_));
 sg13g2_nand2_1 _11283_ (.Y(_03895_),
    .A(net3081),
    .B(net2645));
 sg13g2_xnor2_1 _11284_ (.Y(_03896_),
    .A(net3081),
    .B(net2645));
 sg13g2_nor2_1 _11285_ (.A(_03884_),
    .B(_03891_),
    .Y(_03897_));
 sg13g2_nor2_1 _11286_ (.A(_03883_),
    .B(_03890_),
    .Y(_03898_));
 sg13g2_a221oi_1 _11287_ (.B2(_03897_),
    .C1(_03898_),
    .B1(_03885_),
    .A1(\am_sdr0.cic1.integ2[14] ),
    .Y(_03899_),
    .A2(\am_sdr0.cic1.integ3[11] ));
 sg13g2_and2_1 _11288_ (.A(_03886_),
    .B(_03897_),
    .X(_03900_));
 sg13g2_inv_1 _11289_ (.Y(_03901_),
    .A(_03900_));
 sg13g2_a21oi_1 _11290_ (.A1(_03866_),
    .A2(_03870_),
    .Y(_03902_),
    .B1(_03901_));
 sg13g2_nor2b_1 _11291_ (.A(_03902_),
    .B_N(_03899_),
    .Y(_03903_));
 sg13g2_or2_1 _11292_ (.X(_03904_),
    .B(_03903_),
    .A(_03896_));
 sg13g2_nand2_1 _11293_ (.Y(_03905_),
    .A(net1899),
    .B(_03904_));
 sg13g2_a21oi_1 _11294_ (.A1(_03896_),
    .A2(_03903_),
    .Y(_00637_),
    .B1(_03905_));
 sg13g2_nor2_1 _11295_ (.A(\am_sdr0.cic1.integ2[16] ),
    .B(net1398),
    .Y(_03906_));
 sg13g2_nand2_1 _11296_ (.Y(_03907_),
    .A(\am_sdr0.cic1.integ2[16] ),
    .B(net1398));
 sg13g2_nor2b_1 _11297_ (.A(_03906_),
    .B_N(_03907_),
    .Y(_03908_));
 sg13g2_nand2_1 _11298_ (.Y(_03909_),
    .A(_03895_),
    .B(_03904_));
 sg13g2_o21ai_1 _11299_ (.B1(net1897),
    .Y(_03910_),
    .A1(_03908_),
    .A2(_03909_));
 sg13g2_a21oi_1 _11300_ (.A1(_03908_),
    .A2(_03909_),
    .Y(_00638_),
    .B1(_03910_));
 sg13g2_nand2_1 _11301_ (.Y(_03911_),
    .A(\am_sdr0.cic1.integ2[17] ),
    .B(net2354));
 sg13g2_xor2_1 _11302_ (.B(net3309),
    .A(\am_sdr0.cic1.integ2[17] ),
    .X(_03912_));
 sg13g2_xnor2_1 _11303_ (.Y(_03913_),
    .A(\am_sdr0.cic1.integ2[17] ),
    .B(\am_sdr0.cic1.integ3[14] ));
 sg13g2_o21ai_1 _11304_ (.B1(_03907_),
    .Y(_03914_),
    .A1(_03895_),
    .A2(_03906_));
 sg13g2_nand2b_1 _11305_ (.Y(_03915_),
    .B(_03908_),
    .A_N(_03896_));
 sg13g2_nor2_1 _11306_ (.A(_03903_),
    .B(_03915_),
    .Y(_03916_));
 sg13g2_nor3_1 _11307_ (.A(_03912_),
    .B(_03914_),
    .C(_03916_),
    .Y(_03917_));
 sg13g2_o21ai_1 _11308_ (.B1(_03912_),
    .Y(_03918_),
    .A1(_03914_),
    .A2(_03916_));
 sg13g2_nand2_1 _11309_ (.Y(_03919_),
    .A(net1897),
    .B(_03918_));
 sg13g2_nor2_1 _11310_ (.A(_03917_),
    .B(_03919_),
    .Y(_00639_));
 sg13g2_nor2_1 _11311_ (.A(\am_sdr0.cic1.integ2[18] ),
    .B(\am_sdr0.cic1.integ3[15] ),
    .Y(_03920_));
 sg13g2_xnor2_1 _11312_ (.Y(_03921_),
    .A(\am_sdr0.cic1.integ2[18] ),
    .B(net2176));
 sg13g2_and3_1 _11313_ (.X(_03922_),
    .A(_03911_),
    .B(_03918_),
    .C(_03921_));
 sg13g2_a21oi_1 _11314_ (.A1(_03911_),
    .A2(_03918_),
    .Y(_03923_),
    .B1(_03921_));
 sg13g2_nor3_1 _11315_ (.A(net1874),
    .B(_03922_),
    .C(_03923_),
    .Y(_00640_));
 sg13g2_nor2_1 _11316_ (.A(_03911_),
    .B(_03920_),
    .Y(_03924_));
 sg13g2_a21oi_1 _11317_ (.A1(\am_sdr0.cic1.integ2[18] ),
    .A2(\am_sdr0.cic1.integ3[15] ),
    .Y(_03925_),
    .B1(_03924_));
 sg13g2_nor2_1 _11318_ (.A(_03913_),
    .B(_03921_),
    .Y(_03926_));
 sg13g2_nor2_1 _11319_ (.A(_03899_),
    .B(_03915_),
    .Y(_03927_));
 sg13g2_o21ai_1 _11320_ (.B1(_03926_),
    .Y(_03928_),
    .A1(_03914_),
    .A2(_03927_));
 sg13g2_nand2_1 _11321_ (.Y(_03929_),
    .A(_03925_),
    .B(_03928_));
 sg13g2_or4_1 _11322_ (.A(_03901_),
    .B(_03913_),
    .C(_03915_),
    .D(_03921_),
    .X(_03930_));
 sg13g2_a21oi_1 _11323_ (.A1(_03866_),
    .A2(_03870_),
    .Y(_03931_),
    .B1(_03930_));
 sg13g2_nor2_1 _11324_ (.A(_03929_),
    .B(_03931_),
    .Y(_03932_));
 sg13g2_nand2_1 _11325_ (.Y(_03933_),
    .A(net3087),
    .B(net2157));
 sg13g2_xnor2_1 _11326_ (.Y(_03934_),
    .A(net3087),
    .B(net2157));
 sg13g2_inv_1 _11327_ (.Y(_03935_),
    .A(_03934_));
 sg13g2_o21ai_1 _11328_ (.B1(_03935_),
    .Y(_03936_),
    .A1(_03929_),
    .A2(_03931_));
 sg13g2_nand2_1 _11329_ (.Y(_03937_),
    .A(net1897),
    .B(_03936_));
 sg13g2_a21oi_1 _11330_ (.A1(_03932_),
    .A2(_03934_),
    .Y(_00641_),
    .B1(_03937_));
 sg13g2_xor2_1 _11331_ (.B(net2997),
    .A(net3153),
    .X(_03938_));
 sg13g2_nand2_1 _11332_ (.Y(_03939_),
    .A(_03933_),
    .B(_03936_));
 sg13g2_o21ai_1 _11333_ (.B1(net1897),
    .Y(_03940_),
    .A1(_03938_),
    .A2(_03939_));
 sg13g2_a21oi_1 _11334_ (.A1(_03938_),
    .A2(_03939_),
    .Y(_00642_),
    .B1(_03940_));
 sg13g2_a22oi_1 _11335_ (.Y(_03941_),
    .B1(\am_sdr0.cic1.integ2[20] ),
    .B2(net2997),
    .A2(\am_sdr0.cic1.integ3[16] ),
    .A1(\am_sdr0.cic1.integ2[19] ));
 sg13g2_nand2_1 _11336_ (.Y(_03942_),
    .A(_03936_),
    .B(_03941_));
 sg13g2_o21ai_1 _11337_ (.B1(_03942_),
    .Y(_03943_),
    .A1(\am_sdr0.cic1.integ2[20] ),
    .A2(net2997));
 sg13g2_xnor2_1 _11338_ (.Y(_03944_),
    .A(\am_sdr0.cic1.integ2[21] ),
    .B(net1406));
 sg13g2_a221oi_1 _11339_ (.B2(_03941_),
    .C1(_03944_),
    .B1(_03936_),
    .A1(_01590_),
    .Y(_03945_),
    .A2(_01591_));
 sg13g2_nand2b_1 _11340_ (.Y(_03946_),
    .B(net1897),
    .A_N(_03945_));
 sg13g2_a21oi_1 _11341_ (.A1(net2998),
    .A2(_03944_),
    .Y(_00643_),
    .B1(_03946_));
 sg13g2_a21oi_1 _11342_ (.A1(\am_sdr0.cic1.integ2[21] ),
    .A2(net1406),
    .Y(_03947_),
    .B1(_03945_));
 sg13g2_xnor2_1 _11343_ (.Y(_03948_),
    .A(net2982),
    .B(net1379));
 sg13g2_o21ai_1 _11344_ (.B1(net1897),
    .Y(_03949_),
    .A1(_03947_),
    .A2(_03948_));
 sg13g2_a21oi_1 _11345_ (.A1(_03947_),
    .A2(_03948_),
    .Y(_00644_),
    .B1(_03949_));
 sg13g2_and3_1 _11346_ (.X(_03950_),
    .A(\am_sdr0.cic0.count[0] ),
    .B(\am_sdr0.cic0.count[1] ),
    .C(net1219));
 sg13g2_and2_1 _11347_ (.A(net2033),
    .B(_03950_),
    .X(_03951_));
 sg13g2_and2_1 _11348_ (.A(net1425),
    .B(_03951_),
    .X(_03952_));
 sg13g2_nand2_1 _11349_ (.Y(_03953_),
    .A(net2810),
    .B(_03952_));
 sg13g2_or2_1 _11350_ (.X(_03954_),
    .B(net1410),
    .A(net1252));
 sg13g2_nor3_1 _11351_ (.A(net1885),
    .B(_03953_),
    .C(_03954_),
    .Y(_00839_));
 sg13g2_mux2_1 _11352_ (.A0(\am_sdr0.cic0.integ_sample[0] ),
    .A1(net2523),
    .S(net1543),
    .X(_00645_));
 sg13g2_nand2_1 _11353_ (.Y(_03955_),
    .A(net2290),
    .B(net1543));
 sg13g2_o21ai_1 _11354_ (.B1(_03955_),
    .Y(_00646_),
    .A1(_01302_),
    .A2(net1545));
 sg13g2_nand2_1 _11355_ (.Y(_03956_),
    .A(net1499),
    .B(net1543));
 sg13g2_o21ai_1 _11356_ (.B1(_03956_),
    .Y(_00647_),
    .A1(_01301_),
    .A2(net1543));
 sg13g2_nand2_1 _11357_ (.Y(_03957_),
    .A(net1433),
    .B(net1543));
 sg13g2_o21ai_1 _11358_ (.B1(_03957_),
    .Y(_00648_),
    .A1(_01300_),
    .A2(net1543));
 sg13g2_nand2_1 _11359_ (.Y(_03958_),
    .A(net1501),
    .B(net1543));
 sg13g2_o21ai_1 _11360_ (.B1(_03958_),
    .Y(_00649_),
    .A1(_01299_),
    .A2(net1543));
 sg13g2_nand2_1 _11361_ (.Y(_03959_),
    .A(net2052),
    .B(net1544));
 sg13g2_o21ai_1 _11362_ (.B1(_03959_),
    .Y(_00650_),
    .A1(_01298_),
    .A2(net1544));
 sg13g2_nand2_1 _11363_ (.Y(_03960_),
    .A(net1400),
    .B(net1544));
 sg13g2_o21ai_1 _11364_ (.B1(_03960_),
    .Y(_00651_),
    .A1(_01296_),
    .A2(net1544));
 sg13g2_nand2_1 _11365_ (.Y(_03961_),
    .A(net2055),
    .B(net1544));
 sg13g2_o21ai_1 _11366_ (.B1(_03961_),
    .Y(_00652_),
    .A1(_01295_),
    .A2(net1544));
 sg13g2_nand2_1 _11367_ (.Y(_03962_),
    .A(net1437),
    .B(net1544));
 sg13g2_o21ai_1 _11368_ (.B1(_03962_),
    .Y(_00653_),
    .A1(_01294_),
    .A2(net1544));
 sg13g2_nand2_1 _11369_ (.Y(_03963_),
    .A(net1443),
    .B(net1541));
 sg13g2_o21ai_1 _11370_ (.B1(_03963_),
    .Y(_00654_),
    .A1(_01293_),
    .A2(net1542));
 sg13g2_nand2_1 _11371_ (.Y(_03964_),
    .A(net1512),
    .B(net1541));
 sg13g2_o21ai_1 _11372_ (.B1(_03964_),
    .Y(_00655_),
    .A1(_01291_),
    .A2(net1542));
 sg13g2_nand2_1 _11373_ (.Y(_03965_),
    .A(net2240),
    .B(net1541));
 sg13g2_o21ai_1 _11374_ (.B1(_03965_),
    .Y(_00656_),
    .A1(_01290_),
    .A2(net1541));
 sg13g2_nand2_1 _11375_ (.Y(_03966_),
    .A(net2267),
    .B(net1541));
 sg13g2_o21ai_1 _11376_ (.B1(_03966_),
    .Y(_00657_),
    .A1(_01289_),
    .A2(net1541));
 sg13g2_nand2_1 _11377_ (.Y(_03967_),
    .A(net2205),
    .B(net1541));
 sg13g2_o21ai_1 _11378_ (.B1(_03967_),
    .Y(_00658_),
    .A1(_01288_),
    .A2(net1541));
 sg13g2_nand2_1 _11379_ (.Y(_03968_),
    .A(net2109),
    .B(net1542));
 sg13g2_o21ai_1 _11380_ (.B1(_03968_),
    .Y(_00659_),
    .A1(_01287_),
    .A2(net1542));
 sg13g2_mux2_1 _11381_ (.A0(net2867),
    .A1(\am_sdr0.cic0.integ3[15] ),
    .S(net1542),
    .X(_00660_));
 sg13g2_nand2_1 _11382_ (.Y(_03969_),
    .A(net1518),
    .B(net1540));
 sg13g2_o21ai_1 _11383_ (.B1(_03969_),
    .Y(_00661_),
    .A1(_01285_),
    .A2(net1540));
 sg13g2_nor2_1 _11384_ (.A(net2597),
    .B(net1540),
    .Y(_03970_));
 sg13g2_a21oi_1 _11385_ (.A1(_01589_),
    .A2(net1540),
    .Y(_00662_),
    .B1(_03970_));
 sg13g2_nand2_1 _11386_ (.Y(_03971_),
    .A(net1514),
    .B(net1540));
 sg13g2_o21ai_1 _11387_ (.B1(_03971_),
    .Y(_00663_),
    .A1(_01282_),
    .A2(net1540));
 sg13g2_nand2_1 _11388_ (.Y(_03972_),
    .A(net1309),
    .B(net1540));
 sg13g2_o21ai_1 _11389_ (.B1(_03972_),
    .Y(_00664_),
    .A1(_01281_),
    .A2(net1540));
 sg13g2_o21ai_1 _11390_ (.B1(net1963),
    .Y(_03973_),
    .A1(net1791),
    .A2(\am_sdr0.cic1.x_out[8] ));
 sg13g2_a21oi_1 _11391_ (.A1(net1791),
    .A2(_01338_),
    .Y(_00665_),
    .B1(_03973_));
 sg13g2_o21ai_1 _11392_ (.B1(net1963),
    .Y(_03974_),
    .A1(net1792),
    .A2(\am_sdr0.cic1.x_out[9] ));
 sg13g2_a21oi_1 _11393_ (.A1(net1792),
    .A2(_01337_),
    .Y(_00666_),
    .B1(_03974_));
 sg13g2_o21ai_1 _11394_ (.B1(net1961),
    .Y(_03975_),
    .A1(net1791),
    .A2(\am_sdr0.cic1.x_out[10] ));
 sg13g2_a21oi_1 _11395_ (.A1(net1792),
    .A2(_01336_),
    .Y(_00667_),
    .B1(_03975_));
 sg13g2_o21ai_1 _11396_ (.B1(net1961),
    .Y(_03976_),
    .A1(net1789),
    .A2(\am_sdr0.cic1.x_out[11] ));
 sg13g2_a21oi_1 _11397_ (.A1(net1789),
    .A2(_01335_),
    .Y(_00668_),
    .B1(_03976_));
 sg13g2_o21ai_1 _11398_ (.B1(net1961),
    .Y(_03977_),
    .A1(net1790),
    .A2(\am_sdr0.cic1.x_out[12] ));
 sg13g2_a21oi_1 _11399_ (.A1(net1789),
    .A2(_01334_),
    .Y(_00669_),
    .B1(_03977_));
 sg13g2_o21ai_1 _11400_ (.B1(net1961),
    .Y(_03978_),
    .A1(net1789),
    .A2(\am_sdr0.cic1.x_out[13] ));
 sg13g2_a21oi_1 _11401_ (.A1(net1789),
    .A2(_01333_),
    .Y(_00670_),
    .B1(_03978_));
 sg13g2_o21ai_1 _11402_ (.B1(net1961),
    .Y(_03979_),
    .A1(net1789),
    .A2(\am_sdr0.cic1.x_out[14] ));
 sg13g2_a21oi_1 _11403_ (.A1(net1789),
    .A2(_01332_),
    .Y(_00671_),
    .B1(_03979_));
 sg13g2_o21ai_1 _11404_ (.B1(net1961),
    .Y(_03980_),
    .A1(net1789),
    .A2(\am_sdr0.cic1.x_out[15] ));
 sg13g2_a21oi_1 _11405_ (.A1(net1790),
    .A2(_01331_),
    .Y(_00672_),
    .B1(_03980_));
 sg13g2_nand2b_1 _11406_ (.Y(_03981_),
    .B(net2035),
    .A_N(net2630));
 sg13g2_a21oi_1 _11407_ (.A1(_01382_),
    .A2(net2630),
    .Y(_03982_),
    .B1(net1637));
 sg13g2_nor2_1 _11408_ (.A(net1640),
    .B(net1888),
    .Y(_00781_));
 sg13g2_a221oi_1 _11409_ (.B2(_03982_),
    .C1(net1878),
    .B1(_03981_),
    .A1(net1637),
    .Y(_00673_),
    .A2(_01360_));
 sg13g2_nor2b_1 _11410_ (.A(net2931),
    .B_N(\am_sdr0.cic1.integ_sample[1] ),
    .Y(_03983_));
 sg13g2_xnor2_1 _11411_ (.Y(_03984_),
    .A(net2931),
    .B(net2359));
 sg13g2_xnor2_1 _11412_ (.Y(_03985_),
    .A(_03981_),
    .B(_03984_));
 sg13g2_o21ai_1 _11413_ (.B1(net1919),
    .Y(_03986_),
    .A1(net1776),
    .A2(net2468));
 sg13g2_a21oi_1 _11414_ (.A1(net1776),
    .A2(_03985_),
    .Y(_00674_),
    .B1(_03986_));
 sg13g2_nand2b_1 _11415_ (.Y(_03987_),
    .B(net3301),
    .A_N(\am_sdr0.cic1.comb1_in_del[2] ));
 sg13g2_xor2_1 _11416_ (.B(net2561),
    .A(\am_sdr0.cic1.comb1_in_del[2] ),
    .X(_03988_));
 sg13g2_a21oi_1 _11417_ (.A1(_03981_),
    .A2(_03984_),
    .Y(_03989_),
    .B1(_03983_));
 sg13g2_xnor2_1 _11418_ (.Y(_03990_),
    .A(_03988_),
    .B(_03989_));
 sg13g2_o21ai_1 _11419_ (.B1(net1917),
    .Y(_03991_),
    .A1(net1774),
    .A2(net2492));
 sg13g2_a21oi_1 _11420_ (.A1(net1776),
    .A2(net2932),
    .Y(_00675_),
    .B1(_03991_));
 sg13g2_nor2_1 _11421_ (.A(\am_sdr0.cic1.comb1_in_del[3] ),
    .B(_01379_),
    .Y(_03992_));
 sg13g2_nand2_1 _11422_ (.Y(_03993_),
    .A(\am_sdr0.cic1.comb1_in_del[3] ),
    .B(_01379_));
 sg13g2_nor2b_1 _11423_ (.A(_03992_),
    .B_N(_03993_),
    .Y(_03994_));
 sg13g2_o21ai_1 _11424_ (.B1(_03987_),
    .Y(_03995_),
    .A1(_03988_),
    .A2(_03989_));
 sg13g2_xnor2_1 _11425_ (.Y(_03996_),
    .A(_03994_),
    .B(_03995_));
 sg13g2_o21ai_1 _11426_ (.B1(net1918),
    .Y(_03997_),
    .A1(net1774),
    .A2(net2263));
 sg13g2_a21oi_1 _11427_ (.A1(net1774),
    .A2(_03996_),
    .Y(_00676_),
    .B1(_03997_));
 sg13g2_nor2_1 _11428_ (.A(net2692),
    .B(_01378_),
    .Y(_03998_));
 sg13g2_xor2_1 _11429_ (.B(\am_sdr0.cic1.integ_sample[4] ),
    .A(net2774),
    .X(_03999_));
 sg13g2_a21oi_2 _11430_ (.B1(_03992_),
    .Y(_04000_),
    .A2(_03995_),
    .A1(_03993_));
 sg13g2_nor2_1 _11431_ (.A(_03999_),
    .B(_04000_),
    .Y(_04001_));
 sg13g2_xnor2_1 _11432_ (.Y(_04002_),
    .A(net2775),
    .B(_04000_));
 sg13g2_o21ai_1 _11433_ (.B1(net1917),
    .Y(_04003_),
    .A1(net1774),
    .A2(net2670));
 sg13g2_a21oi_1 _11434_ (.A1(net1774),
    .A2(_04002_),
    .Y(_00677_),
    .B1(_04003_));
 sg13g2_nand2_1 _11435_ (.Y(_04004_),
    .A(\am_sdr0.cic1.comb1_in_del[5] ),
    .B(_01377_));
 sg13g2_xor2_1 _11436_ (.B(net2877),
    .A(\am_sdr0.cic1.comb1_in_del[5] ),
    .X(_04005_));
 sg13g2_nor2_1 _11437_ (.A(_03998_),
    .B(_04001_),
    .Y(_04006_));
 sg13g2_xnor2_1 _11438_ (.Y(_04007_),
    .A(_04005_),
    .B(_04006_));
 sg13g2_o21ai_1 _11439_ (.B1(net1917),
    .Y(_04008_),
    .A1(net1773),
    .A2(net3012));
 sg13g2_a21oi_1 _11440_ (.A1(net1773),
    .A2(_04007_),
    .Y(_00678_),
    .B1(_04008_));
 sg13g2_nor2_1 _11441_ (.A(\am_sdr0.cic1.comb1_in_del[6] ),
    .B(_01375_),
    .Y(_04009_));
 sg13g2_xor2_1 _11442_ (.B(net2965),
    .A(\am_sdr0.cic1.comb1_in_del[6] ),
    .X(_04010_));
 sg13g2_inv_1 _11443_ (.Y(_04011_),
    .A(_04010_));
 sg13g2_a21oi_1 _11444_ (.A1(_01376_),
    .A2(\am_sdr0.cic1.integ_sample[5] ),
    .Y(_04012_),
    .B1(_03998_));
 sg13g2_o21ai_1 _11445_ (.B1(_04012_),
    .Y(_04013_),
    .A1(_03999_),
    .A2(_04000_));
 sg13g2_and3_1 _11446_ (.X(_04014_),
    .A(_04004_),
    .B(_04011_),
    .C(_04013_));
 sg13g2_a21oi_1 _11447_ (.A1(_04004_),
    .A2(_04013_),
    .Y(_04015_),
    .B1(_04011_));
 sg13g2_or2_1 _11448_ (.X(_04016_),
    .B(_04015_),
    .A(_04014_));
 sg13g2_o21ai_1 _11449_ (.B1(net1917),
    .Y(_04017_),
    .A1(net1772),
    .A2(net2732));
 sg13g2_a21oi_1 _11450_ (.A1(net1773),
    .A2(_04016_),
    .Y(_00679_),
    .B1(_04017_));
 sg13g2_nand2b_1 _11451_ (.Y(_04018_),
    .B(\am_sdr0.cic1.integ_sample[7] ),
    .A_N(\am_sdr0.cic1.comb1_in_del[7] ));
 sg13g2_xor2_1 _11452_ (.B(\am_sdr0.cic1.integ_sample[7] ),
    .A(\am_sdr0.cic1.comb1_in_del[7] ),
    .X(_04019_));
 sg13g2_inv_1 _11453_ (.Y(_04020_),
    .A(_04019_));
 sg13g2_o21ai_1 _11454_ (.B1(_04020_),
    .Y(_04021_),
    .A1(_04009_),
    .A2(_04014_));
 sg13g2_or3_1 _11455_ (.A(_04009_),
    .B(_04014_),
    .C(_04020_),
    .X(_04022_));
 sg13g2_nand2_1 _11456_ (.Y(_04023_),
    .A(_04021_),
    .B(_04022_));
 sg13g2_o21ai_1 _11457_ (.B1(net1909),
    .Y(_04024_),
    .A1(net1778),
    .A2(net2442));
 sg13g2_a21oi_1 _11458_ (.A1(net1772),
    .A2(_04023_),
    .Y(_00680_),
    .B1(_04024_));
 sg13g2_nand2_1 _11459_ (.Y(_04025_),
    .A(_04018_),
    .B(_04021_));
 sg13g2_nor2_1 _11460_ (.A(net2700),
    .B(_01373_),
    .Y(_04026_));
 sg13g2_xnor2_1 _11461_ (.Y(_04027_),
    .A(\am_sdr0.cic1.comb1_in_del[8] ),
    .B(net2807));
 sg13g2_inv_1 _11462_ (.Y(_04028_),
    .A(_04027_));
 sg13g2_xnor2_1 _11463_ (.Y(_04029_),
    .A(_04025_),
    .B(net2808));
 sg13g2_o21ai_1 _11464_ (.B1(net1910),
    .Y(_04030_),
    .A1(net1778),
    .A2(net2485));
 sg13g2_a21oi_1 _11465_ (.A1(net1778),
    .A2(_04029_),
    .Y(_00681_),
    .B1(_04030_));
 sg13g2_xor2_1 _11466_ (.B(net2903),
    .A(\am_sdr0.cic1.comb1_in_del[9] ),
    .X(_04031_));
 sg13g2_a21oi_1 _11467_ (.A1(_04025_),
    .A2(_04027_),
    .Y(_04032_),
    .B1(_04026_));
 sg13g2_xnor2_1 _11468_ (.Y(_04033_),
    .A(_04031_),
    .B(_04032_));
 sg13g2_o21ai_1 _11469_ (.B1(net1910),
    .Y(_04034_),
    .A1(net1778),
    .A2(net2950));
 sg13g2_a21oi_1 _11470_ (.A1(net1773),
    .A2(_04033_),
    .Y(_00682_),
    .B1(_04034_));
 sg13g2_nand2b_1 _11471_ (.Y(_04035_),
    .B(\am_sdr0.cic1.integ_sample[10] ),
    .A_N(\am_sdr0.cic1.comb1_in_del[10] ));
 sg13g2_xor2_1 _11472_ (.B(\am_sdr0.cic1.integ_sample[10] ),
    .A(net2920),
    .X(_04036_));
 sg13g2_a21oi_1 _11473_ (.A1(_01371_),
    .A2(\am_sdr0.cic1.integ_sample[9] ),
    .Y(_04037_),
    .B1(_04026_));
 sg13g2_a21oi_1 _11474_ (.A1(\am_sdr0.cic1.comb1_in_del[9] ),
    .A2(_01372_),
    .Y(_04038_),
    .B1(_04037_));
 sg13g2_nor2_1 _11475_ (.A(_04028_),
    .B(_04031_),
    .Y(_04039_));
 sg13g2_a21oi_1 _11476_ (.A1(_04025_),
    .A2(_04039_),
    .Y(_04040_),
    .B1(_04038_));
 sg13g2_xnor2_1 _11477_ (.Y(_04041_),
    .A(_04036_),
    .B(_04040_));
 sg13g2_o21ai_1 _11478_ (.B1(net1909),
    .Y(_04042_),
    .A1(net1770),
    .A2(net2329));
 sg13g2_a21oi_1 _11479_ (.A1(net1764),
    .A2(_04041_),
    .Y(_00683_),
    .B1(_04042_));
 sg13g2_nor2b_1 _11480_ (.A(\am_sdr0.cic1.integ_sample[11] ),
    .B_N(\am_sdr0.cic1.comb1_in_del[11] ),
    .Y(_04043_));
 sg13g2_nand2b_1 _11481_ (.Y(_04044_),
    .B(\am_sdr0.cic1.integ_sample[11] ),
    .A_N(\am_sdr0.cic1.comb1_in_del[11] ));
 sg13g2_nand2b_1 _11482_ (.Y(_04045_),
    .B(_04044_),
    .A_N(_04043_));
 sg13g2_o21ai_1 _11483_ (.B1(_04035_),
    .Y(_04046_),
    .A1(_04036_),
    .A2(_04040_));
 sg13g2_xor2_1 _11484_ (.B(_04046_),
    .A(_04045_),
    .X(_04047_));
 sg13g2_o21ai_1 _11485_ (.B1(net1909),
    .Y(_04048_),
    .A1(net1769),
    .A2(net2863));
 sg13g2_a21oi_1 _11486_ (.A1(net1769),
    .A2(_04047_),
    .Y(_00684_),
    .B1(_04048_));
 sg13g2_xor2_1 _11487_ (.B(\am_sdr0.cic1.integ_sample[12] ),
    .A(\am_sdr0.cic1.comb1_in_del[12] ),
    .X(_04049_));
 sg13g2_nor2_1 _11488_ (.A(_04036_),
    .B(_04045_),
    .Y(_04050_));
 sg13g2_o21ai_1 _11489_ (.B1(_04044_),
    .Y(_04051_),
    .A1(_04035_),
    .A2(_04043_));
 sg13g2_a21o_1 _11490_ (.A2(_04050_),
    .A1(_04038_),
    .B1(_04051_),
    .X(_04052_));
 sg13g2_inv_1 _11491_ (.Y(_04053_),
    .A(_04052_));
 sg13g2_nand2_1 _11492_ (.Y(_04054_),
    .A(_04039_),
    .B(_04050_));
 sg13g2_a21o_1 _11493_ (.A2(_04021_),
    .A1(_04018_),
    .B1(_04054_),
    .X(_04055_));
 sg13g2_nand2_1 _11494_ (.Y(_04056_),
    .A(_04053_),
    .B(_04055_));
 sg13g2_a21oi_1 _11495_ (.A1(_04053_),
    .A2(_04055_),
    .Y(_04057_),
    .B1(_04049_));
 sg13g2_xor2_1 _11496_ (.B(_04056_),
    .A(_04049_),
    .X(_04058_));
 sg13g2_o21ai_1 _11497_ (.B1(net1909),
    .Y(_04059_),
    .A1(net1769),
    .A2(net2964));
 sg13g2_a21oi_1 _11498_ (.A1(net1769),
    .A2(_04058_),
    .Y(_00685_),
    .B1(_04059_));
 sg13g2_nand2_1 _11499_ (.Y(_04060_),
    .A(\am_sdr0.cic1.comb1_in_del[13] ),
    .B(_01367_));
 sg13g2_xor2_1 _11500_ (.B(\am_sdr0.cic1.integ_sample[13] ),
    .A(\am_sdr0.cic1.comb1_in_del[13] ),
    .X(_04061_));
 sg13g2_a21oi_1 _11501_ (.A1(_01368_),
    .A2(\am_sdr0.cic1.integ_sample[12] ),
    .Y(_04062_),
    .B1(_04057_));
 sg13g2_xnor2_1 _11502_ (.Y(_04063_),
    .A(_04061_),
    .B(_04062_));
 sg13g2_o21ai_1 _11503_ (.B1(net1907),
    .Y(_04064_),
    .A1(net1769),
    .A2(net2327));
 sg13g2_a21oi_1 _11504_ (.A1(net1769),
    .A2(_04063_),
    .Y(_00686_),
    .B1(_04064_));
 sg13g2_nand2b_1 _11505_ (.Y(_04065_),
    .B(\am_sdr0.cic1.integ_sample[14] ),
    .A_N(\am_sdr0.cic1.comb1_in_del[14] ));
 sg13g2_xor2_1 _11506_ (.B(\am_sdr0.cic1.integ_sample[14] ),
    .A(\am_sdr0.cic1.comb1_in_del[14] ),
    .X(_04066_));
 sg13g2_nand3_1 _11507_ (.B(\am_sdr0.cic1.integ_sample[12] ),
    .C(_04060_),
    .A(_01368_),
    .Y(_04067_));
 sg13g2_o21ai_1 _11508_ (.B1(_04067_),
    .Y(_04068_),
    .A1(\am_sdr0.cic1.comb1_in_del[13] ),
    .A2(_01367_));
 sg13g2_a21oi_1 _11509_ (.A1(_04057_),
    .A2(_04060_),
    .Y(_04069_),
    .B1(_04068_));
 sg13g2_xnor2_1 _11510_ (.Y(_04070_),
    .A(_04066_),
    .B(_04069_));
 sg13g2_o21ai_1 _11511_ (.B1(net1907),
    .Y(_04071_),
    .A1(net1767),
    .A2(net2398));
 sg13g2_a21oi_1 _11512_ (.A1(net1767),
    .A2(_04070_),
    .Y(_00687_),
    .B1(_04071_));
 sg13g2_nor2b_1 _11513_ (.A(\am_sdr0.cic1.integ_sample[15] ),
    .B_N(\am_sdr0.cic1.comb1_in_del[15] ),
    .Y(_04072_));
 sg13g2_nand2b_1 _11514_ (.Y(_04073_),
    .B(\am_sdr0.cic1.integ_sample[15] ),
    .A_N(\am_sdr0.cic1.comb1_in_del[15] ));
 sg13g2_nand2b_1 _11515_ (.Y(_04074_),
    .B(_04073_),
    .A_N(_04072_));
 sg13g2_o21ai_1 _11516_ (.B1(_04065_),
    .Y(_04075_),
    .A1(_04066_),
    .A2(_04069_));
 sg13g2_xor2_1 _11517_ (.B(_04075_),
    .A(_04074_),
    .X(_04076_));
 sg13g2_o21ai_1 _11518_ (.B1(net1916),
    .Y(_04077_),
    .A1(net1767),
    .A2(net2973));
 sg13g2_a21oi_1 _11519_ (.A1(net1767),
    .A2(_04076_),
    .Y(_00688_),
    .B1(_04077_));
 sg13g2_nor2_1 _11520_ (.A(\am_sdr0.cic1.comb1_in_del[16] ),
    .B(_01364_),
    .Y(_04078_));
 sg13g2_xnor2_1 _11521_ (.Y(_04079_),
    .A(\am_sdr0.cic1.comb1_in_del[16] ),
    .B(\am_sdr0.cic1.integ_sample[16] ));
 sg13g2_inv_1 _11522_ (.Y(_04080_),
    .A(_04079_));
 sg13g2_nor2_1 _11523_ (.A(_04066_),
    .B(_04074_),
    .Y(_04081_));
 sg13g2_nor4_1 _11524_ (.A(_04049_),
    .B(_04061_),
    .C(_04066_),
    .D(_04074_),
    .Y(_04082_));
 sg13g2_or4_1 _11525_ (.A(_04049_),
    .B(_04061_),
    .C(_04066_),
    .D(_04074_),
    .X(_04083_));
 sg13g2_o21ai_1 _11526_ (.B1(_04073_),
    .Y(_04084_),
    .A1(_04065_),
    .A2(_04072_));
 sg13g2_a221oi_1 _11527_ (.B2(_04052_),
    .C1(_04084_),
    .B1(_04082_),
    .A1(_04068_),
    .Y(_04085_),
    .A2(_04081_));
 sg13g2_o21ai_1 _11528_ (.B1(_04085_),
    .Y(_04086_),
    .A1(_04055_),
    .A2(_04083_));
 sg13g2_xnor2_1 _11529_ (.Y(_04087_),
    .A(_04079_),
    .B(_04086_));
 sg13g2_o21ai_1 _11530_ (.B1(net1907),
    .Y(_04088_),
    .A1(net1766),
    .A2(net2773));
 sg13g2_a21oi_1 _11531_ (.A1(net1766),
    .A2(_04087_),
    .Y(_00689_),
    .B1(_04088_));
 sg13g2_nand2_1 _11532_ (.Y(_04089_),
    .A(\am_sdr0.cic1.comb1_in_del[17] ),
    .B(_01363_));
 sg13g2_nor2_1 _11533_ (.A(\am_sdr0.cic1.comb1_in_del[17] ),
    .B(_01363_),
    .Y(_04090_));
 sg13g2_xor2_1 _11534_ (.B(\am_sdr0.cic1.integ_sample[17] ),
    .A(\am_sdr0.cic1.comb1_in_del[17] ),
    .X(_04091_));
 sg13g2_a21oi_1 _11535_ (.A1(_04079_),
    .A2(_04086_),
    .Y(_04092_),
    .B1(_04078_));
 sg13g2_xnor2_1 _11536_ (.Y(_04093_),
    .A(_04091_),
    .B(_04092_));
 sg13g2_o21ai_1 _11537_ (.B1(net1907),
    .Y(_04094_),
    .A1(net1766),
    .A2(net2816));
 sg13g2_a21oi_1 _11538_ (.A1(net1766),
    .A2(_04093_),
    .Y(_00690_),
    .B1(_04094_));
 sg13g2_nand2b_1 _11539_ (.Y(_04095_),
    .B(\am_sdr0.cic1.integ_sample[18] ),
    .A_N(\am_sdr0.cic1.comb1_in_del[18] ));
 sg13g2_xor2_1 _11540_ (.B(\am_sdr0.cic1.integ_sample[18] ),
    .A(net2663),
    .X(_04096_));
 sg13g2_nor2_1 _11541_ (.A(_04080_),
    .B(_04091_),
    .Y(_04097_));
 sg13g2_a221oi_1 _11542_ (.B2(_04086_),
    .C1(_04090_),
    .B1(_04097_),
    .A1(_04078_),
    .Y(_04098_),
    .A2(_04089_));
 sg13g2_xnor2_1 _11543_ (.Y(_04099_),
    .A(_04096_),
    .B(_04098_));
 sg13g2_o21ai_1 _11544_ (.B1(net1907),
    .Y(_04100_),
    .A1(net1766),
    .A2(net2760));
 sg13g2_a21oi_1 _11545_ (.A1(net1766),
    .A2(_04099_),
    .Y(_00691_),
    .B1(_04100_));
 sg13g2_o21ai_1 _11546_ (.B1(_04095_),
    .Y(_04101_),
    .A1(_04096_),
    .A2(_04098_));
 sg13g2_xnor2_1 _11547_ (.Y(_04102_),
    .A(net2690),
    .B(net2141));
 sg13g2_xnor2_1 _11548_ (.Y(_04103_),
    .A(_04101_),
    .B(_04102_));
 sg13g2_o21ai_1 _11549_ (.B1(net1907),
    .Y(_04104_),
    .A1(net1767),
    .A2(net2119));
 sg13g2_a21oi_1 _11550_ (.A1(net1766),
    .A2(net2691),
    .Y(_00692_),
    .B1(_04104_));
 sg13g2_o21ai_1 _11551_ (.B1(net1920),
    .Y(_04105_),
    .A1(net1637),
    .A2(\am_sdr0.cic1.integ_sample[0] ));
 sg13g2_a21oi_1 _11552_ (.A1(net1637),
    .A2(_01382_),
    .Y(_00693_),
    .B1(_04105_));
 sg13g2_o21ai_1 _11553_ (.B1(net1920),
    .Y(_04106_),
    .A1(net1775),
    .A2(\am_sdr0.cic1.comb1_in_del[1] ));
 sg13g2_a21oi_1 _11554_ (.A1(net1775),
    .A2(_01381_),
    .Y(_00694_),
    .B1(_04106_));
 sg13g2_o21ai_1 _11555_ (.B1(net1918),
    .Y(_04107_),
    .A1(net1775),
    .A2(\am_sdr0.cic1.comb1_in_del[2] ));
 sg13g2_a21oi_1 _11556_ (.A1(net1775),
    .A2(_01380_),
    .Y(_00695_),
    .B1(_04107_));
 sg13g2_o21ai_1 _11557_ (.B1(net1918),
    .Y(_04108_),
    .A1(net1775),
    .A2(\am_sdr0.cic1.comb1_in_del[3] ));
 sg13g2_a21oi_1 _11558_ (.A1(net1775),
    .A2(_01379_),
    .Y(_00696_),
    .B1(_04108_));
 sg13g2_o21ai_1 _11559_ (.B1(net1918),
    .Y(_04109_),
    .A1(net1775),
    .A2(net2692));
 sg13g2_a21oi_1 _11560_ (.A1(net1775),
    .A2(_01378_),
    .Y(_00697_),
    .B1(_04109_));
 sg13g2_o21ai_1 _11561_ (.B1(net1918),
    .Y(_04110_),
    .A1(net1772),
    .A2(\am_sdr0.cic1.comb1_in_del[5] ));
 sg13g2_a21oi_1 _11562_ (.A1(net1772),
    .A2(_01377_),
    .Y(_00698_),
    .B1(_04110_));
 sg13g2_o21ai_1 _11563_ (.B1(net1918),
    .Y(_04111_),
    .A1(net1772),
    .A2(\am_sdr0.cic1.comb1_in_del[6] ));
 sg13g2_a21oi_1 _11564_ (.A1(net1772),
    .A2(_01375_),
    .Y(_00699_),
    .B1(_04111_));
 sg13g2_o21ai_1 _11565_ (.B1(net1910),
    .Y(_04112_),
    .A1(net1772),
    .A2(\am_sdr0.cic1.comb1_in_del[7] ));
 sg13g2_a21oi_1 _11566_ (.A1(net1772),
    .A2(_01374_),
    .Y(_00700_),
    .B1(_04112_));
 sg13g2_o21ai_1 _11567_ (.B1(net1910),
    .Y(_04113_),
    .A1(net1773),
    .A2(net2700));
 sg13g2_a21oi_1 _11568_ (.A1(net1773),
    .A2(_01373_),
    .Y(_00701_),
    .B1(_04113_));
 sg13g2_o21ai_1 _11569_ (.B1(net1910),
    .Y(_04114_),
    .A1(net1765),
    .A2(\am_sdr0.cic1.comb1_in_del[9] ));
 sg13g2_a21oi_1 _11570_ (.A1(net1764),
    .A2(_01372_),
    .Y(_00702_),
    .B1(_04114_));
 sg13g2_o21ai_1 _11571_ (.B1(net1910),
    .Y(_04115_),
    .A1(net1764),
    .A2(net2656));
 sg13g2_a21oi_1 _11572_ (.A1(net1764),
    .A2(_01370_),
    .Y(_00703_),
    .B1(_04115_));
 sg13g2_o21ai_1 _11573_ (.B1(net1910),
    .Y(_04116_),
    .A1(net1764),
    .A2(\am_sdr0.cic1.comb1_in_del[11] ));
 sg13g2_a21oi_1 _11574_ (.A1(net1764),
    .A2(_01369_),
    .Y(_00704_),
    .B1(_04116_));
 sg13g2_o21ai_1 _11575_ (.B1(net1908),
    .Y(_04117_),
    .A1(net1638),
    .A2(\am_sdr0.cic1.integ_sample[12] ));
 sg13g2_a21oi_1 _11576_ (.A1(net1638),
    .A2(_01368_),
    .Y(_00705_),
    .B1(_04117_));
 sg13g2_o21ai_1 _11577_ (.B1(net1908),
    .Y(_04118_),
    .A1(net1764),
    .A2(net2930));
 sg13g2_a21oi_1 _11578_ (.A1(net1764),
    .A2(_01367_),
    .Y(_00706_),
    .B1(_04118_));
 sg13g2_o21ai_1 _11579_ (.B1(net1908),
    .Y(_04119_),
    .A1(net1762),
    .A2(\am_sdr0.cic1.comb1_in_del[14] ));
 sg13g2_a21oi_1 _11580_ (.A1(net1762),
    .A2(_01366_),
    .Y(_00707_),
    .B1(_04119_));
 sg13g2_o21ai_1 _11581_ (.B1(net1908),
    .Y(_04120_),
    .A1(net1762),
    .A2(net2411));
 sg13g2_a21oi_1 _11582_ (.A1(net1762),
    .A2(_01365_),
    .Y(_00708_),
    .B1(_04120_));
 sg13g2_o21ai_1 _11583_ (.B1(net1908),
    .Y(_04121_),
    .A1(net1763),
    .A2(net2753));
 sg13g2_a21oi_1 _11584_ (.A1(net1763),
    .A2(_01364_),
    .Y(_00709_),
    .B1(_04121_));
 sg13g2_o21ai_1 _11585_ (.B1(net1907),
    .Y(_04122_),
    .A1(net1763),
    .A2(net2927));
 sg13g2_a21oi_1 _11586_ (.A1(net1762),
    .A2(_01363_),
    .Y(_00710_),
    .B1(_04122_));
 sg13g2_o21ai_1 _11587_ (.B1(net1908),
    .Y(_04123_),
    .A1(net1763),
    .A2(net2663));
 sg13g2_a21oi_1 _11588_ (.A1(net1762),
    .A2(_01362_),
    .Y(_00711_),
    .B1(_04123_));
 sg13g2_o21ai_1 _11589_ (.B1(net1908),
    .Y(_04124_),
    .A1(net1762),
    .A2(\am_sdr0.cic1.comb1_in_del[19] ));
 sg13g2_a21oi_1 _11590_ (.A1(net1762),
    .A2(_01361_),
    .Y(_00712_),
    .B1(_04124_));
 sg13g2_nand2b_1 _11591_ (.Y(_04125_),
    .B(net2458),
    .A_N(net2388));
 sg13g2_a21oi_1 _11592_ (.A1(_01359_),
    .A2(net2388),
    .Y(_04126_),
    .B1(net1637));
 sg13g2_a221oi_1 _11593_ (.B2(_04126_),
    .C1(net1878),
    .B1(_04125_),
    .A1(net1638),
    .Y(_00713_),
    .A2(_01330_));
 sg13g2_nor2b_1 _11594_ (.A(net2763),
    .B_N(\am_sdr0.cic1.comb1[1] ),
    .Y(_04127_));
 sg13g2_xnor2_1 _11595_ (.Y(_04128_),
    .A(net2763),
    .B(net2468));
 sg13g2_xnor2_1 _11596_ (.Y(_04129_),
    .A(_04125_),
    .B(_04128_));
 sg13g2_o21ai_1 _11597_ (.B1(net1923),
    .Y(_04130_),
    .A1(net1782),
    .A2(net2307));
 sg13g2_a21oi_1 _11598_ (.A1(net1780),
    .A2(_04129_),
    .Y(_00714_),
    .B1(_04130_));
 sg13g2_nand2b_1 _11599_ (.Y(_04131_),
    .B(\am_sdr0.cic1.comb1[2] ),
    .A_N(\am_sdr0.cic1.comb2_in_del[2] ));
 sg13g2_xor2_1 _11600_ (.B(\am_sdr0.cic1.comb1[2] ),
    .A(\am_sdr0.cic1.comb2_in_del[2] ),
    .X(_04132_));
 sg13g2_a21oi_1 _11601_ (.A1(_04125_),
    .A2(_04128_),
    .Y(_04133_),
    .B1(_04127_));
 sg13g2_xnor2_1 _11602_ (.Y(_04134_),
    .A(_04132_),
    .B(_04133_));
 sg13g2_o21ai_1 _11603_ (.B1(net1921),
    .Y(_04135_),
    .A1(net1782),
    .A2(net2901));
 sg13g2_a21oi_1 _11604_ (.A1(net1781),
    .A2(_04134_),
    .Y(_00715_),
    .B1(_04135_));
 sg13g2_nor2_1 _11605_ (.A(net2605),
    .B(_01356_),
    .Y(_04136_));
 sg13g2_nand2_1 _11606_ (.Y(_04137_),
    .A(net2566),
    .B(_01356_));
 sg13g2_nor2b_1 _11607_ (.A(_04136_),
    .B_N(_04137_),
    .Y(_04138_));
 sg13g2_o21ai_1 _11608_ (.B1(_04131_),
    .Y(_04139_),
    .A1(_04132_),
    .A2(_04133_));
 sg13g2_xnor2_1 _11609_ (.Y(_04140_),
    .A(_04138_),
    .B(_04139_));
 sg13g2_o21ai_1 _11610_ (.B1(net1922),
    .Y(_04141_),
    .A1(net1781),
    .A2(net2842));
 sg13g2_a21oi_1 _11611_ (.A1(net1781),
    .A2(_04140_),
    .Y(_00716_),
    .B1(_04141_));
 sg13g2_nor2_1 _11612_ (.A(\am_sdr0.cic1.comb2_in_del[4] ),
    .B(_01355_),
    .Y(_04142_));
 sg13g2_xor2_1 _11613_ (.B(net3297),
    .A(\am_sdr0.cic1.comb2_in_del[4] ),
    .X(_04143_));
 sg13g2_a21oi_2 _11614_ (.B1(_04136_),
    .Y(_04144_),
    .A2(_04139_),
    .A1(_04137_));
 sg13g2_nor2_1 _11615_ (.A(_04143_),
    .B(_04144_),
    .Y(_04145_));
 sg13g2_xnor2_1 _11616_ (.Y(_04146_),
    .A(_04143_),
    .B(_04144_));
 sg13g2_o21ai_1 _11617_ (.B1(net1922),
    .Y(_04147_),
    .A1(net1781),
    .A2(net2370));
 sg13g2_a21oi_1 _11618_ (.A1(net1781),
    .A2(_04146_),
    .Y(_00717_),
    .B1(_04147_));
 sg13g2_nor2_1 _11619_ (.A(_01354_),
    .B(\am_sdr0.cic1.comb1[5] ),
    .Y(_04148_));
 sg13g2_xor2_1 _11620_ (.B(\am_sdr0.cic1.comb1[5] ),
    .A(net2583),
    .X(_04149_));
 sg13g2_nor2_1 _11621_ (.A(_04142_),
    .B(_04145_),
    .Y(_04150_));
 sg13g2_xnor2_1 _11622_ (.Y(_04151_),
    .A(_04149_),
    .B(_04150_));
 sg13g2_o21ai_1 _11623_ (.B1(net1921),
    .Y(_04152_),
    .A1(net1796),
    .A2(net2864));
 sg13g2_a21oi_1 _11624_ (.A1(net1781),
    .A2(_04151_),
    .Y(_00718_),
    .B1(_04152_));
 sg13g2_nand2b_1 _11625_ (.Y(_04153_),
    .B(\am_sdr0.cic1.comb1[6] ),
    .A_N(net2882));
 sg13g2_xnor2_1 _11626_ (.Y(_04154_),
    .A(net2608),
    .B(net3311));
 sg13g2_a21oi_1 _11627_ (.A1(_01354_),
    .A2(\am_sdr0.cic1.comb1[5] ),
    .Y(_04155_),
    .B1(_04142_));
 sg13g2_o21ai_1 _11628_ (.B1(_04155_),
    .Y(_04156_),
    .A1(_04143_),
    .A2(_04144_));
 sg13g2_nor2b_1 _11629_ (.A(_04148_),
    .B_N(_04156_),
    .Y(_04157_));
 sg13g2_nand3b_1 _11630_ (.B(_04154_),
    .C(_04156_),
    .Y(_04158_),
    .A_N(_04148_));
 sg13g2_xnor2_1 _11631_ (.Y(_04159_),
    .A(_04154_),
    .B(_04157_));
 sg13g2_o21ai_1 _11632_ (.B1(net1921),
    .Y(_04160_),
    .A1(net1795),
    .A2(net2392));
 sg13g2_a21oi_1 _11633_ (.A1(net1779),
    .A2(_04159_),
    .Y(_00719_),
    .B1(_04160_));
 sg13g2_nand2b_1 _11634_ (.Y(_04161_),
    .B(\am_sdr0.cic1.comb1[7] ),
    .A_N(\am_sdr0.cic1.comb2_in_del[7] ));
 sg13g2_xor2_1 _11635_ (.B(\am_sdr0.cic1.comb1[7] ),
    .A(\am_sdr0.cic1.comb2_in_del[7] ),
    .X(_04162_));
 sg13g2_a21o_1 _11636_ (.A2(_04158_),
    .A1(_04153_),
    .B1(_04162_),
    .X(_04163_));
 sg13g2_nand3_1 _11637_ (.B(_04158_),
    .C(_04162_),
    .A(net2883),
    .Y(_04164_));
 sg13g2_a21oi_1 _11638_ (.A1(_04163_),
    .A2(_04164_),
    .Y(_04165_),
    .B1(net1637));
 sg13g2_o21ai_1 _11639_ (.B1(net1921),
    .Y(_04166_),
    .A1(net1795),
    .A2(net2494));
 sg13g2_nor2_1 _11640_ (.A(_04165_),
    .B(_04166_),
    .Y(_00720_));
 sg13g2_nand2_1 _11641_ (.Y(_04167_),
    .A(_04161_),
    .B(_04163_));
 sg13g2_nor2_1 _11642_ (.A(\am_sdr0.cic1.comb2_in_del[8] ),
    .B(_01351_),
    .Y(_04168_));
 sg13g2_xnor2_1 _11643_ (.Y(_04169_),
    .A(\am_sdr0.cic1.comb2_in_del[8] ),
    .B(\am_sdr0.cic1.comb1[8] ));
 sg13g2_inv_1 _11644_ (.Y(_04170_),
    .A(_04169_));
 sg13g2_xnor2_1 _11645_ (.Y(_04171_),
    .A(_04167_),
    .B(_04169_));
 sg13g2_o21ai_1 _11646_ (.B1(net1913),
    .Y(_04172_),
    .A1(net1794),
    .A2(net2403));
 sg13g2_a21oi_1 _11647_ (.A1(net1779),
    .A2(_04171_),
    .Y(_00721_),
    .B1(_04172_));
 sg13g2_xor2_1 _11648_ (.B(\am_sdr0.cic1.comb1[9] ),
    .A(net3321),
    .X(_04173_));
 sg13g2_a21oi_1 _11649_ (.A1(_04167_),
    .A2(_04169_),
    .Y(_04174_),
    .B1(_04168_));
 sg13g2_xnor2_1 _11650_ (.Y(_04175_),
    .A(_04173_),
    .B(_04174_));
 sg13g2_o21ai_1 _11651_ (.B1(net1913),
    .Y(_04176_),
    .A1(net1794),
    .A2(net2836));
 sg13g2_a21oi_1 _11652_ (.A1(net1779),
    .A2(_04175_),
    .Y(_00722_),
    .B1(_04176_));
 sg13g2_nand2b_1 _11653_ (.Y(_04177_),
    .B(\am_sdr0.cic1.comb1[10] ),
    .A_N(\am_sdr0.cic1.comb2_in_del[10] ));
 sg13g2_xor2_1 _11654_ (.B(\am_sdr0.cic1.comb1[10] ),
    .A(\am_sdr0.cic1.comb2_in_del[10] ),
    .X(_04178_));
 sg13g2_a21oi_1 _11655_ (.A1(_01349_),
    .A2(\am_sdr0.cic1.comb1[9] ),
    .Y(_04179_),
    .B1(_04168_));
 sg13g2_a21oi_1 _11656_ (.A1(\am_sdr0.cic1.comb2_in_del[9] ),
    .A2(_01350_),
    .Y(_04180_),
    .B1(_04179_));
 sg13g2_nor2_1 _11657_ (.A(_04170_),
    .B(_04173_),
    .Y(_04181_));
 sg13g2_a21oi_1 _11658_ (.A1(_04167_),
    .A2(_04181_),
    .Y(_04182_),
    .B1(_04180_));
 sg13g2_xnor2_1 _11659_ (.Y(_04183_),
    .A(_04178_),
    .B(_04182_));
 sg13g2_o21ai_1 _11660_ (.B1(net1913),
    .Y(_04184_),
    .A1(net1787),
    .A2(net2780));
 sg13g2_a21oi_1 _11661_ (.A1(net1770),
    .A2(_04183_),
    .Y(_00723_),
    .B1(_04184_));
 sg13g2_nor2b_1 _11662_ (.A(\am_sdr0.cic1.comb1[11] ),
    .B_N(\am_sdr0.cic1.comb2_in_del[11] ),
    .Y(_04185_));
 sg13g2_nand2b_1 _11663_ (.Y(_04186_),
    .B(\am_sdr0.cic1.comb1[11] ),
    .A_N(\am_sdr0.cic1.comb2_in_del[11] ));
 sg13g2_nand2b_1 _11664_ (.Y(_04187_),
    .B(_04186_),
    .A_N(_04185_));
 sg13g2_o21ai_1 _11665_ (.B1(_04177_),
    .Y(_04188_),
    .A1(_04178_),
    .A2(_04182_));
 sg13g2_xor2_1 _11666_ (.B(_04188_),
    .A(_04187_),
    .X(_04189_));
 sg13g2_o21ai_1 _11667_ (.B1(net1913),
    .Y(_04190_),
    .A1(net1786),
    .A2(net2571));
 sg13g2_a21oi_1 _11668_ (.A1(net1786),
    .A2(_04189_),
    .Y(_00724_),
    .B1(_04190_));
 sg13g2_nand2b_1 _11669_ (.Y(_04191_),
    .B(\am_sdr0.cic1.comb1[12] ),
    .A_N(\am_sdr0.cic1.comb2_in_del[12] ));
 sg13g2_xor2_1 _11670_ (.B(\am_sdr0.cic1.comb1[12] ),
    .A(net3071),
    .X(_04192_));
 sg13g2_nor2_1 _11671_ (.A(_04178_),
    .B(_04187_),
    .Y(_04193_));
 sg13g2_o21ai_1 _11672_ (.B1(_04186_),
    .Y(_04194_),
    .A1(_04177_),
    .A2(_04185_));
 sg13g2_a21o_1 _11673_ (.A2(_04193_),
    .A1(_04180_),
    .B1(_04194_),
    .X(_04195_));
 sg13g2_nand2_1 _11674_ (.Y(_04196_),
    .A(_04181_),
    .B(_04193_));
 sg13g2_a21oi_2 _11675_ (.B1(_04196_),
    .Y(_04197_),
    .A2(_04163_),
    .A1(_04161_));
 sg13g2_nor2_1 _11676_ (.A(_04195_),
    .B(_04197_),
    .Y(_04198_));
 sg13g2_xnor2_1 _11677_ (.Y(_04199_),
    .A(_04192_),
    .B(_04198_));
 sg13g2_o21ai_1 _11678_ (.B1(net1914),
    .Y(_04200_),
    .A1(net1788),
    .A2(net2718));
 sg13g2_a21oi_1 _11679_ (.A1(net1786),
    .A2(_04199_),
    .Y(_00725_),
    .B1(_04200_));
 sg13g2_nor2b_1 _11680_ (.A(\am_sdr0.cic1.comb1[13] ),
    .B_N(\am_sdr0.cic1.comb2_in_del[13] ),
    .Y(_04201_));
 sg13g2_nand2b_1 _11681_ (.Y(_04202_),
    .B(\am_sdr0.cic1.comb1[13] ),
    .A_N(\am_sdr0.cic1.comb2_in_del[13] ));
 sg13g2_nand2b_1 _11682_ (.Y(_04203_),
    .B(_04202_),
    .A_N(_04201_));
 sg13g2_o21ai_1 _11683_ (.B1(_04191_),
    .Y(_04204_),
    .A1(_04192_),
    .A2(_04198_));
 sg13g2_xor2_1 _11684_ (.B(_04204_),
    .A(_04203_),
    .X(_04205_));
 sg13g2_o21ai_1 _11685_ (.B1(net1914),
    .Y(_04206_),
    .A1(net1787),
    .A2(net2335));
 sg13g2_a21oi_1 _11686_ (.A1(net1786),
    .A2(_04205_),
    .Y(_00726_),
    .B1(_04206_));
 sg13g2_nor2_1 _11687_ (.A(\am_sdr0.cic1.comb2_in_del[14] ),
    .B(_01344_),
    .Y(_04207_));
 sg13g2_nand2_1 _11688_ (.Y(_04208_),
    .A(\am_sdr0.cic1.comb2_in_del[14] ),
    .B(_01344_));
 sg13g2_nand2b_2 _11689_ (.Y(_04209_),
    .B(_04208_),
    .A_N(_04207_));
 sg13g2_o21ai_1 _11690_ (.B1(_04202_),
    .Y(_04210_),
    .A1(_04191_),
    .A2(_04201_));
 sg13g2_inv_1 _11691_ (.Y(_04211_),
    .A(_04210_));
 sg13g2_or2_1 _11692_ (.X(_04212_),
    .B(_04203_),
    .A(_04192_));
 sg13g2_o21ai_1 _11693_ (.B1(_04211_),
    .Y(_04213_),
    .A1(_04198_),
    .A2(_04212_));
 sg13g2_xor2_1 _11694_ (.B(_04213_),
    .A(_04209_),
    .X(_04214_));
 sg13g2_o21ai_1 _11695_ (.B1(net1911),
    .Y(_04215_),
    .A1(net1786),
    .A2(net2500));
 sg13g2_a21oi_1 _11696_ (.A1(net1786),
    .A2(_04214_),
    .Y(_00727_),
    .B1(_04215_));
 sg13g2_nand2_1 _11697_ (.Y(_04216_),
    .A(_01343_),
    .B(\am_sdr0.cic1.comb1[15] ));
 sg13g2_xor2_1 _11698_ (.B(\am_sdr0.cic1.comb1[15] ),
    .A(\am_sdr0.cic1.comb2_in_del[15] ),
    .X(_04217_));
 sg13g2_a21oi_1 _11699_ (.A1(_04208_),
    .A2(_04213_),
    .Y(_04218_),
    .B1(_04207_));
 sg13g2_xnor2_1 _11700_ (.Y(_04219_),
    .A(_04217_),
    .B(_04218_));
 sg13g2_o21ai_1 _11701_ (.B1(net1911),
    .Y(_04220_),
    .A1(net1784),
    .A2(net2376));
 sg13g2_a21oi_1 _11702_ (.A1(net1784),
    .A2(_04219_),
    .Y(_00728_),
    .B1(_04220_));
 sg13g2_nor2_1 _11703_ (.A(\am_sdr0.cic1.comb2_in_del[16] ),
    .B(_01342_),
    .Y(_04221_));
 sg13g2_xor2_1 _11704_ (.B(\am_sdr0.cic1.comb1[16] ),
    .A(\am_sdr0.cic1.comb2_in_del[16] ),
    .X(_04222_));
 sg13g2_nor2_1 _11705_ (.A(_04209_),
    .B(_04217_),
    .Y(_04223_));
 sg13g2_nor3_2 _11706_ (.A(_04209_),
    .B(_04212_),
    .C(_04217_),
    .Y(_04224_));
 sg13g2_o21ai_1 _11707_ (.B1(_04207_),
    .Y(_04225_),
    .A1(_01343_),
    .A2(\am_sdr0.cic1.comb1[15] ));
 sg13g2_a22oi_1 _11708_ (.Y(_04226_),
    .B1(_04224_),
    .B2(_04195_),
    .A2(_04223_),
    .A1(_04210_));
 sg13g2_nand3_1 _11709_ (.B(_04225_),
    .C(_04226_),
    .A(_04216_),
    .Y(_04227_));
 sg13g2_a21oi_2 _11710_ (.B1(_04227_),
    .Y(_04228_),
    .A2(_04224_),
    .A1(_04197_));
 sg13g2_nor2_1 _11711_ (.A(_04222_),
    .B(_04228_),
    .Y(_04229_));
 sg13g2_xnor2_1 _11712_ (.Y(_04230_),
    .A(_04222_),
    .B(_04228_));
 sg13g2_o21ai_1 _11713_ (.B1(net1912),
    .Y(_04231_),
    .A1(net1784),
    .A2(net2147));
 sg13g2_a21oi_1 _11714_ (.A1(net1785),
    .A2(_04230_),
    .Y(_00729_),
    .B1(_04231_));
 sg13g2_nand2_1 _11715_ (.Y(_04232_),
    .A(\am_sdr0.cic1.comb2_in_del[17] ),
    .B(_01341_));
 sg13g2_nor2_1 _11716_ (.A(\am_sdr0.cic1.comb2_in_del[17] ),
    .B(_01341_),
    .Y(_04233_));
 sg13g2_xnor2_1 _11717_ (.Y(_04234_),
    .A(\am_sdr0.cic1.comb2_in_del[17] ),
    .B(\am_sdr0.cic1.comb1[17] ));
 sg13g2_nor2_1 _11718_ (.A(_04221_),
    .B(_04229_),
    .Y(_04235_));
 sg13g2_xor2_1 _11719_ (.B(_04235_),
    .A(_04234_),
    .X(_04236_));
 sg13g2_o21ai_1 _11720_ (.B1(net1911),
    .Y(_04237_),
    .A1(net1784),
    .A2(net2256));
 sg13g2_a21oi_1 _11721_ (.A1(net1784),
    .A2(_04236_),
    .Y(_00730_),
    .B1(_04237_));
 sg13g2_nor2_1 _11722_ (.A(\am_sdr0.cic1.comb2_in_del[18] ),
    .B(_01340_),
    .Y(_04238_));
 sg13g2_xnor2_1 _11723_ (.Y(_04239_),
    .A(\am_sdr0.cic1.comb2_in_del[18] ),
    .B(\am_sdr0.cic1.comb1[18] ));
 sg13g2_nand2b_1 _11724_ (.Y(_04240_),
    .B(_04234_),
    .A_N(_04222_));
 sg13g2_a21oi_1 _11725_ (.A1(_04221_),
    .A2(_04232_),
    .Y(_04241_),
    .B1(_04233_));
 sg13g2_o21ai_1 _11726_ (.B1(_04241_),
    .Y(_04242_),
    .A1(_04228_),
    .A2(_04240_));
 sg13g2_xnor2_1 _11727_ (.Y(_04243_),
    .A(net2610),
    .B(_04242_));
 sg13g2_o21ai_1 _11728_ (.B1(net1911),
    .Y(_04244_),
    .A1(net1788),
    .A2(net2145));
 sg13g2_a21oi_1 _11729_ (.A1(net1784),
    .A2(_04243_),
    .Y(_00731_),
    .B1(_04244_));
 sg13g2_a21oi_1 _11730_ (.A1(_04239_),
    .A2(_04242_),
    .Y(_04245_),
    .B1(_04238_));
 sg13g2_xor2_1 _11731_ (.B(net2119),
    .A(net2309),
    .X(_04246_));
 sg13g2_inv_1 _11732_ (.Y(_04247_),
    .A(_04246_));
 sg13g2_nand2b_1 _11733_ (.Y(_04248_),
    .B(_04246_),
    .A_N(_04245_));
 sg13g2_a21oi_1 _11734_ (.A1(_04245_),
    .A2(_04247_),
    .Y(_04249_),
    .B1(net1639));
 sg13g2_a221oi_1 _11735_ (.B2(_04249_),
    .C1(net1878),
    .B1(net2310),
    .A1(_01305_),
    .Y(_00732_),
    .A2(net1639));
 sg13g2_o21ai_1 _11736_ (.B1(net1919),
    .Y(_04250_),
    .A1(net1774),
    .A2(\am_sdr0.cic1.comb2_in_del[0] ));
 sg13g2_a21oi_1 _11737_ (.A1(net1774),
    .A2(_01360_),
    .Y(_00733_),
    .B1(_04250_));
 sg13g2_o21ai_1 _11738_ (.B1(net1919),
    .Y(_04251_),
    .A1(net1782),
    .A2(\am_sdr0.cic1.comb2_in_del[1] ));
 sg13g2_a21oi_1 _11739_ (.A1(net1780),
    .A2(_01358_),
    .Y(_00734_),
    .B1(_04251_));
 sg13g2_o21ai_1 _11740_ (.B1(net1917),
    .Y(_04252_),
    .A1(net1780),
    .A2(\am_sdr0.cic1.comb2_in_del[2] ));
 sg13g2_a21oi_1 _11741_ (.A1(net1774),
    .A2(_01357_),
    .Y(_00735_),
    .B1(_04252_));
 sg13g2_o21ai_1 _11742_ (.B1(net1918),
    .Y(_04253_),
    .A1(net1780),
    .A2(net2566));
 sg13g2_a21oi_1 _11743_ (.A1(net1780),
    .A2(_01356_),
    .Y(_00736_),
    .B1(_04253_));
 sg13g2_o21ai_1 _11744_ (.B1(net1917),
    .Y(_04254_),
    .A1(net1780),
    .A2(\am_sdr0.cic1.comb2_in_del[4] ));
 sg13g2_a21oi_1 _11745_ (.A1(net1780),
    .A2(_01355_),
    .Y(_00737_),
    .B1(_04254_));
 sg13g2_o21ai_1 _11746_ (.B1(net1917),
    .Y(_04255_),
    .A1(net1638),
    .A2(\am_sdr0.cic1.comb1[5] ));
 sg13g2_a21oi_1 _11747_ (.A1(net1637),
    .A2(_01354_),
    .Y(_00738_),
    .B1(_04255_));
 sg13g2_o21ai_1 _11748_ (.B1(net1917),
    .Y(_04256_),
    .A1(net1779),
    .A2(net2608));
 sg13g2_a21oi_1 _11749_ (.A1(net1779),
    .A2(_01353_),
    .Y(_00739_),
    .B1(_04256_));
 sg13g2_o21ai_1 _11750_ (.B1(net1909),
    .Y(_04257_),
    .A1(net1778),
    .A2(\am_sdr0.cic1.comb2_in_del[7] ));
 sg13g2_a21oi_1 _11751_ (.A1(net1778),
    .A2(_01352_),
    .Y(_00740_),
    .B1(_04257_));
 sg13g2_o21ai_1 _11752_ (.B1(net1909),
    .Y(_04258_),
    .A1(net1778),
    .A2(\am_sdr0.cic1.comb2_in_del[8] ));
 sg13g2_a21oi_1 _11753_ (.A1(net1778),
    .A2(_01351_),
    .Y(_00741_),
    .B1(_04258_));
 sg13g2_o21ai_1 _11754_ (.B1(net1913),
    .Y(_04259_),
    .A1(net1779),
    .A2(net2847));
 sg13g2_a21oi_1 _11755_ (.A1(net1779),
    .A2(_01350_),
    .Y(_00742_),
    .B1(_04259_));
 sg13g2_o21ai_1 _11756_ (.B1(net1909),
    .Y(_04260_),
    .A1(net1769),
    .A2(\am_sdr0.cic1.comb2_in_del[10] ));
 sg13g2_a21oi_1 _11757_ (.A1(net1770),
    .A2(_01348_),
    .Y(_00743_),
    .B1(_04260_));
 sg13g2_o21ai_1 _11758_ (.B1(net1909),
    .Y(_04261_),
    .A1(net1770),
    .A2(net2242));
 sg13g2_a21oi_1 _11759_ (.A1(net1769),
    .A2(_01347_),
    .Y(_00744_),
    .B1(_04261_));
 sg13g2_o21ai_1 _11760_ (.B1(net1913),
    .Y(_04262_),
    .A1(net1771),
    .A2(net2648));
 sg13g2_a21oi_1 _11761_ (.A1(net1770),
    .A2(_01346_),
    .Y(_00745_),
    .B1(_04262_));
 sg13g2_o21ai_1 _11762_ (.B1(net1912),
    .Y(_04263_),
    .A1(net1770),
    .A2(\am_sdr0.cic1.comb2_in_del[13] ));
 sg13g2_a21oi_1 _11763_ (.A1(net1770),
    .A2(_01345_),
    .Y(_00746_),
    .B1(_04263_));
 sg13g2_o21ai_1 _11764_ (.B1(net1912),
    .Y(_04264_),
    .A1(net1771),
    .A2(net2563));
 sg13g2_a21oi_1 _11765_ (.A1(net1768),
    .A2(_01344_),
    .Y(_00747_),
    .B1(_04264_));
 sg13g2_o21ai_1 _11766_ (.B1(net1912),
    .Y(_04265_),
    .A1(net1638),
    .A2(\am_sdr0.cic1.comb1[15] ));
 sg13g2_a21oi_1 _11767_ (.A1(net1638),
    .A2(_01343_),
    .Y(_00748_),
    .B1(_04265_));
 sg13g2_o21ai_1 _11768_ (.B1(net1912),
    .Y(_04266_),
    .A1(net1768),
    .A2(net2689));
 sg13g2_a21oi_1 _11769_ (.A1(net1768),
    .A2(_01342_),
    .Y(_00749_),
    .B1(_04266_));
 sg13g2_o21ai_1 _11770_ (.B1(net1912),
    .Y(_04267_),
    .A1(net1768),
    .A2(net2929));
 sg13g2_a21oi_1 _11771_ (.A1(net1768),
    .A2(_01341_),
    .Y(_00750_),
    .B1(_04267_));
 sg13g2_o21ai_1 _11772_ (.B1(net1912),
    .Y(_04268_),
    .A1(net1768),
    .A2(net2609));
 sg13g2_a21oi_1 _11773_ (.A1(net1768),
    .A2(_01340_),
    .Y(_00751_),
    .B1(_04268_));
 sg13g2_o21ai_1 _11774_ (.B1(net1907),
    .Y(_04269_),
    .A1(net1768),
    .A2(\am_sdr0.cic1.comb2_in_del[19] ));
 sg13g2_a21oi_1 _11775_ (.A1(net1766),
    .A2(_01339_),
    .Y(_00752_),
    .B1(_04269_));
 sg13g2_nand2_1 _11776_ (.Y(_04270_),
    .A(\am_sdr0.cic1.comb3_in_del[4] ),
    .B(_01326_));
 sg13g2_nand2b_1 _11777_ (.Y(_04271_),
    .B(\am_sdr0.cic1.comb3_in_del[1] ),
    .A_N(\am_sdr0.cic1.comb2[1] ));
 sg13g2_nand2b_1 _11778_ (.Y(_04272_),
    .B(\am_sdr0.cic1.comb3_in_del[0] ),
    .A_N(\am_sdr0.cic1.comb2[0] ));
 sg13g2_nor2b_1 _11779_ (.A(\am_sdr0.cic1.comb3_in_del[1] ),
    .B_N(\am_sdr0.cic1.comb2[1] ),
    .Y(_04273_));
 sg13g2_a221oi_1 _11780_ (.B2(_04272_),
    .C1(_04273_),
    .B1(_04271_),
    .A1(_01328_),
    .Y(_04274_),
    .A2(\am_sdr0.cic1.comb2[2] ));
 sg13g2_nand2b_1 _11781_ (.Y(_04275_),
    .B(\am_sdr0.cic1.comb3_in_del[3] ),
    .A_N(\am_sdr0.cic1.comb2[3] ));
 sg13g2_o21ai_1 _11782_ (.B1(_04275_),
    .Y(_04276_),
    .A1(_01328_),
    .A2(\am_sdr0.cic1.comb2[2] ));
 sg13g2_a22oi_1 _11783_ (.Y(_04277_),
    .B1(_01327_),
    .B2(\am_sdr0.cic1.comb2[3] ),
    .A2(\am_sdr0.cic1.comb2[4] ),
    .A1(_01325_));
 sg13g2_o21ai_1 _11784_ (.B1(_04277_),
    .Y(_04278_),
    .A1(_04274_),
    .A2(_04276_));
 sg13g2_a22oi_1 _11785_ (.Y(_04279_),
    .B1(_04270_),
    .B2(_04278_),
    .A2(\am_sdr0.cic1.comb2[5] ),
    .A1(_01324_));
 sg13g2_nand2_1 _11786_ (.Y(_04280_),
    .A(\am_sdr0.cic1.comb3_in_del[6] ),
    .B(_01323_));
 sg13g2_o21ai_1 _11787_ (.B1(_04280_),
    .Y(_04281_),
    .A1(_01324_),
    .A2(\am_sdr0.cic1.comb2[5] ));
 sg13g2_a22oi_1 _11788_ (.Y(_04282_),
    .B1(_01322_),
    .B2(\am_sdr0.cic1.comb2[6] ),
    .A2(\am_sdr0.cic1.comb2[7] ),
    .A1(_01320_));
 sg13g2_o21ai_1 _11789_ (.B1(_04282_),
    .Y(_04283_),
    .A1(_04279_),
    .A2(_04281_));
 sg13g2_nand2_1 _11790_ (.Y(_04284_),
    .A(\am_sdr0.cic1.comb3_in_del[11] ),
    .B(_01315_));
 sg13g2_a22oi_1 _11791_ (.Y(_04285_),
    .B1(_01318_),
    .B2(\am_sdr0.cic1.comb2[8] ),
    .A2(\am_sdr0.cic1.comb2[9] ),
    .A1(_01317_));
 sg13g2_nand2b_1 _11792_ (.Y(_04286_),
    .B(\am_sdr0.cic1.comb3_in_del[10] ),
    .A_N(\am_sdr0.cic1.comb2[10] ));
 sg13g2_o21ai_1 _11793_ (.B1(_04286_),
    .Y(_04287_),
    .A1(_01317_),
    .A2(\am_sdr0.cic1.comb2[9] ));
 sg13g2_a22oi_1 _11794_ (.Y(_04288_),
    .B1(_01316_),
    .B2(\am_sdr0.cic1.comb2[10] ),
    .A2(\am_sdr0.cic1.comb2[11] ),
    .A1(_01314_));
 sg13g2_nand3b_1 _11795_ (.B(_04288_),
    .C(_04284_),
    .Y(_04289_),
    .A_N(_04287_));
 sg13g2_a221oi_1 _11796_ (.B2(_01321_),
    .C1(_04289_),
    .B1(\am_sdr0.cic1.comb3_in_del[7] ),
    .A1(\am_sdr0.cic1.comb3_in_del[8] ),
    .Y(_04290_),
    .A2(_01319_));
 sg13g2_and2_1 _11797_ (.A(_04285_),
    .B(_04290_),
    .X(_04291_));
 sg13g2_o21ai_1 _11798_ (.B1(_04288_),
    .Y(_04292_),
    .A1(_04285_),
    .A2(_04287_));
 sg13g2_a22oi_1 _11799_ (.Y(_04293_),
    .B1(_04292_),
    .B2(_04284_),
    .A2(_04291_),
    .A1(_04283_));
 sg13g2_xnor2_1 _11800_ (.Y(_04294_),
    .A(net2367),
    .B(net3326));
 sg13g2_nor2b_1 _11801_ (.A(_04293_),
    .B_N(_04294_),
    .Y(_04295_));
 sg13g2_xor2_1 _11802_ (.B(_04294_),
    .A(_04293_),
    .X(_04296_));
 sg13g2_o21ai_1 _11803_ (.B1(net1963),
    .Y(_04297_),
    .A1(net1792),
    .A2(net1283));
 sg13g2_a21oi_1 _11804_ (.A1(net1791),
    .A2(_04296_),
    .Y(_00753_),
    .B1(_04297_));
 sg13g2_nand2_1 _11805_ (.Y(_04298_),
    .A(\am_sdr0.cic1.comb3_in_del[13] ),
    .B(_01312_));
 sg13g2_xnor2_1 _11806_ (.Y(_04299_),
    .A(\am_sdr0.cic1.comb3_in_del[13] ),
    .B(net2335));
 sg13g2_a21oi_1 _11807_ (.A1(_01313_),
    .A2(\am_sdr0.cic1.comb2[12] ),
    .Y(_04300_),
    .B1(_04295_));
 sg13g2_o21ai_1 _11808_ (.B1(net1791),
    .Y(_04301_),
    .A1(_04299_),
    .A2(_04300_));
 sg13g2_a21oi_1 _11809_ (.A1(net2336),
    .A2(_04300_),
    .Y(_04302_),
    .B1(_04301_));
 sg13g2_o21ai_1 _11810_ (.B1(net1963),
    .Y(_04303_),
    .A1(net1791),
    .A2(net1337));
 sg13g2_nor2_1 _11811_ (.A(net2337),
    .B(_04303_),
    .Y(_00754_));
 sg13g2_nor2_1 _11812_ (.A(net2323),
    .B(_01311_),
    .Y(_04304_));
 sg13g2_xor2_1 _11813_ (.B(\am_sdr0.cic1.comb2[14] ),
    .A(net2323),
    .X(_04305_));
 sg13g2_nand3_1 _11814_ (.B(\am_sdr0.cic1.comb2[12] ),
    .C(_04298_),
    .A(_01313_),
    .Y(_04306_));
 sg13g2_o21ai_1 _11815_ (.B1(_04306_),
    .Y(_04307_),
    .A1(\am_sdr0.cic1.comb3_in_del[13] ),
    .A2(_01312_));
 sg13g2_a21oi_1 _11816_ (.A1(_04295_),
    .A2(_04299_),
    .Y(_04308_),
    .B1(_04307_));
 sg13g2_nor2_1 _11817_ (.A(_04305_),
    .B(_04308_),
    .Y(_04309_));
 sg13g2_xnor2_1 _11818_ (.Y(_04310_),
    .A(net2324),
    .B(_04308_));
 sg13g2_o21ai_1 _11819_ (.B1(net1961),
    .Y(_04311_),
    .A1(net1792),
    .A2(net1241));
 sg13g2_a21oi_1 _11820_ (.A1(net1791),
    .A2(_04310_),
    .Y(_00755_),
    .B1(_04311_));
 sg13g2_nor2_1 _11821_ (.A(net2414),
    .B(_01310_),
    .Y(_04312_));
 sg13g2_nand2_1 _11822_ (.Y(_04313_),
    .A(net2414),
    .B(_01310_));
 sg13g2_nor2b_1 _11823_ (.A(_04312_),
    .B_N(_04313_),
    .Y(_04314_));
 sg13g2_nor2_1 _11824_ (.A(_04304_),
    .B(_04309_),
    .Y(_04315_));
 sg13g2_o21ai_1 _11825_ (.B1(net1791),
    .Y(_04316_),
    .A1(_04314_),
    .A2(_04315_));
 sg13g2_a21oi_1 _11826_ (.A1(_04314_),
    .A2(_04315_),
    .Y(_04317_),
    .B1(_04316_));
 sg13g2_o21ai_1 _11827_ (.B1(net1962),
    .Y(_04318_),
    .A1(net1790),
    .A2(net1226));
 sg13g2_nor2_1 _11828_ (.A(_04317_),
    .B(_04318_),
    .Y(_00756_));
 sg13g2_nor2_1 _11829_ (.A(\am_sdr0.cic1.comb3_in_del[16] ),
    .B(_01309_),
    .Y(_04319_));
 sg13g2_xnor2_1 _11830_ (.Y(_04320_),
    .A(net2269),
    .B(net2147));
 sg13g2_nor2b_1 _11831_ (.A(_04305_),
    .B_N(_04314_),
    .Y(_04321_));
 sg13g2_nand3_1 _11832_ (.B(_04299_),
    .C(_04321_),
    .A(_04294_),
    .Y(_04322_));
 sg13g2_a221oi_1 _11833_ (.B2(_04307_),
    .C1(_04312_),
    .B1(_04321_),
    .A1(_04304_),
    .Y(_04323_),
    .A2(_04313_));
 sg13g2_o21ai_1 _11834_ (.B1(_04323_),
    .Y(_04324_),
    .A1(_04293_),
    .A2(_04322_));
 sg13g2_xnor2_1 _11835_ (.Y(_04325_),
    .A(_04320_),
    .B(_04324_));
 sg13g2_o21ai_1 _11836_ (.B1(net1962),
    .Y(_04326_),
    .A1(net1790),
    .A2(net1366));
 sg13g2_a21oi_1 _11837_ (.A1(net1790),
    .A2(_04325_),
    .Y(_00757_),
    .B1(_04326_));
 sg13g2_a21oi_1 _11838_ (.A1(_04320_),
    .A2(_04324_),
    .Y(_04327_),
    .B1(_04319_));
 sg13g2_nand2b_1 _11839_ (.Y(_04328_),
    .B(\am_sdr0.cic1.comb2[17] ),
    .A_N(\am_sdr0.cic1.comb3_in_del[17] ));
 sg13g2_nor2b_1 _11840_ (.A(net2256),
    .B_N(\am_sdr0.cic1.comb3_in_del[17] ),
    .Y(_04329_));
 sg13g2_xnor2_1 _11841_ (.Y(_04330_),
    .A(net2029),
    .B(\am_sdr0.cic1.comb2[17] ));
 sg13g2_or2_1 _11842_ (.X(_04331_),
    .B(net2030),
    .A(_04327_));
 sg13g2_a21oi_1 _11843_ (.A1(_04327_),
    .A2(net2030),
    .Y(_04332_),
    .B1(net1640));
 sg13g2_a221oi_1 _11844_ (.B2(_04332_),
    .C1(net1888),
    .B1(_04331_),
    .A1(net1640),
    .Y(_00758_),
    .A2(_01333_));
 sg13g2_xnor2_1 _11845_ (.Y(_04333_),
    .A(\am_sdr0.cic1.comb3_in_del[18] ),
    .B(net2145));
 sg13g2_a21oi_1 _11846_ (.A1(_04327_),
    .A2(_04328_),
    .Y(_04334_),
    .B1(net2257));
 sg13g2_nand2_1 _11847_ (.Y(_04335_),
    .A(_04333_),
    .B(_04334_));
 sg13g2_xnor2_1 _11848_ (.Y(_04336_),
    .A(_04333_),
    .B(net2258));
 sg13g2_o21ai_1 _11849_ (.B1(net1961),
    .Y(_04337_),
    .A1(net1790),
    .A2(net1264));
 sg13g2_a21oi_1 _11850_ (.A1(net1790),
    .A2(net2259),
    .Y(_00759_),
    .B1(_04337_));
 sg13g2_o21ai_1 _11851_ (.B1(_04335_),
    .Y(_04338_),
    .A1(\am_sdr0.cic1.comb3_in_del[18] ),
    .A2(_01307_));
 sg13g2_xor2_1 _11852_ (.B(net2061),
    .A(net2178),
    .X(_04339_));
 sg13g2_or2_1 _11853_ (.X(_04340_),
    .B(_04339_),
    .A(_04338_));
 sg13g2_a21oi_1 _11854_ (.A1(_04338_),
    .A2(_04339_),
    .Y(_04341_),
    .B1(net1639));
 sg13g2_a221oi_1 _11855_ (.B2(net2179),
    .C1(net1888),
    .B1(_04340_),
    .A1(net1639),
    .Y(_00760_),
    .A2(_01331_));
 sg13g2_o21ai_1 _11856_ (.B1(net1919),
    .Y(_04342_),
    .A1(net1781),
    .A2(\am_sdr0.cic1.comb3_in_del[0] ));
 sg13g2_a21oi_1 _11857_ (.A1(net1780),
    .A2(_01330_),
    .Y(_00761_),
    .B1(_04342_));
 sg13g2_o21ai_1 _11858_ (.B1(net1923),
    .Y(_04343_),
    .A1(net1782),
    .A2(\am_sdr0.cic1.comb3_in_del[1] ));
 sg13g2_a21oi_1 _11859_ (.A1(net1781),
    .A2(_01329_),
    .Y(_00762_),
    .B1(_04343_));
 sg13g2_o21ai_1 _11860_ (.B1(net1921),
    .Y(_04344_),
    .A1(net1638),
    .A2(\am_sdr0.cic1.comb2[2] ));
 sg13g2_a21oi_1 _11861_ (.A1(net1641),
    .A2(_01328_),
    .Y(_00763_),
    .B1(_04344_));
 sg13g2_o21ai_1 _11862_ (.B1(net1921),
    .Y(_04345_),
    .A1(net1637),
    .A2(\am_sdr0.cic1.comb2[3] ));
 sg13g2_a21oi_1 _11863_ (.A1(net1641),
    .A2(_01327_),
    .Y(_00764_),
    .B1(_04345_));
 sg13g2_o21ai_1 _11864_ (.B1(net1922),
    .Y(_04346_),
    .A1(net1796),
    .A2(\am_sdr0.cic1.comb3_in_del[4] ));
 sg13g2_a21oi_1 _11865_ (.A1(net1796),
    .A2(_01326_),
    .Y(_00765_),
    .B1(_04346_));
 sg13g2_o21ai_1 _11866_ (.B1(net1921),
    .Y(_04347_),
    .A1(net1640),
    .A2(\am_sdr0.cic1.comb2[5] ));
 sg13g2_a21oi_1 _11867_ (.A1(net1640),
    .A2(_01324_),
    .Y(_00766_),
    .B1(_04347_));
 sg13g2_o21ai_1 _11868_ (.B1(net1921),
    .Y(_04348_),
    .A1(net1794),
    .A2(\am_sdr0.cic1.comb3_in_del[6] ));
 sg13g2_a21oi_1 _11869_ (.A1(net1794),
    .A2(_01323_),
    .Y(_00767_),
    .B1(_04348_));
 sg13g2_o21ai_1 _11870_ (.B1(net1925),
    .Y(_04349_),
    .A1(net1794),
    .A2(\am_sdr0.cic1.comb3_in_del[7] ));
 sg13g2_a21oi_1 _11871_ (.A1(net1794),
    .A2(_01321_),
    .Y(_00768_),
    .B1(_04349_));
 sg13g2_o21ai_1 _11872_ (.B1(net1914),
    .Y(_04350_),
    .A1(net1794),
    .A2(\am_sdr0.cic1.comb3_in_del[8] ));
 sg13g2_a21oi_1 _11873_ (.A1(net1794),
    .A2(_01319_),
    .Y(_00769_),
    .B1(_04350_));
 sg13g2_o21ai_1 _11874_ (.B1(net1913),
    .Y(_04351_),
    .A1(net1640),
    .A2(\am_sdr0.cic1.comb2[9] ));
 sg13g2_a21oi_1 _11875_ (.A1(net1640),
    .A2(_01317_),
    .Y(_00770_),
    .B1(_04351_));
 sg13g2_o21ai_1 _11876_ (.B1(net1913),
    .Y(_04352_),
    .A1(net1639),
    .A2(\am_sdr0.cic1.comb2[10] ));
 sg13g2_a21oi_1 _11877_ (.A1(net1639),
    .A2(_01316_),
    .Y(_00771_),
    .B1(_04352_));
 sg13g2_o21ai_1 _11878_ (.B1(net1914),
    .Y(_04353_),
    .A1(net1786),
    .A2(net2427));
 sg13g2_a21oi_1 _11879_ (.A1(net1786),
    .A2(_01315_),
    .Y(_00772_),
    .B1(_04353_));
 sg13g2_o21ai_1 _11880_ (.B1(net1914),
    .Y(_04354_),
    .A1(net1639),
    .A2(net2718));
 sg13g2_a21oi_1 _11881_ (.A1(net1639),
    .A2(_01313_),
    .Y(_00773_),
    .B1(_04354_));
 sg13g2_o21ai_1 _11882_ (.B1(net1914),
    .Y(_04355_),
    .A1(net1787),
    .A2(net2825));
 sg13g2_a21oi_1 _11883_ (.A1(net1787),
    .A2(_01312_),
    .Y(_00774_),
    .B1(_04355_));
 sg13g2_o21ai_1 _11884_ (.B1(net1915),
    .Y(_04356_),
    .A1(net1787),
    .A2(net2323));
 sg13g2_a21oi_1 _11885_ (.A1(net1787),
    .A2(_01311_),
    .Y(_00775_),
    .B1(_04356_));
 sg13g2_o21ai_1 _11886_ (.B1(net1915),
    .Y(_04357_),
    .A1(net1787),
    .A2(net2414));
 sg13g2_a21oi_1 _11887_ (.A1(net1788),
    .A2(_01310_),
    .Y(_00776_),
    .B1(_04357_));
 sg13g2_o21ai_1 _11888_ (.B1(net1911),
    .Y(_04358_),
    .A1(net1785),
    .A2(\am_sdr0.cic1.comb3_in_del[16] ));
 sg13g2_a21oi_1 _11889_ (.A1(net1785),
    .A2(_01309_),
    .Y(_00777_),
    .B1(_04358_));
 sg13g2_o21ai_1 _11890_ (.B1(net1911),
    .Y(_04359_),
    .A1(net1785),
    .A2(net2029));
 sg13g2_a21oi_1 _11891_ (.A1(net1785),
    .A2(_01308_),
    .Y(_00778_),
    .B1(_04359_));
 sg13g2_o21ai_1 _11892_ (.B1(net1911),
    .Y(_04360_),
    .A1(net1785),
    .A2(\am_sdr0.cic1.comb3_in_del[18] ));
 sg13g2_a21oi_1 _11893_ (.A1(net1785),
    .A2(_01307_),
    .Y(_00779_),
    .B1(_04360_));
 sg13g2_o21ai_1 _11894_ (.B1(net1911),
    .Y(_04361_),
    .A1(\am_sdr0.cic1.comb3_in_del[19] ),
    .A2(net1784));
 sg13g2_a21oi_1 _11895_ (.A1(_01305_),
    .A2(net1784),
    .Y(_00780_),
    .B1(_04361_));
 sg13g2_o21ai_1 _11896_ (.B1(net1901),
    .Y(_04362_),
    .A1(_02974_),
    .A2(_02975_));
 sg13g2_nor2_1 _11897_ (.A(_01594_),
    .B(_04362_),
    .Y(_00782_));
 sg13g2_xnor2_1 _11898_ (.Y(_04363_),
    .A(\am_sdr0.cic1.count[0] ),
    .B(net2174));
 sg13g2_nor2_1 _11899_ (.A(_04362_),
    .B(net2175),
    .Y(_00783_));
 sg13g2_a21oi_1 _11900_ (.A1(\am_sdr0.cic1.count[0] ),
    .A2(\am_sdr0.cic1.count[1] ),
    .Y(_04364_),
    .B1(net1202));
 sg13g2_nor3_1 _11901_ (.A(_02971_),
    .B(_04362_),
    .C(net1203),
    .Y(_00784_));
 sg13g2_nor2_1 _11902_ (.A(net1439),
    .B(_02971_),
    .Y(_04365_));
 sg13g2_nor3_1 _11903_ (.A(net1877),
    .B(_02972_),
    .C(net1440),
    .Y(_00785_));
 sg13g2_nor2_1 _11904_ (.A(net1429),
    .B(_02972_),
    .Y(_04366_));
 sg13g2_nor3_1 _11905_ (.A(net1877),
    .B(_02973_),
    .C(net1430),
    .Y(_00786_));
 sg13g2_o21ai_1 _11906_ (.B1(net1901),
    .Y(_04367_),
    .A1(net2857),
    .A2(_02973_));
 sg13g2_nor2b_1 _11907_ (.A(_04367_),
    .B_N(_02974_),
    .Y(_00787_));
 sg13g2_a21oi_1 _11908_ (.A1(\am_sdr0.cic1.count[5] ),
    .A2(_02973_),
    .Y(_04368_),
    .B1(net1372));
 sg13g2_and3_1 _11909_ (.X(_04369_),
    .A(\am_sdr0.cic1.count[5] ),
    .B(net1372),
    .C(_02973_));
 sg13g2_nor3_1 _11910_ (.A(_04362_),
    .B(net1373),
    .C(_04369_),
    .Y(_00788_));
 sg13g2_o21ai_1 _11911_ (.B1(net1901),
    .Y(_04370_),
    .A1(net1208),
    .A2(_04369_));
 sg13g2_a21oi_1 _11912_ (.A1(net1208),
    .A2(_04369_),
    .Y(_00789_),
    .B1(_04370_));
 sg13g2_nand2_1 _11913_ (.Y(_04371_),
    .A(net3122),
    .B(net2185));
 sg13g2_o21ai_1 _11914_ (.B1(net1930),
    .Y(_04372_),
    .A1(\am_sdr0.Q_out[0] ),
    .A2(net2185));
 sg13g2_nor2b_1 _11915_ (.A(net2186),
    .B_N(_04371_),
    .Y(_00790_));
 sg13g2_nand2_1 _11916_ (.Y(_04373_),
    .A(\am_sdr0.Q_out[1] ),
    .B(\am_sdr0.cic1.integ1[1] ));
 sg13g2_xnor2_1 _11917_ (.Y(_04374_),
    .A(\am_sdr0.Q_out[1] ),
    .B(\am_sdr0.cic1.integ1[1] ));
 sg13g2_and2_1 _11918_ (.A(_04371_),
    .B(_04374_),
    .X(_04375_));
 sg13g2_nor2_1 _11919_ (.A(_04371_),
    .B(_04374_),
    .Y(_04376_));
 sg13g2_nor3_1 _11920_ (.A(net1879),
    .B(net3123),
    .C(_04376_),
    .Y(_00791_));
 sg13g2_and2_1 _11921_ (.A(net3084),
    .B(net3282),
    .X(_04377_));
 sg13g2_xnor2_1 _11922_ (.Y(_04378_),
    .A(net3084),
    .B(\am_sdr0.cic1.integ1[2] ));
 sg13g2_inv_1 _11923_ (.Y(_04379_),
    .A(_04378_));
 sg13g2_a21oi_1 _11924_ (.A1(\am_sdr0.Q_out[1] ),
    .A2(\am_sdr0.cic1.integ1[1] ),
    .Y(_04380_),
    .B1(_04376_));
 sg13g2_o21ai_1 _11925_ (.B1(_04373_),
    .Y(_04381_),
    .A1(_04371_),
    .A2(_04374_));
 sg13g2_o21ai_1 _11926_ (.B1(net1904),
    .Y(_04382_),
    .A1(net3085),
    .A2(_04380_));
 sg13g2_a21oi_1 _11927_ (.A1(net3085),
    .A2(_04380_),
    .Y(_00792_),
    .B1(_04382_));
 sg13g2_nand2_1 _11928_ (.Y(_04383_),
    .A(\am_sdr0.Q_out[3] ),
    .B(\am_sdr0.cic1.integ1[3] ));
 sg13g2_xnor2_1 _11929_ (.Y(_04384_),
    .A(net3230),
    .B(\am_sdr0.cic1.integ1[3] ));
 sg13g2_a21oi_1 _11930_ (.A1(_04379_),
    .A2(_04381_),
    .Y(_04385_),
    .B1(_04377_));
 sg13g2_nor2_1 _11931_ (.A(_04384_),
    .B(_04385_),
    .Y(_04386_));
 sg13g2_a21oi_1 _11932_ (.A1(_04384_),
    .A2(_04385_),
    .Y(_04387_),
    .B1(net1877));
 sg13g2_nor2b_1 _11933_ (.A(_04386_),
    .B_N(_04387_),
    .Y(_00793_));
 sg13g2_a21oi_1 _11934_ (.A1(net3230),
    .A2(\am_sdr0.cic1.integ1[3] ),
    .Y(_04388_),
    .B1(_04386_));
 sg13g2_o21ai_1 _11935_ (.B1(_04383_),
    .Y(_04389_),
    .A1(_04384_),
    .A2(_04385_));
 sg13g2_xnor2_1 _11936_ (.Y(_04390_),
    .A(net3057),
    .B(\am_sdr0.cic1.integ1[4] ));
 sg13g2_nor2_1 _11937_ (.A(_04388_),
    .B(_04390_),
    .Y(_04391_));
 sg13g2_a21oi_1 _11938_ (.A1(_04388_),
    .A2(_04390_),
    .Y(_04392_),
    .B1(net1877));
 sg13g2_nor2b_1 _11939_ (.A(_04391_),
    .B_N(_04392_),
    .Y(_00794_));
 sg13g2_nand2_1 _11940_ (.Y(_04393_),
    .A(\am_sdr0.Q_out[5] ),
    .B(\am_sdr0.cic1.integ1[5] ));
 sg13g2_or2_1 _11941_ (.X(_04394_),
    .B(\am_sdr0.cic1.integ1[5] ),
    .A(\am_sdr0.Q_out[5] ));
 sg13g2_nand2_1 _11942_ (.Y(_04395_),
    .A(_04393_),
    .B(_04394_));
 sg13g2_a21oi_1 _11943_ (.A1(net3057),
    .A2(\am_sdr0.cic1.integ1[4] ),
    .Y(_04396_),
    .B1(_04391_));
 sg13g2_o21ai_1 _11944_ (.B1(net1901),
    .Y(_04397_),
    .A1(_04395_),
    .A2(net3058));
 sg13g2_a21oi_1 _11945_ (.A1(_04395_),
    .A2(net3058),
    .Y(_00795_),
    .B1(_04397_));
 sg13g2_nand2_1 _11946_ (.Y(_04398_),
    .A(net3149),
    .B(\am_sdr0.cic1.integ1[6] ));
 sg13g2_xnor2_1 _11947_ (.Y(_04399_),
    .A(net3149),
    .B(\am_sdr0.cic1.integ1[6] ));
 sg13g2_nor2_1 _11948_ (.A(_04390_),
    .B(_04395_),
    .Y(_04400_));
 sg13g2_nand3_1 _11949_ (.B(\am_sdr0.cic1.integ1[4] ),
    .C(_04394_),
    .A(net3057),
    .Y(_04401_));
 sg13g2_nand2_1 _11950_ (.Y(_04402_),
    .A(_04393_),
    .B(_04401_));
 sg13g2_a21oi_1 _11951_ (.A1(_04389_),
    .A2(_04400_),
    .Y(_04403_),
    .B1(_04402_));
 sg13g2_o21ai_1 _11952_ (.B1(net1904),
    .Y(_04404_),
    .A1(_04399_),
    .A2(_04403_));
 sg13g2_a21oi_1 _11953_ (.A1(net3150),
    .A2(_04403_),
    .Y(_00796_),
    .B1(_04404_));
 sg13g2_and2_1 _11954_ (.A(net1662),
    .B(net3197),
    .X(_04405_));
 sg13g2_or2_1 _11955_ (.X(_04406_),
    .B(net3197),
    .A(net1662));
 sg13g2_nand2b_1 _11956_ (.Y(_04407_),
    .B(_04406_),
    .A_N(_04405_));
 sg13g2_o21ai_1 _11957_ (.B1(_04398_),
    .Y(_04408_),
    .A1(_04399_),
    .A2(_04403_));
 sg13g2_nand2b_1 _11958_ (.Y(_04409_),
    .B(_04407_),
    .A_N(_04408_));
 sg13g2_nand2b_1 _11959_ (.Y(_04410_),
    .B(_04408_),
    .A_N(_04407_));
 sg13g2_and3_1 _11960_ (.X(_00797_),
    .A(net1902),
    .B(_04409_),
    .C(_04410_));
 sg13g2_a21oi_1 _11961_ (.A1(_04406_),
    .A2(_04408_),
    .Y(_04411_),
    .B1(_04405_));
 sg13g2_a21o_1 _11962_ (.A2(_04408_),
    .A1(_04406_),
    .B1(_04405_),
    .X(_04412_));
 sg13g2_nand2_1 _11963_ (.Y(_04413_),
    .A(net1660),
    .B(net3285));
 sg13g2_xnor2_1 _11964_ (.Y(_04414_),
    .A(net1660),
    .B(\am_sdr0.cic1.integ1[8] ));
 sg13g2_nand2b_1 _11965_ (.Y(_04415_),
    .B(_04412_),
    .A_N(_04414_));
 sg13g2_nand2_1 _11966_ (.Y(_04416_),
    .A(net1902),
    .B(_04415_));
 sg13g2_a21oi_1 _11967_ (.A1(_04411_),
    .A2(_04414_),
    .Y(_00798_),
    .B1(_04416_));
 sg13g2_xnor2_1 _11968_ (.Y(_04417_),
    .A(net1660),
    .B(net3283));
 sg13g2_a21oi_1 _11969_ (.A1(_04413_),
    .A2(_04415_),
    .Y(_04418_),
    .B1(_04417_));
 sg13g2_and3_1 _11970_ (.X(_04419_),
    .A(_04413_),
    .B(_04415_),
    .C(_04417_));
 sg13g2_nor3_1 _11971_ (.A(net1876),
    .B(_04418_),
    .C(_04419_),
    .Y(_00799_));
 sg13g2_nand2_1 _11972_ (.Y(_04420_),
    .A(net1660),
    .B(\am_sdr0.cic1.integ1[10] ));
 sg13g2_xor2_1 _11973_ (.B(\am_sdr0.cic1.integ1[10] ),
    .A(net1660),
    .X(_04421_));
 sg13g2_xnor2_1 _11974_ (.Y(_04422_),
    .A(net1660),
    .B(\am_sdr0.cic1.integ1[10] ));
 sg13g2_o21ai_1 _11975_ (.B1(net1662),
    .Y(_04423_),
    .A1(\am_sdr0.cic1.integ1[8] ),
    .A2(\am_sdr0.cic1.integ1[9] ));
 sg13g2_o21ai_1 _11976_ (.B1(_04423_),
    .Y(_04424_),
    .A1(_04415_),
    .A2(_04417_));
 sg13g2_nand2_1 _11977_ (.Y(_04425_),
    .A(_04421_),
    .B(_04424_));
 sg13g2_o21ai_1 _11978_ (.B1(net1902),
    .Y(_04426_),
    .A1(_04421_),
    .A2(_04424_));
 sg13g2_nor2b_1 _11979_ (.A(_04426_),
    .B_N(_04425_),
    .Y(_00800_));
 sg13g2_xnor2_1 _11980_ (.Y(_04427_),
    .A(net1660),
    .B(net3237));
 sg13g2_and3_1 _11981_ (.X(_04428_),
    .A(_04420_),
    .B(_04425_),
    .C(_04427_));
 sg13g2_a21oi_1 _11982_ (.A1(_04420_),
    .A2(_04425_),
    .Y(_04429_),
    .B1(_04427_));
 sg13g2_nor3_1 _11983_ (.A(net1876),
    .B(_04428_),
    .C(_04429_),
    .Y(_00801_));
 sg13g2_nand2_1 _11984_ (.Y(_04430_),
    .A(net1661),
    .B(net3218));
 sg13g2_xnor2_1 _11985_ (.Y(_04431_),
    .A(net1661),
    .B(net3325));
 sg13g2_o21ai_1 _11986_ (.B1(net1660),
    .Y(_04432_),
    .A1(\am_sdr0.cic1.integ1[10] ),
    .A2(\am_sdr0.cic1.integ1[11] ));
 sg13g2_nand2_1 _11987_ (.Y(_04433_),
    .A(_04423_),
    .B(_04432_));
 sg13g2_nor4_1 _11988_ (.A(_04414_),
    .B(_04417_),
    .C(_04422_),
    .D(_04427_),
    .Y(_04434_));
 sg13g2_a21oi_1 _11989_ (.A1(_04412_),
    .A2(_04434_),
    .Y(_04435_),
    .B1(_04433_));
 sg13g2_or2_1 _11990_ (.X(_04436_),
    .B(_04435_),
    .A(_04431_));
 sg13g2_a21oi_1 _11991_ (.A1(_04431_),
    .A2(_04435_),
    .Y(_04437_),
    .B1(net1876));
 sg13g2_and2_1 _11992_ (.A(_04436_),
    .B(_04437_),
    .X(_00802_));
 sg13g2_xor2_1 _11993_ (.B(\am_sdr0.cic1.integ1[13] ),
    .A(net1661),
    .X(_04438_));
 sg13g2_nand2_1 _11994_ (.Y(_04439_),
    .A(_04430_),
    .B(_04436_));
 sg13g2_o21ai_1 _11995_ (.B1(net1898),
    .Y(_04440_),
    .A1(_04438_),
    .A2(_04439_));
 sg13g2_a21oi_1 _11996_ (.A1(_04438_),
    .A2(_04439_),
    .Y(_00803_),
    .B1(_04440_));
 sg13g2_nand2_1 _11997_ (.Y(_04441_),
    .A(net1661),
    .B(\am_sdr0.cic1.integ1[14] ));
 sg13g2_xnor2_1 _11998_ (.Y(_04442_),
    .A(net1661),
    .B(net3248));
 sg13g2_o21ai_1 _11999_ (.B1(net1661),
    .Y(_04443_),
    .A1(\am_sdr0.cic1.integ1[12] ),
    .A2(\am_sdr0.cic1.integ1[13] ));
 sg13g2_nand2b_1 _12000_ (.Y(_04444_),
    .B(_04438_),
    .A_N(_04431_));
 sg13g2_nor2_1 _12001_ (.A(_04435_),
    .B(_04444_),
    .Y(_04445_));
 sg13g2_nor2b_1 _12002_ (.A(_04445_),
    .B_N(_04443_),
    .Y(_04446_));
 sg13g2_or2_1 _12003_ (.X(_04447_),
    .B(_04446_),
    .A(_04442_));
 sg13g2_nand2_1 _12004_ (.Y(_04448_),
    .A(net1898),
    .B(_04447_));
 sg13g2_a21oi_1 _12005_ (.A1(_04442_),
    .A2(_04446_),
    .Y(_00804_),
    .B1(_04448_));
 sg13g2_xnor2_1 _12006_ (.Y(_04449_),
    .A(net1661),
    .B(\am_sdr0.cic1.integ1[15] ));
 sg13g2_nand3_1 _12007_ (.B(_04447_),
    .C(_04449_),
    .A(_04441_),
    .Y(_04450_));
 sg13g2_a21o_1 _12008_ (.A2(_04447_),
    .A1(_04441_),
    .B1(_04449_),
    .X(_04451_));
 sg13g2_and3_1 _12009_ (.X(_00805_),
    .A(net1898),
    .B(_04450_),
    .C(_04451_));
 sg13g2_nor3_1 _12010_ (.A(_04442_),
    .B(_04444_),
    .C(_04449_),
    .Y(_04452_));
 sg13g2_and2_1 _12011_ (.A(_04434_),
    .B(_04452_),
    .X(_04453_));
 sg13g2_o21ai_1 _12012_ (.B1(net1661),
    .Y(_04454_),
    .A1(\am_sdr0.cic1.integ1[14] ),
    .A2(\am_sdr0.cic1.integ1[15] ));
 sg13g2_nand4_1 _12013_ (.B(_04432_),
    .C(_04443_),
    .A(_04423_),
    .Y(_04455_),
    .D(_04454_));
 sg13g2_a21oi_2 _12014_ (.B1(_04455_),
    .Y(_04456_),
    .A2(_04453_),
    .A1(_04412_));
 sg13g2_xnor2_1 _12015_ (.Y(_04457_),
    .A(net1658),
    .B(\am_sdr0.cic1.integ1[16] ));
 sg13g2_nor2_1 _12016_ (.A(_04456_),
    .B(_04457_),
    .Y(_04458_));
 sg13g2_a21oi_1 _12017_ (.A1(_04456_),
    .A2(_04457_),
    .Y(_04459_),
    .B1(net1875));
 sg13g2_nor2b_1 _12018_ (.A(_04458_),
    .B_N(_04459_),
    .Y(_00806_));
 sg13g2_xor2_1 _12019_ (.B(\am_sdr0.cic1.integ1[17] ),
    .A(net1659),
    .X(_04460_));
 sg13g2_xnor2_1 _12020_ (.Y(_04461_),
    .A(net1658),
    .B(net3264));
 sg13g2_a21oi_1 _12021_ (.A1(net1658),
    .A2(\am_sdr0.cic1.integ1[16] ),
    .Y(_04462_),
    .B1(_04458_));
 sg13g2_o21ai_1 _12022_ (.B1(net1898),
    .Y(_04463_),
    .A1(_04461_),
    .A2(_04462_));
 sg13g2_a21oi_1 _12023_ (.A1(_04461_),
    .A2(_04462_),
    .Y(_00807_),
    .B1(_04463_));
 sg13g2_and2_1 _12024_ (.A(net1658),
    .B(\am_sdr0.cic1.integ1[18] ),
    .X(_04464_));
 sg13g2_xnor2_1 _12025_ (.Y(_04465_),
    .A(net1658),
    .B(\am_sdr0.cic1.integ1[18] ));
 sg13g2_o21ai_1 _12026_ (.B1(net1658),
    .Y(_04466_),
    .A1(\am_sdr0.cic1.integ1[16] ),
    .A2(\am_sdr0.cic1.integ1[17] ));
 sg13g2_inv_1 _12027_ (.Y(_04467_),
    .A(_04466_));
 sg13g2_a21oi_1 _12028_ (.A1(_04458_),
    .A2(_04460_),
    .Y(_04468_),
    .B1(_04467_));
 sg13g2_nor2_1 _12029_ (.A(_04465_),
    .B(_04468_),
    .Y(_04469_));
 sg13g2_a21oi_1 _12030_ (.A1(_04465_),
    .A2(_04468_),
    .Y(_04470_),
    .B1(net1875));
 sg13g2_nor2b_1 _12031_ (.A(_04469_),
    .B_N(_04470_),
    .Y(_00808_));
 sg13g2_xor2_1 _12032_ (.B(\am_sdr0.cic1.integ1[19] ),
    .A(net1658),
    .X(_04471_));
 sg13g2_or3_1 _12033_ (.A(_04464_),
    .B(_04469_),
    .C(_04471_),
    .X(_04472_));
 sg13g2_o21ai_1 _12034_ (.B1(_04471_),
    .Y(_04473_),
    .A1(_04464_),
    .A2(_04469_));
 sg13g2_and3_1 _12035_ (.X(_00809_),
    .A(net1896),
    .B(_04472_),
    .C(_04473_));
 sg13g2_nor2_1 _12036_ (.A(_04457_),
    .B(_04461_),
    .Y(_04474_));
 sg13g2_nand3b_1 _12037_ (.B(_04471_),
    .C(_04474_),
    .Y(_04475_),
    .A_N(_04465_));
 sg13g2_nor2_1 _12038_ (.A(_04456_),
    .B(_04475_),
    .Y(_04476_));
 sg13g2_o21ai_1 _12039_ (.B1(net1658),
    .Y(_04477_),
    .A1(\am_sdr0.cic1.integ1[18] ),
    .A2(\am_sdr0.cic1.integ1[19] ));
 sg13g2_and2_1 _12040_ (.A(_04466_),
    .B(_04477_),
    .X(_04478_));
 sg13g2_o21ai_1 _12041_ (.B1(_04478_),
    .Y(_04479_),
    .A1(_04456_),
    .A2(_04475_));
 sg13g2_nand2_1 _12042_ (.Y(_04480_),
    .A(net1659),
    .B(\am_sdr0.cic1.integ1[20] ));
 sg13g2_xnor2_1 _12043_ (.Y(_04481_),
    .A(net1659),
    .B(\am_sdr0.cic1.integ1[20] ));
 sg13g2_nand2b_1 _12044_ (.Y(_04482_),
    .B(_04481_),
    .A_N(_04479_));
 sg13g2_nand2b_1 _12045_ (.Y(_04483_),
    .B(_04479_),
    .A_N(_04481_));
 sg13g2_and3_1 _12046_ (.X(_00810_),
    .A(net1906),
    .B(_04482_),
    .C(_04483_));
 sg13g2_xnor2_1 _12047_ (.Y(_04484_),
    .A(net1659),
    .B(net2072));
 sg13g2_nand3_1 _12048_ (.B(_04483_),
    .C(_04484_),
    .A(_04480_),
    .Y(_04485_));
 sg13g2_a21oi_1 _12049_ (.A1(_04480_),
    .A2(_04483_),
    .Y(_04486_),
    .B1(_04484_));
 sg13g2_nand2_1 _12050_ (.Y(_04487_),
    .A(net1906),
    .B(_04485_));
 sg13g2_nor2_1 _12051_ (.A(_04486_),
    .B(_04487_),
    .Y(_00811_));
 sg13g2_nand2_1 _12052_ (.Y(_04488_),
    .A(net1657),
    .B(net3238));
 sg13g2_xnor2_1 _12053_ (.Y(_04489_),
    .A(net1657),
    .B(\am_sdr0.cic1.integ1[22] ));
 sg13g2_o21ai_1 _12054_ (.B1(net1657),
    .Y(_04490_),
    .A1(\am_sdr0.cic1.integ1[20] ),
    .A2(net2072));
 sg13g2_inv_1 _12055_ (.Y(_04491_),
    .A(_04490_));
 sg13g2_nor2_1 _12056_ (.A(_04481_),
    .B(_04484_),
    .Y(_04492_));
 sg13g2_a21oi_1 _12057_ (.A1(_04479_),
    .A2(_04492_),
    .Y(_04493_),
    .B1(_04491_));
 sg13g2_or2_1 _12058_ (.X(_04494_),
    .B(_04493_),
    .A(_04489_));
 sg13g2_a21oi_1 _12059_ (.A1(_04489_),
    .A2(_04493_),
    .Y(_04495_),
    .B1(net1874));
 sg13g2_and2_1 _12060_ (.A(_04494_),
    .B(_04495_),
    .X(_00812_));
 sg13g2_xnor2_1 _12061_ (.Y(_04496_),
    .A(net1657),
    .B(net3118));
 sg13g2_and3_1 _12062_ (.X(_04497_),
    .A(_04488_),
    .B(_04494_),
    .C(_04496_));
 sg13g2_a21oi_1 _12063_ (.A1(_04488_),
    .A2(_04494_),
    .Y(_04498_),
    .B1(_04496_));
 sg13g2_nor3_1 _12064_ (.A(net1874),
    .B(_04497_),
    .C(_04498_),
    .Y(_00813_));
 sg13g2_nor4_1 _12065_ (.A(_04481_),
    .B(_04484_),
    .C(_04489_),
    .D(_04496_),
    .Y(_04499_));
 sg13g2_o21ai_1 _12066_ (.B1(net1657),
    .Y(_04500_),
    .A1(\am_sdr0.cic1.integ1[22] ),
    .A2(\am_sdr0.cic1.integ1[23] ));
 sg13g2_nand3_1 _12067_ (.B(_04490_),
    .C(net3119),
    .A(_04478_),
    .Y(_04501_));
 sg13g2_a21oi_1 _12068_ (.A1(_04476_),
    .A2(_04499_),
    .Y(_04502_),
    .B1(_04501_));
 sg13g2_nand2_1 _12069_ (.Y(_04503_),
    .A(net1657),
    .B(net3034));
 sg13g2_xnor2_1 _12070_ (.Y(_04504_),
    .A(net1657),
    .B(net3034));
 sg13g2_or2_1 _12071_ (.X(_04505_),
    .B(_04504_),
    .A(_04502_));
 sg13g2_nand2_1 _12072_ (.Y(_04506_),
    .A(net1896),
    .B(_04505_));
 sg13g2_a21oi_1 _12073_ (.A1(_04502_),
    .A2(_04504_),
    .Y(_00814_),
    .B1(_04506_));
 sg13g2_xnor2_1 _12074_ (.Y(_04507_),
    .A(net1657),
    .B(net3042));
 sg13g2_and3_1 _12075_ (.X(_04508_),
    .A(_04503_),
    .B(_04505_),
    .C(_04507_));
 sg13g2_a21oi_1 _12076_ (.A1(_04503_),
    .A2(_04505_),
    .Y(_04509_),
    .B1(_04507_));
 sg13g2_nor3_1 _12077_ (.A(net1874),
    .B(_04508_),
    .C(_04509_),
    .Y(_00815_));
 sg13g2_nand2_1 _12078_ (.Y(_04510_),
    .A(\am_sdr0.cic1.integ1[3] ),
    .B(net2196));
 sg13g2_o21ai_1 _12079_ (.B1(net1903),
    .Y(_04511_),
    .A1(\am_sdr0.cic1.integ1[3] ),
    .A2(net2196));
 sg13g2_nor2b_1 _12080_ (.A(net2197),
    .B_N(_04510_),
    .Y(_00816_));
 sg13g2_nand2_1 _12081_ (.Y(_04512_),
    .A(\am_sdr0.cic1.integ1[4] ),
    .B(net2941));
 sg13g2_xnor2_1 _12082_ (.Y(_04513_),
    .A(\am_sdr0.cic1.integ1[4] ),
    .B(net2941));
 sg13g2_o21ai_1 _12083_ (.B1(net1901),
    .Y(_04514_),
    .A1(_04510_),
    .A2(_04513_));
 sg13g2_a21oi_1 _12084_ (.A1(_04510_),
    .A2(net2942),
    .Y(_00817_),
    .B1(_04514_));
 sg13g2_and2_1 _12085_ (.A(\am_sdr0.cic1.integ1[5] ),
    .B(net3175),
    .X(_04515_));
 sg13g2_xor2_1 _12086_ (.B(net3175),
    .A(net3216),
    .X(_04516_));
 sg13g2_o21ai_1 _12087_ (.B1(_04512_),
    .Y(_04517_),
    .A1(_04510_),
    .A2(_04513_));
 sg13g2_nor2_1 _12088_ (.A(_04516_),
    .B(_04517_),
    .Y(_04518_));
 sg13g2_a21oi_1 _12089_ (.A1(_04516_),
    .A2(_04517_),
    .Y(_04519_),
    .B1(net1877));
 sg13g2_nor2b_1 _12090_ (.A(_04518_),
    .B_N(_04519_),
    .Y(_00818_));
 sg13g2_nand2_1 _12091_ (.Y(_04520_),
    .A(\am_sdr0.cic1.integ2[3] ),
    .B(\am_sdr0.cic1.integ1[6] ));
 sg13g2_xnor2_1 _12092_ (.Y(_04521_),
    .A(net2588),
    .B(\am_sdr0.cic1.integ1[6] ));
 sg13g2_a21oi_2 _12093_ (.B1(net3176),
    .Y(_04522_),
    .A2(_04517_),
    .A1(_04516_));
 sg13g2_o21ai_1 _12094_ (.B1(net1904),
    .Y(_04523_),
    .A1(_04521_),
    .A2(_04522_));
 sg13g2_a21oi_1 _12095_ (.A1(_04521_),
    .A2(_04522_),
    .Y(_00819_),
    .B1(_04523_));
 sg13g2_and2_1 _12096_ (.A(\am_sdr0.cic1.integ1[7] ),
    .B(net2976),
    .X(_04524_));
 sg13g2_xor2_1 _12097_ (.B(\am_sdr0.cic1.integ2[4] ),
    .A(\am_sdr0.cic1.integ1[7] ),
    .X(_04525_));
 sg13g2_o21ai_1 _12098_ (.B1(_04520_),
    .Y(_04526_),
    .A1(_04521_),
    .A2(_04522_));
 sg13g2_or2_1 _12099_ (.X(_04527_),
    .B(_04526_),
    .A(_04525_));
 sg13g2_a21oi_1 _12100_ (.A1(_04525_),
    .A2(_04526_),
    .Y(_04528_),
    .B1(net1876));
 sg13g2_and2_1 _12101_ (.A(_04527_),
    .B(_04528_),
    .X(_00820_));
 sg13g2_a21oi_1 _12102_ (.A1(_04525_),
    .A2(_04526_),
    .Y(_04529_),
    .B1(_04524_));
 sg13g2_nor2_1 _12103_ (.A(\am_sdr0.cic1.integ1[8] ),
    .B(net3292),
    .Y(_04530_));
 sg13g2_xnor2_1 _12104_ (.Y(_04531_),
    .A(\am_sdr0.cic1.integ1[8] ),
    .B(net3169));
 sg13g2_o21ai_1 _12105_ (.B1(net1902),
    .Y(_04532_),
    .A1(_04529_),
    .A2(_04531_));
 sg13g2_a21oi_1 _12106_ (.A1(_04529_),
    .A2(net3170),
    .Y(_00821_),
    .B1(_04532_));
 sg13g2_and2_1 _12107_ (.A(net3283),
    .B(net3130),
    .X(_04533_));
 sg13g2_xnor2_1 _12108_ (.Y(_04534_),
    .A(net3283),
    .B(net3130));
 sg13g2_a221oi_1 _12109_ (.B2(_04526_),
    .C1(_04524_),
    .B1(_04525_),
    .A1(\am_sdr0.cic1.integ1[8] ),
    .Y(_04535_),
    .A2(\am_sdr0.cic1.integ2[5] ));
 sg13g2_o21ai_1 _12110_ (.B1(_04534_),
    .Y(_04536_),
    .A1(_04530_),
    .A2(_04535_));
 sg13g2_nor3_2 _12111_ (.A(_04530_),
    .B(_04534_),
    .C(_04535_),
    .Y(_04537_));
 sg13g2_nand2_1 _12112_ (.Y(_04538_),
    .A(net1902),
    .B(_04536_));
 sg13g2_nor2_1 _12113_ (.A(_04537_),
    .B(_04538_),
    .Y(_00822_));
 sg13g2_nand2_1 _12114_ (.Y(_04539_),
    .A(\am_sdr0.cic1.integ1[10] ),
    .B(\am_sdr0.cic1.integ2[7] ));
 sg13g2_xor2_1 _12115_ (.B(\am_sdr0.cic1.integ2[7] ),
    .A(\am_sdr0.cic1.integ1[10] ),
    .X(_04540_));
 sg13g2_nor3_1 _12116_ (.A(_04533_),
    .B(_04537_),
    .C(_04540_),
    .Y(_04541_));
 sg13g2_o21ai_1 _12117_ (.B1(_04540_),
    .Y(_04542_),
    .A1(_04533_),
    .A2(_04537_));
 sg13g2_nand2_1 _12118_ (.Y(_04543_),
    .A(net1902),
    .B(_04542_));
 sg13g2_nor2_1 _12119_ (.A(net3284),
    .B(_04543_),
    .Y(_00823_));
 sg13g2_nand2_1 _12120_ (.Y(_04544_),
    .A(_04539_),
    .B(_04542_));
 sg13g2_nand2_1 _12121_ (.Y(_04545_),
    .A(net3237),
    .B(net3105));
 sg13g2_xor2_1 _12122_ (.B(net3290),
    .A(net3237),
    .X(_04546_));
 sg13g2_inv_1 _12123_ (.Y(_04547_),
    .A(_04546_));
 sg13g2_nand2_1 _12124_ (.Y(_04548_),
    .A(_04544_),
    .B(_04546_));
 sg13g2_o21ai_1 _12125_ (.B1(net1902),
    .Y(_04549_),
    .A1(_04544_),
    .A2(_04546_));
 sg13g2_nor2b_1 _12126_ (.A(_04549_),
    .B_N(_04548_),
    .Y(_00824_));
 sg13g2_nor2_1 _12127_ (.A(\am_sdr0.cic1.integ1[12] ),
    .B(net3243),
    .Y(_04550_));
 sg13g2_nand2_1 _12128_ (.Y(_04551_),
    .A(net3218),
    .B(net3243));
 sg13g2_nand2b_1 _12129_ (.Y(_04552_),
    .B(_04551_),
    .A_N(_04550_));
 sg13g2_and2_1 _12130_ (.A(_04545_),
    .B(_04548_),
    .X(_04553_));
 sg13g2_o21ai_1 _12131_ (.B1(net1902),
    .Y(_04554_),
    .A1(_04552_),
    .A2(_04553_));
 sg13g2_a21oi_1 _12132_ (.A1(net3244),
    .A2(_04553_),
    .Y(_00825_),
    .B1(_04554_));
 sg13g2_nand2_1 _12133_ (.Y(_04555_),
    .A(net3257),
    .B(net3250));
 sg13g2_xnor2_1 _12134_ (.Y(_04556_),
    .A(\am_sdr0.cic1.integ1[13] ),
    .B(\am_sdr0.cic1.integ2[10] ));
 sg13g2_nor2_1 _12135_ (.A(_04547_),
    .B(_04552_),
    .Y(_04557_));
 sg13g2_o21ai_1 _12136_ (.B1(_04551_),
    .Y(_04558_),
    .A1(_04545_),
    .A2(_04550_));
 sg13g2_a21oi_1 _12137_ (.A1(_04544_),
    .A2(_04557_),
    .Y(_04559_),
    .B1(_04558_));
 sg13g2_or2_1 _12138_ (.X(_04560_),
    .B(_04559_),
    .A(_04556_));
 sg13g2_a21oi_1 _12139_ (.A1(_04556_),
    .A2(_04559_),
    .Y(_04561_),
    .B1(net1874));
 sg13g2_and2_1 _12140_ (.A(_04560_),
    .B(_04561_),
    .X(_00826_));
 sg13g2_nor2_1 _12141_ (.A(\am_sdr0.cic1.integ1[14] ),
    .B(\am_sdr0.cic1.integ2[11] ),
    .Y(_04562_));
 sg13g2_xnor2_1 _12142_ (.Y(_04563_),
    .A(\am_sdr0.cic1.integ1[14] ),
    .B(net3227));
 sg13g2_and3_1 _12143_ (.X(_04564_),
    .A(_04555_),
    .B(_04560_),
    .C(_04563_));
 sg13g2_a21oi_1 _12144_ (.A1(_04555_),
    .A2(_04560_),
    .Y(_04565_),
    .B1(_04563_));
 sg13g2_nor3_1 _12145_ (.A(net1874),
    .B(_04564_),
    .C(_04565_),
    .Y(_00827_));
 sg13g2_nand2_1 _12146_ (.Y(_04566_),
    .A(\am_sdr0.cic1.integ1[15] ),
    .B(net3234));
 sg13g2_xor2_1 _12147_ (.B(\am_sdr0.cic1.integ2[12] ),
    .A(\am_sdr0.cic1.integ1[15] ),
    .X(_04567_));
 sg13g2_inv_1 _12148_ (.Y(_04568_),
    .A(_04567_));
 sg13g2_nor2_1 _12149_ (.A(_04556_),
    .B(_04563_),
    .Y(_04569_));
 sg13g2_nor2_1 _12150_ (.A(_04555_),
    .B(_04562_),
    .Y(_04570_));
 sg13g2_a221oi_1 _12151_ (.B2(_04569_),
    .C1(_04570_),
    .B1(_04558_),
    .A1(\am_sdr0.cic1.integ1[14] ),
    .Y(_04571_),
    .A2(\am_sdr0.cic1.integ2[11] ));
 sg13g2_inv_1 _12152_ (.Y(_04572_),
    .A(_04571_));
 sg13g2_nand2_1 _12153_ (.Y(_04573_),
    .A(_04557_),
    .B(_04569_));
 sg13g2_a21oi_2 _12154_ (.B1(_04573_),
    .Y(_04574_),
    .A2(_04542_),
    .A1(_04539_));
 sg13g2_nor3_1 _12155_ (.A(_04567_),
    .B(_04572_),
    .C(_04574_),
    .Y(_04575_));
 sg13g2_o21ai_1 _12156_ (.B1(_04567_),
    .Y(_04576_),
    .A1(_04572_),
    .A2(_04574_));
 sg13g2_nand2_1 _12157_ (.Y(_04577_),
    .A(net1898),
    .B(_04576_));
 sg13g2_nor2_1 _12158_ (.A(_04575_),
    .B(_04577_),
    .Y(_00828_));
 sg13g2_nor2_1 _12159_ (.A(\am_sdr0.cic1.integ1[16] ),
    .B(net3280),
    .Y(_04578_));
 sg13g2_xnor2_1 _12160_ (.Y(_04579_),
    .A(\am_sdr0.cic1.integ1[16] ),
    .B(\am_sdr0.cic1.integ2[13] ));
 sg13g2_and3_1 _12161_ (.X(_04580_),
    .A(net3235),
    .B(_04576_),
    .C(_04579_));
 sg13g2_a21oi_1 _12162_ (.A1(net3235),
    .A2(_04576_),
    .Y(_04581_),
    .B1(_04579_));
 sg13g2_nor3_1 _12163_ (.A(net1875),
    .B(_04580_),
    .C(net3236),
    .Y(_00829_));
 sg13g2_nand2_1 _12164_ (.Y(_04582_),
    .A(net3264),
    .B(net3212));
 sg13g2_xnor2_1 _12165_ (.Y(_04583_),
    .A(net3264),
    .B(net3212));
 sg13g2_a22oi_1 _12166_ (.Y(_04584_),
    .B1(\am_sdr0.cic1.integ2[13] ),
    .B2(\am_sdr0.cic1.integ1[16] ),
    .A2(\am_sdr0.cic1.integ2[12] ),
    .A1(\am_sdr0.cic1.integ1[15] ));
 sg13g2_a21o_1 _12167_ (.A2(_04584_),
    .A1(_04576_),
    .B1(_04578_),
    .X(_04585_));
 sg13g2_or2_1 _12168_ (.X(_04586_),
    .B(_04585_),
    .A(_04583_));
 sg13g2_nand2_1 _12169_ (.Y(_04587_),
    .A(net1898),
    .B(_04586_));
 sg13g2_a21oi_1 _12170_ (.A1(_04583_),
    .A2(_04585_),
    .Y(_00830_),
    .B1(_04587_));
 sg13g2_nor2_1 _12171_ (.A(\am_sdr0.cic1.integ1[18] ),
    .B(\am_sdr0.cic1.integ2[15] ),
    .Y(_04588_));
 sg13g2_xnor2_1 _12172_ (.Y(_04589_),
    .A(\am_sdr0.cic1.integ1[18] ),
    .B(net3273));
 sg13g2_and3_1 _12173_ (.X(_04590_),
    .A(_04582_),
    .B(_04586_),
    .C(_04589_));
 sg13g2_a21oi_1 _12174_ (.A1(_04582_),
    .A2(_04586_),
    .Y(_04591_),
    .B1(_04589_));
 sg13g2_nor3_1 _12175_ (.A(net1874),
    .B(_04590_),
    .C(_04591_),
    .Y(_00831_));
 sg13g2_xnor2_1 _12176_ (.Y(_04592_),
    .A(\am_sdr0.cic1.integ1[19] ),
    .B(\am_sdr0.cic1.integ2[16] ));
 sg13g2_nor4_2 _12177_ (.A(_04568_),
    .B(_04579_),
    .C(_04583_),
    .Y(_04593_),
    .D(_04589_));
 sg13g2_nor2_1 _12178_ (.A(_04582_),
    .B(_04588_),
    .Y(_04594_));
 sg13g2_a21oi_1 _12179_ (.A1(\am_sdr0.cic1.integ1[18] ),
    .A2(\am_sdr0.cic1.integ2[15] ),
    .Y(_04595_),
    .B1(_04594_));
 sg13g2_nor4_1 _12180_ (.A(_04578_),
    .B(_04583_),
    .C(_04584_),
    .D(_04589_),
    .Y(_04596_));
 sg13g2_a21oi_1 _12181_ (.A1(_04572_),
    .A2(_04593_),
    .Y(_04597_),
    .B1(_04596_));
 sg13g2_nand2_1 _12182_ (.Y(_04598_),
    .A(_04595_),
    .B(_04597_));
 sg13g2_a21oi_2 _12183_ (.B1(_04598_),
    .Y(_04599_),
    .A2(_04593_),
    .A1(_04574_));
 sg13g2_nor2_1 _12184_ (.A(_04592_),
    .B(_04599_),
    .Y(_04600_));
 sg13g2_a21oi_1 _12185_ (.A1(_04592_),
    .A2(_04599_),
    .Y(_04601_),
    .B1(net1874));
 sg13g2_nor2b_1 _12186_ (.A(_04600_),
    .B_N(_04601_),
    .Y(_00832_));
 sg13g2_nor2_1 _12187_ (.A(\am_sdr0.cic1.integ1[20] ),
    .B(\am_sdr0.cic1.integ2[17] ),
    .Y(_04602_));
 sg13g2_xnor2_1 _12188_ (.Y(_04603_),
    .A(\am_sdr0.cic1.integ1[20] ),
    .B(\am_sdr0.cic1.integ2[17] ));
 sg13g2_a21oi_1 _12189_ (.A1(net3165),
    .A2(\am_sdr0.cic1.integ2[16] ),
    .Y(_04604_),
    .B1(_04600_));
 sg13g2_o21ai_1 _12190_ (.B1(net1896),
    .Y(_04605_),
    .A1(_04603_),
    .A2(net3166));
 sg13g2_a21oi_1 _12191_ (.A1(_04603_),
    .A2(net3166),
    .Y(_00833_),
    .B1(_04605_));
 sg13g2_and2_1 _12192_ (.A(net2072),
    .B(\am_sdr0.cic1.integ2[18] ),
    .X(_04606_));
 sg13g2_or2_1 _12193_ (.X(_04607_),
    .B(\am_sdr0.cic1.integ2[18] ),
    .A(net2072));
 sg13g2_nand2b_1 _12194_ (.Y(_04608_),
    .B(_04607_),
    .A_N(_04606_));
 sg13g2_nor2_1 _12195_ (.A(_04592_),
    .B(_04603_),
    .Y(_04609_));
 sg13g2_inv_1 _12196_ (.Y(_04610_),
    .A(_04609_));
 sg13g2_a22oi_1 _12197_ (.Y(_04611_),
    .B1(\am_sdr0.cic1.integ2[17] ),
    .B2(\am_sdr0.cic1.integ1[20] ),
    .A2(\am_sdr0.cic1.integ2[16] ),
    .A1(\am_sdr0.cic1.integ1[19] ));
 sg13g2_nor2_1 _12198_ (.A(_04602_),
    .B(_04611_),
    .Y(_04612_));
 sg13g2_inv_1 _12199_ (.Y(_04613_),
    .A(_04612_));
 sg13g2_o21ai_1 _12200_ (.B1(_04613_),
    .Y(_04614_),
    .A1(_04599_),
    .A2(_04610_));
 sg13g2_inv_1 _12201_ (.Y(_04615_),
    .A(_04614_));
 sg13g2_o21ai_1 _12202_ (.B1(net1896),
    .Y(_04616_),
    .A1(_04608_),
    .A2(_04615_));
 sg13g2_a21oi_1 _12203_ (.A1(_04608_),
    .A2(_04615_),
    .Y(_00834_),
    .B1(_04616_));
 sg13g2_and2_1 _12204_ (.A(\am_sdr0.cic1.integ1[22] ),
    .B(\am_sdr0.cic1.integ2[19] ),
    .X(_04617_));
 sg13g2_or2_1 _12205_ (.X(_04618_),
    .B(net3295),
    .A(\am_sdr0.cic1.integ1[22] ));
 sg13g2_nand2b_1 _12206_ (.Y(_04619_),
    .B(_04618_),
    .A_N(_04617_));
 sg13g2_a21oi_1 _12207_ (.A1(_04607_),
    .A2(_04614_),
    .Y(_04620_),
    .B1(net2073));
 sg13g2_o21ai_1 _12208_ (.B1(net1896),
    .Y(_04621_),
    .A1(_04619_),
    .A2(_04620_));
 sg13g2_a21oi_1 _12209_ (.A1(_04619_),
    .A2(_04620_),
    .Y(_00835_),
    .B1(_04621_));
 sg13g2_nor2_1 _12210_ (.A(_04608_),
    .B(_04619_),
    .Y(_04622_));
 sg13g2_nand2_1 _12211_ (.Y(_04623_),
    .A(_04609_),
    .B(_04622_));
 sg13g2_a221oi_1 _12212_ (.B2(_04612_),
    .C1(_04617_),
    .B1(_04622_),
    .A1(_04606_),
    .Y(_04624_),
    .A2(_04618_));
 sg13g2_o21ai_1 _12213_ (.B1(_04624_),
    .Y(_04625_),
    .A1(_04599_),
    .A2(_04623_));
 sg13g2_and2_1 _12214_ (.A(net3118),
    .B(\am_sdr0.cic1.integ2[20] ),
    .X(_04626_));
 sg13g2_xnor2_1 _12215_ (.Y(_04627_),
    .A(net3118),
    .B(\am_sdr0.cic1.integ2[20] ));
 sg13g2_inv_1 _12216_ (.Y(_04628_),
    .A(_04627_));
 sg13g2_o21ai_1 _12217_ (.B1(net1896),
    .Y(_04629_),
    .A1(_04625_),
    .A2(_04628_));
 sg13g2_a21oi_1 _12218_ (.A1(_04625_),
    .A2(_04628_),
    .Y(_00836_),
    .B1(_04629_));
 sg13g2_or2_1 _12219_ (.X(_04630_),
    .B(\am_sdr0.cic1.integ2[21] ),
    .A(\am_sdr0.cic1.integ1[24] ));
 sg13g2_and2_1 _12220_ (.A(\am_sdr0.cic1.integ1[24] ),
    .B(\am_sdr0.cic1.integ2[21] ),
    .X(_04631_));
 sg13g2_xnor2_1 _12221_ (.Y(_04632_),
    .A(net3034),
    .B(net3245));
 sg13g2_a21oi_1 _12222_ (.A1(_04625_),
    .A2(_04628_),
    .Y(_04633_),
    .B1(_04626_));
 sg13g2_o21ai_1 _12223_ (.B1(net1896),
    .Y(_04634_),
    .A1(_04632_),
    .A2(_04633_));
 sg13g2_a21oi_1 _12224_ (.A1(_04632_),
    .A2(_04633_),
    .Y(_00837_),
    .B1(_04634_));
 sg13g2_nor2_1 _12225_ (.A(_04627_),
    .B(_04632_),
    .Y(_04635_));
 sg13g2_a221oi_1 _12226_ (.B2(_04625_),
    .C1(_04631_),
    .B1(_04635_),
    .A1(_04626_),
    .Y(_04636_),
    .A2(_04630_));
 sg13g2_xnor2_1 _12227_ (.Y(_04637_),
    .A(net3042),
    .B(net2982));
 sg13g2_o21ai_1 _12228_ (.B1(net1896),
    .Y(_04638_),
    .A1(_04636_),
    .A2(_04637_));
 sg13g2_a21oi_1 _12229_ (.A1(_04636_),
    .A2(_04637_),
    .Y(_00838_),
    .B1(_04638_));
 sg13g2_nand2_1 _12230_ (.Y(_04639_),
    .A(net2756),
    .B(net2523));
 sg13g2_o21ai_1 _12231_ (.B1(net1937),
    .Y(_04640_),
    .A1(net2756),
    .A2(net2523));
 sg13g2_nor2b_1 _12232_ (.A(_04640_),
    .B_N(_04639_),
    .Y(_00840_));
 sg13g2_nand2_1 _12233_ (.Y(_04641_),
    .A(net2990),
    .B(net2290));
 sg13g2_xnor2_1 _12234_ (.Y(_04642_),
    .A(net2990),
    .B(net2290));
 sg13g2_o21ai_1 _12235_ (.B1(net1937),
    .Y(_04643_),
    .A1(_04639_),
    .A2(_04642_));
 sg13g2_a21oi_1 _12236_ (.A1(_04639_),
    .A2(_04642_),
    .Y(_00841_),
    .B1(_04643_));
 sg13g2_and2_1 _12237_ (.A(\am_sdr0.cic0.integ2[5] ),
    .B(net1499),
    .X(_04644_));
 sg13g2_xor2_1 _12238_ (.B(net1499),
    .A(net3181),
    .X(_04645_));
 sg13g2_o21ai_1 _12239_ (.B1(_04641_),
    .Y(_04646_),
    .A1(_04639_),
    .A2(_04642_));
 sg13g2_nor2_1 _12240_ (.A(_04645_),
    .B(_04646_),
    .Y(_04647_));
 sg13g2_a21oi_1 _12241_ (.A1(_04645_),
    .A2(_04646_),
    .Y(_04648_),
    .B1(net1884));
 sg13g2_nor2b_1 _12242_ (.A(_04647_),
    .B_N(_04648_),
    .Y(_00842_));
 sg13g2_nand2_1 _12243_ (.Y(_04649_),
    .A(\am_sdr0.cic0.integ2[6] ),
    .B(\am_sdr0.cic0.integ3[3] ));
 sg13g2_xnor2_1 _12244_ (.Y(_04650_),
    .A(net3142),
    .B(net1433));
 sg13g2_a21oi_1 _12245_ (.A1(_04645_),
    .A2(_04646_),
    .Y(_04651_),
    .B1(_04644_));
 sg13g2_o21ai_1 _12246_ (.B1(net1950),
    .Y(_04652_),
    .A1(_04650_),
    .A2(_04651_));
 sg13g2_a21oi_1 _12247_ (.A1(_04650_),
    .A2(_04651_),
    .Y(_00843_),
    .B1(_04652_));
 sg13g2_and2_1 _12248_ (.A(\am_sdr0.cic0.integ2[7] ),
    .B(net1501),
    .X(_04653_));
 sg13g2_xor2_1 _12249_ (.B(\am_sdr0.cic0.integ3[4] ),
    .A(\am_sdr0.cic0.integ2[7] ),
    .X(_04654_));
 sg13g2_o21ai_1 _12250_ (.B1(_04649_),
    .Y(_04655_),
    .A1(_04650_),
    .A2(_04651_));
 sg13g2_or2_1 _12251_ (.X(_04656_),
    .B(_04655_),
    .A(_04654_));
 sg13g2_a21oi_1 _12252_ (.A1(_04654_),
    .A2(_04655_),
    .Y(_04657_),
    .B1(net1884));
 sg13g2_and2_1 _12253_ (.A(_04656_),
    .B(_04657_),
    .X(_00844_));
 sg13g2_a21oi_1 _12254_ (.A1(_04654_),
    .A2(_04655_),
    .Y(_04658_),
    .B1(_04653_));
 sg13g2_nor2_1 _12255_ (.A(\am_sdr0.cic0.integ2[8] ),
    .B(net3268),
    .Y(_04659_));
 sg13g2_xnor2_1 _12256_ (.Y(_04660_),
    .A(net3099),
    .B(net2052));
 sg13g2_o21ai_1 _12257_ (.B1(net1950),
    .Y(_04661_),
    .A1(_04658_),
    .A2(_04660_));
 sg13g2_a21oi_1 _12258_ (.A1(_04658_),
    .A2(_04660_),
    .Y(_00845_),
    .B1(_04661_));
 sg13g2_and2_1 _12259_ (.A(net3231),
    .B(net1400),
    .X(_04662_));
 sg13g2_xnor2_1 _12260_ (.Y(_04663_),
    .A(net3231),
    .B(net1400));
 sg13g2_a221oi_1 _12261_ (.B2(_04655_),
    .C1(_04653_),
    .B1(_04654_),
    .A1(\am_sdr0.cic0.integ2[8] ),
    .Y(_04664_),
    .A2(\am_sdr0.cic0.integ3[5] ));
 sg13g2_o21ai_1 _12262_ (.B1(_04663_),
    .Y(_04665_),
    .A1(_04659_),
    .A2(_04664_));
 sg13g2_nor3_2 _12263_ (.A(_04659_),
    .B(_04663_),
    .C(_04664_),
    .Y(_04666_));
 sg13g2_nand2_1 _12264_ (.Y(_04667_),
    .A(net1950),
    .B(_04665_));
 sg13g2_nor2_1 _12265_ (.A(_04666_),
    .B(_04667_),
    .Y(_00846_));
 sg13g2_nand2_2 _12266_ (.Y(_04668_),
    .A(\am_sdr0.cic0.integ2[10] ),
    .B(net3306));
 sg13g2_xor2_1 _12267_ (.B(net2055),
    .A(\am_sdr0.cic0.integ2[10] ),
    .X(_04669_));
 sg13g2_nor3_1 _12268_ (.A(_04662_),
    .B(_04666_),
    .C(net3256),
    .Y(_04670_));
 sg13g2_o21ai_1 _12269_ (.B1(_04669_),
    .Y(_04671_),
    .A1(_04662_),
    .A2(_04666_));
 sg13g2_nand2_1 _12270_ (.Y(_04672_),
    .A(net1942),
    .B(_04671_));
 sg13g2_nor2_1 _12271_ (.A(_04670_),
    .B(_04672_),
    .Y(_00847_));
 sg13g2_nand2_1 _12272_ (.Y(_04673_),
    .A(_04668_),
    .B(_04671_));
 sg13g2_nand2_1 _12273_ (.Y(_04674_),
    .A(\am_sdr0.cic0.integ2[11] ),
    .B(net1437));
 sg13g2_xor2_1 _12274_ (.B(net1437),
    .A(\am_sdr0.cic0.integ2[11] ),
    .X(_04675_));
 sg13g2_inv_1 _12275_ (.Y(_04676_),
    .A(_04675_));
 sg13g2_nand2_1 _12276_ (.Y(_04677_),
    .A(_04673_),
    .B(_04675_));
 sg13g2_o21ai_1 _12277_ (.B1(net1942),
    .Y(_04678_),
    .A1(_04673_),
    .A2(net3263));
 sg13g2_nor2b_1 _12278_ (.A(_04678_),
    .B_N(_04677_),
    .Y(_00848_));
 sg13g2_nor2_1 _12279_ (.A(\am_sdr0.cic0.integ2[12] ),
    .B(net1443),
    .Y(_04679_));
 sg13g2_nand2_1 _12280_ (.Y(_04680_),
    .A(net3207),
    .B(net1443));
 sg13g2_nand2b_1 _12281_ (.Y(_04681_),
    .B(_04680_),
    .A_N(_04679_));
 sg13g2_and2_1 _12282_ (.A(_04674_),
    .B(_04677_),
    .X(_04682_));
 sg13g2_o21ai_1 _12283_ (.B1(net1942),
    .Y(_04683_),
    .A1(_04681_),
    .A2(_04682_));
 sg13g2_a21oi_1 _12284_ (.A1(net3208),
    .A2(_04682_),
    .Y(_00849_),
    .B1(_04683_));
 sg13g2_nand2_1 _12285_ (.Y(_04684_),
    .A(net3126),
    .B(net1512));
 sg13g2_xnor2_1 _12286_ (.Y(_04685_),
    .A(net3126),
    .B(net1512));
 sg13g2_o21ai_1 _12287_ (.B1(_04680_),
    .Y(_04686_),
    .A1(_04674_),
    .A2(_04679_));
 sg13g2_nor2_1 _12288_ (.A(_04676_),
    .B(_04681_),
    .Y(_04687_));
 sg13g2_a21oi_1 _12289_ (.A1(_04673_),
    .A2(_04687_),
    .Y(_04688_),
    .B1(_04686_));
 sg13g2_or2_1 _12290_ (.X(_04689_),
    .B(_04688_),
    .A(_04685_));
 sg13g2_nand2_1 _12291_ (.Y(_04690_),
    .A(net1942),
    .B(_04689_));
 sg13g2_a21oi_1 _12292_ (.A1(_04685_),
    .A2(_04688_),
    .Y(_00850_),
    .B1(_04690_));
 sg13g2_nor2_1 _12293_ (.A(\am_sdr0.cic0.integ2[14] ),
    .B(\am_sdr0.cic0.integ3[11] ),
    .Y(_04691_));
 sg13g2_xnor2_1 _12294_ (.Y(_04692_),
    .A(net3215),
    .B(net2240));
 sg13g2_and3_1 _12295_ (.X(_04693_),
    .A(_04684_),
    .B(_04689_),
    .C(_04692_));
 sg13g2_a21oi_1 _12296_ (.A1(_04684_),
    .A2(_04689_),
    .Y(_04694_),
    .B1(_04692_));
 sg13g2_nor3_1 _12297_ (.A(net1886),
    .B(_04693_),
    .C(_04694_),
    .Y(_00851_));
 sg13g2_nand2_1 _12298_ (.Y(_04695_),
    .A(net3179),
    .B(net2267));
 sg13g2_xor2_1 _12299_ (.B(\am_sdr0.cic0.integ3[12] ),
    .A(\am_sdr0.cic0.integ2[15] ),
    .X(_04696_));
 sg13g2_nor2_1 _12300_ (.A(_04685_),
    .B(_04692_),
    .Y(_04697_));
 sg13g2_nor2_1 _12301_ (.A(_04684_),
    .B(_04691_),
    .Y(_04698_));
 sg13g2_a221oi_1 _12302_ (.B2(_04697_),
    .C1(_04698_),
    .B1(_04686_),
    .A1(\am_sdr0.cic0.integ2[14] ),
    .Y(_04699_),
    .A2(\am_sdr0.cic0.integ3[11] ));
 sg13g2_inv_1 _12303_ (.Y(_04700_),
    .A(_04699_));
 sg13g2_and2_1 _12304_ (.A(_04687_),
    .B(_04697_),
    .X(_04701_));
 sg13g2_inv_1 _12305_ (.Y(_04702_),
    .A(_04701_));
 sg13g2_a21oi_1 _12306_ (.A1(_04668_),
    .A2(_04671_),
    .Y(_04703_),
    .B1(_04702_));
 sg13g2_nor3_1 _12307_ (.A(_04696_),
    .B(_04700_),
    .C(_04703_),
    .Y(_04704_));
 sg13g2_o21ai_1 _12308_ (.B1(_04696_),
    .Y(_04705_),
    .A1(_04700_),
    .A2(_04703_));
 sg13g2_nand2_1 _12309_ (.Y(_04706_),
    .A(net1940),
    .B(_04705_));
 sg13g2_nor2_1 _12310_ (.A(_04704_),
    .B(_04706_),
    .Y(_00852_));
 sg13g2_nor2_1 _12311_ (.A(\am_sdr0.cic0.integ2[16] ),
    .B(\am_sdr0.cic0.integ3[13] ),
    .Y(_04707_));
 sg13g2_xor2_1 _12312_ (.B(net2205),
    .A(\am_sdr0.cic0.integ2[16] ),
    .X(_04708_));
 sg13g2_nand2_1 _12313_ (.Y(_04709_),
    .A(_04695_),
    .B(_04705_));
 sg13g2_o21ai_1 _12314_ (.B1(net1940),
    .Y(_04710_),
    .A1(_04708_),
    .A2(_04709_));
 sg13g2_a21oi_1 _12315_ (.A1(_04708_),
    .A2(_04709_),
    .Y(_00853_),
    .B1(_04710_));
 sg13g2_and2_1 _12316_ (.A(\am_sdr0.cic0.integ2[17] ),
    .B(net3316),
    .X(_04711_));
 sg13g2_xnor2_1 _12317_ (.Y(_04712_),
    .A(\am_sdr0.cic0.integ2[17] ),
    .B(net2109));
 sg13g2_a22oi_1 _12318_ (.Y(_04713_),
    .B1(\am_sdr0.cic0.integ3[13] ),
    .B2(\am_sdr0.cic0.integ2[16] ),
    .A2(\am_sdr0.cic0.integ3[12] ),
    .A1(\am_sdr0.cic0.integ2[15] ));
 sg13g2_nand2_1 _12319_ (.Y(_04714_),
    .A(_04696_),
    .B(_04708_));
 sg13g2_a21o_1 _12320_ (.A2(_04713_),
    .A1(_04705_),
    .B1(_04707_),
    .X(_04715_));
 sg13g2_nor2_1 _12321_ (.A(_04712_),
    .B(_04715_),
    .Y(_04716_));
 sg13g2_a21oi_1 _12322_ (.A1(_04712_),
    .A2(_04715_),
    .Y(_04717_),
    .B1(net1886));
 sg13g2_nor2b_1 _12323_ (.A(_04716_),
    .B_N(_04717_),
    .Y(_00854_));
 sg13g2_nand2_1 _12324_ (.Y(_04718_),
    .A(\am_sdr0.cic0.integ2[18] ),
    .B(\am_sdr0.cic0.integ3[15] ));
 sg13g2_xor2_1 _12325_ (.B(\am_sdr0.cic0.integ3[15] ),
    .A(\am_sdr0.cic0.integ2[18] ),
    .X(_04719_));
 sg13g2_or3_1 _12326_ (.A(_04711_),
    .B(_04716_),
    .C(_04719_),
    .X(_04720_));
 sg13g2_o21ai_1 _12327_ (.B1(_04719_),
    .Y(_04721_),
    .A1(_04711_),
    .A2(_04716_));
 sg13g2_and3_1 _12328_ (.X(_00855_),
    .A(net1940),
    .B(_04720_),
    .C(_04721_));
 sg13g2_nand2_1 _12329_ (.Y(_04722_),
    .A(net3093),
    .B(net1518));
 sg13g2_xnor2_1 _12330_ (.Y(_04723_),
    .A(net3093),
    .B(net1518));
 sg13g2_inv_1 _12331_ (.Y(_04724_),
    .A(_04723_));
 sg13g2_nand2b_1 _12332_ (.Y(_04725_),
    .B(_04719_),
    .A_N(_04712_));
 sg13g2_nor2_1 _12333_ (.A(_04714_),
    .B(_04725_),
    .Y(_04726_));
 sg13g2_o21ai_1 _12334_ (.B1(_04711_),
    .Y(_04727_),
    .A1(\am_sdr0.cic0.integ2[18] ),
    .A2(\am_sdr0.cic0.integ3[15] ));
 sg13g2_nor3_1 _12335_ (.A(_04707_),
    .B(_04713_),
    .C(_04725_),
    .Y(_04728_));
 sg13g2_a21oi_1 _12336_ (.A1(_04700_),
    .A2(_04726_),
    .Y(_04729_),
    .B1(_04728_));
 sg13g2_nand3_1 _12337_ (.B(_04727_),
    .C(_04729_),
    .A(_04718_),
    .Y(_04730_));
 sg13g2_nand2_1 _12338_ (.Y(_04731_),
    .A(_04701_),
    .B(_04726_));
 sg13g2_a21oi_2 _12339_ (.B1(_04731_),
    .Y(_04732_),
    .A2(_04671_),
    .A1(_04668_));
 sg13g2_nor2_1 _12340_ (.A(_04730_),
    .B(_04732_),
    .Y(_04733_));
 sg13g2_o21ai_1 _12341_ (.B1(_04724_),
    .Y(_04734_),
    .A1(_04730_),
    .A2(_04732_));
 sg13g2_nand2_1 _12342_ (.Y(_04735_),
    .A(net1940),
    .B(_04734_));
 sg13g2_a21oi_1 _12343_ (.A1(_04723_),
    .A2(_04733_),
    .Y(_00856_),
    .B1(_04735_));
 sg13g2_xor2_1 _12344_ (.B(net3025),
    .A(net3144),
    .X(_04736_));
 sg13g2_nand2_1 _12345_ (.Y(_04737_),
    .A(_04722_),
    .B(_04734_));
 sg13g2_o21ai_1 _12346_ (.B1(net1920),
    .Y(_04738_),
    .A1(_04736_),
    .A2(_04737_));
 sg13g2_a21oi_1 _12347_ (.A1(_04736_),
    .A2(_04737_),
    .Y(_00857_),
    .B1(_04738_));
 sg13g2_a22oi_1 _12348_ (.Y(_04739_),
    .B1(net3025),
    .B2(\am_sdr0.cic0.integ2[20] ),
    .A2(net1518),
    .A1(\am_sdr0.cic0.integ2[19] ));
 sg13g2_nand2_1 _12349_ (.Y(_04740_),
    .A(_04734_),
    .B(_04739_));
 sg13g2_o21ai_1 _12350_ (.B1(_04740_),
    .Y(_04741_),
    .A1(\am_sdr0.cic0.integ2[20] ),
    .A2(net3025));
 sg13g2_xnor2_1 _12351_ (.Y(_04742_),
    .A(\am_sdr0.cic0.integ2[21] ),
    .B(net1514));
 sg13g2_a221oi_1 _12352_ (.B2(_04739_),
    .C1(_04742_),
    .B1(_04734_),
    .A1(_01588_),
    .Y(_04743_),
    .A2(_01589_));
 sg13g2_nand2b_1 _12353_ (.Y(_04744_),
    .B(net1920),
    .A_N(_04743_));
 sg13g2_a21oi_1 _12354_ (.A1(net3026),
    .A2(_04742_),
    .Y(_00858_),
    .B1(_04744_));
 sg13g2_a21oi_1 _12355_ (.A1(\am_sdr0.cic0.integ2[21] ),
    .A2(net1514),
    .Y(_04745_),
    .B1(_04743_));
 sg13g2_xnor2_1 _12356_ (.Y(_04746_),
    .A(net3019),
    .B(net1309));
 sg13g2_o21ai_1 _12357_ (.B1(net1920),
    .Y(_04747_),
    .A1(_04745_),
    .A2(_04746_));
 sg13g2_a21oi_1 _12358_ (.A1(_04745_),
    .A2(_04746_),
    .Y(_00859_),
    .B1(_04747_));
 sg13g2_nor2b_2 _12359_ (.A(net1341),
    .B_N(\am_sdr0.spi0.state[0] ),
    .Y(_04748_));
 sg13g2_nor3_1 _12360_ (.A(net1884),
    .B(_01569_),
    .C(net1404),
    .Y(_04749_));
 sg13g2_a22oi_1 _12361_ (.Y(_04750_),
    .B1(_04749_),
    .B2(_01194_),
    .A2(net1342),
    .A1(net1952));
 sg13g2_nand2b_1 _12362_ (.Y(_04751_),
    .B(\am_sdr0.spi0.SCK_qq ),
    .A_N(\am_sdr0.spi0.SCK_qqq ));
 sg13g2_a21o_1 _12363_ (.A2(_04751_),
    .A1(\am_sdr0.spi0.state[0] ),
    .B1(_04750_),
    .X(_04752_));
 sg13g2_nand2_1 _12364_ (.Y(_04753_),
    .A(net1302),
    .B(net1615));
 sg13g2_nand2_1 _12365_ (.Y(_04754_),
    .A(\am_sdr0.spi0.shift_reg[0] ),
    .B(net1561));
 sg13g2_o21ai_1 _12366_ (.B1(_04754_),
    .Y(_00860_),
    .A1(net1561),
    .A2(_04753_));
 sg13g2_nand2_1 _12367_ (.Y(_04755_),
    .A(net1470),
    .B(net1615));
 sg13g2_nand2_1 _12368_ (.Y(_04756_),
    .A(net1388),
    .B(net1561));
 sg13g2_o21ai_1 _12369_ (.B1(_04756_),
    .Y(_00861_),
    .A1(net1561),
    .A2(_04755_));
 sg13g2_nand2_1 _12370_ (.Y(_04757_),
    .A(net1388),
    .B(net1615));
 sg13g2_nand2_1 _12371_ (.Y(_04758_),
    .A(net1271),
    .B(net1561));
 sg13g2_o21ai_1 _12372_ (.B1(_04758_),
    .Y(_00862_),
    .A1(net1561),
    .A2(_04757_));
 sg13g2_nand2_1 _12373_ (.Y(_04759_),
    .A(net1271),
    .B(net1615));
 sg13g2_nand2_1 _12374_ (.Y(_04760_),
    .A(net1325),
    .B(net1561));
 sg13g2_o21ai_1 _12375_ (.B1(_04760_),
    .Y(_00863_),
    .A1(net1561),
    .A2(_04759_));
 sg13g2_nand2_1 _12376_ (.Y(_04761_),
    .A(net1325),
    .B(net1615));
 sg13g2_nand2_1 _12377_ (.Y(_04762_),
    .A(net1291),
    .B(net1559));
 sg13g2_o21ai_1 _12378_ (.B1(_04762_),
    .Y(_00864_),
    .A1(net1558),
    .A2(_04761_));
 sg13g2_nand2_1 _12379_ (.Y(_04763_),
    .A(net1291),
    .B(net1614));
 sg13g2_nand2_1 _12380_ (.Y(_04764_),
    .A(net1330),
    .B(net1559));
 sg13g2_o21ai_1 _12381_ (.B1(_04764_),
    .Y(_00865_),
    .A1(net1558),
    .A2(_04763_));
 sg13g2_nand2_1 _12382_ (.Y(_04765_),
    .A(net1330),
    .B(net1614));
 sg13g2_nand2_1 _12383_ (.Y(_04766_),
    .A(net1408),
    .B(net1559));
 sg13g2_o21ai_1 _12384_ (.B1(_04766_),
    .Y(_00866_),
    .A1(net1559),
    .A2(_04765_));
 sg13g2_nand2_1 _12385_ (.Y(_04767_),
    .A(net1408),
    .B(net1614));
 sg13g2_nand2_1 _12386_ (.Y(_04768_),
    .A(net1418),
    .B(net1558));
 sg13g2_o21ai_1 _12387_ (.B1(_04768_),
    .Y(_00867_),
    .A1(net1558),
    .A2(_04767_));
 sg13g2_nand2_1 _12388_ (.Y(_04769_),
    .A(net1418),
    .B(net1614));
 sg13g2_nand2_1 _12389_ (.Y(_04770_),
    .A(net1422),
    .B(net1558));
 sg13g2_o21ai_1 _12390_ (.B1(_04770_),
    .Y(_00868_),
    .A1(net1558),
    .A2(_04769_));
 sg13g2_nand2_1 _12391_ (.Y(_04771_),
    .A(\am_sdr0.spi0.shift_reg[8] ),
    .B(net1614));
 sg13g2_nand2_1 _12392_ (.Y(_04772_),
    .A(net1382),
    .B(net1555));
 sg13g2_o21ai_1 _12393_ (.B1(_04772_),
    .Y(_00869_),
    .A1(net1555),
    .A2(_04771_));
 sg13g2_nand2_1 _12394_ (.Y(_04773_),
    .A(\am_sdr0.spi0.shift_reg[9] ),
    .B(net1612));
 sg13g2_nand2_1 _12395_ (.Y(_04774_),
    .A(net1315),
    .B(net1555));
 sg13g2_o21ai_1 _12396_ (.B1(_04774_),
    .Y(_00870_),
    .A1(net1555),
    .A2(_04773_));
 sg13g2_nand2_1 _12397_ (.Y(_04775_),
    .A(net1315),
    .B(net1612));
 sg13g2_nand2_1 _12398_ (.Y(_04776_),
    .A(net1409),
    .B(net1554));
 sg13g2_o21ai_1 _12399_ (.B1(_04776_),
    .Y(_00871_),
    .A1(net1554),
    .A2(_04775_));
 sg13g2_nand2_1 _12400_ (.Y(_04777_),
    .A(\am_sdr0.spi0.shift_reg[11] ),
    .B(net1613));
 sg13g2_nand2_1 _12401_ (.Y(_04778_),
    .A(net1362),
    .B(net1556));
 sg13g2_o21ai_1 _12402_ (.B1(_04778_),
    .Y(_00872_),
    .A1(net1556),
    .A2(_04777_));
 sg13g2_nand2_1 _12403_ (.Y(_04779_),
    .A(\am_sdr0.spi0.shift_reg[12] ),
    .B(net1613));
 sg13g2_nand2_1 _12404_ (.Y(_04780_),
    .A(net1298),
    .B(net1557));
 sg13g2_o21ai_1 _12405_ (.B1(_04780_),
    .Y(_00873_),
    .A1(net1556),
    .A2(_04779_));
 sg13g2_nand2_1 _12406_ (.Y(_04781_),
    .A(net1298),
    .B(net1613));
 sg13g2_nand2_1 _12407_ (.Y(_04782_),
    .A(net1345),
    .B(net1557));
 sg13g2_o21ai_1 _12408_ (.B1(_04782_),
    .Y(_00874_),
    .A1(net1557),
    .A2(_04781_));
 sg13g2_nand2_1 _12409_ (.Y(_04783_),
    .A(net1345),
    .B(net1613));
 sg13g2_nand2_1 _12410_ (.Y(_04784_),
    .A(net1420),
    .B(net1556));
 sg13g2_o21ai_1 _12411_ (.B1(_04784_),
    .Y(_00875_),
    .A1(net1556),
    .A2(_04783_));
 sg13g2_nand2_1 _12412_ (.Y(_04785_),
    .A(\am_sdr0.spi0.shift_reg[15] ),
    .B(net1613));
 sg13g2_nand2_1 _12413_ (.Y(_04786_),
    .A(net1393),
    .B(net1557));
 sg13g2_o21ai_1 _12414_ (.B1(_04786_),
    .Y(_00876_),
    .A1(net1556),
    .A2(_04785_));
 sg13g2_nand2_1 _12415_ (.Y(_04787_),
    .A(\am_sdr0.spi0.shift_reg[16] ),
    .B(net1614));
 sg13g2_nand2_1 _12416_ (.Y(_04788_),
    .A(net1360),
    .B(net1557));
 sg13g2_o21ai_1 _12417_ (.B1(_04788_),
    .Y(_00877_),
    .A1(net1557),
    .A2(_04787_));
 sg13g2_nand2_1 _12418_ (.Y(_04789_),
    .A(net1360),
    .B(net1613));
 sg13g2_nand2_1 _12419_ (.Y(_04790_),
    .A(net2043),
    .B(net1556));
 sg13g2_o21ai_1 _12420_ (.B1(_04790_),
    .Y(_00878_),
    .A1(net1556),
    .A2(_04789_));
 sg13g2_nand2_1 _12421_ (.Y(_04791_),
    .A(\am_sdr0.spi0.shift_reg[18] ),
    .B(net1612));
 sg13g2_nand2_1 _12422_ (.Y(_04792_),
    .A(net1289),
    .B(net1554));
 sg13g2_o21ai_1 _12423_ (.B1(_04792_),
    .Y(_00879_),
    .A1(net1554),
    .A2(_04791_));
 sg13g2_nand2_1 _12424_ (.Y(_04793_),
    .A(net1289),
    .B(net1612));
 sg13g2_nand2_1 _12425_ (.Y(_04794_),
    .A(net1381),
    .B(net1553));
 sg13g2_o21ai_1 _12426_ (.B1(_04794_),
    .Y(_00880_),
    .A1(net1554),
    .A2(_04793_));
 sg13g2_nand2_1 _12427_ (.Y(_04795_),
    .A(net1381),
    .B(net1612));
 sg13g2_nand2_1 _12428_ (.Y(_04796_),
    .A(net1419),
    .B(net1553));
 sg13g2_o21ai_1 _12429_ (.B1(_04796_),
    .Y(_00881_),
    .A1(net1553),
    .A2(_04795_));
 sg13g2_nand2_1 _12430_ (.Y(_04797_),
    .A(net1419),
    .B(net1612));
 sg13g2_nand2_1 _12431_ (.Y(_04798_),
    .A(net1455),
    .B(net1553));
 sg13g2_o21ai_1 _12432_ (.B1(_04798_),
    .Y(_00882_),
    .A1(net1553),
    .A2(_04797_));
 sg13g2_nand2_1 _12433_ (.Y(_04799_),
    .A(\am_sdr0.spi0.shift_reg[22] ),
    .B(net1612));
 sg13g2_nand2_1 _12434_ (.Y(_04800_),
    .A(net1415),
    .B(net1553));
 sg13g2_o21ai_1 _12435_ (.B1(_04800_),
    .Y(_00883_),
    .A1(net1553),
    .A2(_04799_));
 sg13g2_nand2_1 _12436_ (.Y(_04801_),
    .A(\am_sdr0.spi0.shift_reg[23] ),
    .B(net1612));
 sg13g2_nand2_1 _12437_ (.Y(_04802_),
    .A(net1343),
    .B(net1553));
 sg13g2_o21ai_1 _12438_ (.B1(_04802_),
    .Y(_00884_),
    .A1(net1554),
    .A2(_04801_));
 sg13g2_nand2_1 _12439_ (.Y(_04803_),
    .A(net1343),
    .B(net1613));
 sg13g2_nand2_1 _12440_ (.Y(_04804_),
    .A(net2161),
    .B(net1555));
 sg13g2_o21ai_1 _12441_ (.B1(_04804_),
    .Y(_00885_),
    .A1(net1555),
    .A2(_04803_));
 sg13g2_nand2_1 _12442_ (.Y(_04805_),
    .A(net2161),
    .B(net1614));
 sg13g2_nand2_1 _12443_ (.Y(_04806_),
    .A(net2415),
    .B(net1558));
 sg13g2_o21ai_1 _12444_ (.B1(_04806_),
    .Y(_00886_),
    .A1(net1558),
    .A2(_04805_));
 sg13g2_nand2_1 _12445_ (.Y(_04807_),
    .A(\am_sdr0.spi0.shift_reg[26] ),
    .B(net1615));
 sg13g2_nand2_1 _12446_ (.Y(_04808_),
    .A(net1482),
    .B(net1562));
 sg13g2_o21ai_1 _12447_ (.B1(_04808_),
    .Y(_00887_),
    .A1(net1562),
    .A2(_04807_));
 sg13g2_nand2_1 _12448_ (.Y(_04809_),
    .A(\am_sdr0.spi0.shift_reg[27] ),
    .B(net1615));
 sg13g2_nand2_1 _12449_ (.Y(_04810_),
    .A(net1235),
    .B(net1562));
 sg13g2_o21ai_1 _12450_ (.B1(_04810_),
    .Y(_00888_),
    .A1(net1562),
    .A2(_04809_));
 sg13g2_o21ai_1 _12451_ (.B1(net2013),
    .Y(_04811_),
    .A1(net1729),
    .A2(\am_sdr0.cic0.x_out[8] ));
 sg13g2_a21oi_1 _12452_ (.A1(net1729),
    .A2(_01256_),
    .Y(_00889_),
    .B1(_04811_));
 sg13g2_o21ai_1 _12453_ (.B1(net1948),
    .Y(_04812_),
    .A1(net1728),
    .A2(\am_sdr0.cic0.x_out[9] ));
 sg13g2_a21oi_1 _12454_ (.A1(net1728),
    .A2(_01255_),
    .Y(_00890_),
    .B1(_04812_));
 sg13g2_o21ai_1 _12455_ (.B1(net2005),
    .Y(_04813_),
    .A1(net1713),
    .A2(\am_sdr0.cic0.x_out[10] ));
 sg13g2_a21oi_1 _12456_ (.A1(net1713),
    .A2(_01254_),
    .Y(_00891_),
    .B1(_04813_));
 sg13g2_o21ai_1 _12457_ (.B1(net1948),
    .Y(_04814_),
    .A1(net1713),
    .A2(\am_sdr0.cic0.x_out[11] ));
 sg13g2_a21oi_1 _12458_ (.A1(net1713),
    .A2(_01253_),
    .Y(_00892_),
    .B1(_04814_));
 sg13g2_o21ai_1 _12459_ (.B1(net1945),
    .Y(_04815_),
    .A1(net1712),
    .A2(\am_sdr0.cic0.x_out[12] ));
 sg13g2_a21oi_1 _12460_ (.A1(net1712),
    .A2(_01252_),
    .Y(_00893_),
    .B1(_04815_));
 sg13g2_o21ai_1 _12461_ (.B1(net1946),
    .Y(_04816_),
    .A1(net1715),
    .A2(\am_sdr0.cic0.x_out[13] ));
 sg13g2_a21oi_1 _12462_ (.A1(net1715),
    .A2(_01251_),
    .Y(_00894_),
    .B1(_04816_));
 sg13g2_o21ai_1 _12463_ (.B1(net1925),
    .Y(_04817_),
    .A1(net1709),
    .A2(\am_sdr0.cic0.x_out[14] ));
 sg13g2_a21oi_1 _12464_ (.A1(net1709),
    .A2(_01250_),
    .Y(_00895_),
    .B1(_04817_));
 sg13g2_o21ai_1 _12465_ (.B1(net1924),
    .Y(_04818_),
    .A1(net1709),
    .A2(net1694));
 sg13g2_a21oi_1 _12466_ (.A1(net1709),
    .A2(_01249_),
    .Y(_00896_),
    .B1(_04818_));
 sg13g2_nand2b_1 _12467_ (.Y(_04819_),
    .B(net2121),
    .A_N(net2614));
 sg13g2_a21oi_1 _12468_ (.A1(_01303_),
    .A2(net2614),
    .Y(_04820_),
    .B1(net1645));
 sg13g2_nor2_1 _12469_ (.A(net1643),
    .B(net1884),
    .Y(_01005_));
 sg13g2_a221oi_1 _12470_ (.B2(_04820_),
    .C1(net1884),
    .B1(_04819_),
    .A1(net1645),
    .Y(_00897_),
    .A2(_01280_));
 sg13g2_nor2b_1 _12471_ (.A(net2667),
    .B_N(\am_sdr0.cic0.integ_sample[1] ),
    .Y(_04821_));
 sg13g2_xnor2_1 _12472_ (.Y(_04822_),
    .A(net2667),
    .B(net2922));
 sg13g2_xnor2_1 _12473_ (.Y(_04823_),
    .A(_04819_),
    .B(_04822_));
 sg13g2_o21ai_1 _12474_ (.B1(net1952),
    .Y(_04824_),
    .A1(net1723),
    .A2(net2722));
 sg13g2_a21oi_1 _12475_ (.A1(net1723),
    .A2(_04823_),
    .Y(_00898_),
    .B1(_04824_));
 sg13g2_nand2b_1 _12476_ (.Y(_04825_),
    .B(\am_sdr0.cic0.integ_sample[2] ),
    .A_N(\am_sdr0.cic0.comb1_in_del[2] ));
 sg13g2_xor2_1 _12477_ (.B(net2928),
    .A(\am_sdr0.cic0.comb1_in_del[2] ),
    .X(_04826_));
 sg13g2_a21oi_1 _12478_ (.A1(_04819_),
    .A2(_04822_),
    .Y(_04827_),
    .B1(_04821_));
 sg13g2_xnor2_1 _12479_ (.Y(_04828_),
    .A(_04826_),
    .B(_04827_));
 sg13g2_o21ai_1 _12480_ (.B1(net1953),
    .Y(_04829_),
    .A1(net1723),
    .A2(net2545));
 sg13g2_a21oi_1 _12481_ (.A1(net1723),
    .A2(_04828_),
    .Y(_00899_),
    .B1(_04829_));
 sg13g2_nor2_1 _12482_ (.A(\am_sdr0.cic0.comb1_in_del[3] ),
    .B(_01300_),
    .Y(_04830_));
 sg13g2_nand2_1 _12483_ (.Y(_04831_),
    .A(\am_sdr0.cic0.comb1_in_del[3] ),
    .B(_01300_));
 sg13g2_nand2b_1 _12484_ (.Y(_04832_),
    .B(_04831_),
    .A_N(_04830_));
 sg13g2_o21ai_1 _12485_ (.B1(_04825_),
    .Y(_04833_),
    .A1(_04826_),
    .A2(_04827_));
 sg13g2_xor2_1 _12486_ (.B(_04833_),
    .A(_04832_),
    .X(_04834_));
 sg13g2_o21ai_1 _12487_ (.B1(net1953),
    .Y(_04835_),
    .A1(net1722),
    .A2(net2221));
 sg13g2_a21oi_1 _12488_ (.A1(net1722),
    .A2(_04834_),
    .Y(_00900_),
    .B1(_04835_));
 sg13g2_nor2_1 _12489_ (.A(\am_sdr0.cic0.comb1_in_del[4] ),
    .B(_01299_),
    .Y(_04836_));
 sg13g2_xor2_1 _12490_ (.B(net2738),
    .A(\am_sdr0.cic0.comb1_in_del[4] ),
    .X(_04837_));
 sg13g2_a21oi_1 _12491_ (.A1(_04831_),
    .A2(_04833_),
    .Y(_04838_),
    .B1(_04830_));
 sg13g2_or2_1 _12492_ (.X(_04839_),
    .B(_04838_),
    .A(_04837_));
 sg13g2_xnor2_1 _12493_ (.Y(_04840_),
    .A(_04837_),
    .B(_04838_));
 sg13g2_o21ai_1 _12494_ (.B1(net1950),
    .Y(_04841_),
    .A1(net1722),
    .A2(net2823));
 sg13g2_a21oi_1 _12495_ (.A1(net1721),
    .A2(_04840_),
    .Y(_00901_),
    .B1(_04841_));
 sg13g2_xor2_1 _12496_ (.B(net2626),
    .A(\am_sdr0.cic0.comb1_in_del[5] ),
    .X(_04842_));
 sg13g2_nor2b_1 _12497_ (.A(_04836_),
    .B_N(_04839_),
    .Y(_04843_));
 sg13g2_xnor2_1 _12498_ (.Y(_04844_),
    .A(net2627),
    .B(_04843_));
 sg13g2_o21ai_1 _12499_ (.B1(net1950),
    .Y(_04845_),
    .A1(net1722),
    .A2(net2431));
 sg13g2_a21oi_1 _12500_ (.A1(net1722),
    .A2(net2628),
    .Y(_00902_),
    .B1(_04845_));
 sg13g2_nor2_1 _12501_ (.A(\am_sdr0.cic0.comb1_in_del[6] ),
    .B(_01296_),
    .Y(_04846_));
 sg13g2_xor2_1 _12502_ (.B(net2858),
    .A(net2685),
    .X(_04847_));
 sg13g2_a21oi_1 _12503_ (.A1(_01297_),
    .A2(\am_sdr0.cic0.integ_sample[5] ),
    .Y(_04848_),
    .B1(_04836_));
 sg13g2_a22oi_1 _12504_ (.Y(_04849_),
    .B1(_04839_),
    .B2(_04848_),
    .A2(_01298_),
    .A1(net3324));
 sg13g2_a221oi_1 _12505_ (.B2(_04848_),
    .C1(_04847_),
    .B1(_04839_),
    .A1(\am_sdr0.cic0.comb1_in_del[5] ),
    .Y(_04850_),
    .A2(_01298_));
 sg13g2_xor2_1 _12506_ (.B(_04849_),
    .A(_04847_),
    .X(_04851_));
 sg13g2_o21ai_1 _12507_ (.B1(net1950),
    .Y(_04852_),
    .A1(net1718),
    .A2(net2331));
 sg13g2_a21oi_1 _12508_ (.A1(net1718),
    .A2(_04851_),
    .Y(_00903_),
    .B1(_04852_));
 sg13g2_nand2b_1 _12509_ (.Y(_04853_),
    .B(\am_sdr0.cic0.integ_sample[7] ),
    .A_N(\am_sdr0.cic0.comb1_in_del[7] ));
 sg13g2_xnor2_1 _12510_ (.Y(_04854_),
    .A(\am_sdr0.cic0.comb1_in_del[7] ),
    .B(\am_sdr0.cic0.integ_sample[7] ));
 sg13g2_o21ai_1 _12511_ (.B1(_04854_),
    .Y(_04855_),
    .A1(_04846_),
    .A2(_04850_));
 sg13g2_or3_1 _12512_ (.A(_04846_),
    .B(_04850_),
    .C(_04854_),
    .X(_04856_));
 sg13g2_and2_1 _12513_ (.A(_04855_),
    .B(_04856_),
    .X(_04857_));
 sg13g2_mux2_1 _12514_ (.A0(net2107),
    .A1(_04857_),
    .S(net1718),
    .X(_04858_));
 sg13g2_and2_1 _12515_ (.A(net1953),
    .B(_04858_),
    .X(_00904_));
 sg13g2_nand2_1 _12516_ (.Y(_04859_),
    .A(_04853_),
    .B(_04855_));
 sg13g2_nor2_1 _12517_ (.A(\am_sdr0.cic0.comb1_in_del[8] ),
    .B(_01294_),
    .Y(_04860_));
 sg13g2_xnor2_1 _12518_ (.Y(_04861_),
    .A(\am_sdr0.cic0.comb1_in_del[8] ),
    .B(net2703));
 sg13g2_inv_1 _12519_ (.Y(_04862_),
    .A(_04861_));
 sg13g2_xnor2_1 _12520_ (.Y(_04863_),
    .A(_04859_),
    .B(_04861_));
 sg13g2_o21ai_1 _12521_ (.B1(net1942),
    .Y(_04864_),
    .A1(net1717),
    .A2(net2440));
 sg13g2_a21oi_1 _12522_ (.A1(net1717),
    .A2(_04863_),
    .Y(_00905_),
    .B1(_04864_));
 sg13g2_xor2_1 _12523_ (.B(net2971),
    .A(\am_sdr0.cic0.comb1_in_del[9] ),
    .X(_04865_));
 sg13g2_a21oi_1 _12524_ (.A1(_04859_),
    .A2(_04861_),
    .Y(_04866_),
    .B1(_04860_));
 sg13g2_xnor2_1 _12525_ (.Y(_04867_),
    .A(net2972),
    .B(_04866_));
 sg13g2_o21ai_1 _12526_ (.B1(net1941),
    .Y(_04868_),
    .A1(net1717),
    .A2(net2894));
 sg13g2_a21oi_1 _12527_ (.A1(net1717),
    .A2(_04867_),
    .Y(_00906_),
    .B1(_04868_));
 sg13g2_nand2b_1 _12528_ (.Y(_04869_),
    .B(\am_sdr0.cic0.integ_sample[10] ),
    .A_N(\am_sdr0.cic0.comb1_in_del[10] ));
 sg13g2_xor2_1 _12529_ (.B(\am_sdr0.cic0.integ_sample[10] ),
    .A(\am_sdr0.cic0.comb1_in_del[10] ),
    .X(_04870_));
 sg13g2_a21oi_1 _12530_ (.A1(_01292_),
    .A2(\am_sdr0.cic0.integ_sample[9] ),
    .Y(_04871_),
    .B1(_04860_));
 sg13g2_a21oi_1 _12531_ (.A1(\am_sdr0.cic0.comb1_in_del[9] ),
    .A2(_01293_),
    .Y(_04872_),
    .B1(_04871_));
 sg13g2_nor2_1 _12532_ (.A(_04862_),
    .B(_04865_),
    .Y(_04873_));
 sg13g2_a21oi_1 _12533_ (.A1(_04859_),
    .A2(_04873_),
    .Y(_04874_),
    .B1(_04872_));
 sg13g2_xnor2_1 _12534_ (.Y(_04875_),
    .A(_04870_),
    .B(_04874_));
 sg13g2_o21ai_1 _12535_ (.B1(net1941),
    .Y(_04876_),
    .A1(net1717),
    .A2(net2401));
 sg13g2_a21oi_1 _12536_ (.A1(net1717),
    .A2(_04875_),
    .Y(_00907_),
    .B1(_04876_));
 sg13g2_nor2b_1 _12537_ (.A(\am_sdr0.cic0.integ_sample[11] ),
    .B_N(\am_sdr0.cic0.comb1_in_del[11] ),
    .Y(_04877_));
 sg13g2_nand2b_1 _12538_ (.Y(_04878_),
    .B(\am_sdr0.cic0.integ_sample[11] ),
    .A_N(\am_sdr0.cic0.comb1_in_del[11] ));
 sg13g2_nand2b_1 _12539_ (.Y(_04879_),
    .B(_04878_),
    .A_N(_04877_));
 sg13g2_o21ai_1 _12540_ (.B1(_04869_),
    .Y(_04880_),
    .A1(_04870_),
    .A2(_04874_));
 sg13g2_xor2_1 _12541_ (.B(_04880_),
    .A(_04879_),
    .X(_04881_));
 sg13g2_o21ai_1 _12542_ (.B1(net1941),
    .Y(_04882_),
    .A1(net1704),
    .A2(net2911));
 sg13g2_a21oi_1 _12543_ (.A1(net1704),
    .A2(_04881_),
    .Y(_00908_),
    .B1(_04882_));
 sg13g2_nand2b_1 _12544_ (.Y(_04883_),
    .B(\am_sdr0.cic0.integ_sample[12] ),
    .A_N(\am_sdr0.cic0.comb1_in_del[12] ));
 sg13g2_xor2_1 _12545_ (.B(\am_sdr0.cic0.integ_sample[12] ),
    .A(\am_sdr0.cic0.comb1_in_del[12] ),
    .X(_04884_));
 sg13g2_nor2_1 _12546_ (.A(_04870_),
    .B(_04879_),
    .Y(_04885_));
 sg13g2_o21ai_1 _12547_ (.B1(_04878_),
    .Y(_04886_),
    .A1(_04869_),
    .A2(_04877_));
 sg13g2_a21o_1 _12548_ (.A2(_04885_),
    .A1(_04872_),
    .B1(_04886_),
    .X(_04887_));
 sg13g2_nand2_1 _12549_ (.Y(_04888_),
    .A(_04873_),
    .B(_04885_));
 sg13g2_a21oi_2 _12550_ (.B1(_04888_),
    .Y(_04889_),
    .A2(_04855_),
    .A1(_04853_));
 sg13g2_nor2_1 _12551_ (.A(_04887_),
    .B(_04889_),
    .Y(_04890_));
 sg13g2_xnor2_1 _12552_ (.Y(_04891_),
    .A(_04884_),
    .B(_04890_));
 sg13g2_o21ai_1 _12553_ (.B1(net1941),
    .Y(_04892_),
    .A1(net1704),
    .A2(net3047));
 sg13g2_a21oi_1 _12554_ (.A1(net1706),
    .A2(_04891_),
    .Y(_00909_),
    .B1(_04892_));
 sg13g2_nor2b_1 _12555_ (.A(\am_sdr0.cic0.integ_sample[13] ),
    .B_N(\am_sdr0.cic0.comb1_in_del[13] ),
    .Y(_04893_));
 sg13g2_nand2b_1 _12556_ (.Y(_04894_),
    .B(\am_sdr0.cic0.integ_sample[13] ),
    .A_N(\am_sdr0.cic0.comb1_in_del[13] ));
 sg13g2_nand2b_1 _12557_ (.Y(_04895_),
    .B(_04894_),
    .A_N(_04893_));
 sg13g2_o21ai_1 _12558_ (.B1(_04883_),
    .Y(_04896_),
    .A1(_04884_),
    .A2(_04890_));
 sg13g2_xor2_1 _12559_ (.B(_04896_),
    .A(_04895_),
    .X(_04897_));
 sg13g2_o21ai_1 _12560_ (.B1(net1940),
    .Y(_04898_),
    .A1(net1703),
    .A2(net2694));
 sg13g2_a21oi_1 _12561_ (.A1(net1703),
    .A2(_04897_),
    .Y(_00910_),
    .B1(_04898_));
 sg13g2_nor2_1 _12562_ (.A(\am_sdr0.cic0.comb1_in_del[14] ),
    .B(_01287_),
    .Y(_04899_));
 sg13g2_nand2_1 _12563_ (.Y(_04900_),
    .A(net2916),
    .B(_01287_));
 sg13g2_nand2b_2 _12564_ (.Y(_04901_),
    .B(_04900_),
    .A_N(_04899_));
 sg13g2_o21ai_1 _12565_ (.B1(_04894_),
    .Y(_04902_),
    .A1(_04883_),
    .A2(_04893_));
 sg13g2_inv_1 _12566_ (.Y(_04903_),
    .A(_04902_));
 sg13g2_or2_1 _12567_ (.X(_04904_),
    .B(_04895_),
    .A(_04884_));
 sg13g2_o21ai_1 _12568_ (.B1(_04903_),
    .Y(_04905_),
    .A1(_04890_),
    .A2(_04904_));
 sg13g2_xor2_1 _12569_ (.B(_04905_),
    .A(_04901_),
    .X(_04906_));
 sg13g2_o21ai_1 _12570_ (.B1(net1940),
    .Y(_04907_),
    .A1(net1703),
    .A2(net2472));
 sg13g2_a21oi_1 _12571_ (.A1(net1703),
    .A2(_04906_),
    .Y(_00911_),
    .B1(_04907_));
 sg13g2_nand2_1 _12572_ (.Y(_04908_),
    .A(_01286_),
    .B(\am_sdr0.cic0.integ_sample[15] ));
 sg13g2_xor2_1 _12573_ (.B(\am_sdr0.cic0.integ_sample[15] ),
    .A(\am_sdr0.cic0.comb1_in_del[15] ),
    .X(_04909_));
 sg13g2_a21oi_1 _12574_ (.A1(_04900_),
    .A2(_04905_),
    .Y(_04910_),
    .B1(_04899_));
 sg13g2_xnor2_1 _12575_ (.Y(_04911_),
    .A(_04909_),
    .B(net2917));
 sg13g2_o21ai_1 _12576_ (.B1(net1945),
    .Y(_04912_),
    .A1(net1703),
    .A2(net2743));
 sg13g2_a21oi_1 _12577_ (.A1(net1703),
    .A2(_04911_),
    .Y(_00912_),
    .B1(_04912_));
 sg13g2_nand2b_1 _12578_ (.Y(_04913_),
    .B(net2852),
    .A_N(\am_sdr0.cic0.comb1_in_del[16] ));
 sg13g2_xor2_1 _12579_ (.B(net2852),
    .A(net2555),
    .X(_04914_));
 sg13g2_nor2_1 _12580_ (.A(_04901_),
    .B(_04909_),
    .Y(_04915_));
 sg13g2_nor3_2 _12581_ (.A(_04901_),
    .B(_04904_),
    .C(_04909_),
    .Y(_04916_));
 sg13g2_o21ai_1 _12582_ (.B1(_04899_),
    .Y(_04917_),
    .A1(_01286_),
    .A2(\am_sdr0.cic0.integ_sample[15] ));
 sg13g2_a22oi_1 _12583_ (.Y(_04918_),
    .B1(_04916_),
    .B2(_04887_),
    .A2(_04915_),
    .A1(_04902_));
 sg13g2_nand3_1 _12584_ (.B(_04917_),
    .C(_04918_),
    .A(_04908_),
    .Y(_04919_));
 sg13g2_a21oi_2 _12585_ (.B1(_04919_),
    .Y(_04920_),
    .A2(_04916_),
    .A1(_04889_));
 sg13g2_xnor2_1 _12586_ (.Y(_04921_),
    .A(_04914_),
    .B(_04920_));
 sg13g2_o21ai_1 _12587_ (.B1(net1943),
    .Y(_04922_),
    .A1(net1701),
    .A2(net2272));
 sg13g2_a21oi_1 _12588_ (.A1(net1701),
    .A2(_04921_),
    .Y(_00913_),
    .B1(_04922_));
 sg13g2_xnor2_1 _12589_ (.Y(_04923_),
    .A(\am_sdr0.cic0.comb1_in_del[17] ),
    .B(net2936));
 sg13g2_o21ai_1 _12590_ (.B1(_04913_),
    .Y(_04924_),
    .A1(_04914_),
    .A2(_04920_));
 sg13g2_xnor2_1 _12591_ (.Y(_04925_),
    .A(_04923_),
    .B(_04924_));
 sg13g2_o21ai_1 _12592_ (.B1(net1923),
    .Y(_04926_),
    .A1(net1701),
    .A2(net2748));
 sg13g2_a21oi_1 _12593_ (.A1(net1701),
    .A2(net2937),
    .Y(_00914_),
    .B1(_04926_));
 sg13g2_nor2_1 _12594_ (.A(\am_sdr0.cic0.comb1_in_del[18] ),
    .B(_01282_),
    .Y(_04927_));
 sg13g2_xnor2_1 _12595_ (.Y(_04928_),
    .A(\am_sdr0.cic0.comb1_in_del[18] ),
    .B(net2661));
 sg13g2_nand2b_1 _12596_ (.Y(_04929_),
    .B(_04923_),
    .A_N(_04914_));
 sg13g2_a21oi_1 _12597_ (.A1(\am_sdr0.cic0.comb1_in_del[17] ),
    .A2(_01284_),
    .Y(_04930_),
    .B1(_04913_));
 sg13g2_a21oi_1 _12598_ (.A1(_01283_),
    .A2(\am_sdr0.cic0.integ_sample[17] ),
    .Y(_04931_),
    .B1(_04930_));
 sg13g2_o21ai_1 _12599_ (.B1(_04931_),
    .Y(_04932_),
    .A1(_04920_),
    .A2(_04929_));
 sg13g2_xnor2_1 _12600_ (.Y(_04933_),
    .A(net2662),
    .B(_04932_));
 sg13g2_o21ai_1 _12601_ (.B1(net1919),
    .Y(_04934_),
    .A1(net1700),
    .A2(net2589));
 sg13g2_a21oi_1 _12602_ (.A1(net1700),
    .A2(_04933_),
    .Y(_00915_),
    .B1(_04934_));
 sg13g2_a21oi_1 _12603_ (.A1(_04928_),
    .A2(_04932_),
    .Y(_04935_),
    .B1(_04927_));
 sg13g2_xor2_1 _12604_ (.B(net2287),
    .A(net2682),
    .X(_04936_));
 sg13g2_xnor2_1 _12605_ (.Y(_04937_),
    .A(_04935_),
    .B(_04936_));
 sg13g2_o21ai_1 _12606_ (.B1(net1920),
    .Y(_04938_),
    .A1(net1700),
    .A2(net2123));
 sg13g2_a21oi_1 _12607_ (.A1(net1700),
    .A2(net2683),
    .Y(_00916_),
    .B1(_04938_));
 sg13g2_o21ai_1 _12608_ (.B1(net1952),
    .Y(_04939_),
    .A1(net1645),
    .A2(\am_sdr0.cic0.integ_sample[0] ));
 sg13g2_a21oi_1 _12609_ (.A1(net1645),
    .A2(_01303_),
    .Y(_00917_),
    .B1(_04939_));
 sg13g2_o21ai_1 _12610_ (.B1(net1952),
    .Y(_04940_),
    .A1(net1726),
    .A2(net2667));
 sg13g2_a21oi_1 _12611_ (.A1(net1726),
    .A2(_01302_),
    .Y(_00918_),
    .B1(_04940_));
 sg13g2_o21ai_1 _12612_ (.B1(net1952),
    .Y(_04941_),
    .A1(net1721),
    .A2(\am_sdr0.cic0.comb1_in_del[2] ));
 sg13g2_a21oi_1 _12613_ (.A1(net1721),
    .A2(_01301_),
    .Y(_00919_),
    .B1(_04941_));
 sg13g2_o21ai_1 _12614_ (.B1(net1950),
    .Y(_04942_),
    .A1(net1721),
    .A2(\am_sdr0.cic0.comb1_in_del[3] ));
 sg13g2_a21oi_1 _12615_ (.A1(net1721),
    .A2(_01300_),
    .Y(_00920_),
    .B1(_04942_));
 sg13g2_o21ai_1 _12616_ (.B1(net1950),
    .Y(_04943_),
    .A1(net1721),
    .A2(\am_sdr0.cic0.comb1_in_del[4] ));
 sg13g2_a21oi_1 _12617_ (.A1(net1721),
    .A2(_01299_),
    .Y(_00921_),
    .B1(_04943_));
 sg13g2_o21ai_1 _12618_ (.B1(net1953),
    .Y(_04944_),
    .A1(net1720),
    .A2(net2994));
 sg13g2_a21oi_1 _12619_ (.A1(net1720),
    .A2(_01298_),
    .Y(_00922_),
    .B1(_04944_));
 sg13g2_o21ai_1 _12620_ (.B1(net1953),
    .Y(_04945_),
    .A1(net1716),
    .A2(net2685));
 sg13g2_a21oi_1 _12621_ (.A1(net1716),
    .A2(_01296_),
    .Y(_00923_),
    .B1(_04945_));
 sg13g2_o21ai_1 _12622_ (.B1(net1941),
    .Y(_04946_),
    .A1(net1716),
    .A2(net2624));
 sg13g2_a21oi_1 _12623_ (.A1(net1716),
    .A2(_01295_),
    .Y(_00924_),
    .B1(_04946_));
 sg13g2_o21ai_1 _12624_ (.B1(net1941),
    .Y(_04947_),
    .A1(net1716),
    .A2(net2782));
 sg13g2_a21oi_1 _12625_ (.A1(net1716),
    .A2(_01294_),
    .Y(_00925_),
    .B1(_04947_));
 sg13g2_o21ai_1 _12626_ (.B1(net1942),
    .Y(_04948_),
    .A1(net1716),
    .A2(net2843));
 sg13g2_a21oi_1 _12627_ (.A1(net1716),
    .A2(_01293_),
    .Y(_00926_),
    .B1(_04948_));
 sg13g2_o21ai_1 _12628_ (.B1(net1941),
    .Y(_04949_),
    .A1(net1705),
    .A2(\am_sdr0.cic0.comb1_in_del[10] ));
 sg13g2_a21oi_1 _12629_ (.A1(net1705),
    .A2(_01291_),
    .Y(_00927_),
    .B1(_04949_));
 sg13g2_o21ai_1 _12630_ (.B1(net1941),
    .Y(_04950_),
    .A1(net1705),
    .A2(\am_sdr0.cic0.comb1_in_del[11] ));
 sg13g2_a21oi_1 _12631_ (.A1(net1705),
    .A2(_01290_),
    .Y(_00928_),
    .B1(_04950_));
 sg13g2_o21ai_1 _12632_ (.B1(net1940),
    .Y(_04951_),
    .A1(net1705),
    .A2(net2573));
 sg13g2_a21oi_1 _12633_ (.A1(net1705),
    .A2(_01289_),
    .Y(_00929_),
    .B1(_04951_));
 sg13g2_o21ai_1 _12634_ (.B1(net1940),
    .Y(_04952_),
    .A1(net1705),
    .A2(net2216));
 sg13g2_a21oi_1 _12635_ (.A1(net1705),
    .A2(_01288_),
    .Y(_00930_),
    .B1(_04952_));
 sg13g2_o21ai_1 _12636_ (.B1(net1943),
    .Y(_04953_),
    .A1(net1699),
    .A2(net2462));
 sg13g2_a21oi_1 _12637_ (.A1(net1699),
    .A2(_01287_),
    .Y(_00931_),
    .B1(_04953_));
 sg13g2_o21ai_1 _12638_ (.B1(net1943),
    .Y(_04954_),
    .A1(net1642),
    .A2(\am_sdr0.cic0.integ_sample[15] ));
 sg13g2_a21oi_1 _12639_ (.A1(net1642),
    .A2(_01286_),
    .Y(_00932_),
    .B1(_04954_));
 sg13g2_o21ai_1 _12640_ (.B1(net1919),
    .Y(_04955_),
    .A1(net1702),
    .A2(net2555));
 sg13g2_a21oi_1 _12641_ (.A1(net1702),
    .A2(_01285_),
    .Y(_00933_),
    .B1(_04955_));
 sg13g2_o21ai_1 _12642_ (.B1(net1919),
    .Y(_04956_),
    .A1(net1699),
    .A2(net2638));
 sg13g2_a21oi_1 _12643_ (.A1(net1699),
    .A2(_01284_),
    .Y(_00934_),
    .B1(_04956_));
 sg13g2_o21ai_1 _12644_ (.B1(net1919),
    .Y(_04957_),
    .A1(net1699),
    .A2(net2688));
 sg13g2_a21oi_1 _12645_ (.A1(net1699),
    .A2(_01282_),
    .Y(_00935_),
    .B1(_04957_));
 sg13g2_o21ai_1 _12646_ (.B1(net1920),
    .Y(_04958_),
    .A1(net1699),
    .A2(\am_sdr0.cic0.comb1_in_del[19] ));
 sg13g2_a21oi_1 _12647_ (.A1(net1699),
    .A2(_01281_),
    .Y(_00936_),
    .B1(_04958_));
 sg13g2_nand2b_1 _12648_ (.Y(_04959_),
    .B(net2377),
    .A_N(net2547));
 sg13g2_a21oi_1 _12649_ (.A1(_01279_),
    .A2(net2547),
    .Y(_04960_),
    .B1(net1645));
 sg13g2_a221oi_1 _12650_ (.B2(_04960_),
    .C1(net1885),
    .B1(_04959_),
    .A1(net1645),
    .Y(_00937_),
    .A2(_01248_));
 sg13g2_nor2b_1 _12651_ (.A(net2672),
    .B_N(\am_sdr0.cic0.comb1[1] ),
    .Y(_04961_));
 sg13g2_xnor2_1 _12652_ (.Y(_04962_),
    .A(net2672),
    .B(\am_sdr0.cic0.comb1[1] ));
 sg13g2_xnor2_1 _12653_ (.Y(_04963_),
    .A(_04959_),
    .B(net2723));
 sg13g2_o21ai_1 _12654_ (.B1(net1956),
    .Y(_04964_),
    .A1(net1731),
    .A2(net2074));
 sg13g2_a21oi_1 _12655_ (.A1(net1731),
    .A2(_04963_),
    .Y(_00938_),
    .B1(_04964_));
 sg13g2_nand2b_1 _12656_ (.Y(_04965_),
    .B(\am_sdr0.cic0.comb1[2] ),
    .A_N(\am_sdr0.cic0.comb2_in_del[2] ));
 sg13g2_xor2_1 _12657_ (.B(\am_sdr0.cic0.comb1[2] ),
    .A(\am_sdr0.cic0.comb2_in_del[2] ),
    .X(_04966_));
 sg13g2_a21oi_1 _12658_ (.A1(_04959_),
    .A2(_04962_),
    .Y(_04967_),
    .B1(_04961_));
 sg13g2_xnor2_1 _12659_ (.Y(_04968_),
    .A(_04966_),
    .B(_04967_));
 sg13g2_o21ai_1 _12660_ (.B1(net1956),
    .Y(_04969_),
    .A1(net1731),
    .A2(net2913));
 sg13g2_a21oi_1 _12661_ (.A1(net1731),
    .A2(_04968_),
    .Y(_00939_),
    .B1(_04969_));
 sg13g2_nor2_1 _12662_ (.A(\am_sdr0.cic0.comb2_in_del[3] ),
    .B(_01276_),
    .Y(_04970_));
 sg13g2_nand2_1 _12663_ (.Y(_04971_),
    .A(\am_sdr0.cic0.comb2_in_del[3] ),
    .B(_01276_));
 sg13g2_nor2b_1 _12664_ (.A(_04970_),
    .B_N(_04971_),
    .Y(_04972_));
 sg13g2_o21ai_1 _12665_ (.B1(_04965_),
    .Y(_04973_),
    .A1(_04966_),
    .A2(_04967_));
 sg13g2_xnor2_1 _12666_ (.Y(_04974_),
    .A(_04972_),
    .B(_04973_));
 sg13g2_o21ai_1 _12667_ (.B1(net1956),
    .Y(_04975_),
    .A1(net1732),
    .A2(net2793));
 sg13g2_a21oi_1 _12668_ (.A1(net1732),
    .A2(_04974_),
    .Y(_00940_),
    .B1(_04975_));
 sg13g2_nor2_1 _12669_ (.A(\am_sdr0.cic0.comb2_in_del[4] ),
    .B(_01275_),
    .Y(_04976_));
 sg13g2_xor2_1 _12670_ (.B(\am_sdr0.cic0.comb1[4] ),
    .A(\am_sdr0.cic0.comb2_in_del[4] ),
    .X(_04977_));
 sg13g2_a21oi_2 _12671_ (.B1(_04970_),
    .Y(_04978_),
    .A2(_04973_),
    .A1(_04971_));
 sg13g2_nor2_1 _12672_ (.A(_04977_),
    .B(_04978_),
    .Y(_04979_));
 sg13g2_xnor2_1 _12673_ (.Y(_04980_),
    .A(_04977_),
    .B(_04978_));
 sg13g2_o21ai_1 _12674_ (.B1(net1954),
    .Y(_04981_),
    .A1(net1732),
    .A2(net2399));
 sg13g2_a21oi_1 _12675_ (.A1(net1732),
    .A2(_04980_),
    .Y(_00941_),
    .B1(_04981_));
 sg13g2_nand2b_1 _12676_ (.Y(_04982_),
    .B(net2431),
    .A_N(\am_sdr0.cic0.comb2_in_del[5] ));
 sg13g2_nand2_1 _12677_ (.Y(_04983_),
    .A(\am_sdr0.cic0.comb2_in_del[5] ),
    .B(_01274_));
 sg13g2_nor2_1 _12678_ (.A(_04976_),
    .B(_04979_),
    .Y(_04984_));
 sg13g2_a21oi_1 _12679_ (.A1(_04982_),
    .A2(_04983_),
    .Y(_04985_),
    .B1(_04984_));
 sg13g2_nand3_1 _12680_ (.B(_04983_),
    .C(_04984_),
    .A(_04982_),
    .Y(_04986_));
 sg13g2_nor2_1 _12681_ (.A(net1644),
    .B(_04985_),
    .Y(_04987_));
 sg13g2_a221oi_1 _12682_ (.B2(_04987_),
    .C1(net1884),
    .B1(_04986_),
    .A1(net1644),
    .Y(_00942_),
    .A2(_01242_));
 sg13g2_nand2b_1 _12683_ (.Y(_04988_),
    .B(net2331),
    .A_N(\am_sdr0.cic0.comb2_in_del[6] ));
 sg13g2_xnor2_1 _12684_ (.Y(_04989_),
    .A(\am_sdr0.cic0.comb2_in_del[6] ),
    .B(\am_sdr0.cic0.comb1[6] ));
 sg13g2_nor2b_1 _12685_ (.A(_04976_),
    .B_N(_04982_),
    .Y(_04990_));
 sg13g2_o21ai_1 _12686_ (.B1(_04990_),
    .Y(_04991_),
    .A1(_04977_),
    .A2(_04978_));
 sg13g2_nand3_1 _12687_ (.B(_04989_),
    .C(_04991_),
    .A(_04983_),
    .Y(_04992_));
 sg13g2_a21o_1 _12688_ (.A2(_04991_),
    .A1(_04983_),
    .B1(_04989_),
    .X(_04993_));
 sg13g2_nand2_1 _12689_ (.Y(_04994_),
    .A(_04992_),
    .B(_04993_));
 sg13g2_o21ai_1 _12690_ (.B1(net1958),
    .Y(_04995_),
    .A1(net1732),
    .A2(net2444));
 sg13g2_a21oi_1 _12691_ (.A1(net1732),
    .A2(_04994_),
    .Y(_00943_),
    .B1(_04995_));
 sg13g2_nand2b_1 _12692_ (.Y(_04996_),
    .B(\am_sdr0.cic0.comb1[7] ),
    .A_N(\am_sdr0.cic0.comb2_in_del[7] ));
 sg13g2_xor2_1 _12693_ (.B(\am_sdr0.cic0.comb1[7] ),
    .A(\am_sdr0.cic0.comb2_in_del[7] ),
    .X(_04997_));
 sg13g2_a21o_1 _12694_ (.A2(_04992_),
    .A1(_04988_),
    .B1(_04997_),
    .X(_04998_));
 sg13g2_nand3_1 _12695_ (.B(_04992_),
    .C(_04997_),
    .A(_04988_),
    .Y(_04999_));
 sg13g2_a21oi_1 _12696_ (.A1(_04998_),
    .A2(_04999_),
    .Y(_05000_),
    .B1(net1643));
 sg13g2_o21ai_1 _12697_ (.B1(net1954),
    .Y(_05001_),
    .A1(net1727),
    .A2(net2641));
 sg13g2_nor2_1 _12698_ (.A(_05000_),
    .B(_05001_),
    .Y(_00944_));
 sg13g2_nand2_1 _12699_ (.Y(_05002_),
    .A(_04996_),
    .B(_04998_));
 sg13g2_nor2_1 _12700_ (.A(\am_sdr0.cic0.comb2_in_del[8] ),
    .B(_01271_),
    .Y(_05003_));
 sg13g2_xnor2_1 _12701_ (.Y(_05004_),
    .A(\am_sdr0.cic0.comb2_in_del[8] ),
    .B(\am_sdr0.cic0.comb1[8] ));
 sg13g2_inv_1 _12702_ (.Y(_05005_),
    .A(_05004_));
 sg13g2_xnor2_1 _12703_ (.Y(_05006_),
    .A(_05002_),
    .B(net2441));
 sg13g2_o21ai_1 _12704_ (.B1(net1955),
    .Y(_05007_),
    .A1(net1730),
    .A2(net2319));
 sg13g2_a21oi_1 _12705_ (.A1(net1730),
    .A2(_05006_),
    .Y(_00945_),
    .B1(_05007_));
 sg13g2_xor2_1 _12706_ (.B(\am_sdr0.cic0.comb1[9] ),
    .A(\am_sdr0.cic0.comb2_in_del[9] ),
    .X(_05008_));
 sg13g2_a21oi_1 _12707_ (.A1(_05002_),
    .A2(_05004_),
    .Y(_05009_),
    .B1(_05003_));
 sg13g2_xnor2_1 _12708_ (.Y(_05010_),
    .A(_05008_),
    .B(_05009_));
 sg13g2_o21ai_1 _12709_ (.B1(net1955),
    .Y(_05011_),
    .A1(net1730),
    .A2(net2880));
 sg13g2_a21oi_1 _12710_ (.A1(net1727),
    .A2(_05010_),
    .Y(_00946_),
    .B1(_05011_));
 sg13g2_nand2b_1 _12711_ (.Y(_05012_),
    .B(net3328),
    .A_N(\am_sdr0.cic0.comb2_in_del[10] ));
 sg13g2_xor2_1 _12712_ (.B(net3323),
    .A(\am_sdr0.cic0.comb2_in_del[10] ),
    .X(_05013_));
 sg13g2_a21oi_1 _12713_ (.A1(_01269_),
    .A2(\am_sdr0.cic0.comb1[9] ),
    .Y(_05014_),
    .B1(_05003_));
 sg13g2_a21oi_1 _12714_ (.A1(\am_sdr0.cic0.comb2_in_del[9] ),
    .A2(_01270_),
    .Y(_05015_),
    .B1(_05014_));
 sg13g2_nor2_1 _12715_ (.A(_05005_),
    .B(_05008_),
    .Y(_05016_));
 sg13g2_a21oi_1 _12716_ (.A1(_05002_),
    .A2(_05016_),
    .Y(_05017_),
    .B1(_05015_));
 sg13g2_xnor2_1 _12717_ (.Y(_05018_),
    .A(_05013_),
    .B(_05017_));
 sg13g2_o21ai_1 _12718_ (.B1(net1947),
    .Y(_05019_),
    .A1(net1727),
    .A2(net2212));
 sg13g2_a21oi_1 _12719_ (.A1(net1727),
    .A2(_05018_),
    .Y(_00947_),
    .B1(_05019_));
 sg13g2_nor2b_1 _12720_ (.A(\am_sdr0.cic0.comb1[11] ),
    .B_N(\am_sdr0.cic0.comb2_in_del[11] ),
    .Y(_05020_));
 sg13g2_nand2b_1 _12721_ (.Y(_05021_),
    .B(\am_sdr0.cic0.comb1[11] ),
    .A_N(\am_sdr0.cic0.comb2_in_del[11] ));
 sg13g2_nand2b_1 _12722_ (.Y(_05022_),
    .B(_05021_),
    .A_N(_05020_));
 sg13g2_o21ai_1 _12723_ (.B1(_05012_),
    .Y(_05023_),
    .A1(_05013_),
    .A2(_05017_));
 sg13g2_xor2_1 _12724_ (.B(_05023_),
    .A(_05022_),
    .X(_05024_));
 sg13g2_o21ai_1 _12725_ (.B1(net1947),
    .Y(_05025_),
    .A1(net1727),
    .A2(net2838));
 sg13g2_a21oi_1 _12726_ (.A1(net1727),
    .A2(_05024_),
    .Y(_00948_),
    .B1(_05025_));
 sg13g2_xor2_1 _12727_ (.B(\am_sdr0.cic0.comb1[12] ),
    .A(\am_sdr0.cic0.comb2_in_del[12] ),
    .X(_05026_));
 sg13g2_nor2_1 _12728_ (.A(_05013_),
    .B(_05022_),
    .Y(_05027_));
 sg13g2_o21ai_1 _12729_ (.B1(_05021_),
    .Y(_05028_),
    .A1(_05012_),
    .A2(_05020_));
 sg13g2_a21oi_2 _12730_ (.B1(_05028_),
    .Y(_05029_),
    .A2(_05027_),
    .A1(_05015_));
 sg13g2_nand2_1 _12731_ (.Y(_05030_),
    .A(_05016_),
    .B(_05027_));
 sg13g2_a21o_1 _12732_ (.A2(_04998_),
    .A1(_04996_),
    .B1(_05030_),
    .X(_05031_));
 sg13g2_and3_1 _12733_ (.X(_05032_),
    .A(_05026_),
    .B(_05029_),
    .C(_05031_));
 sg13g2_a21oi_1 _12734_ (.A1(_05029_),
    .A2(_05031_),
    .Y(_05033_),
    .B1(_05026_));
 sg13g2_or2_1 _12735_ (.X(_05034_),
    .B(_05033_),
    .A(_05032_));
 sg13g2_o21ai_1 _12736_ (.B1(net1947),
    .Y(_05035_),
    .A1(net1711),
    .A2(net2684));
 sg13g2_a21oi_1 _12737_ (.A1(net1711),
    .A2(_05034_),
    .Y(_00949_),
    .B1(_05035_));
 sg13g2_nand2_1 _12738_ (.Y(_05036_),
    .A(\am_sdr0.cic0.comb2_in_del[13] ),
    .B(_01265_));
 sg13g2_xor2_1 _12739_ (.B(net2746),
    .A(\am_sdr0.cic0.comb2_in_del[13] ),
    .X(_05037_));
 sg13g2_a21oi_1 _12740_ (.A1(_01266_),
    .A2(\am_sdr0.cic0.comb1[12] ),
    .Y(_05038_),
    .B1(_05033_));
 sg13g2_xnor2_1 _12741_ (.Y(_05039_),
    .A(_05037_),
    .B(_05038_));
 sg13g2_o21ai_1 _12742_ (.B1(net1947),
    .Y(_05040_),
    .A1(net1711),
    .A2(net2092));
 sg13g2_a21oi_1 _12743_ (.A1(net1711),
    .A2(net2747),
    .Y(_00950_),
    .B1(_05040_));
 sg13g2_nand2b_1 _12744_ (.Y(_05041_),
    .B(net2731),
    .A_N(\am_sdr0.cic0.comb2_in_del[14] ));
 sg13g2_xor2_1 _12745_ (.B(\am_sdr0.cic0.comb1[14] ),
    .A(\am_sdr0.cic0.comb2_in_del[14] ),
    .X(_05042_));
 sg13g2_nand3_1 _12746_ (.B(\am_sdr0.cic0.comb1[12] ),
    .C(_05036_),
    .A(_01266_),
    .Y(_05043_));
 sg13g2_o21ai_1 _12747_ (.B1(_05043_),
    .Y(_05044_),
    .A1(\am_sdr0.cic0.comb2_in_del[13] ),
    .A2(_01265_));
 sg13g2_a21oi_1 _12748_ (.A1(_05033_),
    .A2(_05036_),
    .Y(_05045_),
    .B1(_05044_));
 sg13g2_xnor2_1 _12749_ (.Y(_05046_),
    .A(_05042_),
    .B(_05045_));
 sg13g2_o21ai_1 _12750_ (.B1(net1944),
    .Y(_05047_),
    .A1(net1710),
    .A2(net2265));
 sg13g2_a21oi_1 _12751_ (.A1(net1710),
    .A2(_05046_),
    .Y(_00951_),
    .B1(_05047_));
 sg13g2_xor2_1 _12752_ (.B(\am_sdr0.cic0.comb1[15] ),
    .A(\am_sdr0.cic0.comb2_in_del[15] ),
    .X(_05048_));
 sg13g2_o21ai_1 _12753_ (.B1(_05041_),
    .Y(_05049_),
    .A1(_05042_),
    .A2(_05045_));
 sg13g2_xor2_1 _12754_ (.B(_05049_),
    .A(_05048_),
    .X(_05050_));
 sg13g2_o21ai_1 _12755_ (.B1(net1944),
    .Y(_05051_),
    .A1(net1710),
    .A2(net2633));
 sg13g2_a21oi_1 _12756_ (.A1(net1710),
    .A2(_05050_),
    .Y(_00952_),
    .B1(_05051_));
 sg13g2_nand2b_1 _12757_ (.Y(_05052_),
    .B(net2272),
    .A_N(\am_sdr0.cic0.comb2_in_del[16] ));
 sg13g2_xor2_1 _12758_ (.B(net2642),
    .A(\am_sdr0.cic0.comb2_in_del[16] ),
    .X(_05053_));
 sg13g2_nor2_1 _12759_ (.A(_05042_),
    .B(_05048_),
    .Y(_05054_));
 sg13g2_nor4_1 _12760_ (.A(_05026_),
    .B(_05037_),
    .C(_05042_),
    .D(_05048_),
    .Y(_05055_));
 sg13g2_a21oi_1 _12761_ (.A1(\am_sdr0.cic0.comb2_in_del[15] ),
    .A2(_01263_),
    .Y(_05056_),
    .B1(_05041_));
 sg13g2_a221oi_1 _12762_ (.B2(_05054_),
    .C1(_05056_),
    .B1(_05044_),
    .A1(_01262_),
    .Y(_05057_),
    .A2(\am_sdr0.cic0.comb1[15] ));
 sg13g2_nor2b_1 _12763_ (.A(_05055_),
    .B_N(_05057_),
    .Y(_05058_));
 sg13g2_and2_1 _12764_ (.A(_05029_),
    .B(_05057_),
    .X(_05059_));
 sg13g2_a21o_2 _12765_ (.A2(_05059_),
    .A1(_05031_),
    .B1(_05058_),
    .X(_05060_));
 sg13g2_xnor2_1 _12766_ (.Y(_05061_),
    .A(net2643),
    .B(_05060_));
 sg13g2_o21ai_1 _12767_ (.B1(net1944),
    .Y(_05062_),
    .A1(net1707),
    .A2(net2560));
 sg13g2_a21oi_1 _12768_ (.A1(net1707),
    .A2(_05061_),
    .Y(_00953_),
    .B1(_05062_));
 sg13g2_xnor2_1 _12769_ (.Y(_05063_),
    .A(\am_sdr0.cic0.comb2_in_del[17] ),
    .B(net2944));
 sg13g2_o21ai_1 _12770_ (.B1(_05052_),
    .Y(_05064_),
    .A1(_05053_),
    .A2(_05060_));
 sg13g2_xnor2_1 _12771_ (.Y(_05065_),
    .A(_05063_),
    .B(_05064_));
 sg13g2_o21ai_1 _12772_ (.B1(net1944),
    .Y(_05066_),
    .A1(net1707),
    .A2(net2550));
 sg13g2_a21oi_1 _12773_ (.A1(net1707),
    .A2(_05065_),
    .Y(_00954_),
    .B1(_05066_));
 sg13g2_nor2_1 _12774_ (.A(\am_sdr0.cic0.comb2_in_del[18] ),
    .B(_01258_),
    .Y(_05067_));
 sg13g2_xnor2_1 _12775_ (.Y(_05068_),
    .A(net2721),
    .B(net2589));
 sg13g2_nand2b_1 _12776_ (.Y(_05069_),
    .B(_05063_),
    .A_N(_05053_));
 sg13g2_a21oi_1 _12777_ (.A1(\am_sdr0.cic0.comb2_in_del[17] ),
    .A2(_01260_),
    .Y(_05070_),
    .B1(_05052_));
 sg13g2_a21oi_1 _12778_ (.A1(_01259_),
    .A2(\am_sdr0.cic0.comb1[17] ),
    .Y(_05071_),
    .B1(_05070_));
 sg13g2_o21ai_1 _12779_ (.B1(_05071_),
    .Y(_05072_),
    .A1(_05060_),
    .A2(_05069_));
 sg13g2_xnor2_1 _12780_ (.Y(_05073_),
    .A(_05068_),
    .B(_05072_));
 sg13g2_o21ai_1 _12781_ (.B1(net1924),
    .Y(_05074_),
    .A1(net1708),
    .A2(net2201));
 sg13g2_a21oi_1 _12782_ (.A1(net1708),
    .A2(_05073_),
    .Y(_00955_),
    .B1(_05074_));
 sg13g2_a21oi_1 _12783_ (.A1(_05068_),
    .A2(_05072_),
    .Y(_05075_),
    .B1(_05067_));
 sg13g2_xnor2_1 _12784_ (.Y(_05076_),
    .A(net2487),
    .B(net2123));
 sg13g2_or2_1 _12785_ (.X(_05077_),
    .B(_05076_),
    .A(_05075_));
 sg13g2_a21oi_1 _12786_ (.A1(_05075_),
    .A2(_05076_),
    .Y(_05078_),
    .B1(net1642));
 sg13g2_a221oi_1 _12787_ (.B2(_05078_),
    .C1(net1878),
    .B1(net2488),
    .A1(_01222_),
    .Y(_00956_),
    .A2(net1642));
 sg13g2_o21ai_1 _12788_ (.B1(net1956),
    .Y(_05079_),
    .A1(net1724),
    .A2(net2377));
 sg13g2_a21oi_1 _12789_ (.A1(net1724),
    .A2(_01280_),
    .Y(_00957_),
    .B1(_05079_));
 sg13g2_o21ai_1 _12790_ (.B1(net1956),
    .Y(_05080_),
    .A1(net1724),
    .A2(net2672));
 sg13g2_a21oi_1 _12791_ (.A1(net1724),
    .A2(_01278_),
    .Y(_00958_),
    .B1(_05080_));
 sg13g2_o21ai_1 _12792_ (.B1(net1956),
    .Y(_05081_),
    .A1(net1723),
    .A2(\am_sdr0.cic0.comb2_in_del[2] ));
 sg13g2_a21oi_1 _12793_ (.A1(net1723),
    .A2(_01277_),
    .Y(_00959_),
    .B1(_05081_));
 sg13g2_o21ai_1 _12794_ (.B1(net1956),
    .Y(_05082_),
    .A1(net1723),
    .A2(net2572));
 sg13g2_a21oi_1 _12795_ (.A1(net1723),
    .A2(_01276_),
    .Y(_00960_),
    .B1(_05082_));
 sg13g2_o21ai_1 _12796_ (.B1(net1955),
    .Y(_05083_),
    .A1(net1725),
    .A2(net2828));
 sg13g2_a21oi_1 _12797_ (.A1(net1722),
    .A2(_01275_),
    .Y(_00961_),
    .B1(_05083_));
 sg13g2_o21ai_1 _12798_ (.B1(net1955),
    .Y(_05084_),
    .A1(net1722),
    .A2(\am_sdr0.cic0.comb2_in_del[5] ));
 sg13g2_a21oi_1 _12799_ (.A1(net1722),
    .A2(_01274_),
    .Y(_00962_),
    .B1(_05084_));
 sg13g2_o21ai_1 _12800_ (.B1(net1955),
    .Y(_05085_),
    .A1(net1718),
    .A2(\am_sdr0.cic0.comb2_in_del[6] ));
 sg13g2_a21oi_1 _12801_ (.A1(net1718),
    .A2(_01273_),
    .Y(_00963_),
    .B1(_05085_));
 sg13g2_o21ai_1 _12802_ (.B1(net1955),
    .Y(_05086_),
    .A1(net1718),
    .A2(\am_sdr0.cic0.comb2_in_del[7] ));
 sg13g2_a21oi_1 _12803_ (.A1(net1718),
    .A2(_01272_),
    .Y(_00964_),
    .B1(_05086_));
 sg13g2_o21ai_1 _12804_ (.B1(net1955),
    .Y(_05087_),
    .A1(net1719),
    .A2(net2717));
 sg13g2_a21oi_1 _12805_ (.A1(net1718),
    .A2(_01271_),
    .Y(_00965_),
    .B1(_05087_));
 sg13g2_o21ai_1 _12806_ (.B1(net1947),
    .Y(_05088_),
    .A1(net1719),
    .A2(\am_sdr0.cic0.comb2_in_del[9] ));
 sg13g2_a21oi_1 _12807_ (.A1(net1719),
    .A2(_01270_),
    .Y(_00966_),
    .B1(_05088_));
 sg13g2_o21ai_1 _12808_ (.B1(net1947),
    .Y(_05089_),
    .A1(net1717),
    .A2(\am_sdr0.cic0.comb2_in_del[10] ));
 sg13g2_a21oi_1 _12809_ (.A1(net1717),
    .A2(_01268_),
    .Y(_00967_),
    .B1(_05089_));
 sg13g2_o21ai_1 _12810_ (.B1(net1947),
    .Y(_05090_),
    .A1(net1704),
    .A2(net2283));
 sg13g2_a21oi_1 _12811_ (.A1(net1704),
    .A2(_01267_),
    .Y(_00968_),
    .B1(_05090_));
 sg13g2_o21ai_1 _12812_ (.B1(net1947),
    .Y(_05091_),
    .A1(net1642),
    .A2(\am_sdr0.cic0.comb1[12] ));
 sg13g2_a21oi_1 _12813_ (.A1(net1642),
    .A2(_01266_),
    .Y(_00969_),
    .B1(_05091_));
 sg13g2_o21ai_1 _12814_ (.B1(net1945),
    .Y(_05092_),
    .A1(net1703),
    .A2(net2873));
 sg13g2_a21oi_1 _12815_ (.A1(net1703),
    .A2(_01265_),
    .Y(_00970_),
    .B1(_05092_));
 sg13g2_o21ai_1 _12816_ (.B1(net1945),
    .Y(_05093_),
    .A1(net1704),
    .A2(\am_sdr0.cic0.comb2_in_del[14] ));
 sg13g2_a21oi_1 _12817_ (.A1(net1704),
    .A2(_01264_),
    .Y(_00971_),
    .B1(_05093_));
 sg13g2_o21ai_1 _12818_ (.B1(net1944),
    .Y(_05094_),
    .A1(net1710),
    .A2(\am_sdr0.cic0.comb2_in_del[15] ));
 sg13g2_a21oi_1 _12819_ (.A1(net1710),
    .A2(_01263_),
    .Y(_00972_),
    .B1(_05094_));
 sg13g2_o21ai_1 _12820_ (.B1(net1944),
    .Y(_05095_),
    .A1(net1701),
    .A2(\am_sdr0.cic0.comb2_in_del[16] ));
 sg13g2_a21oi_1 _12821_ (.A1(net1701),
    .A2(_01261_),
    .Y(_00973_),
    .B1(_05095_));
 sg13g2_o21ai_1 _12822_ (.B1(net1923),
    .Y(_05096_),
    .A1(net1701),
    .A2(\am_sdr0.cic0.comb2_in_del[17] ));
 sg13g2_a21oi_1 _12823_ (.A1(net1701),
    .A2(_01260_),
    .Y(_00974_),
    .B1(_05096_));
 sg13g2_o21ai_1 _12824_ (.B1(net1923),
    .Y(_05097_),
    .A1(net1700),
    .A2(\am_sdr0.cic0.comb2_in_del[18] ));
 sg13g2_a21oi_1 _12825_ (.A1(net1700),
    .A2(_01258_),
    .Y(_00975_),
    .B1(_05097_));
 sg13g2_o21ai_1 _12826_ (.B1(net1923),
    .Y(_05098_),
    .A1(net1700),
    .A2(\am_sdr0.cic0.comb2_in_del[19] ));
 sg13g2_a21oi_1 _12827_ (.A1(net1700),
    .A2(_01257_),
    .Y(_00976_),
    .B1(_05098_));
 sg13g2_nand2_1 _12828_ (.Y(_05099_),
    .A(\am_sdr0.cic0.comb3_in_del[4] ),
    .B(_01244_));
 sg13g2_nand2b_1 _12829_ (.Y(_05100_),
    .B(\am_sdr0.cic0.comb3_in_del[1] ),
    .A_N(\am_sdr0.cic0.comb2[1] ));
 sg13g2_nand2b_1 _12830_ (.Y(_05101_),
    .B(\am_sdr0.cic0.comb3_in_del[0] ),
    .A_N(\am_sdr0.cic0.comb2[0] ));
 sg13g2_nor2b_1 _12831_ (.A(\am_sdr0.cic0.comb3_in_del[1] ),
    .B_N(\am_sdr0.cic0.comb2[1] ),
    .Y(_05102_));
 sg13g2_a221oi_1 _12832_ (.B2(_05101_),
    .C1(_05102_),
    .B1(_05100_),
    .A1(_01246_),
    .Y(_05103_),
    .A2(\am_sdr0.cic0.comb2[2] ));
 sg13g2_nand2b_1 _12833_ (.Y(_05104_),
    .B(\am_sdr0.cic0.comb3_in_del[3] ),
    .A_N(\am_sdr0.cic0.comb2[3] ));
 sg13g2_o21ai_1 _12834_ (.B1(_05104_),
    .Y(_05105_),
    .A1(_01246_),
    .A2(\am_sdr0.cic0.comb2[2] ));
 sg13g2_a22oi_1 _12835_ (.Y(_05106_),
    .B1(_01245_),
    .B2(\am_sdr0.cic0.comb2[3] ),
    .A2(\am_sdr0.cic0.comb2[4] ),
    .A1(_01243_));
 sg13g2_o21ai_1 _12836_ (.B1(_05106_),
    .Y(_05107_),
    .A1(_05103_),
    .A2(_05105_));
 sg13g2_a22oi_1 _12837_ (.Y(_05108_),
    .B1(_05099_),
    .B2(_05107_),
    .A2(\am_sdr0.cic0.comb2[5] ),
    .A1(_01241_));
 sg13g2_nand2_1 _12838_ (.Y(_05109_),
    .A(\am_sdr0.cic0.comb3_in_del[6] ),
    .B(_01240_));
 sg13g2_o21ai_1 _12839_ (.B1(_05109_),
    .Y(_05110_),
    .A1(_01241_),
    .A2(\am_sdr0.cic0.comb2[5] ));
 sg13g2_a22oi_1 _12840_ (.Y(_05111_),
    .B1(_01239_),
    .B2(\am_sdr0.cic0.comb2[6] ),
    .A2(\am_sdr0.cic0.comb2[7] ),
    .A1(_01237_));
 sg13g2_o21ai_1 _12841_ (.B1(_05111_),
    .Y(_05112_),
    .A1(_05108_),
    .A2(_05110_));
 sg13g2_a22oi_1 _12842_ (.Y(_05113_),
    .B1(\am_sdr0.cic0.comb3_in_del[10] ),
    .B2(_01233_),
    .A2(\am_sdr0.cic0.comb2[11] ),
    .A1(_01231_));
 sg13g2_o21ai_1 _12843_ (.B1(_05113_),
    .Y(_05114_),
    .A1(_01234_),
    .A2(\am_sdr0.cic0.comb2[9] ));
 sg13g2_a22oi_1 _12844_ (.Y(_05115_),
    .B1(_01235_),
    .B2(\am_sdr0.cic0.comb2[8] ),
    .A2(\am_sdr0.cic0.comb2[9] ),
    .A1(_01234_));
 sg13g2_nor2_1 _12845_ (.A(\am_sdr0.cic0.comb3_in_del[10] ),
    .B(_01233_),
    .Y(_05116_));
 sg13g2_a21oi_1 _12846_ (.A1(\am_sdr0.cic0.comb3_in_del[8] ),
    .A2(_01236_),
    .Y(_05117_),
    .B1(_05116_));
 sg13g2_nand2_1 _12847_ (.Y(_05118_),
    .A(\am_sdr0.cic0.comb3_in_del[7] ),
    .B(_01238_));
 sg13g2_nand2_1 _12848_ (.Y(_05119_),
    .A(\am_sdr0.cic0.comb3_in_del[11] ),
    .B(_01232_));
 sg13g2_nand4_1 _12849_ (.B(_05117_),
    .C(_05118_),
    .A(_05115_),
    .Y(_05120_),
    .D(_05119_));
 sg13g2_nor2_1 _12850_ (.A(_05114_),
    .B(_05120_),
    .Y(_05121_));
 sg13g2_a21oi_1 _12851_ (.A1(_01231_),
    .A2(\am_sdr0.cic0.comb2[11] ),
    .Y(_05122_),
    .B1(_05116_));
 sg13g2_o21ai_1 _12852_ (.B1(_05122_),
    .Y(_05123_),
    .A1(_05114_),
    .A2(_05115_));
 sg13g2_a22oi_1 _12853_ (.Y(_05124_),
    .B1(_05123_),
    .B2(_05119_),
    .A2(_05121_),
    .A1(_05112_));
 sg13g2_xor2_1 _12854_ (.B(\am_sdr0.cic0.comb2[12] ),
    .A(net2289),
    .X(_05125_));
 sg13g2_inv_1 _12855_ (.Y(_05126_),
    .A(_05125_));
 sg13g2_nor2_1 _12856_ (.A(_05124_),
    .B(_05125_),
    .Y(_05127_));
 sg13g2_xnor2_1 _12857_ (.Y(_05128_),
    .A(_05124_),
    .B(_05125_));
 sg13g2_o21ai_1 _12858_ (.B1(net1948),
    .Y(_05129_),
    .A1(net1728),
    .A2(net1503));
 sg13g2_a21oi_1 _12859_ (.A1(net1728),
    .A2(_05128_),
    .Y(_00977_),
    .B1(_05129_));
 sg13g2_nand2_1 _12860_ (.Y(_05130_),
    .A(\am_sdr0.cic0.comb3_in_del[13] ),
    .B(_01229_));
 sg13g2_xnor2_1 _12861_ (.Y(_05131_),
    .A(\am_sdr0.cic0.comb3_in_del[13] ),
    .B(net2092));
 sg13g2_a21oi_1 _12862_ (.A1(_01230_),
    .A2(net3298),
    .Y(_05132_),
    .B1(_05127_));
 sg13g2_or2_1 _12863_ (.X(_05133_),
    .B(_05132_),
    .A(_05131_));
 sg13g2_a21oi_1 _12864_ (.A1(_05131_),
    .A2(_05132_),
    .Y(_05134_),
    .B1(net1643));
 sg13g2_a221oi_1 _12865_ (.B2(_05134_),
    .C1(net1886),
    .B1(_05133_),
    .A1(net1643),
    .Y(_00978_),
    .A2(_01255_));
 sg13g2_nand2b_1 _12866_ (.Y(_05135_),
    .B(net2390),
    .A_N(\am_sdr0.cic0.comb3_in_del[14] ));
 sg13g2_inv_1 _12867_ (.Y(_05136_),
    .A(_05135_));
 sg13g2_nand2_1 _12868_ (.Y(_05137_),
    .A(\am_sdr0.cic0.comb3_in_del[14] ),
    .B(_01228_));
 sg13g2_nand2_1 _12869_ (.Y(_05138_),
    .A(_05135_),
    .B(_05137_));
 sg13g2_nand3_1 _12870_ (.B(\am_sdr0.cic0.comb2[12] ),
    .C(_05130_),
    .A(_01230_),
    .Y(_05139_));
 sg13g2_o21ai_1 _12871_ (.B1(_05139_),
    .Y(_05140_),
    .A1(\am_sdr0.cic0.comb3_in_del[13] ),
    .A2(_01229_));
 sg13g2_nand3b_1 _12872_ (.B(_05126_),
    .C(_05131_),
    .Y(_05141_),
    .A_N(_05124_));
 sg13g2_nand2b_1 _12873_ (.Y(_05142_),
    .B(_05141_),
    .A_N(_05140_));
 sg13g2_xor2_1 _12874_ (.B(_05142_),
    .A(_05138_),
    .X(_05143_));
 sg13g2_o21ai_1 _12875_ (.B1(net1948),
    .Y(_05144_),
    .A1(net1712),
    .A2(net1478));
 sg13g2_a21oi_1 _12876_ (.A1(net1712),
    .A2(_05143_),
    .Y(_00979_),
    .B1(_05144_));
 sg13g2_nand2b_1 _12877_ (.Y(_05145_),
    .B(net3300),
    .A_N(net2143));
 sg13g2_nand2_1 _12878_ (.Y(_05146_),
    .A(net2143),
    .B(_01227_));
 sg13g2_a21oi_1 _12879_ (.A1(_05137_),
    .A2(_05142_),
    .Y(_05147_),
    .B1(_05136_));
 sg13g2_a21oi_1 _12880_ (.A1(_05145_),
    .A2(_05146_),
    .Y(_05148_),
    .B1(_05147_));
 sg13g2_nand3_1 _12881_ (.B(_05146_),
    .C(_05147_),
    .A(_05145_),
    .Y(_05149_));
 sg13g2_nor2_1 _12882_ (.A(net1642),
    .B(_05148_),
    .Y(_05150_));
 sg13g2_a221oi_1 _12883_ (.B2(_05150_),
    .C1(net1886),
    .B1(net2144),
    .A1(net1642),
    .Y(_00980_),
    .A2(_01253_));
 sg13g2_nor2_1 _12884_ (.A(net2218),
    .B(_01226_),
    .Y(_05151_));
 sg13g2_xnor2_1 _12885_ (.Y(_05152_),
    .A(\am_sdr0.cic0.comb3_in_del[16] ),
    .B(\am_sdr0.cic0.comb2[16] ));
 sg13g2_nor2b_1 _12886_ (.A(_05137_),
    .B_N(_05145_),
    .Y(_05153_));
 sg13g2_nand2_1 _12887_ (.Y(_05154_),
    .A(_05136_),
    .B(_05146_));
 sg13g2_nand2_1 _12888_ (.Y(_05155_),
    .A(_05145_),
    .B(_05154_));
 sg13g2_nor2_1 _12889_ (.A(_05140_),
    .B(_05155_),
    .Y(_05156_));
 sg13g2_a221oi_1 _12890_ (.B2(_05156_),
    .C1(_05153_),
    .B1(_05141_),
    .A1(net2153),
    .Y(_05157_),
    .A2(_01227_));
 sg13g2_xnor2_1 _12891_ (.Y(_05158_),
    .A(_05152_),
    .B(_05157_));
 sg13g2_o21ai_1 _12892_ (.B1(net1945),
    .Y(_05159_),
    .A1(net1712),
    .A2(net1269));
 sg13g2_a21oi_1 _12893_ (.A1(net1712),
    .A2(net2154),
    .Y(_00981_),
    .B1(_05159_));
 sg13g2_a21oi_1 _12894_ (.A1(_05152_),
    .A2(_05157_),
    .Y(_05160_),
    .B1(_05151_));
 sg13g2_nand2b_1 _12895_ (.Y(_05161_),
    .B(\am_sdr0.cic0.comb2[17] ),
    .A_N(\am_sdr0.cic0.comb3_in_del[17] ));
 sg13g2_nor2b_1 _12896_ (.A(net3303),
    .B_N(\am_sdr0.cic0.comb3_in_del[17] ),
    .Y(_05162_));
 sg13g2_xnor2_1 _12897_ (.Y(_05163_),
    .A(\am_sdr0.cic0.comb3_in_del[17] ),
    .B(\am_sdr0.cic0.comb2[17] ));
 sg13g2_o21ai_1 _12898_ (.B1(net1707),
    .Y(_05164_),
    .A1(_05160_),
    .A2(_05163_));
 sg13g2_a21oi_1 _12899_ (.A1(_05160_),
    .A2(_05163_),
    .Y(_05165_),
    .B1(_05164_));
 sg13g2_o21ai_1 _12900_ (.B1(net1946),
    .Y(_05166_),
    .A1(net1709),
    .A2(net1306));
 sg13g2_nor2_1 _12901_ (.A(net2219),
    .B(_05166_),
    .Y(_00982_));
 sg13g2_nor2_1 _12902_ (.A(\am_sdr0.cic0.comb3_in_del[18] ),
    .B(_01224_),
    .Y(_05167_));
 sg13g2_xnor2_1 _12903_ (.Y(_05168_),
    .A(\am_sdr0.cic0.comb3_in_del[18] ),
    .B(net2201));
 sg13g2_a21oi_1 _12904_ (.A1(_05160_),
    .A2(_05161_),
    .Y(_05169_),
    .B1(_05162_));
 sg13g2_xnor2_1 _12905_ (.Y(_05170_),
    .A(net2202),
    .B(_05169_));
 sg13g2_o21ai_1 _12906_ (.B1(net1924),
    .Y(_05171_),
    .A1(net1709),
    .A2(net1293));
 sg13g2_a21oi_1 _12907_ (.A1(net1708),
    .A2(_05170_),
    .Y(_00983_),
    .B1(_05171_));
 sg13g2_a21oi_1 _12908_ (.A1(_05168_),
    .A2(_05169_),
    .Y(_05172_),
    .B1(_05167_));
 sg13g2_xnor2_1 _12909_ (.Y(_05173_),
    .A(\am_sdr0.cic0.comb3_in_del[19] ),
    .B(net2133));
 sg13g2_or2_1 _12910_ (.X(_05174_),
    .B(net2134),
    .A(_05172_));
 sg13g2_a21oi_1 _12911_ (.A1(_05172_),
    .A2(net2134),
    .Y(_05175_),
    .B1(net1646));
 sg13g2_a221oi_1 _12912_ (.B2(_05175_),
    .C1(net1878),
    .B1(_05174_),
    .A1(net1646),
    .Y(_00984_),
    .A2(_01249_));
 sg13g2_o21ai_1 _12913_ (.B1(net1956),
    .Y(_05176_),
    .A1(net1731),
    .A2(\am_sdr0.cic0.comb3_in_del[0] ));
 sg13g2_a21oi_1 _12914_ (.A1(net1731),
    .A2(_01248_),
    .Y(_00985_),
    .B1(_05176_));
 sg13g2_o21ai_1 _12915_ (.B1(net1957),
    .Y(_05177_),
    .A1(net1731),
    .A2(\am_sdr0.cic0.comb3_in_del[1] ));
 sg13g2_a21oi_1 _12916_ (.A1(net1731),
    .A2(_01247_),
    .Y(_00986_),
    .B1(_05177_));
 sg13g2_o21ai_1 _12917_ (.B1(net1957),
    .Y(_05178_),
    .A1(net1644),
    .A2(\am_sdr0.cic0.comb2[2] ));
 sg13g2_a21oi_1 _12918_ (.A1(net1644),
    .A2(_01246_),
    .Y(_00987_),
    .B1(_05178_));
 sg13g2_o21ai_1 _12919_ (.B1(net1957),
    .Y(_05179_),
    .A1(net1644),
    .A2(\am_sdr0.cic0.comb2[3] ));
 sg13g2_a21oi_1 _12920_ (.A1(net1644),
    .A2(_01245_),
    .Y(_00988_),
    .B1(_05179_));
 sg13g2_o21ai_1 _12921_ (.B1(net1954),
    .Y(_05180_),
    .A1(net1733),
    .A2(net2457));
 sg13g2_a21oi_1 _12922_ (.A1(net1733),
    .A2(_01244_),
    .Y(_00989_),
    .B1(_05180_));
 sg13g2_o21ai_1 _12923_ (.B1(net1954),
    .Y(_05181_),
    .A1(net1733),
    .A2(net2275));
 sg13g2_a21oi_1 _12924_ (.A1(net1733),
    .A2(_01242_),
    .Y(_00990_),
    .B1(_05181_));
 sg13g2_o21ai_1 _12925_ (.B1(net1958),
    .Y(_05182_),
    .A1(net1733),
    .A2(net2417));
 sg13g2_a21oi_1 _12926_ (.A1(net1733),
    .A2(_01240_),
    .Y(_00991_),
    .B1(_05182_));
 sg13g2_o21ai_1 _12927_ (.B1(net1954),
    .Y(_05183_),
    .A1(net1728),
    .A2(net2501));
 sg13g2_a21oi_1 _12928_ (.A1(net1728),
    .A2(_01238_),
    .Y(_00992_),
    .B1(_05183_));
 sg13g2_o21ai_1 _12929_ (.B1(net1954),
    .Y(_05184_),
    .A1(net1729),
    .A2(\am_sdr0.cic0.comb3_in_del[8] ));
 sg13g2_a21oi_1 _12930_ (.A1(net1729),
    .A2(_01236_),
    .Y(_00993_),
    .B1(_05184_));
 sg13g2_o21ai_1 _12931_ (.B1(net1954),
    .Y(_05185_),
    .A1(net1643),
    .A2(\am_sdr0.cic0.comb2[9] ));
 sg13g2_a21oi_1 _12932_ (.A1(net1643),
    .A2(_01234_),
    .Y(_00994_),
    .B1(_05185_));
 sg13g2_o21ai_1 _12933_ (.B1(net1948),
    .Y(_05186_),
    .A1(net1727),
    .A2(net2544));
 sg13g2_a21oi_1 _12934_ (.A1(net1727),
    .A2(_01233_),
    .Y(_00995_),
    .B1(_05186_));
 sg13g2_o21ai_1 _12935_ (.B1(net1954),
    .Y(_05187_),
    .A1(net1728),
    .A2(net2429));
 sg13g2_a21oi_1 _12936_ (.A1(net1728),
    .A2(_01232_),
    .Y(_00996_),
    .B1(_05187_));
 sg13g2_o21ai_1 _12937_ (.B1(net1948),
    .Y(_05188_),
    .A1(net1643),
    .A2(net2684));
 sg13g2_a21oi_1 _12938_ (.A1(net1643),
    .A2(_01230_),
    .Y(_00997_),
    .B1(_05188_));
 sg13g2_o21ai_1 _12939_ (.B1(net1948),
    .Y(_05189_),
    .A1(net1710),
    .A2(net2924));
 sg13g2_a21oi_1 _12940_ (.A1(net1710),
    .A2(_01229_),
    .Y(_00998_),
    .B1(_05189_));
 sg13g2_o21ai_1 _12941_ (.B1(net1948),
    .Y(_05190_),
    .A1(net1711),
    .A2(\am_sdr0.cic0.comb3_in_del[14] ));
 sg13g2_a21oi_1 _12942_ (.A1(net1711),
    .A2(_01228_),
    .Y(_00999_),
    .B1(_05190_));
 sg13g2_o21ai_1 _12943_ (.B1(net1945),
    .Y(_05191_),
    .A1(net1712),
    .A2(net2143));
 sg13g2_a21oi_1 _12944_ (.A1(net1712),
    .A2(_01227_),
    .Y(_01000_),
    .B1(_05191_));
 sg13g2_o21ai_1 _12945_ (.B1(net1944),
    .Y(_05192_),
    .A1(net1707),
    .A2(net2218));
 sg13g2_a21oi_1 _12946_ (.A1(net1707),
    .A2(_01226_),
    .Y(_01001_),
    .B1(_05192_));
 sg13g2_o21ai_1 _12947_ (.B1(net1944),
    .Y(_05193_),
    .A1(net1707),
    .A2(\am_sdr0.cic0.comb3_in_del[17] ));
 sg13g2_a21oi_1 _12948_ (.A1(net1709),
    .A2(_01225_),
    .Y(_01002_),
    .B1(_05193_));
 sg13g2_o21ai_1 _12949_ (.B1(net1923),
    .Y(_05194_),
    .A1(net1708),
    .A2(net2419));
 sg13g2_a21oi_1 _12950_ (.A1(net1708),
    .A2(_01224_),
    .Y(_01003_),
    .B1(_05194_));
 sg13g2_o21ai_1 _12951_ (.B1(net1923),
    .Y(_05195_),
    .A1(net2165),
    .A2(net1708));
 sg13g2_a21oi_1 _12952_ (.A1(_01222_),
    .A2(net1708),
    .Y(_01004_),
    .B1(_05195_));
 sg13g2_o21ai_1 _12953_ (.B1(net1957),
    .Y(_05196_),
    .A1(_03953_),
    .A2(_03954_));
 sg13g2_nor2_1 _12954_ (.A(_01595_),
    .B(_05196_),
    .Y(_01006_));
 sg13g2_xnor2_1 _12955_ (.Y(_05197_),
    .A(\am_sdr0.cic0.count[0] ),
    .B(net2253));
 sg13g2_nor2_1 _12956_ (.A(_05196_),
    .B(net2254),
    .Y(_01007_));
 sg13g2_a21oi_1 _12957_ (.A1(\am_sdr0.cic0.count[0] ),
    .A2(\am_sdr0.cic0.count[1] ),
    .Y(_05198_),
    .B1(net1219));
 sg13g2_nor3_1 _12958_ (.A(_03950_),
    .B(_05196_),
    .C(net1220),
    .Y(_01008_));
 sg13g2_nor2_1 _12959_ (.A(net2033),
    .B(_03950_),
    .Y(_05199_));
 sg13g2_nor3_1 _12960_ (.A(net1885),
    .B(_03951_),
    .C(net2034),
    .Y(_01009_));
 sg13g2_nor2_1 _12961_ (.A(net1425),
    .B(_03951_),
    .Y(_05200_));
 sg13g2_nor3_1 _12962_ (.A(net1885),
    .B(_03952_),
    .C(net1426),
    .Y(_01010_));
 sg13g2_o21ai_1 _12963_ (.B1(net1957),
    .Y(_05201_),
    .A1(net2810),
    .A2(_03952_));
 sg13g2_nor2b_1 _12964_ (.A(_05201_),
    .B_N(_03953_),
    .Y(_01011_));
 sg13g2_a21oi_1 _12965_ (.A1(\am_sdr0.cic0.count[5] ),
    .A2(_03952_),
    .Y(_05202_),
    .B1(net1410));
 sg13g2_and3_1 _12966_ (.X(_05203_),
    .A(\am_sdr0.cic0.count[5] ),
    .B(net1410),
    .C(_03952_));
 sg13g2_nor3_1 _12967_ (.A(_05196_),
    .B(net1411),
    .C(_05203_),
    .Y(_01012_));
 sg13g2_o21ai_1 _12968_ (.B1(net1957),
    .Y(_05204_),
    .A1(net1252),
    .A2(_05203_));
 sg13g2_a21oi_1 _12969_ (.A1(net1252),
    .A2(_05203_),
    .Y(_01013_),
    .B1(_05204_));
 sg13g2_nand2_1 _12970_ (.Y(_05205_),
    .A(net3162),
    .B(net2459));
 sg13g2_o21ai_1 _12971_ (.B1(net1927),
    .Y(_05206_),
    .A1(\am_sdr0.I_out[0] ),
    .A2(net2459));
 sg13g2_nor2b_1 _12972_ (.A(net2460),
    .B_N(_05205_),
    .Y(_01014_));
 sg13g2_nand2_1 _12973_ (.Y(_05207_),
    .A(\am_sdr0.I_out[1] ),
    .B(\am_sdr0.cic0.integ1[1] ));
 sg13g2_xnor2_1 _12974_ (.Y(_05208_),
    .A(net3044),
    .B(\am_sdr0.cic0.integ1[1] ));
 sg13g2_and2_1 _12975_ (.A(_05205_),
    .B(_05208_),
    .X(_05209_));
 sg13g2_nor2_1 _12976_ (.A(_05205_),
    .B(_05208_),
    .Y(_05210_));
 sg13g2_nor3_1 _12977_ (.A(net1879),
    .B(net3163),
    .C(_05210_),
    .Y(_01015_));
 sg13g2_and2_1 _12978_ (.A(net3286),
    .B(\am_sdr0.cic0.integ1[2] ),
    .X(_05211_));
 sg13g2_xnor2_1 _12979_ (.Y(_05212_),
    .A(\am_sdr0.I_out[2] ),
    .B(\am_sdr0.cic0.integ1[2] ));
 sg13g2_inv_1 _12980_ (.Y(_05213_),
    .A(_05212_));
 sg13g2_a21oi_1 _12981_ (.A1(net3044),
    .A2(\am_sdr0.cic0.integ1[1] ),
    .Y(_05214_),
    .B1(_05210_));
 sg13g2_o21ai_1 _12982_ (.B1(_05207_),
    .Y(_05215_),
    .A1(_05205_),
    .A2(_05208_));
 sg13g2_o21ai_1 _12983_ (.B1(net1930),
    .Y(_05216_),
    .A1(_05212_),
    .A2(net3045));
 sg13g2_a21oi_1 _12984_ (.A1(_05212_),
    .A2(net3045),
    .Y(_01016_),
    .B1(_05216_));
 sg13g2_nand2_1 _12985_ (.Y(_05217_),
    .A(\am_sdr0.cic0.integ1[3] ),
    .B(\am_sdr0.I_out[3] ));
 sg13g2_xnor2_1 _12986_ (.Y(_05218_),
    .A(\am_sdr0.cic0.integ1[3] ),
    .B(net3249));
 sg13g2_a21oi_1 _12987_ (.A1(_05213_),
    .A2(_05215_),
    .Y(_05219_),
    .B1(_05211_));
 sg13g2_nor2_1 _12988_ (.A(_05218_),
    .B(_05219_),
    .Y(_05220_));
 sg13g2_a21oi_1 _12989_ (.A1(_05218_),
    .A2(_05219_),
    .Y(_05221_),
    .B1(net1879));
 sg13g2_nor2b_1 _12990_ (.A(_05220_),
    .B_N(_05221_),
    .Y(_01017_));
 sg13g2_a21oi_1 _12991_ (.A1(net2845),
    .A2(net3249),
    .Y(_05222_),
    .B1(_05220_));
 sg13g2_o21ai_1 _12992_ (.B1(_05217_),
    .Y(_05223_),
    .A1(_05218_),
    .A2(_05219_));
 sg13g2_xnor2_1 _12993_ (.Y(_05224_),
    .A(\am_sdr0.cic0.integ1[4] ),
    .B(net3102));
 sg13g2_nor2_1 _12994_ (.A(_05222_),
    .B(_05224_),
    .Y(_05225_));
 sg13g2_a21oi_1 _12995_ (.A1(_05222_),
    .A2(_05224_),
    .Y(_05226_),
    .B1(net1879));
 sg13g2_nor2b_1 _12996_ (.A(_05225_),
    .B_N(_05226_),
    .Y(_01018_));
 sg13g2_nand2_1 _12997_ (.Y(_05227_),
    .A(\am_sdr0.cic0.integ1[5] ),
    .B(\am_sdr0.I_out[5] ));
 sg13g2_or2_1 _12998_ (.X(_05228_),
    .B(\am_sdr0.I_out[5] ),
    .A(\am_sdr0.cic0.integ1[5] ));
 sg13g2_nand2_1 _12999_ (.Y(_05229_),
    .A(_05227_),
    .B(_05228_));
 sg13g2_a21oi_1 _13000_ (.A1(\am_sdr0.cic0.integ1[4] ),
    .A2(net3102),
    .Y(_05230_),
    .B1(_05225_));
 sg13g2_o21ai_1 _13001_ (.B1(net1932),
    .Y(_05231_),
    .A1(_05229_),
    .A2(net3103));
 sg13g2_a21oi_1 _13002_ (.A1(_05229_),
    .A2(net3103),
    .Y(_01019_),
    .B1(_05231_));
 sg13g2_nand2_1 _13003_ (.Y(_05232_),
    .A(\am_sdr0.cic0.integ1[6] ),
    .B(\am_sdr0.I_out[6] ));
 sg13g2_xnor2_1 _13004_ (.Y(_05233_),
    .A(\am_sdr0.cic0.integ1[6] ),
    .B(net3134));
 sg13g2_nor2_1 _13005_ (.A(_05224_),
    .B(_05229_),
    .Y(_05234_));
 sg13g2_nand3_1 _13006_ (.B(net3102),
    .C(_05228_),
    .A(\am_sdr0.cic0.integ1[4] ),
    .Y(_05235_));
 sg13g2_nand2_1 _13007_ (.Y(_05236_),
    .A(_05227_),
    .B(_05235_));
 sg13g2_a21oi_2 _13008_ (.B1(_05236_),
    .Y(_05237_),
    .A2(_05234_),
    .A1(_05223_));
 sg13g2_o21ai_1 _13009_ (.B1(net1936),
    .Y(_05238_),
    .A1(_05233_),
    .A2(_05237_));
 sg13g2_a21oi_1 _13010_ (.A1(net3135),
    .A2(_05237_),
    .Y(_01020_),
    .B1(_05238_));
 sg13g2_and2_1 _13011_ (.A(\am_sdr0.cic0.integ1[7] ),
    .B(net1667),
    .X(_05239_));
 sg13g2_or2_1 _13012_ (.X(_05240_),
    .B(net1667),
    .A(\am_sdr0.cic0.integ1[7] ));
 sg13g2_nand2b_1 _13013_ (.Y(_05241_),
    .B(_05240_),
    .A_N(_05239_));
 sg13g2_o21ai_1 _13014_ (.B1(_05232_),
    .Y(_05242_),
    .A1(_05233_),
    .A2(_05237_));
 sg13g2_nand2b_1 _13015_ (.Y(_05243_),
    .B(_05241_),
    .A_N(_05242_));
 sg13g2_nand2b_1 _13016_ (.Y(_05244_),
    .B(_05242_),
    .A_N(_05241_));
 sg13g2_and3_1 _13017_ (.X(_01021_),
    .A(net1936),
    .B(_05243_),
    .C(_05244_));
 sg13g2_a21oi_1 _13018_ (.A1(_05240_),
    .A2(_05242_),
    .Y(_05245_),
    .B1(_05239_));
 sg13g2_a21o_1 _13019_ (.A2(_05242_),
    .A1(_05240_),
    .B1(_05239_),
    .X(_05246_));
 sg13g2_nand2_1 _13020_ (.Y(_05247_),
    .A(net3269),
    .B(net1666));
 sg13g2_xnor2_1 _13021_ (.Y(_05248_),
    .A(\am_sdr0.cic0.integ1[8] ),
    .B(net1666));
 sg13g2_nand2b_1 _13022_ (.Y(_05249_),
    .B(_05246_),
    .A_N(_05248_));
 sg13g2_nand2_1 _13023_ (.Y(_05250_),
    .A(net1936),
    .B(_05249_));
 sg13g2_a21oi_1 _13024_ (.A1(_05245_),
    .A2(_05248_),
    .Y(_01022_),
    .B1(_05250_));
 sg13g2_xnor2_1 _13025_ (.Y(_05251_),
    .A(\am_sdr0.cic0.integ1[9] ),
    .B(net1667));
 sg13g2_a21oi_1 _13026_ (.A1(_05247_),
    .A2(_05249_),
    .Y(_05252_),
    .B1(_05251_));
 sg13g2_and3_1 _13027_ (.X(_05253_),
    .A(_05247_),
    .B(_05249_),
    .C(_05251_));
 sg13g2_nor3_1 _13028_ (.A(net1881),
    .B(_05252_),
    .C(_05253_),
    .Y(_01023_));
 sg13g2_nand2_1 _13029_ (.Y(_05254_),
    .A(net3213),
    .B(net1666));
 sg13g2_xnor2_1 _13030_ (.Y(_05255_),
    .A(net3213),
    .B(net1666));
 sg13g2_o21ai_1 _13031_ (.B1(net1666),
    .Y(_05256_),
    .A1(\am_sdr0.cic0.integ1[8] ),
    .A2(\am_sdr0.cic0.integ1[9] ));
 sg13g2_o21ai_1 _13032_ (.B1(_05256_),
    .Y(_05257_),
    .A1(_05245_),
    .A2(_05248_));
 sg13g2_o21ai_1 _13033_ (.B1(_05257_),
    .Y(_05258_),
    .A1(\am_sdr0.cic0.integ1[9] ),
    .A2(net1666));
 sg13g2_or2_1 _13034_ (.X(_05259_),
    .B(_05258_),
    .A(_05255_));
 sg13g2_nand2_1 _13035_ (.Y(_05260_),
    .A(net1938),
    .B(_05259_));
 sg13g2_a21oi_1 _13036_ (.A1(_05255_),
    .A2(_05258_),
    .Y(_01024_),
    .B1(_05260_));
 sg13g2_xnor2_1 _13037_ (.Y(_05261_),
    .A(net3246),
    .B(net1666));
 sg13g2_nand3_1 _13038_ (.B(_05259_),
    .C(_05261_),
    .A(_05254_),
    .Y(_05262_));
 sg13g2_a21oi_1 _13039_ (.A1(_05254_),
    .A2(_05259_),
    .Y(_05263_),
    .B1(_05261_));
 sg13g2_nand2_1 _13040_ (.Y(_05264_),
    .A(net1938),
    .B(_05262_));
 sg13g2_nor2_1 _13041_ (.A(_05263_),
    .B(_05264_),
    .Y(_01025_));
 sg13g2_nand2_1 _13042_ (.Y(_05265_),
    .A(net3220),
    .B(net1668));
 sg13g2_xnor2_1 _13043_ (.Y(_05266_),
    .A(\am_sdr0.cic0.integ1[12] ),
    .B(net1668));
 sg13g2_o21ai_1 _13044_ (.B1(net1666),
    .Y(_05267_),
    .A1(\am_sdr0.cic0.integ1[10] ),
    .A2(\am_sdr0.cic0.integ1[11] ));
 sg13g2_nand2_1 _13045_ (.Y(_05268_),
    .A(_05256_),
    .B(_05267_));
 sg13g2_nor4_1 _13046_ (.A(_05248_),
    .B(_05251_),
    .C(_05255_),
    .D(_05261_),
    .Y(_05269_));
 sg13g2_a21oi_1 _13047_ (.A1(_05246_),
    .A2(_05269_),
    .Y(_05270_),
    .B1(_05268_));
 sg13g2_or2_1 _13048_ (.X(_05271_),
    .B(_05270_),
    .A(_05266_));
 sg13g2_a21oi_1 _13049_ (.A1(_05266_),
    .A2(_05270_),
    .Y(_05272_),
    .B1(net1881));
 sg13g2_and2_1 _13050_ (.A(_05271_),
    .B(_05272_),
    .X(_01026_));
 sg13g2_xor2_1 _13051_ (.B(net1668),
    .A(\am_sdr0.cic0.integ1[13] ),
    .X(_05273_));
 sg13g2_nand2_1 _13052_ (.Y(_05274_),
    .A(_05265_),
    .B(_05271_));
 sg13g2_o21ai_1 _13053_ (.B1(net1931),
    .Y(_05275_),
    .A1(_05273_),
    .A2(_05274_));
 sg13g2_a21oi_1 _13054_ (.A1(_05273_),
    .A2(_05274_),
    .Y(_01027_),
    .B1(_05275_));
 sg13g2_nand2_1 _13055_ (.Y(_05276_),
    .A(net3272),
    .B(net1669));
 sg13g2_xnor2_1 _13056_ (.Y(_05277_),
    .A(\am_sdr0.cic0.integ1[14] ),
    .B(net1669));
 sg13g2_o21ai_1 _13057_ (.B1(net1668),
    .Y(_05278_),
    .A1(\am_sdr0.cic0.integ1[12] ),
    .A2(\am_sdr0.cic0.integ1[13] ));
 sg13g2_o21ai_1 _13058_ (.B1(_05278_),
    .Y(_05279_),
    .A1(_05266_),
    .A2(_05270_));
 sg13g2_o21ai_1 _13059_ (.B1(_05279_),
    .Y(_05280_),
    .A1(net3222),
    .A2(net1668));
 sg13g2_or2_1 _13060_ (.X(_05281_),
    .B(_05280_),
    .A(_05277_));
 sg13g2_nand2_1 _13061_ (.Y(_05282_),
    .A(net1931),
    .B(_05281_));
 sg13g2_a21oi_1 _13062_ (.A1(_05277_),
    .A2(_05280_),
    .Y(_01028_),
    .B1(_05282_));
 sg13g2_xnor2_1 _13063_ (.Y(_05283_),
    .A(net3239),
    .B(net1669));
 sg13g2_and3_1 _13064_ (.X(_05284_),
    .A(_05276_),
    .B(_05281_),
    .C(_05283_));
 sg13g2_a21oi_1 _13065_ (.A1(_05276_),
    .A2(_05281_),
    .Y(_05285_),
    .B1(_05283_));
 sg13g2_nor3_1 _13066_ (.A(net1880),
    .B(_05284_),
    .C(_05285_),
    .Y(_01029_));
 sg13g2_nor2b_1 _13067_ (.A(_05266_),
    .B_N(_05273_),
    .Y(_05286_));
 sg13g2_nor2_1 _13068_ (.A(_05277_),
    .B(_05283_),
    .Y(_05287_));
 sg13g2_and3_1 _13069_ (.X(_05288_),
    .A(_05269_),
    .B(_05286_),
    .C(_05287_));
 sg13g2_o21ai_1 _13070_ (.B1(net1668),
    .Y(_05289_),
    .A1(\am_sdr0.cic0.integ1[14] ),
    .A2(\am_sdr0.cic0.integ1[15] ));
 sg13g2_nand4_1 _13071_ (.B(_05267_),
    .C(_05278_),
    .A(_05256_),
    .Y(_05290_),
    .D(_05289_));
 sg13g2_a21oi_2 _13072_ (.B1(_05290_),
    .Y(_05291_),
    .A2(_05288_),
    .A1(_05246_));
 sg13g2_nand2_1 _13073_ (.Y(_05292_),
    .A(\am_sdr0.cic0.integ1[16] ),
    .B(net1664));
 sg13g2_xnor2_1 _13074_ (.Y(_05293_),
    .A(\am_sdr0.cic0.integ1[16] ),
    .B(net1669));
 sg13g2_inv_1 _13075_ (.Y(_05294_),
    .A(_05293_));
 sg13g2_o21ai_1 _13076_ (.B1(net1932),
    .Y(_05295_),
    .A1(_05291_),
    .A2(_05293_));
 sg13g2_a21oi_1 _13077_ (.A1(_05291_),
    .A2(_05293_),
    .Y(_01030_),
    .B1(_05295_));
 sg13g2_or2_1 _13078_ (.X(_05296_),
    .B(net1665),
    .A(\am_sdr0.cic0.integ1[17] ));
 sg13g2_xor2_1 _13079_ (.B(net1665),
    .A(net3278),
    .X(_05297_));
 sg13g2_o21ai_1 _13080_ (.B1(_05292_),
    .Y(_05298_),
    .A1(_05291_),
    .A2(_05293_));
 sg13g2_o21ai_1 _13081_ (.B1(net1930),
    .Y(_05299_),
    .A1(_05297_),
    .A2(_05298_));
 sg13g2_a21oi_1 _13082_ (.A1(_05297_),
    .A2(_05298_),
    .Y(_01031_),
    .B1(_05299_));
 sg13g2_nand2_1 _13083_ (.Y(_05300_),
    .A(net3276),
    .B(net1665));
 sg13g2_xor2_1 _13084_ (.B(net1665),
    .A(net3276),
    .X(_05301_));
 sg13g2_o21ai_1 _13085_ (.B1(net1664),
    .Y(_05302_),
    .A1(\am_sdr0.cic0.integ1[16] ),
    .A2(\am_sdr0.cic0.integ1[17] ));
 sg13g2_o21ai_1 _13086_ (.B1(_05302_),
    .Y(_05303_),
    .A1(_05291_),
    .A2(_05293_));
 sg13g2_a21oi_1 _13087_ (.A1(_05296_),
    .A2(_05303_),
    .Y(_05304_),
    .B1(_05301_));
 sg13g2_nand3_1 _13088_ (.B(_05301_),
    .C(_05303_),
    .A(_05296_),
    .Y(_05305_));
 sg13g2_nand2_1 _13089_ (.Y(_05306_),
    .A(net1930),
    .B(_05305_));
 sg13g2_nor2_1 _13090_ (.A(net3277),
    .B(_05306_),
    .Y(_01032_));
 sg13g2_xor2_1 _13091_ (.B(net1664),
    .A(net3199),
    .X(_05307_));
 sg13g2_nand2_1 _13092_ (.Y(_05308_),
    .A(_05300_),
    .B(_05305_));
 sg13g2_o21ai_1 _13093_ (.B1(net1930),
    .Y(_05309_),
    .A1(_05307_),
    .A2(_05308_));
 sg13g2_a21oi_1 _13094_ (.A1(_05307_),
    .A2(_05308_),
    .Y(_01033_),
    .B1(_05309_));
 sg13g2_nand4_1 _13095_ (.B(_05297_),
    .C(_05301_),
    .A(_05294_),
    .Y(_05310_),
    .D(_05307_));
 sg13g2_nand2_1 _13096_ (.Y(_05311_),
    .A(_05300_),
    .B(_05302_));
 sg13g2_a21oi_1 _13097_ (.A1(\am_sdr0.cic0.integ1[19] ),
    .A2(net1664),
    .Y(_05312_),
    .B1(_05311_));
 sg13g2_o21ai_1 _13098_ (.B1(_05312_),
    .Y(_05313_),
    .A1(_05291_),
    .A2(_05310_));
 sg13g2_nand2_1 _13099_ (.Y(_05314_),
    .A(net3266),
    .B(net1664));
 sg13g2_xnor2_1 _13100_ (.Y(_05315_),
    .A(\am_sdr0.cic0.integ1[20] ),
    .B(net1663));
 sg13g2_nand2b_1 _13101_ (.Y(_05316_),
    .B(_05315_),
    .A_N(_05313_));
 sg13g2_nand2b_1 _13102_ (.Y(_05317_),
    .B(_05313_),
    .A_N(_05315_));
 sg13g2_and3_1 _13103_ (.X(_01034_),
    .A(net1930),
    .B(_05316_),
    .C(_05317_));
 sg13g2_xnor2_1 _13104_ (.Y(_05318_),
    .A(\am_sdr0.cic0.integ1[21] ),
    .B(net1663));
 sg13g2_nand3_1 _13105_ (.B(_05317_),
    .C(_05318_),
    .A(_05314_),
    .Y(_05319_));
 sg13g2_a21oi_1 _13106_ (.A1(_05314_),
    .A2(_05317_),
    .Y(_05320_),
    .B1(_05318_));
 sg13g2_nand2_1 _13107_ (.Y(_05321_),
    .A(net1930),
    .B(_05319_));
 sg13g2_nor2_1 _13108_ (.A(_05320_),
    .B(_05321_),
    .Y(_01035_));
 sg13g2_nand2_1 _13109_ (.Y(_05322_),
    .A(net3217),
    .B(net1663));
 sg13g2_xnor2_1 _13110_ (.Y(_05323_),
    .A(net3217),
    .B(net1664));
 sg13g2_o21ai_1 _13111_ (.B1(net1664),
    .Y(_05324_),
    .A1(\am_sdr0.cic0.integ1[20] ),
    .A2(\am_sdr0.cic0.integ1[21] ));
 sg13g2_inv_1 _13112_ (.Y(_05325_),
    .A(_05324_));
 sg13g2_nor2_1 _13113_ (.A(_05315_),
    .B(_05318_),
    .Y(_05326_));
 sg13g2_a21oi_1 _13114_ (.A1(_05313_),
    .A2(_05326_),
    .Y(_05327_),
    .B1(_05325_));
 sg13g2_or2_1 _13115_ (.X(_05328_),
    .B(_05327_),
    .A(_05323_));
 sg13g2_nand2_1 _13116_ (.Y(_05329_),
    .A(net1930),
    .B(_05328_));
 sg13g2_a21oi_1 _13117_ (.A1(_05323_),
    .A2(_05327_),
    .Y(_01036_),
    .B1(_05329_));
 sg13g2_xnor2_1 _13118_ (.Y(_05330_),
    .A(net3224),
    .B(net1663));
 sg13g2_and3_1 _13119_ (.X(_05331_),
    .A(_05322_),
    .B(_05328_),
    .C(_05330_));
 sg13g2_a21oi_1 _13120_ (.A1(_05322_),
    .A2(_05328_),
    .Y(_05332_),
    .B1(_05330_));
 sg13g2_nor3_1 _13121_ (.A(net1876),
    .B(_05331_),
    .C(_05332_),
    .Y(_01037_));
 sg13g2_or4_1 _13122_ (.A(_05315_),
    .B(_05318_),
    .C(_05323_),
    .D(_05330_),
    .X(_05333_));
 sg13g2_nor3_1 _13123_ (.A(_05291_),
    .B(_05310_),
    .C(_05333_),
    .Y(_05334_));
 sg13g2_o21ai_1 _13124_ (.B1(net1663),
    .Y(_05335_),
    .A1(\am_sdr0.cic0.integ1[22] ),
    .A2(\am_sdr0.cic0.integ1[23] ));
 sg13g2_nand3_1 _13125_ (.B(_05324_),
    .C(_05335_),
    .A(_05312_),
    .Y(_05336_));
 sg13g2_nand2_1 _13126_ (.Y(_05337_),
    .A(net3148),
    .B(net1663));
 sg13g2_xor2_1 _13127_ (.B(net1663),
    .A(net3293),
    .X(_05338_));
 sg13g2_nor3_1 _13128_ (.A(_05334_),
    .B(_05336_),
    .C(_05338_),
    .Y(_05339_));
 sg13g2_o21ai_1 _13129_ (.B1(_05338_),
    .Y(_05340_),
    .A1(_05334_),
    .A2(_05336_));
 sg13g2_nand2_1 _13130_ (.Y(_05341_),
    .A(net1904),
    .B(_05340_));
 sg13g2_nor2_1 _13131_ (.A(net3294),
    .B(_05341_),
    .Y(_01038_));
 sg13g2_xnor2_1 _13132_ (.Y(_05342_),
    .A(net3072),
    .B(net1663));
 sg13g2_and3_1 _13133_ (.X(_05343_),
    .A(_05337_),
    .B(_05340_),
    .C(_05342_));
 sg13g2_a21oi_1 _13134_ (.A1(_05337_),
    .A2(_05340_),
    .Y(_05344_),
    .B1(_05342_));
 sg13g2_nor3_1 _13135_ (.A(net1876),
    .B(_05343_),
    .C(_05344_),
    .Y(_01039_));
 sg13g2_nand2_1 _13136_ (.Y(_05345_),
    .A(net2611),
    .B(net2845));
 sg13g2_o21ai_1 _13137_ (.B1(net1932),
    .Y(_05346_),
    .A1(net2611),
    .A2(\am_sdr0.cic0.integ1[3] ));
 sg13g2_nor2b_1 _13138_ (.A(net2612),
    .B_N(_05345_),
    .Y(_01040_));
 sg13g2_nand2_1 _13139_ (.Y(_05347_),
    .A(net3241),
    .B(\am_sdr0.cic0.integ1[4] ));
 sg13g2_xnor2_1 _13140_ (.Y(_05348_),
    .A(\am_sdr0.cic0.integ2[1] ),
    .B(\am_sdr0.cic0.integ1[4] ));
 sg13g2_o21ai_1 _13141_ (.B1(net1932),
    .Y(_05349_),
    .A1(_05345_),
    .A2(_05348_));
 sg13g2_a21oi_1 _13142_ (.A1(_05345_),
    .A2(_05348_),
    .Y(_01041_),
    .B1(_05349_));
 sg13g2_and2_1 _13143_ (.A(net3202),
    .B(\am_sdr0.cic0.integ1[5] ),
    .X(_05350_));
 sg13g2_xor2_1 _13144_ (.B(\am_sdr0.cic0.integ1[5] ),
    .A(net3202),
    .X(_05351_));
 sg13g2_o21ai_1 _13145_ (.B1(_05347_),
    .Y(_05352_),
    .A1(_05345_),
    .A2(_05348_));
 sg13g2_nor2_1 _13146_ (.A(_05351_),
    .B(_05352_),
    .Y(_05353_));
 sg13g2_a21oi_1 _13147_ (.A1(_05351_),
    .A2(_05352_),
    .Y(_05354_),
    .B1(net1879));
 sg13g2_nor2b_1 _13148_ (.A(net3242),
    .B_N(_05354_),
    .Y(_01042_));
 sg13g2_nand2_1 _13149_ (.Y(_05355_),
    .A(\am_sdr0.cic0.integ2[3] ),
    .B(\am_sdr0.cic0.integ1[6] ));
 sg13g2_xnor2_1 _13150_ (.Y(_05356_),
    .A(net2756),
    .B(\am_sdr0.cic0.integ1[6] ));
 sg13g2_a21oi_2 _13151_ (.B1(net3203),
    .Y(_05357_),
    .A2(_05352_),
    .A1(_05351_));
 sg13g2_o21ai_1 _13152_ (.B1(net1936),
    .Y(_05358_),
    .A1(_05356_),
    .A2(_05357_));
 sg13g2_a21oi_1 _13153_ (.A1(_05356_),
    .A2(_05357_),
    .Y(_01043_),
    .B1(_05358_));
 sg13g2_and2_1 _13154_ (.A(net2990),
    .B(\am_sdr0.cic0.integ1[7] ),
    .X(_05359_));
 sg13g2_xor2_1 _13155_ (.B(\am_sdr0.cic0.integ1[7] ),
    .A(\am_sdr0.cic0.integ2[4] ),
    .X(_05360_));
 sg13g2_o21ai_1 _13156_ (.B1(_05355_),
    .Y(_05361_),
    .A1(_05356_),
    .A2(_05357_));
 sg13g2_or2_1 _13157_ (.X(_05362_),
    .B(_05361_),
    .A(_05360_));
 sg13g2_a21oi_1 _13158_ (.A1(_05360_),
    .A2(_05361_),
    .Y(_05363_),
    .B1(net1881));
 sg13g2_and2_1 _13159_ (.A(_05362_),
    .B(_05363_),
    .X(_01044_));
 sg13g2_a21oi_1 _13160_ (.A1(_05360_),
    .A2(_05361_),
    .Y(_05364_),
    .B1(_05359_));
 sg13g2_nor2_1 _13161_ (.A(\am_sdr0.cic0.integ2[5] ),
    .B(\am_sdr0.cic0.integ1[8] ),
    .Y(_05365_));
 sg13g2_xnor2_1 _13162_ (.Y(_05366_),
    .A(net3181),
    .B(\am_sdr0.cic0.integ1[8] ));
 sg13g2_o21ai_1 _13163_ (.B1(net1936),
    .Y(_05367_),
    .A1(_05364_),
    .A2(_05366_));
 sg13g2_a21oi_1 _13164_ (.A1(_05364_),
    .A2(net3182),
    .Y(_01045_),
    .B1(_05367_));
 sg13g2_and2_1 _13165_ (.A(net3142),
    .B(\am_sdr0.cic0.integ1[9] ),
    .X(_05368_));
 sg13g2_xnor2_1 _13166_ (.Y(_05369_),
    .A(net3307),
    .B(\am_sdr0.cic0.integ1[9] ));
 sg13g2_a221oi_1 _13167_ (.B2(_05361_),
    .C1(_05359_),
    .B1(_05360_),
    .A1(\am_sdr0.cic0.integ2[5] ),
    .Y(_05370_),
    .A2(\am_sdr0.cic0.integ1[8] ));
 sg13g2_o21ai_1 _13168_ (.B1(_05369_),
    .Y(_05371_),
    .A1(_05365_),
    .A2(_05370_));
 sg13g2_nor3_2 _13169_ (.A(_05365_),
    .B(_05369_),
    .C(_05370_),
    .Y(_05372_));
 sg13g2_nand2_1 _13170_ (.Y(_05373_),
    .A(net1938),
    .B(_05371_));
 sg13g2_nor2_1 _13171_ (.A(_05372_),
    .B(_05373_),
    .Y(_01046_));
 sg13g2_nand2_1 _13172_ (.Y(_05374_),
    .A(\am_sdr0.cic0.integ2[7] ),
    .B(\am_sdr0.cic0.integ1[10] ));
 sg13g2_xor2_1 _13173_ (.B(net3288),
    .A(\am_sdr0.cic0.integ2[7] ),
    .X(_05375_));
 sg13g2_nor3_1 _13174_ (.A(_05368_),
    .B(_05372_),
    .C(net3289),
    .Y(_05376_));
 sg13g2_o21ai_1 _13175_ (.B1(_05375_),
    .Y(_05377_),
    .A1(_05368_),
    .A2(_05372_));
 sg13g2_nand2_1 _13176_ (.Y(_05378_),
    .A(net1936),
    .B(_05377_));
 sg13g2_nor2_1 _13177_ (.A(_05376_),
    .B(_05378_),
    .Y(_01047_));
 sg13g2_nand2_1 _13178_ (.Y(_05379_),
    .A(_05374_),
    .B(_05377_));
 sg13g2_nand2_1 _13179_ (.Y(_05380_),
    .A(net3099),
    .B(\am_sdr0.cic0.integ1[11] ));
 sg13g2_xor2_1 _13180_ (.B(net3304),
    .A(\am_sdr0.cic0.integ2[8] ),
    .X(_05381_));
 sg13g2_inv_1 _13181_ (.Y(_05382_),
    .A(_05381_));
 sg13g2_nand2_1 _13182_ (.Y(_05383_),
    .A(_05379_),
    .B(_05381_));
 sg13g2_o21ai_1 _13183_ (.B1(net1936),
    .Y(_05384_),
    .A1(_05379_),
    .A2(net3305));
 sg13g2_nor2b_1 _13184_ (.A(_05384_),
    .B_N(_05383_),
    .Y(_01048_));
 sg13g2_nor2_1 _13185_ (.A(net3231),
    .B(\am_sdr0.cic0.integ1[12] ),
    .Y(_05385_));
 sg13g2_nand2_1 _13186_ (.Y(_05386_),
    .A(net3231),
    .B(net3220));
 sg13g2_nand2b_1 _13187_ (.Y(_05387_),
    .B(_05386_),
    .A_N(_05385_));
 sg13g2_and2_1 _13188_ (.A(_05380_),
    .B(_05383_),
    .X(_05388_));
 sg13g2_o21ai_1 _13189_ (.B1(net1936),
    .Y(_05389_),
    .A1(_05387_),
    .A2(_05388_));
 sg13g2_a21oi_1 _13190_ (.A1(net3232),
    .A2(_05388_),
    .Y(_01049_),
    .B1(_05389_));
 sg13g2_nand2_1 _13191_ (.Y(_05390_),
    .A(net3255),
    .B(net3222));
 sg13g2_xnor2_1 _13192_ (.Y(_05391_),
    .A(\am_sdr0.cic0.integ2[10] ),
    .B(\am_sdr0.cic0.integ1[13] ));
 sg13g2_nor2_1 _13193_ (.A(_05382_),
    .B(_05387_),
    .Y(_05392_));
 sg13g2_o21ai_1 _13194_ (.B1(_05386_),
    .Y(_05393_),
    .A1(_05380_),
    .A2(_05385_));
 sg13g2_a21oi_1 _13195_ (.A1(_05379_),
    .A2(_05392_),
    .Y(_05394_),
    .B1(_05393_));
 sg13g2_or2_1 _13196_ (.X(_05395_),
    .B(_05394_),
    .A(_05391_));
 sg13g2_a21oi_1 _13197_ (.A1(_05391_),
    .A2(_05394_),
    .Y(_05396_),
    .B1(net1879));
 sg13g2_and2_1 _13198_ (.A(_05395_),
    .B(_05396_),
    .X(_01050_));
 sg13g2_nor2_1 _13199_ (.A(\am_sdr0.cic0.integ2[11] ),
    .B(\am_sdr0.cic0.integ1[14] ),
    .Y(_05397_));
 sg13g2_xnor2_1 _13200_ (.Y(_05398_),
    .A(net3262),
    .B(net3272));
 sg13g2_and3_1 _13201_ (.X(_05399_),
    .A(_05390_),
    .B(_05395_),
    .C(_05398_));
 sg13g2_a21oi_1 _13202_ (.A1(_05390_),
    .A2(_05395_),
    .Y(_05400_),
    .B1(_05398_));
 sg13g2_nor3_1 _13203_ (.A(net1879),
    .B(_05399_),
    .C(_05400_),
    .Y(_01051_));
 sg13g2_nand2_1 _13204_ (.Y(_05401_),
    .A(net3207),
    .B(net3239));
 sg13g2_xor2_1 _13205_ (.B(\am_sdr0.cic0.integ1[15] ),
    .A(\am_sdr0.cic0.integ2[12] ),
    .X(_05402_));
 sg13g2_inv_1 _13206_ (.Y(_05403_),
    .A(_05402_));
 sg13g2_nor2_1 _13207_ (.A(_05391_),
    .B(_05398_),
    .Y(_05404_));
 sg13g2_nor2_1 _13208_ (.A(_05390_),
    .B(_05397_),
    .Y(_05405_));
 sg13g2_a221oi_1 _13209_ (.B2(_05404_),
    .C1(_05405_),
    .B1(_05393_),
    .A1(\am_sdr0.cic0.integ2[11] ),
    .Y(_05406_),
    .A2(\am_sdr0.cic0.integ1[14] ));
 sg13g2_inv_1 _13210_ (.Y(_05407_),
    .A(_05406_));
 sg13g2_nand2_1 _13211_ (.Y(_05408_),
    .A(_05392_),
    .B(_05404_));
 sg13g2_a21oi_2 _13212_ (.B1(_05408_),
    .Y(_05409_),
    .A2(_05377_),
    .A1(_05374_));
 sg13g2_nor3_1 _13213_ (.A(_05402_),
    .B(_05407_),
    .C(_05409_),
    .Y(_05410_));
 sg13g2_o21ai_1 _13214_ (.B1(_05402_),
    .Y(_05411_),
    .A1(_05407_),
    .A2(_05409_));
 sg13g2_nand2_1 _13215_ (.Y(_05412_),
    .A(net1931),
    .B(_05411_));
 sg13g2_nor2_1 _13216_ (.A(_05410_),
    .B(_05412_),
    .Y(_01052_));
 sg13g2_nor2_1 _13217_ (.A(net3274),
    .B(\am_sdr0.cic0.integ1[16] ),
    .Y(_05413_));
 sg13g2_xnor2_1 _13218_ (.Y(_05414_),
    .A(\am_sdr0.cic0.integ2[13] ),
    .B(\am_sdr0.cic0.integ1[16] ));
 sg13g2_and3_1 _13219_ (.X(_05415_),
    .A(_05401_),
    .B(_05411_),
    .C(_05414_));
 sg13g2_a21oi_1 _13220_ (.A1(_05401_),
    .A2(_05411_),
    .Y(_05416_),
    .B1(_05414_));
 sg13g2_nor3_1 _13221_ (.A(net1880),
    .B(_05415_),
    .C(net3240),
    .Y(_01053_));
 sg13g2_nand2_1 _13222_ (.Y(_05417_),
    .A(net3215),
    .B(net3278));
 sg13g2_xnor2_1 _13223_ (.Y(_05418_),
    .A(net3215),
    .B(\am_sdr0.cic0.integ1[17] ));
 sg13g2_a22oi_1 _13224_ (.Y(_05419_),
    .B1(\am_sdr0.cic0.integ2[13] ),
    .B2(\am_sdr0.cic0.integ1[16] ),
    .A2(\am_sdr0.cic0.integ1[15] ),
    .A1(\am_sdr0.cic0.integ2[12] ));
 sg13g2_a21o_1 _13225_ (.A2(_05419_),
    .A1(_05411_),
    .B1(_05413_),
    .X(_05420_));
 sg13g2_or2_1 _13226_ (.X(_05421_),
    .B(_05420_),
    .A(_05418_));
 sg13g2_nand2_1 _13227_ (.Y(_05422_),
    .A(net1931),
    .B(_05421_));
 sg13g2_a21oi_1 _13228_ (.A1(_05418_),
    .A2(_05420_),
    .Y(_01054_),
    .B1(_05422_));
 sg13g2_nor2_1 _13229_ (.A(\am_sdr0.cic0.integ2[15] ),
    .B(\am_sdr0.cic0.integ1[18] ),
    .Y(_05423_));
 sg13g2_xnor2_1 _13230_ (.Y(_05424_),
    .A(\am_sdr0.cic0.integ2[15] ),
    .B(net3287));
 sg13g2_and3_1 _13231_ (.X(_05425_),
    .A(_05417_),
    .B(_05421_),
    .C(_05424_));
 sg13g2_a21oi_1 _13232_ (.A1(_05417_),
    .A2(_05421_),
    .Y(_05426_),
    .B1(_05424_));
 sg13g2_nor3_1 _13233_ (.A(net1880),
    .B(_05425_),
    .C(_05426_),
    .Y(_01055_));
 sg13g2_xnor2_1 _13234_ (.Y(_05427_),
    .A(\am_sdr0.cic0.integ2[16] ),
    .B(net3312));
 sg13g2_nor4_2 _13235_ (.A(_05403_),
    .B(_05414_),
    .C(_05418_),
    .Y(_05428_),
    .D(_05424_));
 sg13g2_nor2_1 _13236_ (.A(_05417_),
    .B(_05423_),
    .Y(_05429_));
 sg13g2_a21oi_1 _13237_ (.A1(\am_sdr0.cic0.integ2[15] ),
    .A2(\am_sdr0.cic0.integ1[18] ),
    .Y(_05430_),
    .B1(_05429_));
 sg13g2_nor4_1 _13238_ (.A(_05413_),
    .B(_05418_),
    .C(_05419_),
    .D(_05424_),
    .Y(_05431_));
 sg13g2_a21oi_1 _13239_ (.A1(_05407_),
    .A2(_05428_),
    .Y(_05432_),
    .B1(_05431_));
 sg13g2_nand2_1 _13240_ (.Y(_05433_),
    .A(_05430_),
    .B(_05432_));
 sg13g2_a21oi_2 _13241_ (.B1(_05433_),
    .Y(_05434_),
    .A2(_05428_),
    .A1(_05409_));
 sg13g2_nor2_1 _13242_ (.A(_05427_),
    .B(_05434_),
    .Y(_05435_));
 sg13g2_a21oi_1 _13243_ (.A1(_05427_),
    .A2(_05434_),
    .Y(_05436_),
    .B1(net1879));
 sg13g2_nor2b_1 _13244_ (.A(_05435_),
    .B_N(_05436_),
    .Y(_01056_));
 sg13g2_nor2_1 _13245_ (.A(\am_sdr0.cic0.integ2[17] ),
    .B(\am_sdr0.cic0.integ1[20] ),
    .Y(_05437_));
 sg13g2_xnor2_1 _13246_ (.Y(_05438_),
    .A(\am_sdr0.cic0.integ2[17] ),
    .B(\am_sdr0.cic0.integ1[20] ));
 sg13g2_a21oi_1 _13247_ (.A1(\am_sdr0.cic0.integ2[16] ),
    .A2(net3199),
    .Y(_05439_),
    .B1(_05435_));
 sg13g2_o21ai_1 _13248_ (.B1(net1931),
    .Y(_05440_),
    .A1(_05438_),
    .A2(_05439_));
 sg13g2_a21oi_1 _13249_ (.A1(_05438_),
    .A2(net3200),
    .Y(_01057_),
    .B1(_05440_));
 sg13g2_and2_1 _13250_ (.A(\am_sdr0.cic0.integ2[18] ),
    .B(\am_sdr0.cic0.integ1[21] ),
    .X(_05441_));
 sg13g2_or2_1 _13251_ (.X(_05442_),
    .B(net3291),
    .A(\am_sdr0.cic0.integ2[18] ));
 sg13g2_nand2b_1 _13252_ (.Y(_05443_),
    .B(_05442_),
    .A_N(_05441_));
 sg13g2_nor2_1 _13253_ (.A(_05427_),
    .B(_05438_),
    .Y(_05444_));
 sg13g2_inv_1 _13254_ (.Y(_05445_),
    .A(_05444_));
 sg13g2_a22oi_1 _13255_ (.Y(_05446_),
    .B1(\am_sdr0.cic0.integ2[17] ),
    .B2(\am_sdr0.cic0.integ1[20] ),
    .A2(\am_sdr0.cic0.integ1[19] ),
    .A1(\am_sdr0.cic0.integ2[16] ));
 sg13g2_nor2_1 _13256_ (.A(_05437_),
    .B(_05446_),
    .Y(_05447_));
 sg13g2_inv_1 _13257_ (.Y(_05448_),
    .A(_05447_));
 sg13g2_o21ai_1 _13258_ (.B1(_05448_),
    .Y(_05449_),
    .A1(_05434_),
    .A2(_05445_));
 sg13g2_inv_1 _13259_ (.Y(_05450_),
    .A(_05449_));
 sg13g2_o21ai_1 _13260_ (.B1(net1931),
    .Y(_05451_),
    .A1(_05443_),
    .A2(_05450_));
 sg13g2_a21oi_1 _13261_ (.A1(_05443_),
    .A2(_05450_),
    .Y(_01058_),
    .B1(_05451_));
 sg13g2_and2_1 _13262_ (.A(\am_sdr0.cic0.integ2[19] ),
    .B(net3259),
    .X(_05452_));
 sg13g2_or2_1 _13263_ (.X(_05453_),
    .B(net3259),
    .A(\am_sdr0.cic0.integ2[19] ));
 sg13g2_nand2b_1 _13264_ (.Y(_05454_),
    .B(net3260),
    .A_N(_05452_));
 sg13g2_a21oi_1 _13265_ (.A1(_05442_),
    .A2(_05449_),
    .Y(_05455_),
    .B1(_05441_));
 sg13g2_o21ai_1 _13266_ (.B1(net1931),
    .Y(_05456_),
    .A1(_05454_),
    .A2(_05455_));
 sg13g2_a21oi_1 _13267_ (.A1(_05454_),
    .A2(_05455_),
    .Y(_01059_),
    .B1(_05456_));
 sg13g2_nor2_1 _13268_ (.A(_05443_),
    .B(_05454_),
    .Y(_05457_));
 sg13g2_nand2_1 _13269_ (.Y(_05458_),
    .A(_05444_),
    .B(_05457_));
 sg13g2_a221oi_1 _13270_ (.B2(_05447_),
    .C1(_05452_),
    .B1(_05457_),
    .A1(_05441_),
    .Y(_05459_),
    .A2(_05453_));
 sg13g2_o21ai_1 _13271_ (.B1(_05459_),
    .Y(_05460_),
    .A1(_05434_),
    .A2(_05458_));
 sg13g2_and2_1 _13272_ (.A(net3144),
    .B(\am_sdr0.cic0.integ1[23] ),
    .X(_05461_));
 sg13g2_xnor2_1 _13273_ (.Y(_05462_),
    .A(\am_sdr0.cic0.integ2[20] ),
    .B(net3224));
 sg13g2_inv_1 _13274_ (.Y(_05463_),
    .A(_05462_));
 sg13g2_o21ai_1 _13275_ (.B1(net1904),
    .Y(_05464_),
    .A1(_05460_),
    .A2(_05463_));
 sg13g2_a21oi_1 _13276_ (.A1(_05460_),
    .A2(_05463_),
    .Y(_01060_),
    .B1(_05464_));
 sg13g2_or2_1 _13277_ (.X(_05465_),
    .B(\am_sdr0.cic0.integ1[24] ),
    .A(\am_sdr0.cic0.integ2[21] ));
 sg13g2_and2_1 _13278_ (.A(\am_sdr0.cic0.integ2[21] ),
    .B(net3327),
    .X(_05466_));
 sg13g2_xnor2_1 _13279_ (.Y(_05467_),
    .A(net3205),
    .B(net3148));
 sg13g2_a21oi_1 _13280_ (.A1(_05460_),
    .A2(_05463_),
    .Y(_05468_),
    .B1(_05461_));
 sg13g2_o21ai_1 _13281_ (.B1(net1904),
    .Y(_05469_),
    .A1(_05467_),
    .A2(_05468_));
 sg13g2_a21oi_1 _13282_ (.A1(_05467_),
    .A2(_05468_),
    .Y(_01061_),
    .B1(_05469_));
 sg13g2_nor2_1 _13283_ (.A(_05462_),
    .B(_05467_),
    .Y(_05470_));
 sg13g2_a221oi_1 _13284_ (.B2(_05460_),
    .C1(_05466_),
    .B1(_05470_),
    .A1(_05461_),
    .Y(_05471_),
    .A2(_05465_));
 sg13g2_xnor2_1 _13285_ (.Y(_05472_),
    .A(net3019),
    .B(net3072));
 sg13g2_o21ai_1 _13286_ (.B1(net1904),
    .Y(_05473_),
    .A1(_05471_),
    .A2(_05472_));
 sg13g2_a21oi_1 _13287_ (.A1(_05471_),
    .A2(_05472_),
    .Y(_01062_),
    .B1(_05473_));
 sg13g2_nor2_1 _13288_ (.A(net2116),
    .B(net1530),
    .Y(_05474_));
 sg13g2_a21oi_1 _13289_ (.A1(_01561_),
    .A2(net1530),
    .Y(_01063_),
    .B1(_05474_));
 sg13g2_nor2_1 _13290_ (.A(\am_sdr0.cic3.integ3[1] ),
    .B(net1532),
    .Y(_05475_));
 sg13g2_a21oi_1 _13291_ (.A1(_01559_),
    .A2(net1530),
    .Y(_01064_),
    .B1(_05475_));
 sg13g2_nor2_1 _13292_ (.A(\am_sdr0.cic3.integ3[2] ),
    .B(net1532),
    .Y(_05476_));
 sg13g2_a21oi_1 _13293_ (.A1(_01558_),
    .A2(net1530),
    .Y(_01065_),
    .B1(_05476_));
 sg13g2_nor2_1 _13294_ (.A(\am_sdr0.cic3.integ3[3] ),
    .B(net1530),
    .Y(_05477_));
 sg13g2_a21oi_1 _13295_ (.A1(_01557_),
    .A2(net1530),
    .Y(_01066_),
    .B1(_05477_));
 sg13g2_nor2_1 _13296_ (.A(\am_sdr0.cic3.integ3[4] ),
    .B(net1531),
    .Y(_05478_));
 sg13g2_a21oi_1 _13297_ (.A1(_01556_),
    .A2(net1531),
    .Y(_01067_),
    .B1(_05478_));
 sg13g2_nor2_1 _13298_ (.A(net2765),
    .B(net1531),
    .Y(_05479_));
 sg13g2_a21oi_1 _13299_ (.A1(_01555_),
    .A2(net1530),
    .Y(_01068_),
    .B1(_05479_));
 sg13g2_nor2_1 _13300_ (.A(net2478),
    .B(net1531),
    .Y(_05480_));
 sg13g2_a21oi_1 _13301_ (.A1(_01553_),
    .A2(net1530),
    .Y(_01069_),
    .B1(_05480_));
 sg13g2_nor2_1 _13302_ (.A(\am_sdr0.cic3.integ3[7] ),
    .B(net1533),
    .Y(_05481_));
 sg13g2_a21oi_1 _13303_ (.A1(_01552_),
    .A2(net1533),
    .Y(_01070_),
    .B1(_05481_));
 sg13g2_nor2_1 _13304_ (.A(\am_sdr0.cic3.integ3[8] ),
    .B(net1533),
    .Y(_05482_));
 sg13g2_a21oi_1 _13305_ (.A1(_01551_),
    .A2(net1533),
    .Y(_01071_),
    .B1(_05482_));
 sg13g2_nor2_1 _13306_ (.A(net2405),
    .B(net1536),
    .Y(_05483_));
 sg13g2_a21oi_1 _13307_ (.A1(_01550_),
    .A2(net1533),
    .Y(_01072_),
    .B1(_05483_));
 sg13g2_nor2_1 _13308_ (.A(\am_sdr0.cic3.integ3[10] ),
    .B(net1533),
    .Y(_05484_));
 sg13g2_a21oi_1 _13309_ (.A1(_01548_),
    .A2(net1533),
    .Y(_01073_),
    .B1(_05484_));
 sg13g2_nor2_1 _13310_ (.A(\am_sdr0.cic3.integ3[11] ),
    .B(net1533),
    .Y(_05485_));
 sg13g2_a21oi_1 _13311_ (.A1(_01547_),
    .A2(net1535),
    .Y(_01074_),
    .B1(_05485_));
 sg13g2_nor2_1 _13312_ (.A(\am_sdr0.cic3.integ3[12] ),
    .B(net1535),
    .Y(_05486_));
 sg13g2_a21oi_1 _13313_ (.A1(_01546_),
    .A2(net1535),
    .Y(_01075_),
    .B1(_05486_));
 sg13g2_nor2_1 _13314_ (.A(net2787),
    .B(net1535),
    .Y(_05487_));
 sg13g2_a21oi_1 _13315_ (.A1(_01545_),
    .A2(net1535),
    .Y(_01076_),
    .B1(_05487_));
 sg13g2_nor2_1 _13316_ (.A(net2279),
    .B(net1535),
    .Y(_05488_));
 sg13g2_a21oi_1 _13317_ (.A1(_01544_),
    .A2(net1536),
    .Y(_01077_),
    .B1(_05488_));
 sg13g2_nor2_1 _13318_ (.A(net2733),
    .B(net1535),
    .Y(_05489_));
 sg13g2_a21oi_1 _13319_ (.A1(_01543_),
    .A2(net1535),
    .Y(_01078_),
    .B1(_05489_));
 sg13g2_nor2_1 _13320_ (.A(net2517),
    .B(net1534),
    .Y(_05490_));
 sg13g2_a21oi_1 _13321_ (.A1(_01541_),
    .A2(net1534),
    .Y(_01079_),
    .B1(_05490_));
 sg13g2_nor2_1 _13322_ (.A(net2791),
    .B(net1534),
    .Y(_05491_));
 sg13g2_a21oi_1 _13323_ (.A1(_01540_),
    .A2(net1534),
    .Y(_01080_),
    .B1(_05491_));
 sg13g2_nor2_1 _13324_ (.A(net2230),
    .B(net1534),
    .Y(_05492_));
 sg13g2_a21oi_1 _13325_ (.A1(_01539_),
    .A2(net1534),
    .Y(_01081_),
    .B1(_05492_));
 sg13g2_nor2_1 _13326_ (.A(\am_sdr0.cic3.integ3[19] ),
    .B(net1534),
    .Y(_05493_));
 sg13g2_a21oi_1 _13327_ (.A1(_01538_),
    .A2(net1534),
    .Y(_01082_),
    .B1(_05493_));
 sg13g2_and2_1 _13328_ (.A(net1937),
    .B(net2800),
    .X(_01083_));
 sg13g2_and2_1 _13329_ (.A(net1951),
    .B(net1),
    .X(_01084_));
 sg13g2_and2_1 _13330_ (.A(net1938),
    .B(net1205),
    .X(_01085_));
 sg13g2_and2_1 _13331_ (.A(net1927),
    .B(net1189),
    .X(_01086_));
 sg13g2_and2_1 _13332_ (.A(net1927),
    .B(net1184),
    .X(_01087_));
 sg13g2_and2_1 _13333_ (.A(net1927),
    .B(net1188),
    .X(_01088_));
 sg13g2_and2_1 _13334_ (.A(net1901),
    .B(net1190),
    .X(_01089_));
 sg13g2_and2_1 _13335_ (.A(net1905),
    .B(net1178),
    .X(_01090_));
 sg13g2_and2_1 _13336_ (.A(net1905),
    .B(net1187),
    .X(_01091_));
 sg13g2_and2_1 _13337_ (.A(net1901),
    .B(net1185),
    .X(_01092_));
 sg13g2_and2_1 _13338_ (.A(net1901),
    .B(net1182),
    .X(_01093_));
 sg13g2_and2_1 _13339_ (.A(net1927),
    .B(net1186),
    .X(_01094_));
 sg13g2_and2_1 _13340_ (.A(net1933),
    .B(net1180),
    .X(_01095_));
 sg13g2_and2_1 _13341_ (.A(net1927),
    .B(net1193),
    .X(_01096_));
 sg13g2_and2_1 _13342_ (.A(net1927),
    .B(net1194),
    .X(_01097_));
 sg13g2_and2_1 _13343_ (.A(net1929),
    .B(net1214),
    .X(_01098_));
 sg13g2_and2_1 _13344_ (.A(net1928),
    .B(net1177),
    .X(_01099_));
 sg13g2_and2_1 _13345_ (.A(net1929),
    .B(net1191),
    .X(_01100_));
 sg13g2_and2_1 _13346_ (.A(net1929),
    .B(net1192),
    .X(_01101_));
 sg13g2_nand4_1 _13347_ (.B(net2025),
    .C(_01573_),
    .A(net1174),
    .Y(_05494_),
    .D(net1602));
 sg13g2_o21ai_1 _13348_ (.B1(net1175),
    .Y(_01102_),
    .A1(_01564_),
    .A2(_00173_));
 sg13g2_o21ai_1 _13349_ (.B1(_01937_),
    .Y(_01103_),
    .A1(_01573_),
    .A2(_00173_));
 sg13g2_and2_1 _13350_ (.A(net1951),
    .B(net2),
    .X(_01104_));
 sg13g2_and2_1 _13351_ (.A(net1952),
    .B(net1195),
    .X(_01105_));
 sg13g2_and2_1 _13352_ (.A(net1952),
    .B(net1183),
    .X(_01106_));
 sg13g2_nor2_2 _13353_ (.A(_01194_),
    .B(net1357),
    .Y(_05495_));
 sg13g2_a21oi_1 _13354_ (.A1(net1470),
    .A2(net1598),
    .Y(_05496_),
    .B1(net1884));
 sg13g2_o21ai_1 _13355_ (.B1(_05496_),
    .Y(_01107_),
    .A1(_01221_),
    .A2(net1598));
 sg13g2_a21oi_1 _13356_ (.A1(net1388),
    .A2(net1598),
    .Y(_05497_),
    .B1(net1881));
 sg13g2_o21ai_1 _13357_ (.B1(_05497_),
    .Y(_01108_),
    .A1(_01220_),
    .A2(net1598));
 sg13g2_o21ai_1 _13358_ (.B1(net1938),
    .Y(_05498_),
    .A1(\am_sdr0.nco0.phase_inc[2] ),
    .A2(net1598));
 sg13g2_a21oi_1 _13359_ (.A1(_01219_),
    .A2(net1598),
    .Y(_01109_),
    .B1(_05498_));
 sg13g2_a21oi_1 _13360_ (.A1(net1325),
    .A2(net1598),
    .Y(_05499_),
    .B1(net1883));
 sg13g2_o21ai_1 _13361_ (.B1(_05499_),
    .Y(_01110_),
    .A1(_01218_),
    .A2(net1597));
 sg13g2_o21ai_1 _13362_ (.B1(net1937),
    .Y(_05500_),
    .A1(\am_sdr0.nco0.phase_inc[4] ),
    .A2(net1597));
 sg13g2_a21oi_1 _13363_ (.A1(_01217_),
    .A2(net1597),
    .Y(_01111_),
    .B1(_05500_));
 sg13g2_a21oi_1 _13364_ (.A1(net1330),
    .A2(net1597),
    .Y(_05501_),
    .B1(net1883));
 sg13g2_o21ai_1 _13365_ (.B1(_05501_),
    .Y(_01112_),
    .A1(_01216_),
    .A2(net1597));
 sg13g2_a21oi_1 _13366_ (.A1(net1408),
    .A2(net1597),
    .Y(_05502_),
    .B1(net1881));
 sg13g2_o21ai_1 _13367_ (.B1(_05502_),
    .Y(_01113_),
    .A1(_01215_),
    .A2(net1597));
 sg13g2_a21oi_1 _13368_ (.A1(net1418),
    .A2(net1597),
    .Y(_05503_),
    .B1(net1881));
 sg13g2_o21ai_1 _13369_ (.B1(_05503_),
    .Y(_01114_),
    .A1(_01214_),
    .A2(net1595));
 sg13g2_o21ai_1 _13370_ (.B1(net1935),
    .Y(_05504_),
    .A1(net1506),
    .A2(net1593));
 sg13g2_a21oi_1 _13371_ (.A1(_01213_),
    .A2(net1593),
    .Y(_01115_),
    .B1(_05504_));
 sg13g2_a21oi_1 _13372_ (.A1(net1382),
    .A2(net1593),
    .Y(_05505_),
    .B1(net1882));
 sg13g2_o21ai_1 _13373_ (.B1(_05505_),
    .Y(_01116_),
    .A1(_01212_),
    .A2(net1593));
 sg13g2_o21ai_1 _13374_ (.B1(net1934),
    .Y(_05506_),
    .A1(net1391),
    .A2(net1592));
 sg13g2_a21oi_1 _13375_ (.A1(_01211_),
    .A2(net1592),
    .Y(_01117_),
    .B1(_05506_));
 sg13g2_o21ai_1 _13376_ (.B1(net1934),
    .Y(_05507_),
    .A1(net1507),
    .A2(net1594));
 sg13g2_a21oi_1 _13377_ (.A1(_01210_),
    .A2(net1594),
    .Y(_01118_),
    .B1(_05507_));
 sg13g2_a21oi_1 _13378_ (.A1(net1362),
    .A2(net1596),
    .Y(_05508_),
    .B1(net1882));
 sg13g2_o21ai_1 _13379_ (.B1(_05508_),
    .Y(_01119_),
    .A1(_01209_),
    .A2(net1595));
 sg13g2_o21ai_1 _13380_ (.B1(net1939),
    .Y(_05509_),
    .A1(net1354),
    .A2(net1596));
 sg13g2_a21oi_1 _13381_ (.A1(_01208_),
    .A2(net1595),
    .Y(_01120_),
    .B1(_05509_));
 sg13g2_o21ai_1 _13382_ (.B1(net1939),
    .Y(_05510_),
    .A1(\am_sdr0.nco0.phase_inc[14] ),
    .A2(net1595));
 sg13g2_a21oi_1 _13383_ (.A1(_01207_),
    .A2(net1595),
    .Y(_01121_),
    .B1(_05510_));
 sg13g2_o21ai_1 _13384_ (.B1(net1935),
    .Y(_05511_),
    .A1(\am_sdr0.nco0.phase_inc[15] ),
    .A2(net1595));
 sg13g2_a21oi_1 _13385_ (.A1(_01206_),
    .A2(net1594),
    .Y(_01122_),
    .B1(_05511_));
 sg13g2_a21oi_1 _13386_ (.A1(net1393),
    .A2(net1595),
    .Y(_05512_),
    .B1(net1882));
 sg13g2_o21ai_1 _13387_ (.B1(_05512_),
    .Y(_01123_),
    .A1(_01205_),
    .A2(net1594));
 sg13g2_a21oi_1 _13388_ (.A1(net1360),
    .A2(net1594),
    .Y(_05513_),
    .B1(net1882));
 sg13g2_o21ai_1 _13389_ (.B1(_05513_),
    .Y(_01124_),
    .A1(_01204_),
    .A2(net1594));
 sg13g2_o21ai_1 _13390_ (.B1(net1934),
    .Y(_05514_),
    .A1(\am_sdr0.nco0.phase_inc[18] ),
    .A2(net1594));
 sg13g2_a21oi_1 _13391_ (.A1(_01203_),
    .A2(net1594),
    .Y(_01125_),
    .B1(_05514_));
 sg13g2_o21ai_1 _13392_ (.B1(net1934),
    .Y(_05515_),
    .A1(net1481),
    .A2(net1592));
 sg13g2_a21oi_1 _13393_ (.A1(_01202_),
    .A2(net1592),
    .Y(_01126_),
    .B1(_05515_));
 sg13g2_a21oi_1 _13394_ (.A1(net1381),
    .A2(net1592),
    .Y(_05516_),
    .B1(net1882));
 sg13g2_o21ai_1 _13395_ (.B1(_05516_),
    .Y(_01127_),
    .A1(_01201_),
    .A2(net1593));
 sg13g2_o21ai_1 _13396_ (.B1(net1928),
    .Y(_05517_),
    .A1(net1454),
    .A2(net1591));
 sg13g2_a21oi_1 _13397_ (.A1(_01200_),
    .A2(net1591),
    .Y(_01128_),
    .B1(_05517_));
 sg13g2_o21ai_1 _13398_ (.B1(net1928),
    .Y(_05518_),
    .A1(net2129),
    .A2(net1591));
 sg13g2_a21oi_1 _13399_ (.A1(_01199_),
    .A2(net1591),
    .Y(_01129_),
    .B1(_05518_));
 sg13g2_o21ai_1 _13400_ (.B1(net1928),
    .Y(_05519_),
    .A1(net1417),
    .A2(net1591));
 sg13g2_a21oi_1 _13401_ (.A1(_01197_),
    .A2(net1591),
    .Y(_01130_),
    .B1(_05519_));
 sg13g2_o21ai_1 _13402_ (.B1(net1928),
    .Y(_05520_),
    .A1(net2220),
    .A2(net1592));
 sg13g2_a21oi_1 _13403_ (.A1(_01196_),
    .A2(net1592),
    .Y(_01131_),
    .B1(_05520_));
 sg13g2_o21ai_1 _13404_ (.B1(net1929),
    .Y(_05521_),
    .A1(net2537),
    .A2(net1591));
 sg13g2_a21oi_1 _13405_ (.A1(_01195_),
    .A2(net1591),
    .Y(_01132_),
    .B1(_05521_));
 sg13g2_a21oi_1 _13406_ (.A1(_01569_),
    .A2(net1404),
    .Y(_01133_),
    .B1(_04750_));
 sg13g2_and4_1 _13407_ (.A(net1951),
    .B(_01569_),
    .C(net1404),
    .D(net1615),
    .X(_01134_));
 sg13g2_o21ai_1 _13408_ (.B1(net1958),
    .Y(_05522_),
    .A1(net3051),
    .A2(_05495_));
 sg13g2_a21oi_1 _13409_ (.A1(_01193_),
    .A2(net1599),
    .Y(_01135_),
    .B1(_05522_));
 sg13g2_a21oi_1 _13410_ (.A1(net1482),
    .A2(net1599),
    .Y(_05523_),
    .B1(net1884));
 sg13g2_o21ai_1 _13411_ (.B1(_05523_),
    .Y(_01136_),
    .A1(_01192_),
    .A2(net1599));
 sg13g2_o21ai_1 _13412_ (.B1(net1957),
    .Y(_05524_),
    .A1(net2644),
    .A2(net1599));
 sg13g2_a21oi_1 _13413_ (.A1(_01191_),
    .A2(net1599),
    .Y(_01137_),
    .B1(_05524_));
 sg13g2_nand2_1 _13414_ (.Y(_05525_),
    .A(net2054),
    .B(net2136));
 sg13g2_o21ai_1 _13415_ (.B1(net1937),
    .Y(_05526_),
    .A1(net2054),
    .A2(net2136));
 sg13g2_nor2b_1 _13416_ (.A(_05526_),
    .B_N(_05525_),
    .Y(_01138_));
 sg13g2_nand2_1 _13417_ (.Y(_05527_),
    .A(\am_sdr0.nco0.phase_inc[1] ),
    .B(\am_sdr0.nco0.phase[1] ));
 sg13g2_xnor2_1 _13418_ (.Y(_05528_),
    .A(net3168),
    .B(net3066));
 sg13g2_and2_1 _13419_ (.A(_05525_),
    .B(_05528_),
    .X(_05529_));
 sg13g2_nor2_1 _13420_ (.A(_05525_),
    .B(_05528_),
    .Y(_05530_));
 sg13g2_nor3_1 _13421_ (.A(net1883),
    .B(_05529_),
    .C(_05530_),
    .Y(_01139_));
 sg13g2_and2_1 _13422_ (.A(\am_sdr0.nco0.phase_inc[2] ),
    .B(\am_sdr0.nco0.phase[2] ),
    .X(_05531_));
 sg13g2_xnor2_1 _13423_ (.Y(_05532_),
    .A(\am_sdr0.nco0.phase_inc[2] ),
    .B(\am_sdr0.nco0.phase[2] ));
 sg13g2_inv_1 _13424_ (.Y(_05533_),
    .A(_05532_));
 sg13g2_a21oi_1 _13425_ (.A1(net2554),
    .A2(net3066),
    .Y(_05534_),
    .B1(_05530_));
 sg13g2_o21ai_1 _13426_ (.B1(_05527_),
    .Y(_05535_),
    .A1(_05525_),
    .A2(_05528_));
 sg13g2_o21ai_1 _13427_ (.B1(net1938),
    .Y(_05536_),
    .A1(_05532_),
    .A2(_05534_));
 sg13g2_a21oi_1 _13428_ (.A1(_05532_),
    .A2(_05534_),
    .Y(_01140_),
    .B1(_05536_));
 sg13g2_nand2_1 _13429_ (.Y(_05537_),
    .A(\am_sdr0.nco0.phase_inc[3] ),
    .B(\am_sdr0.nco0.phase[3] ));
 sg13g2_xnor2_1 _13430_ (.Y(_05538_),
    .A(net3281),
    .B(net3247));
 sg13g2_a21oi_1 _13431_ (.A1(_05533_),
    .A2(_05535_),
    .Y(_05539_),
    .B1(_05531_));
 sg13g2_nor2_1 _13432_ (.A(_05538_),
    .B(_05539_),
    .Y(_05540_));
 sg13g2_a21oi_1 _13433_ (.A1(_05538_),
    .A2(_05539_),
    .Y(_05541_),
    .B1(net1881));
 sg13g2_nor2b_1 _13434_ (.A(_05540_),
    .B_N(_05541_),
    .Y(_01141_));
 sg13g2_a21oi_1 _13435_ (.A1(net2745),
    .A2(net3247),
    .Y(_05542_),
    .B1(_05540_));
 sg13g2_o21ai_1 _13436_ (.B1(_05537_),
    .Y(_05543_),
    .A1(_05538_),
    .A2(_05539_));
 sg13g2_xnor2_1 _13437_ (.Y(_05544_),
    .A(\am_sdr0.nco0.phase_inc[4] ),
    .B(net3108));
 sg13g2_nor2_1 _13438_ (.A(_05542_),
    .B(_05544_),
    .Y(_05545_));
 sg13g2_a21oi_1 _13439_ (.A1(_05542_),
    .A2(_05544_),
    .Y(_05546_),
    .B1(net1881));
 sg13g2_nor2b_1 _13440_ (.A(_05545_),
    .B_N(_05546_),
    .Y(_01142_));
 sg13g2_nand2_1 _13441_ (.Y(_05547_),
    .A(net2193),
    .B(\am_sdr0.nco0.phase[5] ));
 sg13g2_or2_1 _13442_ (.X(_05548_),
    .B(\am_sdr0.nco0.phase[5] ),
    .A(net2193));
 sg13g2_nand2_1 _13443_ (.Y(_05549_),
    .A(_05547_),
    .B(_05548_));
 sg13g2_a21oi_1 _13444_ (.A1(\am_sdr0.nco0.phase_inc[4] ),
    .A2(net3108),
    .Y(_05550_),
    .B1(_05545_));
 sg13g2_o21ai_1 _13445_ (.B1(net1937),
    .Y(_05551_),
    .A1(_05549_),
    .A2(net3109));
 sg13g2_a21oi_1 _13446_ (.A1(_05549_),
    .A2(net3109),
    .Y(_01143_),
    .B1(_05551_));
 sg13g2_nand2_1 _13447_ (.Y(_05552_),
    .A(\am_sdr0.nco0.phase_inc[6] ),
    .B(\am_sdr0.nco0.phase[6] ));
 sg13g2_xnor2_1 _13448_ (.Y(_05553_),
    .A(net2244),
    .B(net3095));
 sg13g2_nor2_1 _13449_ (.A(_05544_),
    .B(_05549_),
    .Y(_05554_));
 sg13g2_nand3_1 _13450_ (.B(\am_sdr0.nco0.phase[4] ),
    .C(_05548_),
    .A(\am_sdr0.nco0.phase_inc[4] ),
    .Y(_05555_));
 sg13g2_nand2_1 _13451_ (.Y(_05556_),
    .A(_05547_),
    .B(_05555_));
 sg13g2_a21oi_2 _13452_ (.B1(_05556_),
    .Y(_05557_),
    .A2(_05554_),
    .A1(_05543_));
 sg13g2_o21ai_1 _13453_ (.B1(net1937),
    .Y(_05558_),
    .A1(_05553_),
    .A2(_05557_));
 sg13g2_a21oi_1 _13454_ (.A1(_05553_),
    .A2(_05557_),
    .Y(_01144_),
    .B1(_05558_));
 sg13g2_o21ai_1 _13455_ (.B1(_05552_),
    .Y(_05559_),
    .A1(_05553_),
    .A2(_05557_));
 sg13g2_and2_1 _13456_ (.A(net2091),
    .B(\am_sdr0.nco0.phase[7] ),
    .X(_05560_));
 sg13g2_or2_1 _13457_ (.X(_05561_),
    .B(\am_sdr0.nco0.phase[7] ),
    .A(\am_sdr0.nco0.phase_inc[7] ));
 sg13g2_nand2b_1 _13458_ (.Y(_05562_),
    .B(_05561_),
    .A_N(_05560_));
 sg13g2_nand2b_1 _13459_ (.Y(_05563_),
    .B(_05562_),
    .A_N(_05559_));
 sg13g2_nand2b_1 _13460_ (.Y(_05564_),
    .B(_05559_),
    .A_N(_05562_));
 sg13g2_and3_1 _13461_ (.X(_01145_),
    .A(net1937),
    .B(_05563_),
    .C(_05564_));
 sg13g2_a21oi_2 _13462_ (.B1(_05560_),
    .Y(_05565_),
    .A2(_05561_),
    .A1(_05559_));
 sg13g2_nand2_1 _13463_ (.Y(_05566_),
    .A(net1506),
    .B(net3082));
 sg13g2_xnor2_1 _13464_ (.Y(_05567_),
    .A(net1506),
    .B(net3082));
 sg13g2_or2_1 _13465_ (.X(_05568_),
    .B(_05567_),
    .A(_05565_));
 sg13g2_nand2_1 _13466_ (.Y(_05569_),
    .A(net1934),
    .B(_05568_));
 sg13g2_a21oi_1 _13467_ (.A1(_05565_),
    .A2(_05567_),
    .Y(_01146_),
    .B1(_05569_));
 sg13g2_nor2_1 _13468_ (.A(net2076),
    .B(net3184),
    .Y(_05570_));
 sg13g2_nand2_1 _13469_ (.Y(_05571_),
    .A(net2076),
    .B(net3184));
 sg13g2_nand2b_1 _13470_ (.Y(_05572_),
    .B(_05571_),
    .A_N(_05570_));
 sg13g2_and3_1 _13471_ (.X(_05573_),
    .A(_05566_),
    .B(_05568_),
    .C(_05572_));
 sg13g2_a21oi_1 _13472_ (.A1(_05566_),
    .A2(_05568_),
    .Y(_05574_),
    .B1(_05572_));
 sg13g2_nor3_1 _13473_ (.A(net1882),
    .B(_05573_),
    .C(_05574_),
    .Y(_01147_));
 sg13g2_nand2_1 _13474_ (.Y(_05575_),
    .A(net1391),
    .B(net3073));
 sg13g2_xnor2_1 _13475_ (.Y(_05576_),
    .A(net1391),
    .B(net3073));
 sg13g2_o21ai_1 _13476_ (.B1(_05571_),
    .Y(_05577_),
    .A1(_05566_),
    .A2(_05570_));
 sg13g2_nor2_1 _13477_ (.A(_05567_),
    .B(_05572_),
    .Y(_05578_));
 sg13g2_nor2b_1 _13478_ (.A(_05565_),
    .B_N(_05578_),
    .Y(_05579_));
 sg13g2_nor2_1 _13479_ (.A(_05577_),
    .B(_05579_),
    .Y(_05580_));
 sg13g2_or2_1 _13480_ (.X(_05581_),
    .B(_05580_),
    .A(_05576_));
 sg13g2_nand2_1 _13481_ (.Y(_05582_),
    .A(net1934),
    .B(_05581_));
 sg13g2_a21oi_1 _13482_ (.A1(_05576_),
    .A2(_05580_),
    .Y(_01148_),
    .B1(_05582_));
 sg13g2_nor2_1 _13483_ (.A(\am_sdr0.nco0.phase_inc[11] ),
    .B(\am_sdr0.nco0.phase[11] ),
    .Y(_05583_));
 sg13g2_xnor2_1 _13484_ (.Y(_05584_),
    .A(net1507),
    .B(net3196));
 sg13g2_nand3_1 _13485_ (.B(_05581_),
    .C(_05584_),
    .A(_05575_),
    .Y(_05585_));
 sg13g2_a21oi_1 _13486_ (.A1(_05575_),
    .A2(_05581_),
    .Y(_05586_),
    .B1(_05584_));
 sg13g2_nand2_1 _13487_ (.Y(_05587_),
    .A(net1934),
    .B(_05585_));
 sg13g2_nor2_1 _13488_ (.A(_05586_),
    .B(_05587_),
    .Y(_01149_));
 sg13g2_nand2_1 _13489_ (.Y(_05588_),
    .A(net2439),
    .B(net3210));
 sg13g2_xnor2_1 _13490_ (.Y(_05589_),
    .A(net2439),
    .B(net3210));
 sg13g2_nor2_1 _13491_ (.A(_05576_),
    .B(_05584_),
    .Y(_05590_));
 sg13g2_nor2_1 _13492_ (.A(_05575_),
    .B(_05583_),
    .Y(_05591_));
 sg13g2_a221oi_1 _13493_ (.B2(_05590_),
    .C1(_05591_),
    .B1(_05577_),
    .A1(\am_sdr0.nco0.phase_inc[11] ),
    .Y(_05592_),
    .A2(\am_sdr0.nco0.phase[11] ));
 sg13g2_nand2_1 _13494_ (.Y(_05593_),
    .A(_05578_),
    .B(_05590_));
 sg13g2_o21ai_1 _13495_ (.B1(_05592_),
    .Y(_05594_),
    .A1(_05565_),
    .A2(_05593_));
 sg13g2_nand2b_1 _13496_ (.Y(_05595_),
    .B(_05589_),
    .A_N(_05594_));
 sg13g2_nand2b_1 _13497_ (.Y(_05596_),
    .B(_05594_),
    .A_N(_05589_));
 sg13g2_and3_1 _13498_ (.X(_01150_),
    .A(net1935),
    .B(_05595_),
    .C(_05596_));
 sg13g2_nor2_1 _13499_ (.A(\am_sdr0.nco0.phase_inc[13] ),
    .B(\am_sdr0.nco0.phase[13] ),
    .Y(_05597_));
 sg13g2_nand2_1 _13500_ (.Y(_05598_),
    .A(net1354),
    .B(\am_sdr0.nco0.phase[13] ));
 sg13g2_nand2b_1 _13501_ (.Y(_05599_),
    .B(_05598_),
    .A_N(_05597_));
 sg13g2_nand3_1 _13502_ (.B(_05596_),
    .C(_05599_),
    .A(_05588_),
    .Y(_05600_));
 sg13g2_a21oi_1 _13503_ (.A1(_05588_),
    .A2(_05596_),
    .Y(_05601_),
    .B1(_05599_));
 sg13g2_nand2_1 _13504_ (.Y(_05602_),
    .A(net1935),
    .B(_05600_));
 sg13g2_nor2_1 _13505_ (.A(_05601_),
    .B(_05602_),
    .Y(_01151_));
 sg13g2_nand2_1 _13506_ (.Y(_05603_),
    .A(\am_sdr0.nco0.phase_inc[14] ),
    .B(net3115));
 sg13g2_xnor2_1 _13507_ (.Y(_05604_),
    .A(\am_sdr0.nco0.phase_inc[14] ),
    .B(net3115));
 sg13g2_o21ai_1 _13508_ (.B1(_05598_),
    .Y(_05605_),
    .A1(_05588_),
    .A2(_05597_));
 sg13g2_nor2_1 _13509_ (.A(_05589_),
    .B(_05599_),
    .Y(_05606_));
 sg13g2_a21oi_1 _13510_ (.A1(_05594_),
    .A2(_05606_),
    .Y(_05607_),
    .B1(_05605_));
 sg13g2_or2_1 _13511_ (.X(_05608_),
    .B(_05607_),
    .A(_05604_));
 sg13g2_nand2_1 _13512_ (.Y(_05609_),
    .A(net1935),
    .B(_05608_));
 sg13g2_a21oi_1 _13513_ (.A1(net3116),
    .A2(_05607_),
    .Y(_01152_),
    .B1(_05609_));
 sg13g2_nor2_1 _13514_ (.A(\am_sdr0.nco0.phase_inc[15] ),
    .B(\am_sdr0.nco0.phase[15] ),
    .Y(_05610_));
 sg13g2_xnor2_1 _13515_ (.Y(_05611_),
    .A(\am_sdr0.nco0.phase_inc[15] ),
    .B(net3191));
 sg13g2_and3_1 _13516_ (.X(_05612_),
    .A(_05603_),
    .B(_05608_),
    .C(_05611_));
 sg13g2_a21oi_1 _13517_ (.A1(_05603_),
    .A2(_05608_),
    .Y(_05613_),
    .B1(net3192));
 sg13g2_nor3_1 _13518_ (.A(net1882),
    .B(_05612_),
    .C(net3193),
    .Y(_01153_));
 sg13g2_nor2_1 _13519_ (.A(_05604_),
    .B(_05611_),
    .Y(_05614_));
 sg13g2_nand2_1 _13520_ (.Y(_05615_),
    .A(_05606_),
    .B(_05614_));
 sg13g2_or2_1 _13521_ (.X(_05616_),
    .B(_05615_),
    .A(_05593_));
 sg13g2_nor2_1 _13522_ (.A(_05603_),
    .B(_05610_),
    .Y(_05617_));
 sg13g2_a21oi_1 _13523_ (.A1(\am_sdr0.nco0.phase_inc[15] ),
    .A2(\am_sdr0.nco0.phase[15] ),
    .Y(_05618_),
    .B1(_05617_));
 sg13g2_o21ai_1 _13524_ (.B1(_05618_),
    .Y(_05619_),
    .A1(_05592_),
    .A2(_05615_));
 sg13g2_a21oi_1 _13525_ (.A1(_05605_),
    .A2(_05614_),
    .Y(_05620_),
    .B1(_05619_));
 sg13g2_o21ai_1 _13526_ (.B1(_05620_),
    .Y(_05621_),
    .A1(_05565_),
    .A2(_05616_));
 sg13g2_nand2_1 _13527_ (.Y(_05622_),
    .A(net2498),
    .B(net3229));
 sg13g2_xnor2_1 _13528_ (.Y(_05623_),
    .A(net2498),
    .B(net3229));
 sg13g2_nand2b_1 _13529_ (.Y(_05624_),
    .B(_05623_),
    .A_N(_05621_));
 sg13g2_nand2b_1 _13530_ (.Y(_05625_),
    .B(_05621_),
    .A_N(_05623_));
 sg13g2_and3_1 _13531_ (.X(_01154_),
    .A(net1935),
    .B(_05624_),
    .C(_05625_));
 sg13g2_nor2_1 _13532_ (.A(\am_sdr0.nco0.phase_inc[17] ),
    .B(\am_sdr0.nco0.phase[17] ),
    .Y(_05626_));
 sg13g2_nand2_1 _13533_ (.Y(_05627_),
    .A(net2093),
    .B(\am_sdr0.nco0.phase[17] ));
 sg13g2_nand2b_1 _13534_ (.Y(_05628_),
    .B(_05627_),
    .A_N(_05626_));
 sg13g2_nand3_1 _13535_ (.B(_05625_),
    .C(_05628_),
    .A(_05622_),
    .Y(_05629_));
 sg13g2_a21o_1 _13536_ (.A2(_05625_),
    .A1(_05622_),
    .B1(_05628_),
    .X(_05630_));
 sg13g2_and3_1 _13537_ (.X(_01155_),
    .A(net1935),
    .B(_05629_),
    .C(_05630_));
 sg13g2_nand2_1 _13538_ (.Y(_05631_),
    .A(\am_sdr0.nco0.phase_inc[18] ),
    .B(net3031));
 sg13g2_xnor2_1 _13539_ (.Y(_05632_),
    .A(\am_sdr0.nco0.phase_inc[18] ),
    .B(net3031));
 sg13g2_o21ai_1 _13540_ (.B1(_05627_),
    .Y(_05633_),
    .A1(_05622_),
    .A2(_05626_));
 sg13g2_nor2_1 _13541_ (.A(_05623_),
    .B(_05628_),
    .Y(_05634_));
 sg13g2_a21oi_1 _13542_ (.A1(_05621_),
    .A2(_05634_),
    .Y(_05635_),
    .B1(_05633_));
 sg13g2_or2_1 _13543_ (.X(_05636_),
    .B(_05635_),
    .A(_05632_));
 sg13g2_nand2_1 _13544_ (.Y(_05637_),
    .A(net1934),
    .B(_05636_));
 sg13g2_a21oi_1 _13545_ (.A1(net3032),
    .A2(_05635_),
    .Y(_01156_),
    .B1(_05637_));
 sg13g2_nor2_1 _13546_ (.A(\am_sdr0.nco0.phase_inc[19] ),
    .B(\am_sdr0.nco0.phase[19] ),
    .Y(_05638_));
 sg13g2_xnor2_1 _13547_ (.Y(_05639_),
    .A(net1481),
    .B(net3188));
 sg13g2_and3_1 _13548_ (.X(_05640_),
    .A(_05631_),
    .B(_05636_),
    .C(_05639_));
 sg13g2_a21oi_1 _13549_ (.A1(_05631_),
    .A2(_05636_),
    .Y(_05641_),
    .B1(_05639_));
 sg13g2_nor3_1 _13550_ (.A(net1882),
    .B(_05640_),
    .C(net3189),
    .Y(_01157_));
 sg13g2_nor2_1 _13551_ (.A(_05632_),
    .B(_05639_),
    .Y(_05642_));
 sg13g2_and2_1 _13552_ (.A(_05634_),
    .B(_05642_),
    .X(_05643_));
 sg13g2_a22oi_1 _13553_ (.Y(_05644_),
    .B1(_05633_),
    .B2(_05642_),
    .A2(\am_sdr0.nco0.phase[19] ),
    .A1(\am_sdr0.nco0.phase_inc[19] ));
 sg13g2_o21ai_1 _13554_ (.B1(_05644_),
    .Y(_05645_),
    .A1(_05631_),
    .A2(_05638_));
 sg13g2_a21oi_2 _13555_ (.B1(_05645_),
    .Y(_05646_),
    .A2(_05643_),
    .A1(_05621_));
 sg13g2_a21o_1 _13556_ (.A2(_05643_),
    .A1(_05621_),
    .B1(_05645_),
    .X(_05647_));
 sg13g2_nand2_1 _13557_ (.Y(_05648_),
    .A(net2557),
    .B(net3090));
 sg13g2_xnor2_1 _13558_ (.Y(_05649_),
    .A(net2557),
    .B(net3090));
 sg13g2_nand2b_1 _13559_ (.Y(_05650_),
    .B(_05647_),
    .A_N(_05649_));
 sg13g2_nand2_1 _13560_ (.Y(_05651_),
    .A(net1928),
    .B(_05650_));
 sg13g2_a21oi_1 _13561_ (.A1(_05646_),
    .A2(_05649_),
    .Y(_01158_),
    .B1(_05651_));
 sg13g2_nor2_1 _13562_ (.A(net1454),
    .B(net3174),
    .Y(_05652_));
 sg13g2_nand2_1 _13563_ (.Y(_05653_),
    .A(net1454),
    .B(net3174));
 sg13g2_nand2b_1 _13564_ (.Y(_05654_),
    .B(_05653_),
    .A_N(_05652_));
 sg13g2_nand3_1 _13565_ (.B(_05650_),
    .C(_05654_),
    .A(_05648_),
    .Y(_05655_));
 sg13g2_a21oi_1 _13566_ (.A1(_05648_),
    .A2(_05650_),
    .Y(_05656_),
    .B1(_05654_));
 sg13g2_nand2_1 _13567_ (.Y(_05657_),
    .A(net1929),
    .B(_05655_));
 sg13g2_nor2_1 _13568_ (.A(_05656_),
    .B(_05657_),
    .Y(_01159_));
 sg13g2_nand2_1 _13569_ (.Y(_05658_),
    .A(net2129),
    .B(net3018));
 sg13g2_xnor2_1 _13570_ (.Y(_05659_),
    .A(net2129),
    .B(net1654));
 sg13g2_nor2_1 _13571_ (.A(_05649_),
    .B(_05654_),
    .Y(_05660_));
 sg13g2_o21ai_1 _13572_ (.B1(_05653_),
    .Y(_05661_),
    .A1(_05648_),
    .A2(_05652_));
 sg13g2_a21oi_1 _13573_ (.A1(_05647_),
    .A2(_05660_),
    .Y(_05662_),
    .B1(_05661_));
 sg13g2_or2_1 _13574_ (.X(_05663_),
    .B(_05662_),
    .A(_05659_));
 sg13g2_nand2_1 _13575_ (.Y(_05664_),
    .A(net1928),
    .B(_05663_));
 sg13g2_a21oi_1 _13576_ (.A1(_05659_),
    .A2(_05662_),
    .Y(_01160_),
    .B1(_05664_));
 sg13g2_xnor2_1 _13577_ (.Y(_05665_),
    .A(\am_sdr0.nco0.phase_inc[23] ),
    .B(net1653));
 sg13g2_nand3_1 _13578_ (.B(_05663_),
    .C(_05665_),
    .A(_05658_),
    .Y(_05666_));
 sg13g2_a21o_1 _13579_ (.A2(_05663_),
    .A1(_05658_),
    .B1(_05665_),
    .X(_05667_));
 sg13g2_and3_1 _13580_ (.X(_01161_),
    .A(net1927),
    .B(_05666_),
    .C(_05667_));
 sg13g2_and2_1 _13581_ (.A(net2220),
    .B(net2130),
    .X(_05668_));
 sg13g2_xor2_1 _13582_ (.B(net2130),
    .A(net2220),
    .X(_05669_));
 sg13g2_nor2_1 _13583_ (.A(_05659_),
    .B(_05665_),
    .Y(_05670_));
 sg13g2_nand2_1 _13584_ (.Y(_05671_),
    .A(_05660_),
    .B(_05670_));
 sg13g2_a21oi_1 _13585_ (.A1(_01198_),
    .A2(_01575_),
    .Y(_05672_),
    .B1(_05658_));
 sg13g2_a221oi_1 _13586_ (.B2(_05670_),
    .C1(_05672_),
    .B1(_05661_),
    .A1(\am_sdr0.nco0.phase_inc[23] ),
    .Y(_05673_),
    .A2(\am_sdr0.nco0.phase[23] ));
 sg13g2_o21ai_1 _13587_ (.B1(_05673_),
    .Y(_05674_),
    .A1(_05646_),
    .A2(_05671_));
 sg13g2_nor2_1 _13588_ (.A(_05669_),
    .B(_05674_),
    .Y(_05675_));
 sg13g2_a21oi_1 _13589_ (.A1(_05669_),
    .A2(_05674_),
    .Y(_05676_),
    .B1(net1880));
 sg13g2_nor2b_1 _13590_ (.A(_05675_),
    .B_N(_05676_),
    .Y(_01162_));
 sg13g2_a21oi_1 _13591_ (.A1(_05669_),
    .A2(_05674_),
    .Y(_05677_),
    .B1(_05668_));
 sg13g2_xnor2_1 _13592_ (.Y(_05678_),
    .A(net2537),
    .B(net1650));
 sg13g2_o21ai_1 _13593_ (.B1(net1928),
    .Y(_05679_),
    .A1(_05677_),
    .A2(_05678_));
 sg13g2_a21oi_1 _13594_ (.A1(_05677_),
    .A2(_05678_),
    .Y(_01163_),
    .B1(_05679_));
 sg13g2_and2_1 _13595_ (.A(net1951),
    .B(net4),
    .X(_01164_));
 sg13g2_and2_1 _13596_ (.A(net1951),
    .B(net1181),
    .X(_01165_));
 sg13g2_and2_1 _13597_ (.A(net1951),
    .B(net1404),
    .X(_01166_));
 sg13g2_and2_1 _13598_ (.A(net1951),
    .B(net3),
    .X(_01167_));
 sg13g2_nand2_1 _13599_ (.Y(_05680_),
    .A(_01188_),
    .B(\am_sdr0.count[1] ));
 sg13g2_nor2b_1 _13600_ (.A(\am_sdr0.count[0] ),
    .B_N(\am_sdr0.am0.demod_out[8] ),
    .Y(_05681_));
 sg13g2_nor2_1 _13601_ (.A(_01188_),
    .B(\am_sdr0.count[1] ),
    .Y(_05682_));
 sg13g2_a221oi_1 _13602_ (.B2(_05681_),
    .C1(_05682_),
    .B1(_05680_),
    .A1(\am_sdr0.am0.demod_out[10] ),
    .Y(_05683_),
    .A2(_01587_));
 sg13g2_a221oi_1 _13603_ (.B2(_01186_),
    .C1(_05683_),
    .B1(\am_sdr0.count[2] ),
    .A1(_01184_),
    .Y(_05684_),
    .A2(\am_sdr0.count[3] ));
 sg13g2_a221oi_1 _13604_ (.B2(\am_sdr0.am0.demod_out[11] ),
    .C1(_05684_),
    .B1(_01586_),
    .A1(\am_sdr0.am0.demod_out[12] ),
    .Y(_05685_),
    .A2(_01585_));
 sg13g2_a221oi_1 _13605_ (.B2(_01182_),
    .C1(_05685_),
    .B1(\am_sdr0.count[4] ),
    .A1(_01180_),
    .Y(_05686_),
    .A2(\am_sdr0.count[5] ));
 sg13g2_a21oi_1 _13606_ (.A1(\am_sdr0.am0.demod_out[13] ),
    .A2(_01584_),
    .Y(_05687_),
    .B1(_05686_));
 sg13g2_a21oi_1 _13607_ (.A1(_01178_),
    .A2(net1870),
    .Y(_05688_),
    .B1(_05687_));
 sg13g2_a221oi_1 _13608_ (.B2(\am_sdr0.am0.demod_out[14] ),
    .C1(_05688_),
    .B1(_01583_),
    .A1(\am_sdr0.am0.demod_out[15] ),
    .Y(_05689_),
    .A2(net1621));
 sg13g2_nor2_1 _13609_ (.A(\am_sdr0.am0.demod_out[15] ),
    .B(net1621),
    .Y(_05690_));
 sg13g2_or2_1 _13610_ (.X(_05691_),
    .B(\am_sdr0.gain_spi[0] ),
    .A(\am_sdr0.gain_spi[1] ));
 sg13g2_nor4_1 _13611_ (.A(\am_sdr0.gain_spi[2] ),
    .B(_05689_),
    .C(_05690_),
    .D(_05691_),
    .Y(_05692_));
 sg13g2_nor2_1 _13612_ (.A(net1647),
    .B(_01586_),
    .Y(_05693_));
 sg13g2_nand2_1 _13613_ (.Y(_05694_),
    .A(\am_sdr0.am0.demod_out[8] ),
    .B(_01587_));
 sg13g2_a22oi_1 _13614_ (.Y(_05695_),
    .B1(_01586_),
    .B2(net1647),
    .A2(_01585_),
    .A1(\am_sdr0.am0.demod_out[10] ));
 sg13g2_o21ai_1 _13615_ (.B1(_05695_),
    .Y(_05696_),
    .A1(_05693_),
    .A2(_05694_));
 sg13g2_a22oi_1 _13616_ (.Y(_05697_),
    .B1(\am_sdr0.count[4] ),
    .B2(_01186_),
    .A2(\am_sdr0.count[5] ),
    .A1(_01184_));
 sg13g2_a22oi_1 _13617_ (.Y(_05698_),
    .B1(_05696_),
    .B2(_05697_),
    .A2(_01584_),
    .A1(\am_sdr0.am0.demod_out[11] ));
 sg13g2_a21oi_1 _13618_ (.A1(_01182_),
    .A2(net1870),
    .Y(_05699_),
    .B1(_05698_));
 sg13g2_a221oi_1 _13619_ (.B2(\am_sdr0.am0.demod_out[12] ),
    .C1(_05699_),
    .B1(_01583_),
    .A1(\am_sdr0.am0.demod_out[13] ),
    .Y(_05700_),
    .A2(net1621));
 sg13g2_nand2_1 _13620_ (.Y(_05701_),
    .A(_01180_),
    .B(\am_sdr0.count[7] ));
 sg13g2_nand3_1 _13621_ (.B(_00046_),
    .C(_05701_),
    .A(\am_sdr0.gain_spi[1] ),
    .Y(_05702_));
 sg13g2_or3_1 _13622_ (.A(\am_sdr0.gain_spi[0] ),
    .B(_05700_),
    .C(_05702_),
    .X(_05703_));
 sg13g2_a22oi_1 _13623_ (.Y(_05704_),
    .B1(_01586_),
    .B2(\am_sdr0.am0.demod_out[8] ),
    .A2(_01585_),
    .A1(net1647));
 sg13g2_a221oi_1 _13624_ (.B2(_01188_),
    .C1(_05704_),
    .B1(\am_sdr0.count[4] ),
    .A1(_01186_),
    .Y(_05705_),
    .A2(\am_sdr0.count[5] ));
 sg13g2_nand2_1 _13625_ (.Y(_05706_),
    .A(\am_sdr0.gain_spi[1] ),
    .B(\am_sdr0.gain_spi[0] ));
 sg13g2_or2_1 _13626_ (.X(_05707_),
    .B(_05706_),
    .A(\am_sdr0.gain_spi[2] ));
 sg13g2_a221oi_1 _13627_ (.B2(\am_sdr0.am0.demod_out[10] ),
    .C1(_05705_),
    .B1(_01584_),
    .A1(\am_sdr0.am0.demod_out[11] ),
    .Y(_05708_),
    .A2(_01583_));
 sg13g2_a221oi_1 _13628_ (.B2(_01184_),
    .C1(_05708_),
    .B1(net1870),
    .A1(_01182_),
    .Y(_05709_),
    .A2(\am_sdr0.count[7] ));
 sg13g2_a21oi_1 _13629_ (.A1(\am_sdr0.am0.demod_out[12] ),
    .A2(net1621),
    .Y(_05710_),
    .B1(_05709_));
 sg13g2_o21ai_1 _13630_ (.B1(_05703_),
    .Y(_05711_),
    .A1(_05707_),
    .A2(_05710_));
 sg13g2_nand2b_1 _13631_ (.Y(_05712_),
    .B(\am_sdr0.am0.demod_out[8] ),
    .A_N(\am_sdr0.count[1] ));
 sg13g2_a21oi_1 _13632_ (.A1(_01188_),
    .A2(\am_sdr0.count[2] ),
    .Y(_05713_),
    .B1(_05712_));
 sg13g2_a221oi_1 _13633_ (.B2(net1647),
    .C1(_05713_),
    .B1(_01587_),
    .A1(\am_sdr0.am0.demod_out[10] ),
    .Y(_05714_),
    .A2(_01586_));
 sg13g2_a221oi_1 _13634_ (.B2(_01186_),
    .C1(_05714_),
    .B1(\am_sdr0.count[3] ),
    .A1(_01184_),
    .Y(_05715_),
    .A2(\am_sdr0.count[4] ));
 sg13g2_a221oi_1 _13635_ (.B2(\am_sdr0.am0.demod_out[11] ),
    .C1(_05715_),
    .B1(_01585_),
    .A1(\am_sdr0.am0.demod_out[12] ),
    .Y(_05716_),
    .A2(_01584_));
 sg13g2_a221oi_1 _13636_ (.B2(_01182_),
    .C1(_05716_),
    .B1(\am_sdr0.count[5] ),
    .A1(_01180_),
    .Y(_05717_),
    .A2(net1870));
 sg13g2_a221oi_1 _13637_ (.B2(\am_sdr0.am0.demod_out[13] ),
    .C1(_05717_),
    .B1(_01583_),
    .A1(\am_sdr0.am0.demod_out[14] ),
    .Y(_05718_),
    .A2(net1621));
 sg13g2_a21oi_1 _13638_ (.A1(_01178_),
    .A2(\am_sdr0.count[7] ),
    .Y(_05719_),
    .B1(_05718_));
 sg13g2_nand4_1 _13639_ (.B(\am_sdr0.gain_spi[0] ),
    .C(net2480),
    .A(_01192_),
    .Y(_05720_),
    .D(_05719_));
 sg13g2_nor2_1 _13640_ (.A(net1647),
    .B(_01584_),
    .Y(_05721_));
 sg13g2_nand2_1 _13641_ (.Y(_05722_),
    .A(\am_sdr0.am0.demod_out[8] ),
    .B(_01585_));
 sg13g2_a22oi_1 _13642_ (.Y(_05723_),
    .B1(_01584_),
    .B2(net1647),
    .A2(_01583_),
    .A1(\am_sdr0.am0.demod_out[10] ));
 sg13g2_o21ai_1 _13643_ (.B1(_05723_),
    .Y(_05724_),
    .A1(_05721_),
    .A2(_05722_));
 sg13g2_a22oi_1 _13644_ (.Y(_05725_),
    .B1(net1870),
    .B2(_01186_),
    .A2(\am_sdr0.count[7] ),
    .A1(_01184_));
 sg13g2_a22oi_1 _13645_ (.Y(_05726_),
    .B1(_05724_),
    .B2(_05725_),
    .A2(_01582_),
    .A1(\am_sdr0.am0.demod_out[11] ));
 sg13g2_nor3_1 _13646_ (.A(net2480),
    .B(_05691_),
    .C(_05726_),
    .Y(_05727_));
 sg13g2_nand2_1 _13647_ (.Y(_05728_),
    .A(net2480),
    .B(_05706_));
 sg13g2_and3_1 _13648_ (.X(_05729_),
    .A(_05691_),
    .B(_05707_),
    .C(_05728_));
 sg13g2_nor4_1 _13649_ (.A(_05692_),
    .B(_05711_),
    .C(_05727_),
    .D(_05729_),
    .Y(_05730_));
 sg13g2_a22oi_1 _13650_ (.Y(_05731_),
    .B1(_01584_),
    .B2(\am_sdr0.am0.demod_out[8] ),
    .A2(_01583_),
    .A1(net1647));
 sg13g2_a221oi_1 _13651_ (.B2(_01188_),
    .C1(_05731_),
    .B1(\am_sdr0.count[6] ),
    .A1(_01186_),
    .Y(_05732_),
    .A2(\am_sdr0.count[7] ));
 sg13g2_a21oi_1 _13652_ (.A1(\am_sdr0.am0.demod_out[10] ),
    .A2(net1621),
    .Y(_05733_),
    .B1(_05732_));
 sg13g2_a221oi_1 _13653_ (.B2(_05729_),
    .C1(net1891),
    .B1(_05733_),
    .A1(net2481),
    .Y(_01168_),
    .A2(_05730_));
 sg13g2_a22oi_1 _13654_ (.Y(_05734_),
    .B1(net1616),
    .B2(net2301),
    .A2(net1617),
    .A1(net2582));
 sg13g2_inv_1 _13655_ (.Y(_01169_),
    .A(_05734_));
 sg13g2_a22oi_1 _13656_ (.Y(_05735_),
    .B1(net1616),
    .B2(\am_sdr0.am0.q[1] ),
    .A2(net1617),
    .A1(net1402));
 sg13g2_inv_1 _13657_ (.Y(_01170_),
    .A(net1403));
 sg13g2_a22oi_1 _13658_ (.Y(_05736_),
    .B1(net1616),
    .B2(net2127),
    .A2(net1617),
    .A1(\am_sdr0.am0.demod_out[10] ));
 sg13g2_inv_1 _13659_ (.Y(_01171_),
    .A(net2128));
 sg13g2_a22oi_1 _13660_ (.Y(_05737_),
    .B1(net1616),
    .B2(net1522),
    .A2(net1617),
    .A1(\am_sdr0.am0.demod_out[11] ));
 sg13g2_inv_1 _13661_ (.Y(_01172_),
    .A(net1523));
 sg13g2_a22oi_1 _13662_ (.Y(_05738_),
    .B1(net1616),
    .B2(net2168),
    .A2(net1617),
    .A1(\am_sdr0.am0.demod_out[12] ));
 sg13g2_inv_1 _13663_ (.Y(_01173_),
    .A(net2169));
 sg13g2_a22oi_1 _13664_ (.Y(_05739_),
    .B1(net1616),
    .B2(net1488),
    .A2(net1617),
    .A1(net2101));
 sg13g2_inv_1 _13665_ (.Y(_01174_),
    .A(_05739_));
 sg13g2_a22oi_1 _13666_ (.Y(_05740_),
    .B1(net1616),
    .B2(net1435),
    .A2(net1617),
    .A1(net2047));
 sg13g2_inv_1 _13667_ (.Y(_01175_),
    .A(_05740_));
 sg13g2_a22oi_1 _13668_ (.Y(_05741_),
    .B1(net1616),
    .B2(net1323),
    .A2(net1617),
    .A1(net1371));
 sg13g2_inv_1 _13669_ (.Y(_01176_),
    .A(_05741_));
 sg13g2_dfrbp_1 _13670_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net29),
    .D(net1259),
    .Q_N(_06799_),
    .Q(\am_sdr0.am0.state[0] ));
 sg13g2_dfrbp_1 _13671_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net30),
    .D(_00019_),
    .Q_N(_06800_),
    .Q(\am_sdr0.am0.state[1] ));
 sg13g2_dfrbp_1 _13672_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net31),
    .D(_00020_),
    .Q_N(_06801_),
    .Q(\am_sdr0.am0.state[2] ));
 sg13g2_dfrbp_1 _13673_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net32),
    .D(_00015_),
    .Q_N(_06802_),
    .Q(\am_sdr0.am0.state[3] ));
 sg13g2_dfrbp_1 _13674_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net33),
    .D(net1274),
    .Q_N(_06803_),
    .Q(\am_sdr0.am0.state[4] ));
 sg13g2_dfrbp_1 _13675_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net93),
    .D(_00017_),
    .Q_N(_06804_),
    .Q(\am_sdr0.am0.state[5] ));
 sg13g2_dfrbp_1 _13676_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net28),
    .D(_00021_),
    .Q_N(_06798_),
    .Q(\am_sdr0.am0.state[6] ));
 sg13g2_dfrbp_1 _13677_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net132),
    .D(_00079_),
    .Q_N(_00078_),
    .Q(\am_sdr0.am0.m_count[0] ));
 sg13g2_dfrbp_1 _13678_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net130),
    .D(net2164),
    .Q_N(_06797_),
    .Q(\am_sdr0.am0.m_count[1] ));
 sg13g2_dfrbp_1 _13679_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net128),
    .D(_00081_),
    .Q_N(_06796_),
    .Q(\am_sdr0.am0.m_count[2] ));
 sg13g2_dfrbp_1 _13680_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net126),
    .D(_00082_),
    .Q_N(_06795_),
    .Q(\am_sdr0.am0.m_count[3] ));
 sg13g2_dfrbp_1 _13681_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net124),
    .D(_00083_),
    .Q_N(_06794_),
    .Q(\am_sdr0.am0.multB[0] ));
 sg13g2_dfrbp_1 _13682_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net115),
    .D(net2049),
    .Q_N(_06793_),
    .Q(\am_sdr0.am0.multB[1] ));
 sg13g2_dfrbp_1 _13683_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net114),
    .D(net1494),
    .Q_N(_06792_),
    .Q(\am_sdr0.am0.multB[2] ));
 sg13g2_dfrbp_1 _13684_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net113),
    .D(net1521),
    .Q_N(_06791_),
    .Q(\am_sdr0.am0.multB[3] ));
 sg13g2_dfrbp_1 _13685_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net112),
    .D(net1511),
    .Q_N(_06790_),
    .Q(\am_sdr0.am0.multB[4] ));
 sg13g2_dfrbp_1 _13686_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net111),
    .D(net2038),
    .Q_N(_06789_),
    .Q(\am_sdr0.am0.multB[5] ));
 sg13g2_dfrbp_1 _13687_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net110),
    .D(net1428),
    .Q_N(_06788_),
    .Q(\am_sdr0.am0.multB[6] ));
 sg13g2_dfrbp_1 _13688_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net109),
    .D(_00090_),
    .Q_N(_06787_),
    .Q(\am_sdr0.am0.multB[7] ));
 sg13g2_dfrbp_1 _13689_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net108),
    .D(_00091_),
    .Q_N(_06786_),
    .Q(\am_sdr0.am0.multA[0] ));
 sg13g2_dfrbp_1 _13690_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net107),
    .D(net3114),
    .Q_N(_00058_),
    .Q(\am_sdr0.am0.multA[1] ));
 sg13g2_dfrbp_1 _13691_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net106),
    .D(net2926),
    .Q_N(_00060_),
    .Q(\am_sdr0.am0.multA[2] ));
 sg13g2_dfrbp_1 _13692_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net105),
    .D(net2830),
    .Q_N(_00061_),
    .Q(\am_sdr0.am0.multA[3] ));
 sg13g2_dfrbp_1 _13693_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net104),
    .D(net2910),
    .Q_N(_00063_),
    .Q(\am_sdr0.am0.multA[4] ));
 sg13g2_dfrbp_1 _13694_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net103),
    .D(net2906),
    .Q_N(_00064_),
    .Q(\am_sdr0.am0.multA[5] ));
 sg13g2_dfrbp_1 _13695_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net102),
    .D(net2832),
    .Q_N(_00065_),
    .Q(\am_sdr0.am0.multA[6] ));
 sg13g2_dfrbp_1 _13696_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net101),
    .D(net2679),
    .Q_N(_00066_),
    .Q(\am_sdr0.am0.multA[7] ));
 sg13g2_dfrbp_1 _13697_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net100),
    .D(_00099_),
    .Q_N(_00067_),
    .Q(\am_sdr0.am0.multA[8] ));
 sg13g2_dfrbp_1 _13698_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net92),
    .D(_00100_),
    .Q_N(_00068_),
    .Q(\am_sdr0.am0.multA[9] ));
 sg13g2_dfrbp_1 _13699_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net91),
    .D(_00101_),
    .Q_N(_00069_),
    .Q(\am_sdr0.am0.multA[10] ));
 sg13g2_dfrbp_1 _13700_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net90),
    .D(net2986),
    .Q_N(_06785_),
    .Q(\am_sdr0.am0.multA[11] ));
 sg13g2_dfrbp_1 _13701_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net89),
    .D(_00103_),
    .Q_N(_06784_),
    .Q(\am_sdr0.am0.multA[12] ));
 sg13g2_dfrbp_1 _13702_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net88),
    .D(_00104_),
    .Q_N(_00070_),
    .Q(\am_sdr0.am0.multA[13] ));
 sg13g2_dfrbp_1 _13703_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net87),
    .D(net2698),
    .Q_N(_00071_),
    .Q(\am_sdr0.am0.multA[14] ));
 sg13g2_dfrbp_1 _13704_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net86),
    .D(_00106_),
    .Q_N(_00072_),
    .Q(\am_sdr0.am0.multA[15] ));
 sg13g2_dfrbp_1 _13705_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net85),
    .D(_00107_),
    .Q_N(_06783_),
    .Q(\am_sdr0.am0.multA[16] ));
 sg13g2_dfrbp_1 _13706_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net84),
    .D(net1432),
    .Q_N(_06782_),
    .Q(\am_sdr0.am0.sum[0] ));
 sg13g2_dfrbp_1 _13707_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net82),
    .D(_00109_),
    .Q_N(_06781_),
    .Q(\am_sdr0.am0.sum[1] ));
 sg13g2_dfrbp_1 _13708_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net80),
    .D(net2278),
    .Q_N(_00059_),
    .Q(\am_sdr0.am0.sum[2] ));
 sg13g2_dfrbp_1 _13709_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net78),
    .D(_00111_),
    .Q_N(_06780_),
    .Q(\am_sdr0.am0.sum[3] ));
 sg13g2_dfrbp_1 _13710_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net76),
    .D(_00112_),
    .Q_N(_00062_),
    .Q(\am_sdr0.am0.sum[4] ));
 sg13g2_dfrbp_1 _13711_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net74),
    .D(_00113_),
    .Q_N(_06779_),
    .Q(\am_sdr0.am0.sum[5] ));
 sg13g2_dfrbp_1 _13712_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net72),
    .D(_00114_),
    .Q_N(_06778_),
    .Q(\am_sdr0.am0.sum[6] ));
 sg13g2_dfrbp_1 _13713_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net70),
    .D(_00115_),
    .Q_N(_06777_),
    .Q(\am_sdr0.am0.sum[7] ));
 sg13g2_dfrbp_1 _13714_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net68),
    .D(net2248),
    .Q_N(_06776_),
    .Q(\am_sdr0.am0.sum[8] ));
 sg13g2_dfrbp_1 _13715_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net66),
    .D(_00117_),
    .Q_N(_06775_),
    .Q(\am_sdr0.am0.sum[9] ));
 sg13g2_dfrbp_1 _13716_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net64),
    .D(_00118_),
    .Q_N(_06774_),
    .Q(\am_sdr0.am0.sum[10] ));
 sg13g2_dfrbp_1 _13717_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net62),
    .D(net2471),
    .Q_N(_06773_),
    .Q(\am_sdr0.am0.sum[11] ));
 sg13g2_dfrbp_1 _13718_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net60),
    .D(_00120_),
    .Q_N(_06772_),
    .Q(\am_sdr0.am0.sum[12] ));
 sg13g2_dfrbp_1 _13719_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net58),
    .D(_00121_),
    .Q_N(_06771_),
    .Q(\am_sdr0.am0.sum[13] ));
 sg13g2_dfrbp_1 _13720_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net56),
    .D(_00122_),
    .Q_N(_06770_),
    .Q(\am_sdr0.am0.sum[14] ));
 sg13g2_dfrbp_1 _13721_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net54),
    .D(_00123_),
    .Q_N(_06769_),
    .Q(\am_sdr0.am0.sum[15] ));
 sg13g2_dfrbp_1 _13722_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net52),
    .D(_00124_),
    .Q_N(_06768_),
    .Q(\am_sdr0.am0.sum[16] ));
 sg13g2_dfrbp_1 _13723_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net50),
    .D(net1171),
    .Q_N(_00077_),
    .Q(\am_sdr0.am0.count2[0] ));
 sg13g2_dfrbp_1 _13724_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net48),
    .D(net3006),
    .Q_N(_06767_),
    .Q(\am_sdr0.am0.count2[1] ));
 sg13g2_dfrbp_1 _13725_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net46),
    .D(net1255),
    .Q_N(_06766_),
    .Q(\am_sdr0.am0.count2[2] ));
 sg13g2_dfrbp_1 _13726_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net44),
    .D(net2098),
    .Q_N(_06765_),
    .Q(\am_sdr0.am0.count2[3] ));
 sg13g2_dfrbp_1 _13727_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net42),
    .D(_00129_),
    .Q_N(_06764_),
    .Q(\am_sdr0.am0.r[0] ));
 sg13g2_dfrbp_1 _13728_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net40),
    .D(_00130_),
    .Q_N(_06763_),
    .Q(\am_sdr0.am0.r[1] ));
 sg13g2_dfrbp_1 _13729_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net38),
    .D(_00131_),
    .Q_N(_06762_),
    .Q(\am_sdr0.am0.r[2] ));
 sg13g2_dfrbp_1 _13730_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net36),
    .D(_00132_),
    .Q_N(_06761_),
    .Q(\am_sdr0.am0.r[3] ));
 sg13g2_dfrbp_1 _13731_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net34),
    .D(_00133_),
    .Q_N(_06760_),
    .Q(\am_sdr0.am0.r[4] ));
 sg13g2_dfrbp_1 _13732_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1162),
    .D(_00134_),
    .Q_N(_06759_),
    .Q(\am_sdr0.am0.r[5] ));
 sg13g2_dfrbp_1 _13733_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1160),
    .D(_00135_),
    .Q_N(_06758_),
    .Q(\am_sdr0.am0.r[6] ));
 sg13g2_dfrbp_1 _13734_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1158),
    .D(_00136_),
    .Q_N(_06757_),
    .Q(\am_sdr0.am0.r[7] ));
 sg13g2_dfrbp_1 _13735_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net94),
    .D(_00137_),
    .Q_N(_00022_),
    .Q(\am_sdr0.am0.r[9] ));
 sg13g2_dfrbp_1 _13736_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net95),
    .D(_00008_),
    .Q_N(_06805_),
    .Q(\am_sdr0.mix0.sin_in[0] ));
 sg13g2_dfrbp_1 _13737_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net96),
    .D(_00009_),
    .Q_N(_06806_),
    .Q(\am_sdr0.mix0.sin_in[1] ));
 sg13g2_dfrbp_1 _13738_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net97),
    .D(_00010_),
    .Q_N(_06807_),
    .Q(\am_sdr0.mix0.sin_in[2] ));
 sg13g2_dfrbp_1 _13739_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net98),
    .D(_00011_),
    .Q_N(_06808_),
    .Q(\am_sdr0.mix0.sin_in[3] ));
 sg13g2_dfrbp_1 _13740_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net99),
    .D(_00012_),
    .Q_N(_06809_),
    .Q(\am_sdr0.mix0.sin_in[4] ));
 sg13g2_dfrbp_1 _13741_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net116),
    .D(_00013_),
    .Q_N(_06810_),
    .Q(\am_sdr0.mix0.sin_in[5] ));
 sg13g2_dfrbp_1 _13742_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1156),
    .D(_00014_),
    .Q_N(_06756_),
    .Q(\am_sdr0.mix0.sin_in[6] ));
 sg13g2_dfrbp_1 _13743_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1154),
    .D(_00138_),
    .Q_N(_06755_),
    .Q(\am_sdr0.am0.a[0] ));
 sg13g2_dfrbp_1 _13744_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1152),
    .D(_00139_),
    .Q_N(_06754_),
    .Q(\am_sdr0.am0.a[1] ));
 sg13g2_dfrbp_1 _13745_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1150),
    .D(net1387),
    .Q_N(_06753_),
    .Q(\am_sdr0.am0.a[2] ));
 sg13g2_dfrbp_1 _13746_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1149),
    .D(net1459),
    .Q_N(_06752_),
    .Q(\am_sdr0.am0.a[3] ));
 sg13g2_dfrbp_1 _13747_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1148),
    .D(net2028),
    .Q_N(_06751_),
    .Q(\am_sdr0.am0.a[4] ));
 sg13g2_dfrbp_1 _13748_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1147),
    .D(net1457),
    .Q_N(_06750_),
    .Q(\am_sdr0.am0.a[5] ));
 sg13g2_dfrbp_1 _13749_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1146),
    .D(net1509),
    .Q_N(_06749_),
    .Q(\am_sdr0.am0.a[6] ));
 sg13g2_dfrbp_1 _13750_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1145),
    .D(net1492),
    .Q_N(_06748_),
    .Q(\am_sdr0.am0.a[7] ));
 sg13g2_dfrbp_1 _13751_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1144),
    .D(net1414),
    .Q_N(_06747_),
    .Q(\am_sdr0.am0.a[8] ));
 sg13g2_dfrbp_1 _13752_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1143),
    .D(net1449),
    .Q_N(_06746_),
    .Q(\am_sdr0.am0.a[9] ));
 sg13g2_dfrbp_1 _13753_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1142),
    .D(net1318),
    .Q_N(_06745_),
    .Q(\am_sdr0.am0.a[10] ));
 sg13g2_dfrbp_1 _13754_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1141),
    .D(_00149_),
    .Q_N(_06744_),
    .Q(\am_sdr0.am0.a[11] ));
 sg13g2_dfrbp_1 _13755_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1140),
    .D(net1359),
    .Q_N(_06743_),
    .Q(\am_sdr0.am0.a[12] ));
 sg13g2_dfrbp_1 _13756_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1139),
    .D(_00151_),
    .Q_N(_06742_),
    .Q(\am_sdr0.am0.a[13] ));
 sg13g2_dfrbp_1 _13757_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1138),
    .D(_00152_),
    .Q_N(_06741_),
    .Q(\am_sdr0.am0.a[14] ));
 sg13g2_dfrbp_1 _13758_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net117),
    .D(_00153_),
    .Q_N(_06811_),
    .Q(\am_sdr0.am0.a[15] ));
 sg13g2_dfrbp_1 _13759_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net118),
    .D(_00000_),
    .Q_N(_06812_),
    .Q(\am_sdr0.cos[0] ));
 sg13g2_dfrbp_1 _13760_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net119),
    .D(_00001_),
    .Q_N(_06813_),
    .Q(\am_sdr0.cos[1] ));
 sg13g2_dfrbp_1 _13761_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net120),
    .D(_00002_),
    .Q_N(_06814_),
    .Q(\am_sdr0.cos[2] ));
 sg13g2_dfrbp_1 _13762_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net121),
    .D(net2410),
    .Q_N(_06815_),
    .Q(\am_sdr0.cos[3] ));
 sg13g2_dfrbp_1 _13763_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net122),
    .D(_00004_),
    .Q_N(_06816_),
    .Q(\am_sdr0.cos[4] ));
 sg13g2_dfrbp_1 _13764_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net123),
    .D(_00005_),
    .Q_N(_06817_),
    .Q(\am_sdr0.cos[5] ));
 sg13g2_dfrbp_1 _13765_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1033),
    .D(_00006_),
    .Q_N(_06818_),
    .Q(\am_sdr0.cos[6] ));
 sg13g2_dfrbp_1 _13766_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1137),
    .D(net1527),
    .Q_N(_06740_),
    .Q(\am_sdr0.cos[7] ));
 sg13g2_dfrbp_1 _13767_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1136),
    .D(_00154_),
    .Q_N(_06739_),
    .Q(\am_sdr0.mix0.sin_in[7] ));
 sg13g2_dfrbp_1 _13768_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1135),
    .D(_00155_),
    .Q_N(_06738_),
    .Q(\am_sdr0.spi0.MOSI_qq ));
 sg13g2_dfrbp_1 _13769_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1134),
    .D(_00156_),
    .Q_N(_00076_),
    .Q(\am_sdr0.count[0] ));
 sg13g2_dfrbp_1 _13770_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1133),
    .D(net2434),
    .Q_N(_06737_),
    .Q(\am_sdr0.count[1] ));
 sg13g2_dfrbp_1 _13771_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1132),
    .D(net2528),
    .Q_N(_06736_),
    .Q(\am_sdr0.count[2] ));
 sg13g2_dfrbp_1 _13772_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1131),
    .D(_00159_),
    .Q_N(_06735_),
    .Q(\am_sdr0.count[3] ));
 sg13g2_dfrbp_1 _13773_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1130),
    .D(_00160_),
    .Q_N(_06734_),
    .Q(\am_sdr0.count[4] ));
 sg13g2_dfrbp_1 _13774_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1129),
    .D(_00161_),
    .Q_N(_06733_),
    .Q(\am_sdr0.count[5] ));
 sg13g2_dfrbp_1 _13775_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1128),
    .D(_00162_),
    .Q_N(_06732_),
    .Q(\am_sdr0.count[6] ));
 sg13g2_dfrbp_1 _13776_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1127),
    .D(_00163_),
    .Q_N(_06731_),
    .Q(\am_sdr0.count[7] ));
 sg13g2_dfrbp_1 _13777_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1126),
    .D(net1173),
    .Q_N(_06730_),
    .Q(\am_sdr0.am0.q[0] ));
 sg13g2_dfrbp_1 _13778_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1124),
    .D(_00165_),
    .Q_N(_06729_),
    .Q(\am_sdr0.am0.q[1] ));
 sg13g2_dfrbp_1 _13779_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1122),
    .D(_00166_),
    .Q_N(_06728_),
    .Q(\am_sdr0.am0.q[2] ));
 sg13g2_dfrbp_1 _13780_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1120),
    .D(_00167_),
    .Q_N(_06727_),
    .Q(\am_sdr0.am0.q[3] ));
 sg13g2_dfrbp_1 _13781_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1118),
    .D(_00168_),
    .Q_N(_06726_),
    .Q(\am_sdr0.am0.q[4] ));
 sg13g2_dfrbp_1 _13782_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1116),
    .D(_00169_),
    .Q_N(_06725_),
    .Q(\am_sdr0.am0.q[5] ));
 sg13g2_dfrbp_1 _13783_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1114),
    .D(_00170_),
    .Q_N(_06724_),
    .Q(\am_sdr0.am0.q[6] ));
 sg13g2_dfrbp_1 _13784_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1112),
    .D(_00171_),
    .Q_N(_06723_),
    .Q(\am_sdr0.am0.q[7] ));
 sg13g2_dfrbp_1 _13785_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1110),
    .D(net2456),
    .Q_N(_06722_),
    .Q(\am_sdr0.am0.sqrt_state[0] ));
 sg13g2_dfrbp_1 _13786_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1108),
    .D(_00173_),
    .Q_N(_06721_),
    .Q(\am_sdr0.am0.sqrt_state[1] ));
 sg13g2_dfrbp_1 _13787_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1106),
    .D(net1473),
    .Q_N(_06720_),
    .Q(\am_sdr0.am0.sqrt_done ));
 sg13g2_dfrbp_1 _13788_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1105),
    .D(_00175_),
    .Q_N(_06719_),
    .Q(\am_sdr0.am0.left[0] ));
 sg13g2_dfrbp_1 _13789_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1103),
    .D(_00176_),
    .Q_N(_06718_),
    .Q(\am_sdr0.am0.left[1] ));
 sg13g2_dfrbp_1 _13790_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1101),
    .D(_00177_),
    .Q_N(_06717_),
    .Q(\am_sdr0.am0.left[2] ));
 sg13g2_dfrbp_1 _13791_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1099),
    .D(_00178_),
    .Q_N(_06716_),
    .Q(\am_sdr0.am0.left[3] ));
 sg13g2_dfrbp_1 _13792_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1097),
    .D(_00179_),
    .Q_N(_06715_),
    .Q(\am_sdr0.am0.left[4] ));
 sg13g2_dfrbp_1 _13793_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1095),
    .D(_00180_),
    .Q_N(_00051_),
    .Q(\am_sdr0.am0.left[5] ));
 sg13g2_dfrbp_1 _13794_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1093),
    .D(_00181_),
    .Q_N(_06714_),
    .Q(\am_sdr0.am0.left[6] ));
 sg13g2_dfrbp_1 _13795_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1091),
    .D(_00182_),
    .Q_N(_06713_),
    .Q(\am_sdr0.am0.left[7] ));
 sg13g2_dfrbp_1 _13796_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1089),
    .D(_00183_),
    .Q_N(_00056_),
    .Q(\am_sdr0.am0.left[8] ));
 sg13g2_dfrbp_1 _13797_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1087),
    .D(_00184_),
    .Q_N(_06712_),
    .Q(\am_sdr0.am0.left[9] ));
 sg13g2_dfrbp_1 _13798_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1085),
    .D(_00185_),
    .Q_N(_06711_),
    .Q(\am_sdr0.am0.right[0] ));
 sg13g2_dfrbp_1 _13799_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1083),
    .D(_00186_),
    .Q_N(_00047_),
    .Q(\am_sdr0.am0.right[1] ));
 sg13g2_dfrbp_1 _13800_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1081),
    .D(_00187_),
    .Q_N(_00048_),
    .Q(\am_sdr0.am0.right[2] ));
 sg13g2_dfrbp_1 _13801_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1079),
    .D(_00188_),
    .Q_N(_00049_),
    .Q(\am_sdr0.am0.right[3] ));
 sg13g2_dfrbp_1 _13802_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1077),
    .D(_00189_),
    .Q_N(_00050_),
    .Q(\am_sdr0.am0.right[4] ));
 sg13g2_dfrbp_1 _13803_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1075),
    .D(_00190_),
    .Q_N(_00052_),
    .Q(\am_sdr0.am0.right[5] ));
 sg13g2_dfrbp_1 _13804_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1073),
    .D(_00191_),
    .Q_N(_00053_),
    .Q(\am_sdr0.am0.right[6] ));
 sg13g2_dfrbp_1 _13805_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1071),
    .D(_00192_),
    .Q_N(_00054_),
    .Q(\am_sdr0.am0.right[7] ));
 sg13g2_dfrbp_1 _13806_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1069),
    .D(_00193_),
    .Q_N(_00057_),
    .Q(\am_sdr0.am0.right[8] ));
 sg13g2_dfrbp_1 _13807_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1067),
    .D(_00194_),
    .Q_N(_00055_),
    .Q(\am_sdr0.am0.right[9] ));
 sg13g2_dfrbp_1 _13808_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1065),
    .D(_00195_),
    .Q_N(_06710_),
    .Q(\am_sdr0.cic3.sample ));
 sg13g2_dfrbp_1 _13809_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1064),
    .D(_00196_),
    .Q_N(_06709_),
    .Q(\am_sdr0.cic2.integ_sample[0] ));
 sg13g2_dfrbp_1 _13810_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1063),
    .D(_00197_),
    .Q_N(_06708_),
    .Q(\am_sdr0.cic2.integ_sample[1] ));
 sg13g2_dfrbp_1 _13811_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1062),
    .D(_00198_),
    .Q_N(_06707_),
    .Q(\am_sdr0.cic2.integ_sample[2] ));
 sg13g2_dfrbp_1 _13812_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1061),
    .D(net2138),
    .Q_N(_06706_),
    .Q(\am_sdr0.cic2.integ_sample[3] ));
 sg13g2_dfrbp_1 _13813_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1060),
    .D(net2448),
    .Q_N(_06705_),
    .Q(\am_sdr0.cic2.integ_sample[4] ));
 sg13g2_dfrbp_1 _13814_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1059),
    .D(net2812),
    .Q_N(_06704_),
    .Q(\am_sdr0.cic2.integ_sample[5] ));
 sg13g2_dfrbp_1 _13815_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1058),
    .D(_00202_),
    .Q_N(_06703_),
    .Q(\am_sdr0.cic2.integ_sample[6] ));
 sg13g2_dfrbp_1 _13816_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1057),
    .D(_00203_),
    .Q_N(_06702_),
    .Q(\am_sdr0.cic2.integ_sample[7] ));
 sg13g2_dfrbp_1 _13817_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1056),
    .D(_00204_),
    .Q_N(_06701_),
    .Q(\am_sdr0.cic2.integ_sample[8] ));
 sg13g2_dfrbp_1 _13818_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1055),
    .D(_00205_),
    .Q_N(_06700_),
    .Q(\am_sdr0.cic2.integ_sample[9] ));
 sg13g2_dfrbp_1 _13819_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1054),
    .D(_00206_),
    .Q_N(_06699_),
    .Q(\am_sdr0.cic2.integ_sample[10] ));
 sg13g2_dfrbp_1 _13820_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1053),
    .D(_00207_),
    .Q_N(_06698_),
    .Q(\am_sdr0.cic2.integ_sample[11] ));
 sg13g2_dfrbp_1 _13821_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1052),
    .D(net2357),
    .Q_N(_06697_),
    .Q(\am_sdr0.cic2.integ_sample[12] ));
 sg13g2_dfrbp_1 _13822_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1051),
    .D(net2850),
    .Q_N(_06696_),
    .Q(\am_sdr0.cic2.integ_sample[13] ));
 sg13g2_dfrbp_1 _13823_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1050),
    .D(net1385),
    .Q_N(_06695_),
    .Q(\am_sdr0.cic2.integ_sample[14] ));
 sg13g2_dfrbp_1 _13824_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1049),
    .D(net2227),
    .Q_N(_06694_),
    .Q(\am_sdr0.cic2.integ_sample[15] ));
 sg13g2_dfrbp_1 _13825_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1032),
    .D(net2297),
    .Q_N(_06693_),
    .Q(\am_sdr0.cic2.integ_sample[16] ));
 sg13g2_dfrbp_1 _13826_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1031),
    .D(net2235),
    .Q_N(_06692_),
    .Q(\am_sdr0.cic2.integ_sample[17] ));
 sg13g2_dfrbp_1 _13827_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1030),
    .D(net2343),
    .Q_N(_06691_),
    .Q(\am_sdr0.cic2.integ_sample[18] ));
 sg13g2_dfrbp_1 _13828_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1029),
    .D(_00215_),
    .Q_N(_06690_),
    .Q(\am_sdr0.cic2.integ_sample[19] ));
 sg13g2_dfrbp_1 _13829_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1028),
    .D(net1517),
    .Q_N(_06689_),
    .Q(\am_sdr0.am0.Q_in[0] ));
 sg13g2_dfrbp_1 _13830_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1026),
    .D(net2150),
    .Q_N(_06688_),
    .Q(\am_sdr0.am0.Q_in[1] ));
 sg13g2_dfrbp_1 _13831_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1024),
    .D(net1453),
    .Q_N(_06687_),
    .Q(\am_sdr0.am0.Q_in[2] ));
 sg13g2_dfrbp_1 _13832_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1022),
    .D(net1463),
    .Q_N(_06686_),
    .Q(\am_sdr0.am0.Q_in[3] ));
 sg13g2_dfrbp_1 _13833_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1020),
    .D(net1320),
    .Q_N(_06685_),
    .Q(\am_sdr0.am0.Q_in[4] ));
 sg13g2_dfrbp_1 _13834_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1018),
    .D(net1350),
    .Q_N(_06684_),
    .Q(\am_sdr0.am0.Q_in[5] ));
 sg13g2_dfrbp_1 _13835_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1016),
    .D(net1356),
    .Q_N(_06683_),
    .Q(\am_sdr0.am0.Q_in[6] ));
 sg13g2_dfrbp_1 _13836_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1014),
    .D(net1333),
    .Q_N(_06682_),
    .Q(\am_sdr0.am0.Q_in[7] ));
 sg13g2_dfrbp_1 _13837_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1012),
    .D(_00224_),
    .Q_N(_06681_),
    .Q(\am_sdr0.cic3.comb1[0] ));
 sg13g2_dfrbp_1 _13838_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1010),
    .D(_00225_),
    .Q_N(_06680_),
    .Q(\am_sdr0.cic3.comb1[1] ));
 sg13g2_dfrbp_1 _13839_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1008),
    .D(_00226_),
    .Q_N(_06679_),
    .Q(\am_sdr0.cic3.comb1[2] ));
 sg13g2_dfrbp_1 _13840_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1006),
    .D(_00227_),
    .Q_N(_06678_),
    .Q(\am_sdr0.cic3.comb1[3] ));
 sg13g2_dfrbp_1 _13841_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1004),
    .D(_00228_),
    .Q_N(_06677_),
    .Q(\am_sdr0.cic3.comb1[4] ));
 sg13g2_dfrbp_1 _13842_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1002),
    .D(net2893),
    .Q_N(_06676_),
    .Q(\am_sdr0.cic3.comb1[5] ));
 sg13g2_dfrbp_1 _13843_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1000),
    .D(_00230_),
    .Q_N(_06675_),
    .Q(\am_sdr0.cic3.comb1[6] ));
 sg13g2_dfrbp_1 _13844_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net998),
    .D(_00231_),
    .Q_N(_06674_),
    .Q(\am_sdr0.cic3.comb1[7] ));
 sg13g2_dfrbp_1 _13845_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net996),
    .D(_00232_),
    .Q_N(_06673_),
    .Q(\am_sdr0.cic3.comb1[8] ));
 sg13g2_dfrbp_1 _13846_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net994),
    .D(_00233_),
    .Q_N(_06672_),
    .Q(\am_sdr0.cic3.comb1[9] ));
 sg13g2_dfrbp_1 _13847_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net992),
    .D(_00234_),
    .Q_N(_06671_),
    .Q(\am_sdr0.cic3.comb1[10] ));
 sg13g2_dfrbp_1 _13848_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net990),
    .D(_00235_),
    .Q_N(_06670_),
    .Q(\am_sdr0.cic3.comb1[11] ));
 sg13g2_dfrbp_1 _13849_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net988),
    .D(_00236_),
    .Q_N(_06669_),
    .Q(\am_sdr0.cic3.comb1[12] ));
 sg13g2_dfrbp_1 _13850_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net986),
    .D(_00237_),
    .Q_N(_06668_),
    .Q(\am_sdr0.cic3.comb1[13] ));
 sg13g2_dfrbp_1 _13851_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net984),
    .D(_00238_),
    .Q_N(_06667_),
    .Q(\am_sdr0.cic3.comb1[14] ));
 sg13g2_dfrbp_1 _13852_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net982),
    .D(_00239_),
    .Q_N(_06666_),
    .Q(\am_sdr0.cic3.comb1[15] ));
 sg13g2_dfrbp_1 _13853_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net980),
    .D(_00240_),
    .Q_N(_06665_),
    .Q(\am_sdr0.cic3.comb1[16] ));
 sg13g2_dfrbp_1 _13854_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net978),
    .D(net2737),
    .Q_N(_06664_),
    .Q(\am_sdr0.cic3.comb1[17] ));
 sg13g2_dfrbp_1 _13855_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net976),
    .D(_00242_),
    .Q_N(_06663_),
    .Q(\am_sdr0.cic3.comb1[18] ));
 sg13g2_dfrbp_1 _13856_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net974),
    .D(_00243_),
    .Q_N(_06662_),
    .Q(\am_sdr0.cic3.comb1[19] ));
 sg13g2_dfrbp_1 _13857_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net972),
    .D(_00244_),
    .Q_N(_06661_),
    .Q(\am_sdr0.cic3.comb1_in_del[0] ));
 sg13g2_dfrbp_1 _13858_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net970),
    .D(net2373),
    .Q_N(_06660_),
    .Q(\am_sdr0.cic3.comb1_in_del[1] ));
 sg13g2_dfrbp_1 _13859_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net968),
    .D(_00246_),
    .Q_N(_06659_),
    .Q(\am_sdr0.cic3.comb1_in_del[2] ));
 sg13g2_dfrbp_1 _13860_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net966),
    .D(_00247_),
    .Q_N(_06658_),
    .Q(\am_sdr0.cic3.comb1_in_del[3] ));
 sg13g2_dfrbp_1 _13861_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net964),
    .D(_00248_),
    .Q_N(_06657_),
    .Q(\am_sdr0.cic3.comb1_in_del[4] ));
 sg13g2_dfrbp_1 _13862_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net962),
    .D(_00249_),
    .Q_N(_06656_),
    .Q(\am_sdr0.cic3.comb1_in_del[5] ));
 sg13g2_dfrbp_1 _13863_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net960),
    .D(_00250_),
    .Q_N(_06655_),
    .Q(\am_sdr0.cic3.comb1_in_del[6] ));
 sg13g2_dfrbp_1 _13864_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net958),
    .D(_00251_),
    .Q_N(_06654_),
    .Q(\am_sdr0.cic3.comb1_in_del[7] ));
 sg13g2_dfrbp_1 _13865_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net956),
    .D(_00252_),
    .Q_N(_06653_),
    .Q(\am_sdr0.cic3.comb1_in_del[8] ));
 sg13g2_dfrbp_1 _13866_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net954),
    .D(_00253_),
    .Q_N(_06652_),
    .Q(\am_sdr0.cic3.comb1_in_del[9] ));
 sg13g2_dfrbp_1 _13867_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net952),
    .D(_00254_),
    .Q_N(_06651_),
    .Q(\am_sdr0.cic3.comb1_in_del[10] ));
 sg13g2_dfrbp_1 _13868_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net950),
    .D(_00255_),
    .Q_N(_06650_),
    .Q(\am_sdr0.cic3.comb1_in_del[11] ));
 sg13g2_dfrbp_1 _13869_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net948),
    .D(_00256_),
    .Q_N(_06649_),
    .Q(\am_sdr0.cic3.comb1_in_del[12] ));
 sg13g2_dfrbp_1 _13870_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net946),
    .D(net2940),
    .Q_N(_06648_),
    .Q(\am_sdr0.cic3.comb1_in_del[13] ));
 sg13g2_dfrbp_1 _13871_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net944),
    .D(net2681),
    .Q_N(_06647_),
    .Q(\am_sdr0.cic3.comb1_in_del[14] ));
 sg13g2_dfrbp_1 _13872_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net942),
    .D(net2814),
    .Q_N(_06646_),
    .Q(\am_sdr0.cic3.comb1_in_del[15] ));
 sg13g2_dfrbp_1 _13873_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net940),
    .D(net2622),
    .Q_N(_06645_),
    .Q(\am_sdr0.cic3.comb1_in_del[16] ));
 sg13g2_dfrbp_1 _13874_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net938),
    .D(net2888),
    .Q_N(_06644_),
    .Q(\am_sdr0.cic3.comb1_in_del[17] ));
 sg13g2_dfrbp_1 _13875_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net936),
    .D(net2477),
    .Q_N(_06643_),
    .Q(\am_sdr0.cic3.comb1_in_del[18] ));
 sg13g2_dfrbp_1 _13876_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net934),
    .D(_00263_),
    .Q_N(_06642_),
    .Q(\am_sdr0.cic3.comb1_in_del[19] ));
 sg13g2_dfrbp_1 _13877_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net932),
    .D(_00264_),
    .Q_N(_06641_),
    .Q(\am_sdr0.cic3.comb2[0] ));
 sg13g2_dfrbp_1 _13878_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net930),
    .D(_00265_),
    .Q_N(_06640_),
    .Q(\am_sdr0.cic3.comb2[1] ));
 sg13g2_dfrbp_1 _13879_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net928),
    .D(net2860),
    .Q_N(_06639_),
    .Q(\am_sdr0.cic3.comb2[2] ));
 sg13g2_dfrbp_1 _13880_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net926),
    .D(_00267_),
    .Q_N(_06638_),
    .Q(\am_sdr0.cic3.comb2[3] ));
 sg13g2_dfrbp_1 _13881_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net924),
    .D(_00268_),
    .Q_N(_06637_),
    .Q(\am_sdr0.cic3.comb2[4] ));
 sg13g2_dfrbp_1 _13882_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net922),
    .D(_00269_),
    .Q_N(_06636_),
    .Q(\am_sdr0.cic3.comb2[5] ));
 sg13g2_dfrbp_1 _13883_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net920),
    .D(net2771),
    .Q_N(_06635_),
    .Q(\am_sdr0.cic3.comb2[6] ));
 sg13g2_dfrbp_1 _13884_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net918),
    .D(_00271_),
    .Q_N(_06634_),
    .Q(\am_sdr0.cic3.comb2[7] ));
 sg13g2_dfrbp_1 _13885_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net916),
    .D(_00272_),
    .Q_N(_06633_),
    .Q(\am_sdr0.cic3.comb2[8] ));
 sg13g2_dfrbp_1 _13886_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net914),
    .D(net2651),
    .Q_N(_06632_),
    .Q(\am_sdr0.cic3.comb2[9] ));
 sg13g2_dfrbp_1 _13887_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net912),
    .D(_00274_),
    .Q_N(_06631_),
    .Q(\am_sdr0.cic3.comb2[10] ));
 sg13g2_dfrbp_1 _13888_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net910),
    .D(_00275_),
    .Q_N(_06630_),
    .Q(\am_sdr0.cic3.comb2[11] ));
 sg13g2_dfrbp_1 _13889_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net908),
    .D(_00276_),
    .Q_N(_06629_),
    .Q(\am_sdr0.cic3.comb2[12] ));
 sg13g2_dfrbp_1 _13890_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net906),
    .D(_00277_),
    .Q_N(_06628_),
    .Q(\am_sdr0.cic3.comb2[13] ));
 sg13g2_dfrbp_1 _13891_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net904),
    .D(_00278_),
    .Q_N(_06627_),
    .Q(\am_sdr0.cic3.comb2[14] ));
 sg13g2_dfrbp_1 _13892_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net902),
    .D(net2886),
    .Q_N(_06626_),
    .Q(\am_sdr0.cic3.comb2[15] ));
 sg13g2_dfrbp_1 _13893_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net900),
    .D(_00280_),
    .Q_N(_06625_),
    .Q(\am_sdr0.cic3.comb2[16] ));
 sg13g2_dfrbp_1 _13894_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net898),
    .D(_00281_),
    .Q_N(_06624_),
    .Q(\am_sdr0.cic3.comb2[17] ));
 sg13g2_dfrbp_1 _13895_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net896),
    .D(_00282_),
    .Q_N(_06623_),
    .Q(\am_sdr0.cic3.comb2[18] ));
 sg13g2_dfrbp_1 _13896_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net894),
    .D(_00283_),
    .Q_N(_06622_),
    .Q(\am_sdr0.cic3.comb2[19] ));
 sg13g2_dfrbp_1 _13897_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net892),
    .D(net2261),
    .Q_N(_06621_),
    .Q(\am_sdr0.cic3.comb2_in_del[0] ));
 sg13g2_dfrbp_1 _13898_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net890),
    .D(net2348),
    .Q_N(_06620_),
    .Q(\am_sdr0.cic3.comb2_in_del[1] ));
 sg13g2_dfrbp_1 _13899_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net888),
    .D(net2239),
    .Q_N(_06619_),
    .Q(\am_sdr0.cic3.comb2_in_del[2] ));
 sg13g2_dfrbp_1 _13900_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net886),
    .D(net2534),
    .Q_N(_06618_),
    .Q(\am_sdr0.cic3.comb2_in_del[3] ));
 sg13g2_dfrbp_1 _13901_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net884),
    .D(_00288_),
    .Q_N(_06617_),
    .Q(\am_sdr0.cic3.comb2_in_del[4] ));
 sg13g2_dfrbp_1 _13902_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net882),
    .D(_00289_),
    .Q_N(_06616_),
    .Q(\am_sdr0.cic3.comb2_in_del[5] ));
 sg13g2_dfrbp_1 _13903_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net880),
    .D(net2720),
    .Q_N(_06615_),
    .Q(\am_sdr0.cic3.comb2_in_del[6] ));
 sg13g2_dfrbp_1 _13904_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net878),
    .D(net2576),
    .Q_N(_06614_),
    .Q(\am_sdr0.cic3.comb2_in_del[7] ));
 sg13g2_dfrbp_1 _13905_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net876),
    .D(net2666),
    .Q_N(_06613_),
    .Q(\am_sdr0.cic3.comb2_in_del[8] ));
 sg13g2_dfrbp_1 _13906_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net874),
    .D(net2777),
    .Q_N(_06612_),
    .Q(\am_sdr0.cic3.comb2_in_del[9] ));
 sg13g2_dfrbp_1 _13907_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net872),
    .D(net2380),
    .Q_N(_06611_),
    .Q(\am_sdr0.cic3.comb2_in_del[10] ));
 sg13g2_dfrbp_1 _13908_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net870),
    .D(net2237),
    .Q_N(_06610_),
    .Q(\am_sdr0.cic3.comb2_in_del[11] ));
 sg13g2_dfrbp_1 _13909_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net868),
    .D(_00296_),
    .Q_N(_06609_),
    .Q(\am_sdr0.cic3.comb2_in_del[12] ));
 sg13g2_dfrbp_1 _13910_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net866),
    .D(net2541),
    .Q_N(_06608_),
    .Q(\am_sdr0.cic3.comb2_in_del[13] ));
 sg13g2_dfrbp_1 _13911_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net864),
    .D(net2322),
    .Q_N(_06607_),
    .Q(\am_sdr0.cic3.comb2_in_del[14] ));
 sg13g2_dfrbp_1 _13912_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net862),
    .D(net2759),
    .Q_N(_06606_),
    .Q(\am_sdr0.cic3.comb2_in_del[15] ));
 sg13g2_dfrbp_1 _13913_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net860),
    .D(net2366),
    .Q_N(_06605_),
    .Q(\am_sdr0.cic3.comb2_in_del[16] ));
 sg13g2_dfrbp_1 _13914_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net858),
    .D(_00301_),
    .Q_N(_06604_),
    .Q(\am_sdr0.cic3.comb2_in_del[17] ));
 sg13g2_dfrbp_1 _13915_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net856),
    .D(net2364),
    .Q_N(_06603_),
    .Q(\am_sdr0.cic3.comb2_in_del[18] ));
 sg13g2_dfrbp_1 _13916_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net854),
    .D(net2436),
    .Q_N(_06602_),
    .Q(\am_sdr0.cic3.comb2_in_del[19] ));
 sg13g2_dfrbp_1 _13917_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net852),
    .D(_00304_),
    .Q_N(_06601_),
    .Q(\am_sdr0.cic3.comb3[12] ));
 sg13g2_dfrbp_1 _13918_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net850),
    .D(_00305_),
    .Q_N(_06600_),
    .Q(\am_sdr0.cic3.comb3[13] ));
 sg13g2_dfrbp_1 _13919_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net848),
    .D(_00306_),
    .Q_N(_06599_),
    .Q(\am_sdr0.cic3.comb3[14] ));
 sg13g2_dfrbp_1 _13920_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net846),
    .D(_00307_),
    .Q_N(_06598_),
    .Q(\am_sdr0.cic3.comb3[15] ));
 sg13g2_dfrbp_1 _13921_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net844),
    .D(_00308_),
    .Q_N(_06597_),
    .Q(\am_sdr0.cic3.comb3[16] ));
 sg13g2_dfrbp_1 _13922_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net842),
    .D(_00309_),
    .Q_N(_06596_),
    .Q(\am_sdr0.cic3.comb3[17] ));
 sg13g2_dfrbp_1 _13923_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net840),
    .D(_00310_),
    .Q_N(_06595_),
    .Q(\am_sdr0.cic3.comb3[18] ));
 sg13g2_dfrbp_1 _13924_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net838),
    .D(_00311_),
    .Q_N(_06594_),
    .Q(\am_sdr0.cic3.comb3[19] ));
 sg13g2_dfrbp_1 _13925_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net836),
    .D(net1529),
    .Q_N(_06593_),
    .Q(\am_sdr0.cic3.comb3_in_del[0] ));
 sg13g2_dfrbp_1 _13926_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net834),
    .D(net2046),
    .Q_N(_06592_),
    .Q(\am_sdr0.cic3.comb3_in_del[1] ));
 sg13g2_dfrbp_1 _13927_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net832),
    .D(net2090),
    .Q_N(_06591_),
    .Q(\am_sdr0.cic3.comb3_in_del[2] ));
 sg13g2_dfrbp_1 _13928_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net830),
    .D(_00315_),
    .Q_N(_06590_),
    .Q(\am_sdr0.cic3.comb3_in_del[3] ));
 sg13g2_dfrbp_1 _13929_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net828),
    .D(net2229),
    .Q_N(_06589_),
    .Q(\am_sdr0.cic3.comb3_in_del[4] ));
 sg13g2_dfrbp_1 _13930_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net826),
    .D(net2233),
    .Q_N(_06588_),
    .Q(\am_sdr0.cic3.comb3_in_del[5] ));
 sg13g2_dfrbp_1 _13931_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net824),
    .D(net2200),
    .Q_N(_06587_),
    .Q(\am_sdr0.cic3.comb3_in_del[6] ));
 sg13g2_dfrbp_1 _13932_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net822),
    .D(net2156),
    .Q_N(_06586_),
    .Q(\am_sdr0.cic3.comb3_in_del[7] ));
 sg13g2_dfrbp_1 _13933_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net820),
    .D(net2211),
    .Q_N(_06585_),
    .Q(\am_sdr0.cic3.comb3_in_del[8] ));
 sg13g2_dfrbp_1 _13934_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net818),
    .D(net2182),
    .Q_N(_06584_),
    .Q(\am_sdr0.cic3.comb3_in_del[9] ));
 sg13g2_dfrbp_1 _13935_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net816),
    .D(net2295),
    .Q_N(_06583_),
    .Q(\am_sdr0.cic3.comb3_in_del[10] ));
 sg13g2_dfrbp_1 _13936_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net814),
    .D(net2214),
    .Q_N(_06582_),
    .Q(\am_sdr0.cic3.comb3_in_del[11] ));
 sg13g2_dfrbp_1 _13937_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net812),
    .D(net2271),
    .Q_N(_06581_),
    .Q(\am_sdr0.cic3.comb3_in_del[12] ));
 sg13g2_dfrbp_1 _13938_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net810),
    .D(_00325_),
    .Q_N(_06580_),
    .Q(\am_sdr0.cic3.comb3_in_del[13] ));
 sg13g2_dfrbp_1 _13939_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net808),
    .D(_00326_),
    .Q_N(_06579_),
    .Q(\am_sdr0.cic3.comb3_in_del[14] ));
 sg13g2_dfrbp_1 _13940_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net806),
    .D(net2286),
    .Q_N(_06578_),
    .Q(\am_sdr0.cic3.comb3_in_del[15] ));
 sg13g2_dfrbp_1 _13941_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net804),
    .D(net2491),
    .Q_N(_06577_),
    .Q(\am_sdr0.cic3.comb3_in_del[16] ));
 sg13g2_dfrbp_1 _13942_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net802),
    .D(net2204),
    .Q_N(_06576_),
    .Q(\am_sdr0.cic3.comb3_in_del[17] ));
 sg13g2_dfrbp_1 _13943_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net800),
    .D(_00330_),
    .Q_N(_06575_),
    .Q(\am_sdr0.cic3.comb3_in_del[18] ));
 sg13g2_dfrbp_1 _13944_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net798),
    .D(net2192),
    .Q_N(_06574_),
    .Q(\am_sdr0.cic3.comb3_in_del[19] ));
 sg13g2_dfrbp_1 _13945_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net796),
    .D(_00332_),
    .Q_N(_06573_),
    .Q(\am_sdr0.cic3.count[0] ));
 sg13g2_dfrbp_1 _13946_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net794),
    .D(net1245),
    .Q_N(_06572_),
    .Q(\am_sdr0.cic3.count[1] ));
 sg13g2_dfrbp_1 _13947_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net792),
    .D(_00334_),
    .Q_N(_06571_),
    .Q(\am_sdr0.cic3.count[2] ));
 sg13g2_dfrbp_1 _13948_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net790),
    .D(_00335_),
    .Q_N(_06570_),
    .Q(\am_sdr0.cic3.count[3] ));
 sg13g2_dfrbp_1 _13949_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net788),
    .D(_00336_),
    .Q_N(_06569_),
    .Q(\am_sdr0.cic3.count[4] ));
 sg13g2_dfrbp_1 _13950_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net786),
    .D(_00337_),
    .Q_N(_06568_),
    .Q(\am_sdr0.cic3.count[5] ));
 sg13g2_dfrbp_1 _13951_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net784),
    .D(net2096),
    .Q_N(_06567_),
    .Q(\am_sdr0.cic3.count[6] ));
 sg13g2_dfrbp_1 _13952_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net782),
    .D(net1376),
    .Q_N(_06566_),
    .Q(\am_sdr0.cic3.count[7] ));
 sg13g2_dfrbp_1 _13953_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net780),
    .D(net1279),
    .Q_N(_06565_),
    .Q(\am_sdr0.cic3.integ1[0] ));
 sg13g2_dfrbp_1 _13954_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net778),
    .D(net2806),
    .Q_N(_06564_),
    .Q(\am_sdr0.cic3.integ1[1] ));
 sg13g2_dfrbp_1 _13955_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net776),
    .D(_00342_),
    .Q_N(_06563_),
    .Q(\am_sdr0.cic3.integ1[2] ));
 sg13g2_dfrbp_1 _13956_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net774),
    .D(net3036),
    .Q_N(_06562_),
    .Q(\am_sdr0.cic3.integ1[3] ));
 sg13g2_dfrbp_1 _13957_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net772),
    .D(_00344_),
    .Q_N(_06561_),
    .Q(\am_sdr0.cic3.integ1[4] ));
 sg13g2_dfrbp_1 _13958_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net770),
    .D(_00345_),
    .Q_N(_06560_),
    .Q(\am_sdr0.cic3.integ1[5] ));
 sg13g2_dfrbp_1 _13959_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net768),
    .D(_00346_),
    .Q_N(_06559_),
    .Q(\am_sdr0.cic3.integ1[6] ));
 sg13g2_dfrbp_1 _13960_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net766),
    .D(net3112),
    .Q_N(_06558_),
    .Q(\am_sdr0.cic3.integ1[7] ));
 sg13g2_dfrbp_1 _13961_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net764),
    .D(_00348_),
    .Q_N(_06557_),
    .Q(\am_sdr0.cic3.integ1[8] ));
 sg13g2_dfrbp_1 _13962_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net762),
    .D(_00349_),
    .Q_N(_06556_),
    .Q(\am_sdr0.cic3.integ1[9] ));
 sg13g2_dfrbp_1 _13963_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net760),
    .D(_00350_),
    .Q_N(_06555_),
    .Q(\am_sdr0.cic3.integ1[10] ));
 sg13g2_dfrbp_1 _13964_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net758),
    .D(_00351_),
    .Q_N(_06554_),
    .Q(\am_sdr0.cic3.integ1[11] ));
 sg13g2_dfrbp_1 _13965_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net756),
    .D(_00352_),
    .Q_N(_06553_),
    .Q(\am_sdr0.cic3.integ1[12] ));
 sg13g2_dfrbp_1 _13966_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net754),
    .D(_00353_),
    .Q_N(_06552_),
    .Q(\am_sdr0.cic3.integ1[13] ));
 sg13g2_dfrbp_1 _13967_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net752),
    .D(_00354_),
    .Q_N(_06551_),
    .Q(\am_sdr0.cic3.integ1[14] ));
 sg13g2_dfrbp_1 _13968_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net750),
    .D(_00355_),
    .Q_N(_06550_),
    .Q(\am_sdr0.cic3.integ1[15] ));
 sg13g2_dfrbp_1 _13969_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net748),
    .D(_00356_),
    .Q_N(_06549_),
    .Q(\am_sdr0.cic3.integ1[16] ));
 sg13g2_dfrbp_1 _13970_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net746),
    .D(_00357_),
    .Q_N(_06548_),
    .Q(\am_sdr0.cic3.integ1[17] ));
 sg13g2_dfrbp_1 _13971_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net744),
    .D(_00358_),
    .Q_N(_06547_),
    .Q(\am_sdr0.cic3.integ1[18] ));
 sg13g2_dfrbp_1 _13972_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net742),
    .D(_00359_),
    .Q_N(_06546_),
    .Q(\am_sdr0.cic3.integ1[19] ));
 sg13g2_dfrbp_1 _13973_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net740),
    .D(_00360_),
    .Q_N(_06545_),
    .Q(\am_sdr0.cic3.integ1[20] ));
 sg13g2_dfrbp_1 _13974_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net738),
    .D(_00361_),
    .Q_N(_06544_),
    .Q(\am_sdr0.cic3.integ1[21] ));
 sg13g2_dfrbp_1 _13975_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net736),
    .D(_00362_),
    .Q_N(_06543_),
    .Q(\am_sdr0.cic3.integ1[22] ));
 sg13g2_dfrbp_1 _13976_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net734),
    .D(_00363_),
    .Q_N(_06542_),
    .Q(\am_sdr0.cic3.integ1[23] ));
 sg13g2_dfrbp_1 _13977_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net732),
    .D(_00364_),
    .Q_N(_06541_),
    .Q(\am_sdr0.cic3.integ1[24] ));
 sg13g2_dfrbp_1 _13978_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net730),
    .D(_00365_),
    .Q_N(_06540_),
    .Q(\am_sdr0.cic3.integ1[25] ));
 sg13g2_dfrbp_1 _13979_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net728),
    .D(_00366_),
    .Q_N(_06539_),
    .Q(\am_sdr0.cic3.integ2[0] ));
 sg13g2_dfrbp_1 _13980_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net726),
    .D(_00367_),
    .Q_N(_06538_),
    .Q(\am_sdr0.cic3.integ2[1] ));
 sg13g2_dfrbp_1 _13981_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net724),
    .D(net2653),
    .Q_N(_06537_),
    .Q(\am_sdr0.cic3.integ2[2] ));
 sg13g2_dfrbp_1 _13982_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net722),
    .D(_00369_),
    .Q_N(_06536_),
    .Q(\am_sdr0.cic3.integ2[3] ));
 sg13g2_dfrbp_1 _13983_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net720),
    .D(_00370_),
    .Q_N(_06535_),
    .Q(\am_sdr0.cic3.integ2[4] ));
 sg13g2_dfrbp_1 _13984_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net718),
    .D(_00371_),
    .Q_N(_06534_),
    .Q(\am_sdr0.cic3.integ2[5] ));
 sg13g2_dfrbp_1 _13985_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net716),
    .D(_00372_),
    .Q_N(_06533_),
    .Q(\am_sdr0.cic3.integ2[6] ));
 sg13g2_dfrbp_1 _13986_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net714),
    .D(_00373_),
    .Q_N(_06532_),
    .Q(\am_sdr0.cic3.integ2[7] ));
 sg13g2_dfrbp_1 _13987_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net712),
    .D(_00374_),
    .Q_N(_06531_),
    .Q(\am_sdr0.cic3.integ2[8] ));
 sg13g2_dfrbp_1 _13988_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net710),
    .D(_00375_),
    .Q_N(_06530_),
    .Q(\am_sdr0.cic3.integ2[9] ));
 sg13g2_dfrbp_1 _13989_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net708),
    .D(_00376_),
    .Q_N(_06529_),
    .Q(\am_sdr0.cic3.integ2[10] ));
 sg13g2_dfrbp_1 _13990_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net706),
    .D(_00377_),
    .Q_N(_06528_),
    .Q(\am_sdr0.cic3.integ2[11] ));
 sg13g2_dfrbp_1 _13991_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net704),
    .D(_00378_),
    .Q_N(_06527_),
    .Q(\am_sdr0.cic3.integ2[12] ));
 sg13g2_dfrbp_1 _13992_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net702),
    .D(_00379_),
    .Q_N(_06526_),
    .Q(\am_sdr0.cic3.integ2[13] ));
 sg13g2_dfrbp_1 _13993_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net700),
    .D(_00380_),
    .Q_N(_06525_),
    .Q(\am_sdr0.cic3.integ2[14] ));
 sg13g2_dfrbp_1 _13994_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net698),
    .D(_00381_),
    .Q_N(_06524_),
    .Q(\am_sdr0.cic3.integ2[15] ));
 sg13g2_dfrbp_1 _13995_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net696),
    .D(_00382_),
    .Q_N(_06523_),
    .Q(\am_sdr0.cic3.integ2[16] ));
 sg13g2_dfrbp_1 _13996_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net694),
    .D(_00383_),
    .Q_N(_06522_),
    .Q(\am_sdr0.cic3.integ2[17] ));
 sg13g2_dfrbp_1 _13997_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net692),
    .D(_00384_),
    .Q_N(_06521_),
    .Q(\am_sdr0.cic3.integ2[18] ));
 sg13g2_dfrbp_1 _13998_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net690),
    .D(_00385_),
    .Q_N(_06520_),
    .Q(\am_sdr0.cic3.integ2[19] ));
 sg13g2_dfrbp_1 _13999_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net688),
    .D(_00386_),
    .Q_N(_06519_),
    .Q(\am_sdr0.cic3.integ2[20] ));
 sg13g2_dfrbp_1 _14000_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net686),
    .D(_00387_),
    .Q_N(_06518_),
    .Q(\am_sdr0.cic3.integ2[21] ));
 sg13g2_dfrbp_1 _14001_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net684),
    .D(_00388_),
    .Q_N(_06517_),
    .Q(\am_sdr0.cic3.integ2[22] ));
 sg13g2_dfrbp_1 _14002_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net682),
    .D(_00389_),
    .Q_N(_06516_),
    .Q(\am_sdr0.cic3.integ3[0] ));
 sg13g2_dfrbp_1 _14003_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net680),
    .D(_00390_),
    .Q_N(_06515_),
    .Q(\am_sdr0.cic3.integ3[1] ));
 sg13g2_dfrbp_1 _14004_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net678),
    .D(net2975),
    .Q_N(_06514_),
    .Q(\am_sdr0.cic3.integ3[2] ));
 sg13g2_dfrbp_1 _14005_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net676),
    .D(_00392_),
    .Q_N(_06513_),
    .Q(\am_sdr0.cic3.integ3[3] ));
 sg13g2_dfrbp_1 _14006_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net674),
    .D(_00393_),
    .Q_N(_06512_),
    .Q(\am_sdr0.cic3.integ3[4] ));
 sg13g2_dfrbp_1 _14007_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net672),
    .D(_00394_),
    .Q_N(_06511_),
    .Q(\am_sdr0.cic3.integ3[5] ));
 sg13g2_dfrbp_1 _14008_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net670),
    .D(_00395_),
    .Q_N(_06510_),
    .Q(\am_sdr0.cic3.integ3[6] ));
 sg13g2_dfrbp_1 _14009_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net668),
    .D(_00396_),
    .Q_N(_06509_),
    .Q(\am_sdr0.cic3.integ3[7] ));
 sg13g2_dfrbp_1 _14010_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net666),
    .D(_00397_),
    .Q_N(_06508_),
    .Q(\am_sdr0.cic3.integ3[8] ));
 sg13g2_dfrbp_1 _14011_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net664),
    .D(_00398_),
    .Q_N(_06507_),
    .Q(\am_sdr0.cic3.integ3[9] ));
 sg13g2_dfrbp_1 _14012_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net662),
    .D(_00399_),
    .Q_N(_06506_),
    .Q(\am_sdr0.cic3.integ3[10] ));
 sg13g2_dfrbp_1 _14013_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net660),
    .D(net2960),
    .Q_N(_06505_),
    .Q(\am_sdr0.cic3.integ3[11] ));
 sg13g2_dfrbp_1 _14014_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net658),
    .D(_00401_),
    .Q_N(_06504_),
    .Q(\am_sdr0.cic3.integ3[12] ));
 sg13g2_dfrbp_1 _14015_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net656),
    .D(_00402_),
    .Q_N(_06503_),
    .Q(\am_sdr0.cic3.integ3[13] ));
 sg13g2_dfrbp_1 _14016_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net654),
    .D(_00403_),
    .Q_N(_06502_),
    .Q(\am_sdr0.cic3.integ3[14] ));
 sg13g2_dfrbp_1 _14017_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net652),
    .D(_00404_),
    .Q_N(_06501_),
    .Q(\am_sdr0.cic3.integ3[15] ));
 sg13g2_dfrbp_1 _14018_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net650),
    .D(_00405_),
    .Q_N(_06500_),
    .Q(\am_sdr0.cic3.integ3[16] ));
 sg13g2_dfrbp_1 _14019_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net648),
    .D(_00406_),
    .Q_N(_06499_),
    .Q(\am_sdr0.cic3.integ3[17] ));
 sg13g2_dfrbp_1 _14020_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net646),
    .D(_00407_),
    .Q_N(_06498_),
    .Q(\am_sdr0.cic3.integ3[18] ));
 sg13g2_dfrbp_1 _14021_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net644),
    .D(net2875),
    .Q_N(_06497_),
    .Q(\am_sdr0.cic3.integ3[19] ));
 sg13g2_dfrbp_1 _14022_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net642),
    .D(net1539),
    .Q_N(_06496_),
    .Q(\am_sdr0.cic2.sample ));
 sg13g2_dfrbp_1 _14023_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net641),
    .D(_00410_),
    .Q_N(_06495_),
    .Q(\am_sdr0.am0.load_tick ));
 sg13g2_dfrbp_1 _14024_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net640),
    .D(net2408),
    .Q_N(_06494_),
    .Q(\am_sdr0.cic1.integ_sample[0] ));
 sg13g2_dfrbp_1 _14025_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net639),
    .D(net1390),
    .Q_N(_06493_),
    .Q(\am_sdr0.cic1.integ_sample[1] ));
 sg13g2_dfrbp_1 _14026_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net638),
    .D(net2082),
    .Q_N(_06492_),
    .Q(\am_sdr0.cic1.integ_sample[2] ));
 sg13g2_dfrbp_1 _14027_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net637),
    .D(net2071),
    .Q_N(_06491_),
    .Q(\am_sdr0.cic1.integ_sample[3] ));
 sg13g2_dfrbp_1 _14028_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net636),
    .D(net2160),
    .Q_N(_06490_),
    .Q(\am_sdr0.cic1.integ_sample[4] ));
 sg13g2_dfrbp_1 _14029_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net635),
    .D(net2086),
    .Q_N(_06489_),
    .Q(\am_sdr0.cic1.integ_sample[5] ));
 sg13g2_dfrbp_1 _14030_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net634),
    .D(net1335),
    .Q_N(_06488_),
    .Q(\am_sdr0.cic1.integ_sample[6] ));
 sg13g2_dfrbp_1 _14031_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net633),
    .D(net1442),
    .Q_N(_06487_),
    .Q(\am_sdr0.cic1.integ_sample[7] ));
 sg13g2_dfrbp_1 _14032_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net632),
    .D(net1477),
    .Q_N(_06486_),
    .Q(\am_sdr0.cic1.integ_sample[8] ));
 sg13g2_dfrbp_1 _14033_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net631),
    .D(net1424),
    .Q_N(_06485_),
    .Q(\am_sdr0.cic1.integ_sample[9] ));
 sg13g2_dfrbp_1 _14034_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net630),
    .D(net1498),
    .Q_N(_06484_),
    .Q(\am_sdr0.cic1.integ_sample[10] ));
 sg13g2_dfrbp_1 _14035_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net629),
    .D(net2115),
    .Q_N(_06483_),
    .Q(\am_sdr0.cic1.integ_sample[11] ));
 sg13g2_dfrbp_1 _14036_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net628),
    .D(net2646),
    .Q_N(_06482_),
    .Q(\am_sdr0.cic1.integ_sample[12] ));
 sg13g2_dfrbp_1 _14037_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net627),
    .D(net1399),
    .Q_N(_06481_),
    .Q(\am_sdr0.cic1.integ_sample[13] ));
 sg13g2_dfrbp_1 _14038_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net626),
    .D(net2355),
    .Q_N(_06480_),
    .Q(\am_sdr0.cic1.integ_sample[14] ));
 sg13g2_dfrbp_1 _14039_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net625),
    .D(net2177),
    .Q_N(_06479_),
    .Q(\am_sdr0.cic1.integ_sample[15] ));
 sg13g2_dfrbp_1 _14040_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net624),
    .D(net2158),
    .Q_N(_06478_),
    .Q(\am_sdr0.cic1.integ_sample[16] ));
 sg13g2_dfrbp_1 _14041_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net623),
    .D(net2352),
    .Q_N(_06477_),
    .Q(\am_sdr0.cic1.integ_sample[17] ));
 sg13g2_dfrbp_1 _14042_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net622),
    .D(net1407),
    .Q_N(_06476_),
    .Q(\am_sdr0.cic1.integ_sample[18] ));
 sg13g2_dfrbp_1 _14043_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net621),
    .D(net1380),
    .Q_N(_06475_),
    .Q(\am_sdr0.cic1.integ_sample[19] ));
 sg13g2_dfrbp_1 _14044_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net620),
    .D(net1232),
    .Q_N(_06474_),
    .Q(\am_sdr0.am0.I_in[0] ));
 sg13g2_dfrbp_1 _14045_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net618),
    .D(net1370),
    .Q_N(_06473_),
    .Q(\am_sdr0.am0.I_in[1] ));
 sg13g2_dfrbp_1 _14046_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net616),
    .D(net1296),
    .Q_N(_06472_),
    .Q(\am_sdr0.am0.I_in[2] ));
 sg13g2_dfrbp_1 _14047_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net614),
    .D(net1451),
    .Q_N(_06471_),
    .Q(\am_sdr0.am0.I_in[3] ));
 sg13g2_dfrbp_1 _14048_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net612),
    .D(net1263),
    .Q_N(_06470_),
    .Q(\am_sdr0.am0.I_in[4] ));
 sg13g2_dfrbp_1 _14049_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net610),
    .D(net1286),
    .Q_N(_06469_),
    .Q(\am_sdr0.am0.I_in[5] ));
 sg13g2_dfrbp_1 _14050_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net608),
    .D(net1247),
    .Q_N(_06468_),
    .Q(\am_sdr0.am0.I_in[6] ));
 sg13g2_dfrbp_1 _14051_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net606),
    .D(net1288),
    .Q_N(_06467_),
    .Q(\am_sdr0.am0.I_in[7] ));
 sg13g2_dfrbp_1 _14052_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net604),
    .D(_00439_),
    .Q_N(_06466_),
    .Q(\am_sdr0.cic2.comb1[0] ));
 sg13g2_dfrbp_1 _14053_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net602),
    .D(_00440_),
    .Q_N(_06465_),
    .Q(\am_sdr0.cic2.comb1[1] ));
 sg13g2_dfrbp_1 _14054_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net600),
    .D(_00441_),
    .Q_N(_06464_),
    .Q(\am_sdr0.cic2.comb1[2] ));
 sg13g2_dfrbp_1 _14055_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net598),
    .D(_00442_),
    .Q_N(_06463_),
    .Q(\am_sdr0.cic2.comb1[3] ));
 sg13g2_dfrbp_1 _14056_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net596),
    .D(_00443_),
    .Q_N(_06462_),
    .Q(\am_sdr0.cic2.comb1[4] ));
 sg13g2_dfrbp_1 _14057_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net594),
    .D(_00444_),
    .Q_N(_06461_),
    .Q(\am_sdr0.cic2.comb1[5] ));
 sg13g2_dfrbp_1 _14058_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net592),
    .D(_00445_),
    .Q_N(_06460_),
    .Q(\am_sdr0.cic2.comb1[6] ));
 sg13g2_dfrbp_1 _14059_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net590),
    .D(_00446_),
    .Q_N(_06459_),
    .Q(\am_sdr0.cic2.comb1[7] ));
 sg13g2_dfrbp_1 _14060_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net588),
    .D(_00447_),
    .Q_N(_06458_),
    .Q(\am_sdr0.cic2.comb1[8] ));
 sg13g2_dfrbp_1 _14061_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net586),
    .D(_00448_),
    .Q_N(_06457_),
    .Q(\am_sdr0.cic2.comb1[9] ));
 sg13g2_dfrbp_1 _14062_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net584),
    .D(_00449_),
    .Q_N(_06456_),
    .Q(\am_sdr0.cic2.comb1[10] ));
 sg13g2_dfrbp_1 _14063_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net582),
    .D(_00450_),
    .Q_N(_06455_),
    .Q(\am_sdr0.cic2.comb1[11] ));
 sg13g2_dfrbp_1 _14064_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net580),
    .D(_00451_),
    .Q_N(_06454_),
    .Q(\am_sdr0.cic2.comb1[12] ));
 sg13g2_dfrbp_1 _14065_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net578),
    .D(_00452_),
    .Q_N(_06453_),
    .Q(\am_sdr0.cic2.comb1[13] ));
 sg13g2_dfrbp_1 _14066_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net576),
    .D(_00453_),
    .Q_N(_06452_),
    .Q(\am_sdr0.cic2.comb1[14] ));
 sg13g2_dfrbp_1 _14067_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net574),
    .D(_00454_),
    .Q_N(_06451_),
    .Q(\am_sdr0.cic2.comb1[15] ));
 sg13g2_dfrbp_1 _14068_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net572),
    .D(_00455_),
    .Q_N(_06450_),
    .Q(\am_sdr0.cic2.comb1[16] ));
 sg13g2_dfrbp_1 _14069_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net570),
    .D(net2660),
    .Q_N(_06449_),
    .Q(\am_sdr0.cic2.comb1[17] ));
 sg13g2_dfrbp_1 _14070_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net568),
    .D(_00457_),
    .Q_N(_06448_),
    .Q(\am_sdr0.cic2.comb1[18] ));
 sg13g2_dfrbp_1 _14071_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net566),
    .D(_00458_),
    .Q_N(_06447_),
    .Q(\am_sdr0.cic2.comb1[19] ));
 sg13g2_dfrbp_1 _14072_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net564),
    .D(net2069),
    .Q_N(_06446_),
    .Q(\am_sdr0.cic2.comb1_in_del[0] ));
 sg13g2_dfrbp_1 _14073_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net562),
    .D(net2454),
    .Q_N(_06445_),
    .Q(\am_sdr0.cic2.comb1_in_del[1] ));
 sg13g2_dfrbp_1 _14074_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net560),
    .D(net2600),
    .Q_N(_06444_),
    .Q(\am_sdr0.cic2.comb1_in_del[2] ));
 sg13g2_dfrbp_1 _14075_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net558),
    .D(_00462_),
    .Q_N(_06443_),
    .Q(\am_sdr0.cic2.comb1_in_del[3] ));
 sg13g2_dfrbp_1 _14076_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net556),
    .D(net2565),
    .Q_N(_06442_),
    .Q(\am_sdr0.cic2.comb1_in_del[4] ));
 sg13g2_dfrbp_1 _14077_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net554),
    .D(net2655),
    .Q_N(_06441_),
    .Q(\am_sdr0.cic2.comb1_in_del[5] ));
 sg13g2_dfrbp_1 _14078_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net552),
    .D(net2375),
    .Q_N(_06440_),
    .Q(\am_sdr0.cic2.comb1_in_del[6] ));
 sg13g2_dfrbp_1 _14079_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net550),
    .D(net2397),
    .Q_N(_06439_),
    .Q(\am_sdr0.cic2.comb1_in_del[7] ));
 sg13g2_dfrbp_1 _14080_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net548),
    .D(net2152),
    .Q_N(_06438_),
    .Q(\am_sdr0.cic2.comb1_in_del[8] ));
 sg13g2_dfrbp_1 _14081_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net546),
    .D(net2362),
    .Q_N(_06437_),
    .Q(\am_sdr0.cic2.comb1_in_del[9] ));
 sg13g2_dfrbp_1 _14082_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net544),
    .D(net2078),
    .Q_N(_06436_),
    .Q(\am_sdr0.cic2.comb1_in_del[10] ));
 sg13g2_dfrbp_1 _14083_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net542),
    .D(net2067),
    .Q_N(_06435_),
    .Q(\am_sdr0.cic2.comb1_in_del[11] ));
 sg13g2_dfrbp_1 _14084_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net540),
    .D(_00471_),
    .Q_N(_06434_),
    .Q(\am_sdr0.cic2.comb1_in_del[12] ));
 sg13g2_dfrbp_1 _14085_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net538),
    .D(net2617),
    .Q_N(_06433_),
    .Q(\am_sdr0.cic2.comb1_in_del[13] ));
 sg13g2_dfrbp_1 _14086_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net536),
    .D(_00473_),
    .Q_N(_06432_),
    .Q(\am_sdr0.cic2.comb1_in_del[14] ));
 sg13g2_dfrbp_1 _14087_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net534),
    .D(_00474_),
    .Q_N(_06431_),
    .Q(\am_sdr0.cic2.comb1_in_del[15] ));
 sg13g2_dfrbp_1 _14088_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net532),
    .D(_00475_),
    .Q_N(_06430_),
    .Q(\am_sdr0.cic2.comb1_in_del[16] ));
 sg13g2_dfrbp_1 _14089_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net530),
    .D(_00476_),
    .Q_N(_06429_),
    .Q(\am_sdr0.cic2.comb1_in_del[17] ));
 sg13g2_dfrbp_1 _14090_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net528),
    .D(_00477_),
    .Q_N(_06428_),
    .Q(\am_sdr0.cic2.comb1_in_del[18] ));
 sg13g2_dfrbp_1 _14091_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net526),
    .D(net1487),
    .Q_N(_06427_),
    .Q(\am_sdr0.cic2.comb1_in_del[19] ));
 sg13g2_dfrbp_1 _14092_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net524),
    .D(net2385),
    .Q_N(_06426_),
    .Q(\am_sdr0.cic2.comb2[0] ));
 sg13g2_dfrbp_1 _14093_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net522),
    .D(_00480_),
    .Q_N(_06425_),
    .Q(\am_sdr0.cic2.comb2[1] ));
 sg13g2_dfrbp_1 _14094_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net520),
    .D(net2872),
    .Q_N(_06424_),
    .Q(\am_sdr0.cic2.comb2[2] ));
 sg13g2_dfrbp_1 _14095_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net518),
    .D(_00482_),
    .Q_N(_06423_),
    .Q(\am_sdr0.cic2.comb2[3] ));
 sg13g2_dfrbp_1 _14096_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net516),
    .D(_00483_),
    .Q_N(_06422_),
    .Q(\am_sdr0.cic2.comb2[4] ));
 sg13g2_dfrbp_1 _14097_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net514),
    .D(_00484_),
    .Q_N(_06421_),
    .Q(\am_sdr0.cic2.comb2[5] ));
 sg13g2_dfrbp_1 _14098_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net512),
    .D(_00485_),
    .Q_N(_06420_),
    .Q(\am_sdr0.cic2.comb2[6] ));
 sg13g2_dfrbp_1 _14099_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net510),
    .D(net2786),
    .Q_N(_06419_),
    .Q(\am_sdr0.cic2.comb2[7] ));
 sg13g2_dfrbp_1 _14100_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net508),
    .D(_00487_),
    .Q_N(_06418_),
    .Q(\am_sdr0.cic2.comb2[8] ));
 sg13g2_dfrbp_1 _14101_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net506),
    .D(_00488_),
    .Q_N(_06417_),
    .Q(\am_sdr0.cic2.comb2[9] ));
 sg13g2_dfrbp_1 _14102_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net504),
    .D(_00489_),
    .Q_N(_06416_),
    .Q(\am_sdr0.cic2.comb2[10] ));
 sg13g2_dfrbp_1 _14103_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net502),
    .D(_00490_),
    .Q_N(_06415_),
    .Q(\am_sdr0.cic2.comb2[11] ));
 sg13g2_dfrbp_1 _14104_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net500),
    .D(_00491_),
    .Q_N(_06414_),
    .Q(\am_sdr0.cic2.comb2[12] ));
 sg13g2_dfrbp_1 _14105_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net498),
    .D(_00492_),
    .Q_N(_06413_),
    .Q(\am_sdr0.cic2.comb2[13] ));
 sg13g2_dfrbp_1 _14106_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net496),
    .D(_00493_),
    .Q_N(_06412_),
    .Q(\am_sdr0.cic2.comb2[14] ));
 sg13g2_dfrbp_1 _14107_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net494),
    .D(_00494_),
    .Q_N(_06411_),
    .Q(\am_sdr0.cic2.comb2[15] ));
 sg13g2_dfrbp_1 _14108_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net492),
    .D(_00495_),
    .Q_N(_06410_),
    .Q(\am_sdr0.cic2.comb2[16] ));
 sg13g2_dfrbp_1 _14109_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net490),
    .D(_00496_),
    .Q_N(_06409_),
    .Q(\am_sdr0.cic2.comb2[17] ));
 sg13g2_dfrbp_1 _14110_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net488),
    .D(_00497_),
    .Q_N(_06408_),
    .Q(\am_sdr0.cic2.comb2[18] ));
 sg13g2_dfrbp_1 _14111_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net486),
    .D(_00498_),
    .Q_N(_06407_),
    .Q(\am_sdr0.cic2.comb2[19] ));
 sg13g2_dfrbp_1 _14112_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net484),
    .D(_00499_),
    .Q_N(_06406_),
    .Q(\am_sdr0.cic2.comb2_in_del[0] ));
 sg13g2_dfrbp_1 _14113_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net482),
    .D(net2313),
    .Q_N(_06405_),
    .Q(\am_sdr0.cic2.comb2_in_del[1] ));
 sg13g2_dfrbp_1 _14114_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net480),
    .D(net2421),
    .Q_N(_06404_),
    .Q(\am_sdr0.cic2.comb2_in_del[2] ));
 sg13g2_dfrbp_1 _14115_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net478),
    .D(net2516),
    .Q_N(_06403_),
    .Q(\am_sdr0.cic2.comb2_in_del[3] ));
 sg13g2_dfrbp_1 _14116_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net476),
    .D(net2223),
    .Q_N(_06402_),
    .Q(\am_sdr0.cic2.comb2_in_del[4] ));
 sg13g2_dfrbp_1 _14117_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net474),
    .D(net2387),
    .Q_N(_06401_),
    .Q(\am_sdr0.cic2.comb2_in_del[5] ));
 sg13g2_dfrbp_1 _14118_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net472),
    .D(net2395),
    .Q_N(_06400_),
    .Q(\am_sdr0.cic2.comb2_in_del[6] ));
 sg13g2_dfrbp_1 _14119_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net470),
    .D(net2521),
    .Q_N(_06399_),
    .Q(\am_sdr0.cic2.comb2_in_del[7] ));
 sg13g2_dfrbp_1 _14120_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net468),
    .D(_00507_),
    .Q_N(_06398_),
    .Q(\am_sdr0.cic2.comb2_in_del[8] ));
 sg13g2_dfrbp_1 _14121_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net466),
    .D(net2282),
    .Q_N(_06397_),
    .Q(\am_sdr0.cic2.comb2_in_del[9] ));
 sg13g2_dfrbp_1 _14122_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net464),
    .D(net2497),
    .Q_N(_06396_),
    .Q(\am_sdr0.cic2.comb2_in_del[10] ));
 sg13g2_dfrbp_1 _14123_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net462),
    .D(net2252),
    .Q_N(_06395_),
    .Q(\am_sdr0.cic2.comb2_in_del[11] ));
 sg13g2_dfrbp_1 _14124_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net460),
    .D(_00511_),
    .Q_N(_06394_),
    .Q(\am_sdr0.cic2.comb2_in_del[12] ));
 sg13g2_dfrbp_1 _14125_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net458),
    .D(_00512_),
    .Q_N(_06393_),
    .Q(\am_sdr0.cic2.comb2_in_del[13] ));
 sg13g2_dfrbp_1 _14126_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net456),
    .D(net2568),
    .Q_N(_06392_),
    .Q(\am_sdr0.cic2.comb2_in_del[14] ));
 sg13g2_dfrbp_1 _14127_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net454),
    .D(net2856),
    .Q_N(_06391_),
    .Q(\am_sdr0.cic2.comb2_in_del[15] ));
 sg13g2_dfrbp_1 _14128_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net452),
    .D(net2632),
    .Q_N(_06390_),
    .Q(\am_sdr0.cic2.comb2_in_del[16] ));
 sg13g2_dfrbp_1 _14129_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net450),
    .D(_00516_),
    .Q_N(_06389_),
    .Q(\am_sdr0.cic2.comb2_in_del[17] ));
 sg13g2_dfrbp_1 _14130_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net448),
    .D(net2246),
    .Q_N(_06388_),
    .Q(\am_sdr0.cic2.comb2_in_del[18] ));
 sg13g2_dfrbp_1 _14131_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net446),
    .D(net2316),
    .Q_N(_06387_),
    .Q(\am_sdr0.cic2.comb2_in_del[19] ));
 sg13g2_dfrbp_1 _14132_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net444),
    .D(_00519_),
    .Q_N(_06386_),
    .Q(\am_sdr0.cic2.comb3[12] ));
 sg13g2_dfrbp_1 _14133_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net442),
    .D(_00520_),
    .Q_N(_06385_),
    .Q(\am_sdr0.cic2.comb3[13] ));
 sg13g2_dfrbp_1 _14134_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net440),
    .D(_00521_),
    .Q_N(_06384_),
    .Q(\am_sdr0.cic2.comb3[14] ));
 sg13g2_dfrbp_1 _14135_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net438),
    .D(_00522_),
    .Q_N(_06383_),
    .Q(\am_sdr0.cic2.comb3[15] ));
 sg13g2_dfrbp_1 _14136_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net436),
    .D(_00523_),
    .Q_N(_06382_),
    .Q(\am_sdr0.cic2.comb3[16] ));
 sg13g2_dfrbp_1 _14137_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net434),
    .D(net2042),
    .Q_N(_06381_),
    .Q(\am_sdr0.cic2.comb3[17] ));
 sg13g2_dfrbp_1 _14138_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net432),
    .D(_00525_),
    .Q_N(_06380_),
    .Q(\am_sdr0.cic2.comb3[18] ));
 sg13g2_dfrbp_1 _14139_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net430),
    .D(net2060),
    .Q_N(_06379_),
    .Q(\am_sdr0.cic2.comb3[19] ));
 sg13g2_dfrbp_1 _14140_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net428),
    .D(net1467),
    .Q_N(_06378_),
    .Q(\am_sdr0.cic2.comb3_in_del[0] ));
 sg13g2_dfrbp_1 _14141_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net426),
    .D(net2084),
    .Q_N(_06377_),
    .Q(\am_sdr0.cic2.comb3_in_del[1] ));
 sg13g2_dfrbp_1 _14142_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net424),
    .D(net2112),
    .Q_N(_06376_),
    .Q(\am_sdr0.cic2.comb3_in_del[2] ));
 sg13g2_dfrbp_1 _14143_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net422),
    .D(net2126),
    .Q_N(_06375_),
    .Q(\am_sdr0.cic2.comb3_in_del[3] ));
 sg13g2_dfrbp_1 _14144_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net420),
    .D(net2530),
    .Q_N(_06374_),
    .Q(\am_sdr0.cic2.comb3_in_del[4] ));
 sg13g2_dfrbp_1 _14145_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net418),
    .D(net2382),
    .Q_N(_06373_),
    .Q(\am_sdr0.cic2.comb3_in_del[5] ));
 sg13g2_dfrbp_1 _14146_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net416),
    .D(net2250),
    .Q_N(_06372_),
    .Q(\am_sdr0.cic2.comb3_in_del[6] ));
 sg13g2_dfrbp_1 _14147_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net414),
    .D(net2586),
    .Q_N(_06371_),
    .Q(\am_sdr0.cic2.comb3_in_del[7] ));
 sg13g2_dfrbp_1 _14148_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net412),
    .D(net2326),
    .Q_N(_06370_),
    .Q(\am_sdr0.cic2.comb3_in_del[8] ));
 sg13g2_dfrbp_1 _14149_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net410),
    .D(net2173),
    .Q_N(_06369_),
    .Q(\am_sdr0.cic2.comb3_in_del[9] ));
 sg13g2_dfrbp_1 _14150_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net408),
    .D(net2334),
    .Q_N(_06368_),
    .Q(\am_sdr0.cic2.comb3_in_del[10] ));
 sg13g2_dfrbp_1 _14151_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net406),
    .D(net2512),
    .Q_N(_06367_),
    .Q(\am_sdr0.cic2.comb3_in_del[11] ));
 sg13g2_dfrbp_1 _14152_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net404),
    .D(_00539_),
    .Q_N(_06366_),
    .Q(\am_sdr0.cic2.comb3_in_del[12] ));
 sg13g2_dfrbp_1 _14153_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net402),
    .D(_00540_),
    .Q_N(_06365_),
    .Q(\am_sdr0.cic2.comb3_in_del[13] ));
 sg13g2_dfrbp_1 _14154_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net400),
    .D(_00541_),
    .Q_N(_06364_),
    .Q(\am_sdr0.cic2.comb3_in_del[14] ));
 sg13g2_dfrbp_1 _14155_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net398),
    .D(_00542_),
    .Q_N(_06363_),
    .Q(\am_sdr0.cic2.comb3_in_del[15] ));
 sg13g2_dfrbp_1 _14156_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net396),
    .D(_00543_),
    .Q_N(_06362_),
    .Q(\am_sdr0.cic2.comb3_in_del[16] ));
 sg13g2_dfrbp_1 _14157_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net394),
    .D(_00544_),
    .Q_N(_06361_),
    .Q(\am_sdr0.cic2.comb3_in_del[17] ));
 sg13g2_dfrbp_1 _14158_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net392),
    .D(_00545_),
    .Q_N(_06360_),
    .Q(\am_sdr0.cic2.comb3_in_del[18] ));
 sg13g2_dfrbp_1 _14159_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net390),
    .D(_00546_),
    .Q_N(_06359_),
    .Q(\am_sdr0.cic2.comb3_in_del[19] ));
 sg13g2_dfrbp_1 _14160_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net388),
    .D(_00547_),
    .Q_N(_06358_),
    .Q(\am_sdr0.cic2.count[0] ));
 sg13g2_dfrbp_1 _14161_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net386),
    .D(net1230),
    .Q_N(_06357_),
    .Q(\am_sdr0.cic2.count[1] ));
 sg13g2_dfrbp_1 _14162_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net384),
    .D(_00549_),
    .Q_N(_06356_),
    .Q(\am_sdr0.cic2.count[2] ));
 sg13g2_dfrbp_1 _14163_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net382),
    .D(_00550_),
    .Q_N(_06355_),
    .Q(\am_sdr0.cic2.count[3] ));
 sg13g2_dfrbp_1 _14164_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net380),
    .D(_00551_),
    .Q_N(_06354_),
    .Q(\am_sdr0.cic2.count[4] ));
 sg13g2_dfrbp_1 _14165_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net378),
    .D(_00552_),
    .Q_N(_06353_),
    .Q(\am_sdr0.cic2.count[5] ));
 sg13g2_dfrbp_1 _14166_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net376),
    .D(net2065),
    .Q_N(_06352_),
    .Q(\am_sdr0.cic2.count[6] ));
 sg13g2_dfrbp_1 _14167_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net374),
    .D(net1329),
    .Q_N(_06351_),
    .Q(\am_sdr0.cic2.count[7] ));
 sg13g2_dfrbp_1 _14168_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net372),
    .D(net1282),
    .Q_N(_06350_),
    .Q(\am_sdr0.cic2.integ1[0] ));
 sg13g2_dfrbp_1 _14169_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net370),
    .D(net2841),
    .Q_N(_06349_),
    .Q(\am_sdr0.cic2.integ1[1] ));
 sg13g2_dfrbp_1 _14170_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net368),
    .D(net2803),
    .Q_N(_06348_),
    .Q(\am_sdr0.cic2.integ1[2] ));
 sg13g2_dfrbp_1 _14171_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net366),
    .D(net2962),
    .Q_N(_06347_),
    .Q(\am_sdr0.cic2.integ1[3] ));
 sg13g2_dfrbp_1 _14172_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net364),
    .D(_00559_),
    .Q_N(_06346_),
    .Q(\am_sdr0.cic2.integ1[4] ));
 sg13g2_dfrbp_1 _14173_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net362),
    .D(net2979),
    .Q_N(_06345_),
    .Q(\am_sdr0.cic2.integ1[5] ));
 sg13g2_dfrbp_1 _14174_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net360),
    .D(_00561_),
    .Q_N(_06344_),
    .Q(\am_sdr0.cic2.integ1[6] ));
 sg13g2_dfrbp_1 _14175_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net358),
    .D(net3003),
    .Q_N(_06343_),
    .Q(\am_sdr0.cic2.integ1[7] ));
 sg13g2_dfrbp_1 _14176_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net356),
    .D(_00563_),
    .Q_N(_06342_),
    .Q(\am_sdr0.cic2.integ1[8] ));
 sg13g2_dfrbp_1 _14177_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net354),
    .D(_00564_),
    .Q_N(_06341_),
    .Q(\am_sdr0.cic2.integ1[9] ));
 sg13g2_dfrbp_1 _14178_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net352),
    .D(_00565_),
    .Q_N(_06340_),
    .Q(\am_sdr0.cic2.integ1[10] ));
 sg13g2_dfrbp_1 _14179_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net350),
    .D(_00566_),
    .Q_N(_06339_),
    .Q(\am_sdr0.cic2.integ1[11] ));
 sg13g2_dfrbp_1 _14180_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net348),
    .D(_00567_),
    .Q_N(_06338_),
    .Q(\am_sdr0.cic2.integ1[12] ));
 sg13g2_dfrbp_1 _14181_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net346),
    .D(_00568_),
    .Q_N(_06337_),
    .Q(\am_sdr0.cic2.integ1[13] ));
 sg13g2_dfrbp_1 _14182_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net344),
    .D(_00569_),
    .Q_N(_06336_),
    .Q(\am_sdr0.cic2.integ1[14] ));
 sg13g2_dfrbp_1 _14183_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net342),
    .D(_00570_),
    .Q_N(_06335_),
    .Q(\am_sdr0.cic2.integ1[15] ));
 sg13g2_dfrbp_1 _14184_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net340),
    .D(_00571_),
    .Q_N(_06334_),
    .Q(\am_sdr0.cic2.integ1[16] ));
 sg13g2_dfrbp_1 _14185_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net338),
    .D(_00572_),
    .Q_N(_06333_),
    .Q(\am_sdr0.cic2.integ1[17] ));
 sg13g2_dfrbp_1 _14186_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net336),
    .D(_00573_),
    .Q_N(_06332_),
    .Q(\am_sdr0.cic2.integ1[18] ));
 sg13g2_dfrbp_1 _14187_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net334),
    .D(_00574_),
    .Q_N(_06331_),
    .Q(\am_sdr0.cic2.integ1[19] ));
 sg13g2_dfrbp_1 _14188_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net332),
    .D(_00575_),
    .Q_N(_06330_),
    .Q(\am_sdr0.cic2.integ1[20] ));
 sg13g2_dfrbp_1 _14189_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net330),
    .D(_00576_),
    .Q_N(_06329_),
    .Q(\am_sdr0.cic2.integ1[21] ));
 sg13g2_dfrbp_1 _14190_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net328),
    .D(_00577_),
    .Q_N(_06328_),
    .Q(\am_sdr0.cic2.integ1[22] ));
 sg13g2_dfrbp_1 _14191_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net326),
    .D(_00578_),
    .Q_N(_06327_),
    .Q(\am_sdr0.cic2.integ1[23] ));
 sg13g2_dfrbp_1 _14192_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net324),
    .D(_00579_),
    .Q_N(_06326_),
    .Q(\am_sdr0.cic2.integ1[24] ));
 sg13g2_dfrbp_1 _14193_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net322),
    .D(_00580_),
    .Q_N(_06325_),
    .Q(\am_sdr0.cic2.integ1[25] ));
 sg13g2_dfrbp_1 _14194_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net320),
    .D(_00581_),
    .Q_N(_06324_),
    .Q(\am_sdr0.cic2.integ2[0] ));
 sg13g2_dfrbp_1 _14195_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net318),
    .D(_00582_),
    .Q_N(_06323_),
    .Q(\am_sdr0.cic2.integ2[1] ));
 sg13g2_dfrbp_1 _14196_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net316),
    .D(net2716),
    .Q_N(_06322_),
    .Q(\am_sdr0.cic2.integ2[2] ));
 sg13g2_dfrbp_1 _14197_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net314),
    .D(_00584_),
    .Q_N(_06321_),
    .Q(\am_sdr0.cic2.integ2[3] ));
 sg13g2_dfrbp_1 _14198_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net312),
    .D(net3173),
    .Q_N(_06320_),
    .Q(\am_sdr0.cic2.integ2[4] ));
 sg13g2_dfrbp_1 _14199_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net310),
    .D(_00586_),
    .Q_N(_06319_),
    .Q(\am_sdr0.cic2.integ2[5] ));
 sg13g2_dfrbp_1 _14200_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net308),
    .D(_00587_),
    .Q_N(_06318_),
    .Q(\am_sdr0.cic2.integ2[6] ));
 sg13g2_dfrbp_1 _14201_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net306),
    .D(_00588_),
    .Q_N(_06317_),
    .Q(\am_sdr0.cic2.integ2[7] ));
 sg13g2_dfrbp_1 _14202_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net304),
    .D(_00589_),
    .Q_N(_06316_),
    .Q(\am_sdr0.cic2.integ2[8] ));
 sg13g2_dfrbp_1 _14203_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net302),
    .D(_00590_),
    .Q_N(_06315_),
    .Q(\am_sdr0.cic2.integ2[9] ));
 sg13g2_dfrbp_1 _14204_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net300),
    .D(_00591_),
    .Q_N(_06314_),
    .Q(\am_sdr0.cic2.integ2[10] ));
 sg13g2_dfrbp_1 _14205_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net298),
    .D(_00592_),
    .Q_N(_06313_),
    .Q(\am_sdr0.cic2.integ2[11] ));
 sg13g2_dfrbp_1 _14206_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net296),
    .D(_00593_),
    .Q_N(_06312_),
    .Q(\am_sdr0.cic2.integ2[12] ));
 sg13g2_dfrbp_1 _14207_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net294),
    .D(_00594_),
    .Q_N(_06311_),
    .Q(\am_sdr0.cic2.integ2[13] ));
 sg13g2_dfrbp_1 _14208_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net292),
    .D(_00595_),
    .Q_N(_06310_),
    .Q(\am_sdr0.cic2.integ2[14] ));
 sg13g2_dfrbp_1 _14209_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net290),
    .D(_00596_),
    .Q_N(_06309_),
    .Q(\am_sdr0.cic2.integ2[15] ));
 sg13g2_dfrbp_1 _14210_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net288),
    .D(_00597_),
    .Q_N(_06308_),
    .Q(\am_sdr0.cic2.integ2[16] ));
 sg13g2_dfrbp_1 _14211_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net286),
    .D(_00598_),
    .Q_N(_06307_),
    .Q(\am_sdr0.cic2.integ2[17] ));
 sg13g2_dfrbp_1 _14212_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net284),
    .D(_00599_),
    .Q_N(_06306_),
    .Q(\am_sdr0.cic2.integ2[18] ));
 sg13g2_dfrbp_1 _14213_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net282),
    .D(_00600_),
    .Q_N(_06305_),
    .Q(\am_sdr0.cic2.integ2[19] ));
 sg13g2_dfrbp_1 _14214_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net280),
    .D(_00601_),
    .Q_N(_06304_),
    .Q(\am_sdr0.cic2.integ2[20] ));
 sg13g2_dfrbp_1 _14215_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net278),
    .D(_00602_),
    .Q_N(_06303_),
    .Q(\am_sdr0.cic2.integ2[21] ));
 sg13g2_dfrbp_1 _14216_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net276),
    .D(_00603_),
    .Q_N(_06302_),
    .Q(\am_sdr0.cic2.integ2[22] ));
 sg13g2_dfrbp_1 _14217_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net274),
    .D(_00604_),
    .Q_N(_06301_),
    .Q(\am_sdr0.cic2.integ3[0] ));
 sg13g2_dfrbp_1 _14218_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net272),
    .D(_00605_),
    .Q_N(_06300_),
    .Q(\am_sdr0.cic2.integ3[1] ));
 sg13g2_dfrbp_1 _14219_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net270),
    .D(_00606_),
    .Q_N(_06299_),
    .Q(\am_sdr0.cic2.integ3[2] ));
 sg13g2_dfrbp_1 _14220_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net268),
    .D(_00607_),
    .Q_N(_06298_),
    .Q(\am_sdr0.cic2.integ3[3] ));
 sg13g2_dfrbp_1 _14221_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net266),
    .D(_00608_),
    .Q_N(_06297_),
    .Q(\am_sdr0.cic2.integ3[4] ));
 sg13g2_dfrbp_1 _14222_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net264),
    .D(_00609_),
    .Q_N(_06296_),
    .Q(\am_sdr0.cic2.integ3[5] ));
 sg13g2_dfrbp_1 _14223_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net262),
    .D(_00610_),
    .Q_N(_06295_),
    .Q(\am_sdr0.cic2.integ3[6] ));
 sg13g2_dfrbp_1 _14224_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net260),
    .D(_00611_),
    .Q_N(_06294_),
    .Q(\am_sdr0.cic2.integ3[7] ));
 sg13g2_dfrbp_1 _14225_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net258),
    .D(_00612_),
    .Q_N(_06293_),
    .Q(\am_sdr0.cic2.integ3[8] ));
 sg13g2_dfrbp_1 _14226_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net256),
    .D(_00613_),
    .Q_N(_06292_),
    .Q(\am_sdr0.cic2.integ3[9] ));
 sg13g2_dfrbp_1 _14227_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net254),
    .D(_00614_),
    .Q_N(_06291_),
    .Q(\am_sdr0.cic2.integ3[10] ));
 sg13g2_dfrbp_1 _14228_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net252),
    .D(_00615_),
    .Q_N(_06290_),
    .Q(\am_sdr0.cic2.integ3[11] ));
 sg13g2_dfrbp_1 _14229_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net250),
    .D(_00616_),
    .Q_N(_06289_),
    .Q(\am_sdr0.cic2.integ3[12] ));
 sg13g2_dfrbp_1 _14230_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net248),
    .D(net2988),
    .Q_N(_06288_),
    .Q(\am_sdr0.cic2.integ3[13] ));
 sg13g2_dfrbp_1 _14231_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net246),
    .D(_00618_),
    .Q_N(_06287_),
    .Q(\am_sdr0.cic2.integ3[14] ));
 sg13g2_dfrbp_1 _14232_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net244),
    .D(net3022),
    .Q_N(_06286_),
    .Q(\am_sdr0.cic2.integ3[15] ));
 sg13g2_dfrbp_1 _14233_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net242),
    .D(_00620_),
    .Q_N(_06285_),
    .Q(\am_sdr0.cic2.integ3[16] ));
 sg13g2_dfrbp_1 _14234_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net240),
    .D(net2970),
    .Q_N(_06284_),
    .Q(\am_sdr0.cic2.integ3[17] ));
 sg13g2_dfrbp_1 _14235_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net238),
    .D(_00622_),
    .Q_N(_06283_),
    .Q(\am_sdr0.cic2.integ3[18] ));
 sg13g2_dfrbp_1 _14236_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net236),
    .D(_00623_),
    .Q_N(_06282_),
    .Q(\am_sdr0.cic2.integ3[19] ));
 sg13g2_dfrbp_1 _14237_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net234),
    .D(net1546),
    .Q_N(_06281_),
    .Q(\am_sdr0.cic1.sample ));
 sg13g2_dfrbp_1 _14238_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net233),
    .D(_00625_),
    .Q_N(_06280_),
    .Q(\am_sdr0.cic1.integ3[0] ));
 sg13g2_dfrbp_1 _14239_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net232),
    .D(_00626_),
    .Q_N(_06279_),
    .Q(\am_sdr0.cic1.integ3[1] ));
 sg13g2_dfrbp_1 _14240_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net231),
    .D(_00627_),
    .Q_N(_06278_),
    .Q(\am_sdr0.cic1.integ3[2] ));
 sg13g2_dfrbp_1 _14241_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net230),
    .D(net3131),
    .Q_N(_06277_),
    .Q(\am_sdr0.cic1.integ3[3] ));
 sg13g2_dfrbp_1 _14242_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net229),
    .D(_00629_),
    .Q_N(_06276_),
    .Q(\am_sdr0.cic1.integ3[4] ));
 sg13g2_dfrbp_1 _14243_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net228),
    .D(net3106),
    .Q_N(_06275_),
    .Q(\am_sdr0.cic1.integ3[5] ));
 sg13g2_dfrbp_1 _14244_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net227),
    .D(net3254),
    .Q_N(_06274_),
    .Q(\am_sdr0.cic1.integ3[6] ));
 sg13g2_dfrbp_1 _14245_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net226),
    .D(_00632_),
    .Q_N(_06273_),
    .Q(\am_sdr0.cic1.integ3[7] ));
 sg13g2_dfrbp_1 _14246_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net225),
    .D(_00633_),
    .Q_N(_06272_),
    .Q(\am_sdr0.cic1.integ3[8] ));
 sg13g2_dfrbp_1 _14247_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net224),
    .D(net3228),
    .Q_N(_06271_),
    .Q(\am_sdr0.cic1.integ3[9] ));
 sg13g2_dfrbp_1 _14248_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net223),
    .D(_00635_),
    .Q_N(_06270_),
    .Q(\am_sdr0.cic1.integ3[10] ));
 sg13g2_dfrbp_1 _14249_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net222),
    .D(_00636_),
    .Q_N(_06269_),
    .Q(\am_sdr0.cic1.integ3[11] ));
 sg13g2_dfrbp_1 _14250_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net221),
    .D(_00637_),
    .Q_N(_06268_),
    .Q(\am_sdr0.cic1.integ3[12] ));
 sg13g2_dfrbp_1 _14251_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net220),
    .D(_00638_),
    .Q_N(_06267_),
    .Q(\am_sdr0.cic1.integ3[13] ));
 sg13g2_dfrbp_1 _14252_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net219),
    .D(_00639_),
    .Q_N(_06266_),
    .Q(\am_sdr0.cic1.integ3[14] ));
 sg13g2_dfrbp_1 _14253_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net218),
    .D(_00640_),
    .Q_N(_06265_),
    .Q(\am_sdr0.cic1.integ3[15] ));
 sg13g2_dfrbp_1 _14254_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net217),
    .D(net3088),
    .Q_N(_06264_),
    .Q(\am_sdr0.cic1.integ3[16] ));
 sg13g2_dfrbp_1 _14255_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net216),
    .D(_00642_),
    .Q_N(_06263_),
    .Q(\am_sdr0.cic1.integ3[17] ));
 sg13g2_dfrbp_1 _14256_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net215),
    .D(net2999),
    .Q_N(_06262_),
    .Q(\am_sdr0.cic1.integ3[18] ));
 sg13g2_dfrbp_1 _14257_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net214),
    .D(net2983),
    .Q_N(_06261_),
    .Q(\am_sdr0.cic1.integ3[19] ));
 sg13g2_dfrbp_1 _14258_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net213),
    .D(net2524),
    .Q_N(_06260_),
    .Q(\am_sdr0.cic0.integ_sample[0] ));
 sg13g2_dfrbp_1 _14259_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net212),
    .D(net2291),
    .Q_N(_06259_),
    .Q(\am_sdr0.cic0.integ_sample[1] ));
 sg13g2_dfrbp_1 _14260_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net211),
    .D(net1500),
    .Q_N(_06258_),
    .Q(\am_sdr0.cic0.integ_sample[2] ));
 sg13g2_dfrbp_1 _14261_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net210),
    .D(net1434),
    .Q_N(_06257_),
    .Q(\am_sdr0.cic0.integ_sample[3] ));
 sg13g2_dfrbp_1 _14262_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net209),
    .D(net1502),
    .Q_N(_06256_),
    .Q(\am_sdr0.cic0.integ_sample[4] ));
 sg13g2_dfrbp_1 _14263_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net208),
    .D(net2053),
    .Q_N(_06255_),
    .Q(\am_sdr0.cic0.integ_sample[5] ));
 sg13g2_dfrbp_1 _14264_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net207),
    .D(net1401),
    .Q_N(_06254_),
    .Q(\am_sdr0.cic0.integ_sample[6] ));
 sg13g2_dfrbp_1 _14265_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net206),
    .D(net2056),
    .Q_N(_06253_),
    .Q(\am_sdr0.cic0.integ_sample[7] ));
 sg13g2_dfrbp_1 _14266_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net205),
    .D(net1438),
    .Q_N(_06252_),
    .Q(\am_sdr0.cic0.integ_sample[8] ));
 sg13g2_dfrbp_1 _14267_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net204),
    .D(net1444),
    .Q_N(_06251_),
    .Q(\am_sdr0.cic0.integ_sample[9] ));
 sg13g2_dfrbp_1 _14268_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net203),
    .D(net1513),
    .Q_N(_06250_),
    .Q(\am_sdr0.cic0.integ_sample[10] ));
 sg13g2_dfrbp_1 _14269_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net202),
    .D(net2241),
    .Q_N(_06249_),
    .Q(\am_sdr0.cic0.integ_sample[11] ));
 sg13g2_dfrbp_1 _14270_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net201),
    .D(net2268),
    .Q_N(_06248_),
    .Q(\am_sdr0.cic0.integ_sample[12] ));
 sg13g2_dfrbp_1 _14271_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net200),
    .D(net2206),
    .Q_N(_06247_),
    .Q(\am_sdr0.cic0.integ_sample[13] ));
 sg13g2_dfrbp_1 _14272_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net199),
    .D(net2110),
    .Q_N(_06246_),
    .Q(\am_sdr0.cic0.integ_sample[14] ));
 sg13g2_dfrbp_1 _14273_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net198),
    .D(net2868),
    .Q_N(_06245_),
    .Q(\am_sdr0.cic0.integ_sample[15] ));
 sg13g2_dfrbp_1 _14274_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net197),
    .D(net1519),
    .Q_N(_06244_),
    .Q(\am_sdr0.cic0.integ_sample[16] ));
 sg13g2_dfrbp_1 _14275_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net196),
    .D(net2598),
    .Q_N(_06243_),
    .Q(\am_sdr0.cic0.integ_sample[17] ));
 sg13g2_dfrbp_1 _14276_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net195),
    .D(net1515),
    .Q_N(_06242_),
    .Q(\am_sdr0.cic0.integ_sample[18] ));
 sg13g2_dfrbp_1 _14277_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net194),
    .D(net1310),
    .Q_N(_06241_),
    .Q(\am_sdr0.cic0.integ_sample[19] ));
 sg13g2_dfrbp_1 _14278_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net193),
    .D(net1284),
    .Q_N(_06240_),
    .Q(\am_sdr0.cic1.x_out[8] ));
 sg13g2_dfrbp_1 _14279_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net191),
    .D(net1338),
    .Q_N(_06239_),
    .Q(\am_sdr0.cic1.x_out[9] ));
 sg13g2_dfrbp_1 _14280_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net189),
    .D(net1242),
    .Q_N(_06238_),
    .Q(\am_sdr0.cic1.x_out[10] ));
 sg13g2_dfrbp_1 _14281_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net187),
    .D(net1227),
    .Q_N(_06237_),
    .Q(\am_sdr0.cic1.x_out[11] ));
 sg13g2_dfrbp_1 _14282_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net185),
    .D(net1367),
    .Q_N(_06236_),
    .Q(\am_sdr0.cic1.x_out[12] ));
 sg13g2_dfrbp_1 _14283_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net183),
    .D(net1348),
    .Q_N(_06235_),
    .Q(\am_sdr0.cic1.x_out[13] ));
 sg13g2_dfrbp_1 _14284_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net181),
    .D(net1265),
    .Q_N(_06234_),
    .Q(\am_sdr0.cic1.x_out[14] ));
 sg13g2_dfrbp_1 _14285_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net179),
    .D(net1485),
    .Q_N(_06233_),
    .Q(\am_sdr0.cic1.x_out[15] ));
 sg13g2_dfrbp_1 _14286_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net177),
    .D(_00673_),
    .Q_N(_06232_),
    .Q(\am_sdr0.cic1.comb1[0] ));
 sg13g2_dfrbp_1 _14287_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net175),
    .D(_00674_),
    .Q_N(_06231_),
    .Q(\am_sdr0.cic1.comb1[1] ));
 sg13g2_dfrbp_1 _14288_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net173),
    .D(_00675_),
    .Q_N(_06230_),
    .Q(\am_sdr0.cic1.comb1[2] ));
 sg13g2_dfrbp_1 _14289_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net171),
    .D(_00676_),
    .Q_N(_06229_),
    .Q(\am_sdr0.cic1.comb1[3] ));
 sg13g2_dfrbp_1 _14290_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net169),
    .D(_00677_),
    .Q_N(_06228_),
    .Q(\am_sdr0.cic1.comb1[4] ));
 sg13g2_dfrbp_1 _14291_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net167),
    .D(net3013),
    .Q_N(_06227_),
    .Q(\am_sdr0.cic1.comb1[5] ));
 sg13g2_dfrbp_1 _14292_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net165),
    .D(_00679_),
    .Q_N(_06226_),
    .Q(\am_sdr0.cic1.comb1[6] ));
 sg13g2_dfrbp_1 _14293_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net163),
    .D(_00680_),
    .Q_N(_06225_),
    .Q(\am_sdr0.cic1.comb1[7] ));
 sg13g2_dfrbp_1 _14294_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net161),
    .D(_00681_),
    .Q_N(_06224_),
    .Q(\am_sdr0.cic1.comb1[8] ));
 sg13g2_dfrbp_1 _14295_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net159),
    .D(net2951),
    .Q_N(_06223_),
    .Q(\am_sdr0.cic1.comb1[9] ));
 sg13g2_dfrbp_1 _14296_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net157),
    .D(_00683_),
    .Q_N(_06222_),
    .Q(\am_sdr0.cic1.comb1[10] ));
 sg13g2_dfrbp_1 _14297_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net155),
    .D(_00684_),
    .Q_N(_06221_),
    .Q(\am_sdr0.cic1.comb1[11] ));
 sg13g2_dfrbp_1 _14298_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net153),
    .D(_00685_),
    .Q_N(_06220_),
    .Q(\am_sdr0.cic1.comb1[12] ));
 sg13g2_dfrbp_1 _14299_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net151),
    .D(_00686_),
    .Q_N(_06219_),
    .Q(\am_sdr0.cic1.comb1[13] ));
 sg13g2_dfrbp_1 _14300_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net149),
    .D(_00687_),
    .Q_N(_06218_),
    .Q(\am_sdr0.cic1.comb1[14] ));
 sg13g2_dfrbp_1 _14301_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net147),
    .D(_00688_),
    .Q_N(_06217_),
    .Q(\am_sdr0.cic1.comb1[15] ));
 sg13g2_dfrbp_1 _14302_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net145),
    .D(_00689_),
    .Q_N(_06216_),
    .Q(\am_sdr0.cic1.comb1[16] ));
 sg13g2_dfrbp_1 _14303_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net143),
    .D(net2817),
    .Q_N(_06215_),
    .Q(\am_sdr0.cic1.comb1[17] ));
 sg13g2_dfrbp_1 _14304_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net141),
    .D(_00691_),
    .Q_N(_06214_),
    .Q(\am_sdr0.cic1.comb1[18] ));
 sg13g2_dfrbp_1 _14305_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net139),
    .D(_00692_),
    .Q_N(_06213_),
    .Q(\am_sdr0.cic1.comb1[19] ));
 sg13g2_dfrbp_1 _14306_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net137),
    .D(net2036),
    .Q_N(_06212_),
    .Q(\am_sdr0.cic1.comb1_in_del[0] ));
 sg13g2_dfrbp_1 _14307_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net135),
    .D(net2360),
    .Q_N(_06211_),
    .Q(\am_sdr0.cic1.comb1_in_del[1] ));
 sg13g2_dfrbp_1 _14308_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net133),
    .D(net2562),
    .Q_N(_06210_),
    .Q(\am_sdr0.cic1.comb1_in_del[2] ));
 sg13g2_dfrbp_1 _14309_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net129),
    .D(net2594),
    .Q_N(_06209_),
    .Q(\am_sdr0.cic1.comb1_in_del[3] ));
 sg13g2_dfrbp_1 _14310_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net125),
    .D(net2693),
    .Q_N(_06208_),
    .Q(\am_sdr0.cic1.comb1_in_del[4] ));
 sg13g2_dfrbp_1 _14311_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net81),
    .D(net2878),
    .Q_N(_06207_),
    .Q(\am_sdr0.cic1.comb1_in_del[5] ));
 sg13g2_dfrbp_1 _14312_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net77),
    .D(net2752),
    .Q_N(_06206_),
    .Q(\am_sdr0.cic1.comb1_in_del[6] ));
 sg13g2_dfrbp_1 _14313_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net73),
    .D(net2570),
    .Q_N(_06205_),
    .Q(\am_sdr0.cic1.comb1_in_del[7] ));
 sg13g2_dfrbp_1 _14314_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net69),
    .D(net2701),
    .Q_N(_06204_),
    .Q(\am_sdr0.cic1.comb1_in_del[8] ));
 sg13g2_dfrbp_1 _14315_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net65),
    .D(net2904),
    .Q_N(_06203_),
    .Q(\am_sdr0.cic1.comb1_in_del[9] ));
 sg13g2_dfrbp_1 _14316_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net61),
    .D(net2657),
    .Q_N(_06202_),
    .Q(\am_sdr0.cic1.comb1_in_del[10] ));
 sg13g2_dfrbp_1 _14317_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net57),
    .D(net2299),
    .Q_N(_06201_),
    .Q(\am_sdr0.cic1.comb1_in_del[11] ));
 sg13g2_dfrbp_1 _14318_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net53),
    .D(net2714),
    .Q_N(_06200_),
    .Q(\am_sdr0.cic1.comb1_in_del[12] ));
 sg13g2_dfrbp_1 _14319_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net49),
    .D(_00706_),
    .Q_N(_06199_),
    .Q(\am_sdr0.cic1.comb1_in_del[13] ));
 sg13g2_dfrbp_1 _14320_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net45),
    .D(net2580),
    .Q_N(_06198_),
    .Q(\am_sdr0.cic1.comb1_in_del[14] ));
 sg13g2_dfrbp_1 _14321_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net41),
    .D(net2412),
    .Q_N(_06197_),
    .Q(\am_sdr0.cic1.comb1_in_del[15] ));
 sg13g2_dfrbp_1 _14322_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net37),
    .D(net2754),
    .Q_N(_06196_),
    .Q(\am_sdr0.cic1.comb1_in_del[16] ));
 sg13g2_dfrbp_1 _14323_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net27),
    .D(_00710_),
    .Q_N(_06195_),
    .Q(\am_sdr0.cic1.comb1_in_del[17] ));
 sg13g2_dfrbp_1 _14324_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1159),
    .D(net2664),
    .Q_N(_06194_),
    .Q(\am_sdr0.cic1.comb1_in_del[18] ));
 sg13g2_dfrbp_1 _14325_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1155),
    .D(net2142),
    .Q_N(_06193_),
    .Q(\am_sdr0.cic1.comb1_in_del[19] ));
 sg13g2_dfrbp_1 _14326_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1151),
    .D(_00713_),
    .Q_N(_06192_),
    .Q(\am_sdr0.cic1.comb2[0] ));
 sg13g2_dfrbp_1 _14327_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1123),
    .D(_00714_),
    .Q_N(_06191_),
    .Q(\am_sdr0.cic1.comb2[1] ));
 sg13g2_dfrbp_1 _14328_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1119),
    .D(net2902),
    .Q_N(_06190_),
    .Q(\am_sdr0.cic1.comb2[2] ));
 sg13g2_dfrbp_1 _14329_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1115),
    .D(_00716_),
    .Q_N(_06189_),
    .Q(\am_sdr0.cic1.comb2[3] ));
 sg13g2_dfrbp_1 _14330_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1111),
    .D(_00717_),
    .Q_N(_06188_),
    .Q(\am_sdr0.cic1.comb2[4] ));
 sg13g2_dfrbp_1 _14331_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1107),
    .D(net2865),
    .Q_N(_06187_),
    .Q(\am_sdr0.cic1.comb2[5] ));
 sg13g2_dfrbp_1 _14332_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1102),
    .D(_00719_),
    .Q_N(_06186_),
    .Q(\am_sdr0.cic1.comb2[6] ));
 sg13g2_dfrbp_1 _14333_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1098),
    .D(_00720_),
    .Q_N(_06185_),
    .Q(\am_sdr0.cic1.comb2[7] ));
 sg13g2_dfrbp_1 _14334_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1094),
    .D(_00721_),
    .Q_N(_06184_),
    .Q(\am_sdr0.cic1.comb2[8] ));
 sg13g2_dfrbp_1 _14335_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1090),
    .D(_00722_),
    .Q_N(_06183_),
    .Q(\am_sdr0.cic1.comb2[9] ));
 sg13g2_dfrbp_1 _14336_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1086),
    .D(_00723_),
    .Q_N(_06182_),
    .Q(\am_sdr0.cic1.comb2[10] ));
 sg13g2_dfrbp_1 _14337_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1082),
    .D(_00724_),
    .Q_N(_06181_),
    .Q(\am_sdr0.cic1.comb2[11] ));
 sg13g2_dfrbp_1 _14338_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1078),
    .D(_00725_),
    .Q_N(_06180_),
    .Q(\am_sdr0.cic1.comb2[12] ));
 sg13g2_dfrbp_1 _14339_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1074),
    .D(_00726_),
    .Q_N(_06179_),
    .Q(\am_sdr0.cic1.comb2[13] ));
 sg13g2_dfrbp_1 _14340_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1070),
    .D(_00727_),
    .Q_N(_06178_),
    .Q(\am_sdr0.cic1.comb2[14] ));
 sg13g2_dfrbp_1 _14341_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1066),
    .D(_00728_),
    .Q_N(_06177_),
    .Q(\am_sdr0.cic1.comb2[15] ));
 sg13g2_dfrbp_1 _14342_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1025),
    .D(_00729_),
    .Q_N(_06176_),
    .Q(\am_sdr0.cic1.comb2[16] ));
 sg13g2_dfrbp_1 _14343_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1021),
    .D(_00730_),
    .Q_N(_06175_),
    .Q(\am_sdr0.cic1.comb2[17] ));
 sg13g2_dfrbp_1 _14344_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1017),
    .D(_00731_),
    .Q_N(_06174_),
    .Q(\am_sdr0.cic1.comb2[18] ));
 sg13g2_dfrbp_1 _14345_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1013),
    .D(net2311),
    .Q_N(_06173_),
    .Q(\am_sdr0.cic1.comb2[19] ));
 sg13g2_dfrbp_1 _14346_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1009),
    .D(net2389),
    .Q_N(_06172_),
    .Q(\am_sdr0.cic1.comb2_in_del[0] ));
 sg13g2_dfrbp_1 _14347_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1005),
    .D(net2469),
    .Q_N(_06171_),
    .Q(\am_sdr0.cic1.comb2_in_del[1] ));
 sg13g2_dfrbp_1 _14348_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1001),
    .D(net2493),
    .Q_N(_06170_),
    .Q(\am_sdr0.cic1.comb2_in_del[2] ));
 sg13g2_dfrbp_1 _14349_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net997),
    .D(_00736_),
    .Q_N(_06169_),
    .Q(\am_sdr0.cic1.comb2_in_del[3] ));
 sg13g2_dfrbp_1 _14350_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net993),
    .D(net2671),
    .Q_N(_06168_),
    .Q(\am_sdr0.cic1.comb2_in_del[4] ));
 sg13g2_dfrbp_1 _14351_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net989),
    .D(net2584),
    .Q_N(_06167_),
    .Q(\am_sdr0.cic1.comb2_in_del[5] ));
 sg13g2_dfrbp_1 _14352_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net985),
    .D(_00739_),
    .Q_N(_06166_),
    .Q(\am_sdr0.cic1.comb2_in_del[6] ));
 sg13g2_dfrbp_1 _14353_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net981),
    .D(net2443),
    .Q_N(_06165_),
    .Q(\am_sdr0.cic1.comb2_in_del[7] ));
 sg13g2_dfrbp_1 _14354_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net977),
    .D(net2486),
    .Q_N(_06164_),
    .Q(\am_sdr0.cic1.comb2_in_del[8] ));
 sg13g2_dfrbp_1 _14355_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net973),
    .D(net2848),
    .Q_N(_06163_),
    .Q(\am_sdr0.cic1.comb2_in_del[9] ));
 sg13g2_dfrbp_1 _14356_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net969),
    .D(net2330),
    .Q_N(_06162_),
    .Q(\am_sdr0.cic1.comb2_in_del[10] ));
 sg13g2_dfrbp_1 _14357_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net965),
    .D(net2243),
    .Q_N(_06161_),
    .Q(\am_sdr0.cic1.comb2_in_del[11] ));
 sg13g2_dfrbp_1 _14358_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net961),
    .D(net2649),
    .Q_N(_06160_),
    .Q(\am_sdr0.cic1.comb2_in_del[12] ));
 sg13g2_dfrbp_1 _14359_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net957),
    .D(net2328),
    .Q_N(_06159_),
    .Q(\am_sdr0.cic1.comb2_in_del[13] ));
 sg13g2_dfrbp_1 _14360_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net953),
    .D(_00747_),
    .Q_N(_06158_),
    .Q(\am_sdr0.cic1.comb2_in_del[14] ));
 sg13g2_dfrbp_1 _14361_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net949),
    .D(net2607),
    .Q_N(_06157_),
    .Q(\am_sdr0.cic1.comb2_in_del[15] ));
 sg13g2_dfrbp_1 _14362_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net945),
    .D(_00749_),
    .Q_N(_06156_),
    .Q(\am_sdr0.cic1.comb2_in_del[16] ));
 sg13g2_dfrbp_1 _14363_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net941),
    .D(_00750_),
    .Q_N(_06155_),
    .Q(\am_sdr0.cic1.comb2_in_del[17] ));
 sg13g2_dfrbp_1 _14364_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net937),
    .D(_00751_),
    .Q_N(_06154_),
    .Q(\am_sdr0.cic1.comb2_in_del[18] ));
 sg13g2_dfrbp_1 _14365_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net933),
    .D(net2120),
    .Q_N(_06153_),
    .Q(\am_sdr0.cic1.comb2_in_del[19] ));
 sg13g2_dfrbp_1 _14366_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net929),
    .D(_00753_),
    .Q_N(_06152_),
    .Q(\am_sdr0.cic1.comb3[12] ));
 sg13g2_dfrbp_1 _14367_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net925),
    .D(_00754_),
    .Q_N(_06151_),
    .Q(\am_sdr0.cic1.comb3[13] ));
 sg13g2_dfrbp_1 _14368_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net921),
    .D(_00755_),
    .Q_N(_06150_),
    .Q(\am_sdr0.cic1.comb3[14] ));
 sg13g2_dfrbp_1 _14369_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net917),
    .D(_00756_),
    .Q_N(_06149_),
    .Q(\am_sdr0.cic1.comb3[15] ));
 sg13g2_dfrbp_1 _14370_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net913),
    .D(_00757_),
    .Q_N(_06148_),
    .Q(\am_sdr0.cic1.comb3[16] ));
 sg13g2_dfrbp_1 _14371_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net909),
    .D(net2031),
    .Q_N(_06147_),
    .Q(\am_sdr0.cic1.comb3[17] ));
 sg13g2_dfrbp_1 _14372_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net905),
    .D(_00759_),
    .Q_N(_06146_),
    .Q(\am_sdr0.cic1.comb3[18] ));
 sg13g2_dfrbp_1 _14373_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net901),
    .D(net2180),
    .Q_N(_06145_),
    .Q(\am_sdr0.cic1.comb3[19] ));
 sg13g2_dfrbp_1 _14374_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net897),
    .D(net2167),
    .Q_N(_06144_),
    .Q(\am_sdr0.cic1.comb3_in_del[0] ));
 sg13g2_dfrbp_1 _14375_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net893),
    .D(net2308),
    .Q_N(_06143_),
    .Q(\am_sdr0.cic1.comb3_in_del[1] ));
 sg13g2_dfrbp_1 _14376_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net889),
    .D(net2190),
    .Q_N(_06142_),
    .Q(\am_sdr0.cic1.comb3_in_del[2] ));
 sg13g2_dfrbp_1 _14377_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net885),
    .D(net2184),
    .Q_N(_06141_),
    .Q(\am_sdr0.cic1.comb3_in_del[3] ));
 sg13g2_dfrbp_1 _14378_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net881),
    .D(net2371),
    .Q_N(_06140_),
    .Q(\am_sdr0.cic1.comb3_in_del[4] ));
 sg13g2_dfrbp_1 _14379_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net877),
    .D(net2103),
    .Q_N(_06139_),
    .Q(\am_sdr0.cic1.comb3_in_del[5] ));
 sg13g2_dfrbp_1 _14380_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net873),
    .D(net2393),
    .Q_N(_06138_),
    .Q(\am_sdr0.cic1.comb3_in_del[6] ));
 sg13g2_dfrbp_1 _14381_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net869),
    .D(net2495),
    .Q_N(_06137_),
    .Q(\am_sdr0.cic1.comb3_in_del[7] ));
 sg13g2_dfrbp_1 _14382_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net865),
    .D(net2404),
    .Q_N(_06136_),
    .Q(\am_sdr0.cic1.comb3_in_del[8] ));
 sg13g2_dfrbp_1 _14383_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net861),
    .D(net2208),
    .Q_N(_06135_),
    .Q(\am_sdr0.cic1.comb3_in_del[9] ));
 sg13g2_dfrbp_1 _14384_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net857),
    .D(net2088),
    .Q_N(_06134_),
    .Q(\am_sdr0.cic1.comb3_in_del[10] ));
 sg13g2_dfrbp_1 _14385_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net853),
    .D(net2428),
    .Q_N(_06133_),
    .Q(\am_sdr0.cic1.comb3_in_del[11] ));
 sg13g2_dfrbp_1 _14386_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net849),
    .D(_00773_),
    .Q_N(_06132_),
    .Q(\am_sdr0.cic1.comb3_in_del[12] ));
 sg13g2_dfrbp_1 _14387_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net845),
    .D(_00774_),
    .Q_N(_06131_),
    .Q(\am_sdr0.cic1.comb3_in_del[13] ));
 sg13g2_dfrbp_1 _14388_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net841),
    .D(_00775_),
    .Q_N(_06130_),
    .Q(\am_sdr0.cic1.comb3_in_del[14] ));
 sg13g2_dfrbp_1 _14389_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net837),
    .D(_00776_),
    .Q_N(_06129_),
    .Q(\am_sdr0.cic1.comb3_in_del[15] ));
 sg13g2_dfrbp_1 _14390_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net833),
    .D(net2148),
    .Q_N(_06128_),
    .Q(\am_sdr0.cic1.comb3_in_del[16] ));
 sg13g2_dfrbp_1 _14391_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net829),
    .D(_00778_),
    .Q_N(_06127_),
    .Q(\am_sdr0.cic1.comb3_in_del[17] ));
 sg13g2_dfrbp_1 _14392_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net825),
    .D(net2146),
    .Q_N(_06126_),
    .Q(\am_sdr0.cic1.comb3_in_del[18] ));
 sg13g2_dfrbp_1 _14393_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net821),
    .D(net2062),
    .Q_N(_06125_),
    .Q(\am_sdr0.cic1.comb3_in_del[19] ));
 sg13g2_dfrbp_1 _14394_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net817),
    .D(_00781_),
    .Q_N(_06124_),
    .Q(\am_sdr0.cic1.out_tick ));
 sg13g2_dfrbp_1 _14395_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net815),
    .D(_00782_),
    .Q_N(_00075_),
    .Q(\am_sdr0.cic1.count[0] ));
 sg13g2_dfrbp_1 _14396_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net813),
    .D(_00783_),
    .Q_N(_06123_),
    .Q(\am_sdr0.cic1.count[1] ));
 sg13g2_dfrbp_1 _14397_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net811),
    .D(net1204),
    .Q_N(_06122_),
    .Q(\am_sdr0.cic1.count[2] ));
 sg13g2_dfrbp_1 _14398_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net809),
    .D(_00785_),
    .Q_N(_06121_),
    .Q(\am_sdr0.cic1.count[3] ));
 sg13g2_dfrbp_1 _14399_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net807),
    .D(_00786_),
    .Q_N(_06120_),
    .Q(\am_sdr0.cic1.count[4] ));
 sg13g2_dfrbp_1 _14400_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net805),
    .D(_00787_),
    .Q_N(_06119_),
    .Q(\am_sdr0.cic1.count[5] ));
 sg13g2_dfrbp_1 _14401_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net803),
    .D(net1374),
    .Q_N(_06118_),
    .Q(\am_sdr0.cic1.count[6] ));
 sg13g2_dfrbp_1 _14402_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net801),
    .D(net1209),
    .Q_N(_06117_),
    .Q(\am_sdr0.cic1.count[7] ));
 sg13g2_dfrbp_1 _14403_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net799),
    .D(net2187),
    .Q_N(_06116_),
    .Q(\am_sdr0.cic1.integ1[0] ));
 sg13g2_dfrbp_1 _14404_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net797),
    .D(net3124),
    .Q_N(_06115_),
    .Q(\am_sdr0.cic1.integ1[1] ));
 sg13g2_dfrbp_1 _14405_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net795),
    .D(net3086),
    .Q_N(_06114_),
    .Q(\am_sdr0.cic1.integ1[2] ));
 sg13g2_dfrbp_1 _14406_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net793),
    .D(_00793_),
    .Q_N(_06113_),
    .Q(\am_sdr0.cic1.integ1[3] ));
 sg13g2_dfrbp_1 _14407_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net791),
    .D(_00794_),
    .Q_N(_06112_),
    .Q(\am_sdr0.cic1.integ1[4] ));
 sg13g2_dfrbp_1 _14408_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net789),
    .D(net3059),
    .Q_N(_06111_),
    .Q(\am_sdr0.cic1.integ1[5] ));
 sg13g2_dfrbp_1 _14409_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net787),
    .D(net3151),
    .Q_N(_06110_),
    .Q(\am_sdr0.cic1.integ1[6] ));
 sg13g2_dfrbp_1 _14410_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net785),
    .D(_00797_),
    .Q_N(_06109_),
    .Q(\am_sdr0.cic1.integ1[7] ));
 sg13g2_dfrbp_1 _14411_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net783),
    .D(net3198),
    .Q_N(_06108_),
    .Q(\am_sdr0.cic1.integ1[8] ));
 sg13g2_dfrbp_1 _14412_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net781),
    .D(_00799_),
    .Q_N(_06107_),
    .Q(\am_sdr0.cic1.integ1[9] ));
 sg13g2_dfrbp_1 _14413_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net779),
    .D(_00800_),
    .Q_N(_06106_),
    .Q(\am_sdr0.cic1.integ1[10] ));
 sg13g2_dfrbp_1 _14414_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net777),
    .D(_00801_),
    .Q_N(_06105_),
    .Q(\am_sdr0.cic1.integ1[11] ));
 sg13g2_dfrbp_1 _14415_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net775),
    .D(_00802_),
    .Q_N(_06104_),
    .Q(\am_sdr0.cic1.integ1[12] ));
 sg13g2_dfrbp_1 _14416_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net773),
    .D(net3219),
    .Q_N(_06103_),
    .Q(\am_sdr0.cic1.integ1[13] ));
 sg13g2_dfrbp_1 _14417_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net771),
    .D(_00804_),
    .Q_N(_06102_),
    .Q(\am_sdr0.cic1.integ1[14] ));
 sg13g2_dfrbp_1 _14418_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net769),
    .D(_00805_),
    .Q_N(_06101_),
    .Q(\am_sdr0.cic1.integ1[15] ));
 sg13g2_dfrbp_1 _14419_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net767),
    .D(_00806_),
    .Q_N(_06100_),
    .Q(\am_sdr0.cic1.integ1[16] ));
 sg13g2_dfrbp_1 _14420_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net765),
    .D(net3265),
    .Q_N(_06099_),
    .Q(\am_sdr0.cic1.integ1[17] ));
 sg13g2_dfrbp_1 _14421_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net763),
    .D(_00808_),
    .Q_N(_06098_),
    .Q(\am_sdr0.cic1.integ1[18] ));
 sg13g2_dfrbp_1 _14422_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net761),
    .D(_00809_),
    .Q_N(_06097_),
    .Q(\am_sdr0.cic1.integ1[19] ));
 sg13g2_dfrbp_1 _14423_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net759),
    .D(_00810_),
    .Q_N(_06096_),
    .Q(\am_sdr0.cic1.integ1[20] ));
 sg13g2_dfrbp_1 _14424_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net757),
    .D(_00811_),
    .Q_N(_06095_),
    .Q(\am_sdr0.cic1.integ1[21] ));
 sg13g2_dfrbp_1 _14425_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net755),
    .D(_00812_),
    .Q_N(_06094_),
    .Q(\am_sdr0.cic1.integ1[22] ));
 sg13g2_dfrbp_1 _14426_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net753),
    .D(_00813_),
    .Q_N(_06093_),
    .Q(\am_sdr0.cic1.integ1[23] ));
 sg13g2_dfrbp_1 _14427_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net751),
    .D(_00814_),
    .Q_N(_06092_),
    .Q(\am_sdr0.cic1.integ1[24] ));
 sg13g2_dfrbp_1 _14428_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net749),
    .D(_00815_),
    .Q_N(_06091_),
    .Q(\am_sdr0.cic1.integ1[25] ));
 sg13g2_dfrbp_1 _14429_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net747),
    .D(_00816_),
    .Q_N(_06090_),
    .Q(\am_sdr0.cic1.integ2[0] ));
 sg13g2_dfrbp_1 _14430_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net745),
    .D(net2943),
    .Q_N(_06089_),
    .Q(\am_sdr0.cic1.integ2[1] ));
 sg13g2_dfrbp_1 _14431_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net743),
    .D(_00818_),
    .Q_N(_06088_),
    .Q(\am_sdr0.cic1.integ2[2] ));
 sg13g2_dfrbp_1 _14432_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net741),
    .D(net3177),
    .Q_N(_06087_),
    .Q(\am_sdr0.cic1.integ2[3] ));
 sg13g2_dfrbp_1 _14433_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net739),
    .D(_00820_),
    .Q_N(_06086_),
    .Q(\am_sdr0.cic1.integ2[4] ));
 sg13g2_dfrbp_1 _14434_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net737),
    .D(net3171),
    .Q_N(_06085_),
    .Q(\am_sdr0.cic1.integ2[5] ));
 sg13g2_dfrbp_1 _14435_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net735),
    .D(_00822_),
    .Q_N(_06084_),
    .Q(\am_sdr0.cic1.integ2[6] ));
 sg13g2_dfrbp_1 _14436_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net733),
    .D(_00823_),
    .Q_N(_06083_),
    .Q(\am_sdr0.cic1.integ2[7] ));
 sg13g2_dfrbp_1 _14437_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net731),
    .D(_00824_),
    .Q_N(_06082_),
    .Q(\am_sdr0.cic1.integ2[8] ));
 sg13g2_dfrbp_1 _14438_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net729),
    .D(_00825_),
    .Q_N(_06081_),
    .Q(\am_sdr0.cic1.integ2[9] ));
 sg13g2_dfrbp_1 _14439_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net727),
    .D(_00826_),
    .Q_N(_06080_),
    .Q(\am_sdr0.cic1.integ2[10] ));
 sg13g2_dfrbp_1 _14440_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net725),
    .D(net3258),
    .Q_N(_06079_),
    .Q(\am_sdr0.cic1.integ2[11] ));
 sg13g2_dfrbp_1 _14441_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net723),
    .D(_00828_),
    .Q_N(_06078_),
    .Q(\am_sdr0.cic1.integ2[12] ));
 sg13g2_dfrbp_1 _14442_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net721),
    .D(_00829_),
    .Q_N(_06077_),
    .Q(\am_sdr0.cic1.integ2[13] ));
 sg13g2_dfrbp_1 _14443_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net719),
    .D(_00830_),
    .Q_N(_06076_),
    .Q(\am_sdr0.cic1.integ2[14] ));
 sg13g2_dfrbp_1 _14444_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net717),
    .D(_00831_),
    .Q_N(_06075_),
    .Q(\am_sdr0.cic1.integ2[15] ));
 sg13g2_dfrbp_1 _14445_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net715),
    .D(_00832_),
    .Q_N(_06074_),
    .Q(\am_sdr0.cic1.integ2[16] ));
 sg13g2_dfrbp_1 _14446_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net713),
    .D(net3167),
    .Q_N(_06073_),
    .Q(\am_sdr0.cic1.integ2[17] ));
 sg13g2_dfrbp_1 _14447_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net711),
    .D(_00834_),
    .Q_N(_06072_),
    .Q(\am_sdr0.cic1.integ2[18] ));
 sg13g2_dfrbp_1 _14448_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net709),
    .D(_00835_),
    .Q_N(_06071_),
    .Q(\am_sdr0.cic1.integ2[19] ));
 sg13g2_dfrbp_1 _14449_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net707),
    .D(_00836_),
    .Q_N(_06070_),
    .Q(\am_sdr0.cic1.integ2[20] ));
 sg13g2_dfrbp_1 _14450_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net705),
    .D(_00837_),
    .Q_N(_06069_),
    .Q(\am_sdr0.cic1.integ2[21] ));
 sg13g2_dfrbp_1 _14451_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net703),
    .D(net3043),
    .Q_N(_06068_),
    .Q(\am_sdr0.cic1.integ2[22] ));
 sg13g2_dfrbp_1 _14452_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net701),
    .D(net1545),
    .Q_N(_06067_),
    .Q(\am_sdr0.cic0.sample ));
 sg13g2_dfrbp_1 _14453_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net699),
    .D(_00840_),
    .Q_N(_06066_),
    .Q(\am_sdr0.cic0.integ3[0] ));
 sg13g2_dfrbp_1 _14454_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net697),
    .D(_00841_),
    .Q_N(_06065_),
    .Q(\am_sdr0.cic0.integ3[1] ));
 sg13g2_dfrbp_1 _14455_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net695),
    .D(_00842_),
    .Q_N(_06064_),
    .Q(\am_sdr0.cic0.integ3[2] ));
 sg13g2_dfrbp_1 _14456_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net693),
    .D(net3143),
    .Q_N(_06063_),
    .Q(\am_sdr0.cic0.integ3[3] ));
 sg13g2_dfrbp_1 _14457_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net691),
    .D(_00844_),
    .Q_N(_06062_),
    .Q(\am_sdr0.cic0.integ3[4] ));
 sg13g2_dfrbp_1 _14458_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net689),
    .D(net3100),
    .Q_N(_06061_),
    .Q(\am_sdr0.cic0.integ3[5] ));
 sg13g2_dfrbp_1 _14459_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net687),
    .D(_00846_),
    .Q_N(_06060_),
    .Q(\am_sdr0.cic0.integ3[6] ));
 sg13g2_dfrbp_1 _14460_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net685),
    .D(_00847_),
    .Q_N(_06059_),
    .Q(\am_sdr0.cic0.integ3[7] ));
 sg13g2_dfrbp_1 _14461_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net683),
    .D(_00848_),
    .Q_N(_06058_),
    .Q(\am_sdr0.cic0.integ3[8] ));
 sg13g2_dfrbp_1 _14462_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net681),
    .D(net3209),
    .Q_N(_06057_),
    .Q(\am_sdr0.cic0.integ3[9] ));
 sg13g2_dfrbp_1 _14463_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net679),
    .D(_00850_),
    .Q_N(_06056_),
    .Q(\am_sdr0.cic0.integ3[10] ));
 sg13g2_dfrbp_1 _14464_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net677),
    .D(_00851_),
    .Q_N(_06055_),
    .Q(\am_sdr0.cic0.integ3[11] ));
 sg13g2_dfrbp_1 _14465_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net675),
    .D(_00852_),
    .Q_N(_06054_),
    .Q(\am_sdr0.cic0.integ3[12] ));
 sg13g2_dfrbp_1 _14466_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net673),
    .D(net3180),
    .Q_N(_06053_),
    .Q(\am_sdr0.cic0.integ3[13] ));
 sg13g2_dfrbp_1 _14467_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net671),
    .D(_00854_),
    .Q_N(_06052_),
    .Q(\am_sdr0.cic0.integ3[14] ));
 sg13g2_dfrbp_1 _14468_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net669),
    .D(_00855_),
    .Q_N(_06051_),
    .Q(\am_sdr0.cic0.integ3[15] ));
 sg13g2_dfrbp_1 _14469_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net667),
    .D(net3094),
    .Q_N(_06050_),
    .Q(\am_sdr0.cic0.integ3[16] ));
 sg13g2_dfrbp_1 _14470_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net665),
    .D(_00857_),
    .Q_N(_06049_),
    .Q(\am_sdr0.cic0.integ3[17] ));
 sg13g2_dfrbp_1 _14471_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net663),
    .D(net3027),
    .Q_N(_06048_),
    .Q(\am_sdr0.cic0.integ3[18] ));
 sg13g2_dfrbp_1 _14472_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net661),
    .D(net3020),
    .Q_N(_06047_),
    .Q(\am_sdr0.cic0.integ3[19] ));
 sg13g2_dfrbp_1 _14473_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net659),
    .D(net1303),
    .Q_N(_06046_),
    .Q(\am_sdr0.spi0.shift_reg[0] ));
 sg13g2_dfrbp_1 _14474_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net655),
    .D(_00861_),
    .Q_N(_06045_),
    .Q(\am_sdr0.spi0.shift_reg[1] ));
 sg13g2_dfrbp_1 _14475_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net651),
    .D(_00862_),
    .Q_N(_06044_),
    .Q(\am_sdr0.spi0.shift_reg[2] ));
 sg13g2_dfrbp_1 _14476_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net647),
    .D(_00863_),
    .Q_N(_06043_),
    .Q(\am_sdr0.spi0.shift_reg[3] ));
 sg13g2_dfrbp_1 _14477_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net643),
    .D(_00864_),
    .Q_N(_06042_),
    .Q(\am_sdr0.spi0.shift_reg[4] ));
 sg13g2_dfrbp_1 _14478_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net617),
    .D(net1331),
    .Q_N(_06041_),
    .Q(\am_sdr0.spi0.shift_reg[5] ));
 sg13g2_dfrbp_1 _14479_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net613),
    .D(_00866_),
    .Q_N(_06040_),
    .Q(\am_sdr0.spi0.shift_reg[6] ));
 sg13g2_dfrbp_1 _14480_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net609),
    .D(_00867_),
    .Q_N(_06039_),
    .Q(\am_sdr0.spi0.shift_reg[7] ));
 sg13g2_dfrbp_1 _14481_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net605),
    .D(_00868_),
    .Q_N(_06038_),
    .Q(\am_sdr0.spi0.shift_reg[8] ));
 sg13g2_dfrbp_1 _14482_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net601),
    .D(net1383),
    .Q_N(_06037_),
    .Q(\am_sdr0.spi0.shift_reg[9] ));
 sg13g2_dfrbp_1 _14483_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net597),
    .D(net1316),
    .Q_N(_06036_),
    .Q(\am_sdr0.spi0.shift_reg[10] ));
 sg13g2_dfrbp_1 _14484_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net593),
    .D(_00871_),
    .Q_N(_06035_),
    .Q(\am_sdr0.spi0.shift_reg[11] ));
 sg13g2_dfrbp_1 _14485_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net589),
    .D(net1363),
    .Q_N(_06034_),
    .Q(\am_sdr0.spi0.shift_reg[12] ));
 sg13g2_dfrbp_1 _14486_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net585),
    .D(net1299),
    .Q_N(_06033_),
    .Q(\am_sdr0.spi0.shift_reg[13] ));
 sg13g2_dfrbp_1 _14487_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net581),
    .D(_00874_),
    .Q_N(_06032_),
    .Q(\am_sdr0.spi0.shift_reg[14] ));
 sg13g2_dfrbp_1 _14488_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net577),
    .D(_00875_),
    .Q_N(_06031_),
    .Q(\am_sdr0.spi0.shift_reg[15] ));
 sg13g2_dfrbp_1 _14489_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net573),
    .D(net1394),
    .Q_N(_06030_),
    .Q(\am_sdr0.spi0.shift_reg[16] ));
 sg13g2_dfrbp_1 _14490_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net569),
    .D(net1361),
    .Q_N(_06029_),
    .Q(\am_sdr0.spi0.shift_reg[17] ));
 sg13g2_dfrbp_1 _14491_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net565),
    .D(_00878_),
    .Q_N(_06028_),
    .Q(\am_sdr0.spi0.shift_reg[18] ));
 sg13g2_dfrbp_1 _14492_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net561),
    .D(net1290),
    .Q_N(_06027_),
    .Q(\am_sdr0.spi0.shift_reg[19] ));
 sg13g2_dfrbp_1 _14493_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net557),
    .D(_00880_),
    .Q_N(_06026_),
    .Q(\am_sdr0.spi0.shift_reg[20] ));
 sg13g2_dfrbp_1 _14494_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net553),
    .D(_00881_),
    .Q_N(_06025_),
    .Q(\am_sdr0.spi0.shift_reg[21] ));
 sg13g2_dfrbp_1 _14495_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net549),
    .D(_00882_),
    .Q_N(_06024_),
    .Q(\am_sdr0.spi0.shift_reg[22] ));
 sg13g2_dfrbp_1 _14496_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net545),
    .D(net1416),
    .Q_N(_06023_),
    .Q(\am_sdr0.spi0.shift_reg[23] ));
 sg13g2_dfrbp_1 _14497_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net541),
    .D(net1344),
    .Q_N(_06022_),
    .Q(\am_sdr0.spi0.shift_reg[24] ));
 sg13g2_dfrbp_1 _14498_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net537),
    .D(_00885_),
    .Q_N(_06021_),
    .Q(\am_sdr0.spi0.shift_reg[25] ));
 sg13g2_dfrbp_1 _14499_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net533),
    .D(_00886_),
    .Q_N(_06020_),
    .Q(\am_sdr0.spi0.shift_reg[26] ));
 sg13g2_dfrbp_1 _14500_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net529),
    .D(net1483),
    .Q_N(_06019_),
    .Q(\am_sdr0.spi0.shift_reg[27] ));
 sg13g2_dfrbp_1 _14501_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net525),
    .D(net1236),
    .Q_N(_06018_),
    .Q(\am_sdr0.spi0.shift_reg[28] ));
 sg13g2_dfrbp_1 _14502_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net521),
    .D(net1504),
    .Q_N(_06017_),
    .Q(\am_sdr0.cic0.x_out[8] ));
 sg13g2_dfrbp_1 _14503_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net517),
    .D(net1340),
    .Q_N(_06016_),
    .Q(\am_sdr0.cic0.x_out[9] ));
 sg13g2_dfrbp_1 _14504_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net513),
    .D(net1479),
    .Q_N(_06015_),
    .Q(\am_sdr0.cic0.x_out[10] ));
 sg13g2_dfrbp_1 _14505_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net509),
    .D(net1496),
    .Q_N(_06014_),
    .Q(\am_sdr0.cic0.x_out[11] ));
 sg13g2_dfrbp_1 _14506_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net505),
    .D(net1270),
    .Q_N(_06013_),
    .Q(\am_sdr0.cic0.x_out[12] ));
 sg13g2_dfrbp_1 _14507_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net501),
    .D(net1307),
    .Q_N(_06012_),
    .Q(\am_sdr0.cic0.x_out[13] ));
 sg13g2_dfrbp_1 _14508_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net497),
    .D(net1294),
    .Q_N(_06011_),
    .Q(\am_sdr0.cic0.x_out[14] ));
 sg13g2_dfrbp_1 _14509_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net493),
    .D(_00896_),
    .Q_N(_06010_),
    .Q(\am_sdr0.cic0.x_out[15] ));
 sg13g2_dfrbp_1 _14510_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net489),
    .D(_00897_),
    .Q_N(_06009_),
    .Q(\am_sdr0.cic0.comb1[0] ));
 sg13g2_dfrbp_1 _14511_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net485),
    .D(_00898_),
    .Q_N(_06008_),
    .Q(\am_sdr0.cic0.comb1[1] ));
 sg13g2_dfrbp_1 _14512_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net481),
    .D(_00899_),
    .Q_N(_06007_),
    .Q(\am_sdr0.cic0.comb1[2] ));
 sg13g2_dfrbp_1 _14513_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net477),
    .D(_00900_),
    .Q_N(_06006_),
    .Q(\am_sdr0.cic0.comb1[3] ));
 sg13g2_dfrbp_1 _14514_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net473),
    .D(net2824),
    .Q_N(_06005_),
    .Q(\am_sdr0.cic0.comb1[4] ));
 sg13g2_dfrbp_1 _14515_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net469),
    .D(_00902_),
    .Q_N(_06004_),
    .Q(\am_sdr0.cic0.comb1[5] ));
 sg13g2_dfrbp_1 _14516_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net465),
    .D(_00903_),
    .Q_N(_06003_),
    .Q(\am_sdr0.cic0.comb1[6] ));
 sg13g2_dfrbp_1 _14517_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net461),
    .D(_00904_),
    .Q_N(_06002_),
    .Q(\am_sdr0.cic0.comb1[7] ));
 sg13g2_dfrbp_1 _14518_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net457),
    .D(_00905_),
    .Q_N(_06001_),
    .Q(\am_sdr0.cic0.comb1[8] ));
 sg13g2_dfrbp_1 _14519_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net453),
    .D(_00906_),
    .Q_N(_06000_),
    .Q(\am_sdr0.cic0.comb1[9] ));
 sg13g2_dfrbp_1 _14520_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net449),
    .D(_00907_),
    .Q_N(_05999_),
    .Q(\am_sdr0.cic0.comb1[10] ));
 sg13g2_dfrbp_1 _14521_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net445),
    .D(_00908_),
    .Q_N(_05998_),
    .Q(\am_sdr0.cic0.comb1[11] ));
 sg13g2_dfrbp_1 _14522_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net441),
    .D(net3048),
    .Q_N(_05997_),
    .Q(\am_sdr0.cic0.comb1[12] ));
 sg13g2_dfrbp_1 _14523_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net437),
    .D(net2695),
    .Q_N(_05996_),
    .Q(\am_sdr0.cic0.comb1[13] ));
 sg13g2_dfrbp_1 _14524_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net433),
    .D(_00911_),
    .Q_N(_05995_),
    .Q(\am_sdr0.cic0.comb1[14] ));
 sg13g2_dfrbp_1 _14525_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net429),
    .D(_00912_),
    .Q_N(_05994_),
    .Q(\am_sdr0.cic0.comb1[15] ));
 sg13g2_dfrbp_1 _14526_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net425),
    .D(_00913_),
    .Q_N(_05993_),
    .Q(\am_sdr0.cic0.comb1[16] ));
 sg13g2_dfrbp_1 _14527_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net421),
    .D(_00914_),
    .Q_N(_05992_),
    .Q(\am_sdr0.cic0.comb1[17] ));
 sg13g2_dfrbp_1 _14528_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net417),
    .D(_00915_),
    .Q_N(_05991_),
    .Q(\am_sdr0.cic0.comb1[18] ));
 sg13g2_dfrbp_1 _14529_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net413),
    .D(_00916_),
    .Q_N(_05990_),
    .Q(\am_sdr0.cic0.comb1[19] ));
 sg13g2_dfrbp_1 _14530_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net409),
    .D(net2122),
    .Q_N(_05989_),
    .Q(\am_sdr0.cic0.comb1_in_del[0] ));
 sg13g2_dfrbp_1 _14531_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net405),
    .D(net2668),
    .Q_N(_05988_),
    .Q(\am_sdr0.cic0.comb1_in_del[1] ));
 sg13g2_dfrbp_1 _14532_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net401),
    .D(net2706),
    .Q_N(_05987_),
    .Q(\am_sdr0.cic0.comb1_in_del[2] ));
 sg13g2_dfrbp_1 _14533_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net397),
    .D(net2465),
    .Q_N(_05986_),
    .Q(\am_sdr0.cic0.comb1_in_del[3] ));
 sg13g2_dfrbp_1 _14534_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net393),
    .D(net2739),
    .Q_N(_05985_),
    .Q(\am_sdr0.cic0.comb1_in_del[4] ));
 sg13g2_dfrbp_1 _14535_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net389),
    .D(_00922_),
    .Q_N(_05984_),
    .Q(\am_sdr0.cic0.comb1_in_del[5] ));
 sg13g2_dfrbp_1 _14536_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net385),
    .D(net2686),
    .Q_N(_05983_),
    .Q(\am_sdr0.cic0.comb1_in_del[6] ));
 sg13g2_dfrbp_1 _14537_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net381),
    .D(net2625),
    .Q_N(_05982_),
    .Q(\am_sdr0.cic0.comb1_in_del[7] ));
 sg13g2_dfrbp_1 _14538_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net377),
    .D(_00925_),
    .Q_N(_05981_),
    .Q(\am_sdr0.cic0.comb1_in_del[8] ));
 sg13g2_dfrbp_1 _14539_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net373),
    .D(net2844),
    .Q_N(_05980_),
    .Q(\am_sdr0.cic0.comb1_in_del[9] ));
 sg13g2_dfrbp_1 _14540_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net369),
    .D(net2637),
    .Q_N(_05979_),
    .Q(\am_sdr0.cic0.comb1_in_del[10] ));
 sg13g2_dfrbp_1 _14541_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net365),
    .D(net2293),
    .Q_N(_05978_),
    .Q(\am_sdr0.cic0.comb1_in_del[11] ));
 sg13g2_dfrbp_1 _14542_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net361),
    .D(net2574),
    .Q_N(_05977_),
    .Q(\am_sdr0.cic0.comb1_in_del[12] ));
 sg13g2_dfrbp_1 _14543_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net357),
    .D(net2217),
    .Q_N(_05976_),
    .Q(\am_sdr0.cic0.comb1_in_del[13] ));
 sg13g2_dfrbp_1 _14544_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net353),
    .D(net2463),
    .Q_N(_05975_),
    .Q(\am_sdr0.cic0.comb1_in_del[14] ));
 sg13g2_dfrbp_1 _14545_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net349),
    .D(net2710),
    .Q_N(_05974_),
    .Q(\am_sdr0.cic0.comb1_in_del[15] ));
 sg13g2_dfrbp_1 _14546_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net345),
    .D(net2556),
    .Q_N(_05973_),
    .Q(\am_sdr0.cic0.comb1_in_del[16] ));
 sg13g2_dfrbp_1 _14547_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net341),
    .D(_00934_),
    .Q_N(_05972_),
    .Q(\am_sdr0.cic0.comb1_in_del[17] ));
 sg13g2_dfrbp_1 _14548_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net337),
    .D(_00935_),
    .Q_N(_05971_),
    .Q(\am_sdr0.cic0.comb1_in_del[18] ));
 sg13g2_dfrbp_1 _14549_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net333),
    .D(net2288),
    .Q_N(_05970_),
    .Q(\am_sdr0.cic0.comb1_in_del[19] ));
 sg13g2_dfrbp_1 _14550_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net329),
    .D(_00937_),
    .Q_N(_05969_),
    .Q(\am_sdr0.cic0.comb2[0] ));
 sg13g2_dfrbp_1 _14551_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net325),
    .D(_00938_),
    .Q_N(_05968_),
    .Q(\am_sdr0.cic0.comb2[1] ));
 sg13g2_dfrbp_1 _14552_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net321),
    .D(net2914),
    .Q_N(_05967_),
    .Q(\am_sdr0.cic0.comb2[2] ));
 sg13g2_dfrbp_1 _14553_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net317),
    .D(_00940_),
    .Q_N(_05966_),
    .Q(\am_sdr0.cic0.comb2[3] ));
 sg13g2_dfrbp_1 _14554_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net313),
    .D(net2400),
    .Q_N(_05965_),
    .Q(\am_sdr0.cic0.comb2[4] ));
 sg13g2_dfrbp_1 _14555_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net309),
    .D(net2712),
    .Q_N(_05964_),
    .Q(\am_sdr0.cic0.comb2[5] ));
 sg13g2_dfrbp_1 _14556_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net305),
    .D(_00943_),
    .Q_N(_05963_),
    .Q(\am_sdr0.cic0.comb2[6] ));
 sg13g2_dfrbp_1 _14557_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net301),
    .D(_00944_),
    .Q_N(_05962_),
    .Q(\am_sdr0.cic0.comb2[7] ));
 sg13g2_dfrbp_1 _14558_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net297),
    .D(_00945_),
    .Q_N(_05961_),
    .Q(\am_sdr0.cic0.comb2[8] ));
 sg13g2_dfrbp_1 _14559_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net293),
    .D(net2881),
    .Q_N(_05960_),
    .Q(\am_sdr0.cic0.comb2[9] ));
 sg13g2_dfrbp_1 _14560_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net289),
    .D(_00947_),
    .Q_N(_05959_),
    .Q(\am_sdr0.cic0.comb2[10] ));
 sg13g2_dfrbp_1 _14561_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net285),
    .D(_00948_),
    .Q_N(_05958_),
    .Q(\am_sdr0.cic0.comb2[11] ));
 sg13g2_dfrbp_1 _14562_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net281),
    .D(_00949_),
    .Q_N(_05957_),
    .Q(\am_sdr0.cic0.comb2[12] ));
 sg13g2_dfrbp_1 _14563_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net277),
    .D(_00950_),
    .Q_N(_05956_),
    .Q(\am_sdr0.cic0.comb2[13] ));
 sg13g2_dfrbp_1 _14564_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net273),
    .D(_00951_),
    .Q_N(_05955_),
    .Q(\am_sdr0.cic0.comb2[14] ));
 sg13g2_dfrbp_1 _14565_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net269),
    .D(_00952_),
    .Q_N(_05954_),
    .Q(\am_sdr0.cic0.comb2[15] ));
 sg13g2_dfrbp_1 _14566_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net265),
    .D(_00953_),
    .Q_N(_05953_),
    .Q(\am_sdr0.cic0.comb2[16] ));
 sg13g2_dfrbp_1 _14567_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net261),
    .D(_00954_),
    .Q_N(_05952_),
    .Q(\am_sdr0.cic0.comb2[17] ));
 sg13g2_dfrbp_1 _14568_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net257),
    .D(_00955_),
    .Q_N(_05951_),
    .Q(\am_sdr0.cic0.comb2[18] ));
 sg13g2_dfrbp_1 _14569_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net253),
    .D(net2489),
    .Q_N(_05950_),
    .Q(\am_sdr0.cic0.comb2[19] ));
 sg13g2_dfrbp_1 _14570_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net249),
    .D(net2378),
    .Q_N(_05949_),
    .Q(\am_sdr0.cic0.comb2_in_del[0] ));
 sg13g2_dfrbp_1 _14571_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net245),
    .D(net2673),
    .Q_N(_05948_),
    .Q(\am_sdr0.cic0.comb2_in_del[1] ));
 sg13g2_dfrbp_1 _14572_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net241),
    .D(net2546),
    .Q_N(_05947_),
    .Q(\am_sdr0.cic0.comb2_in_del[2] ));
 sg13g2_dfrbp_1 _14573_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net237),
    .D(_00960_),
    .Q_N(_05946_),
    .Q(\am_sdr0.cic0.comb2_in_del[3] ));
 sg13g2_dfrbp_1 _14574_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net192),
    .D(_00961_),
    .Q_N(_05945_),
    .Q(\am_sdr0.cic0.comb2_in_del[4] ));
 sg13g2_dfrbp_1 _14575_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net188),
    .D(net2432),
    .Q_N(_05944_),
    .Q(\am_sdr0.cic0.comb2_in_del[5] ));
 sg13g2_dfrbp_1 _14576_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net184),
    .D(net2332),
    .Q_N(_05943_),
    .Q(\am_sdr0.cic0.comb2_in_del[6] ));
 sg13g2_dfrbp_1 _14577_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net180),
    .D(net2108),
    .Q_N(_05942_),
    .Q(\am_sdr0.cic0.comb2_in_del[7] ));
 sg13g2_dfrbp_1 _14578_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net176),
    .D(_00965_),
    .Q_N(_05941_),
    .Q(\am_sdr0.cic0.comb2_in_del[8] ));
 sg13g2_dfrbp_1 _14579_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net172),
    .D(net2895),
    .Q_N(_05940_),
    .Q(\am_sdr0.cic0.comb2_in_del[9] ));
 sg13g2_dfrbp_1 _14580_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net168),
    .D(net2402),
    .Q_N(_05939_),
    .Q(\am_sdr0.cic0.comb2_in_del[10] ));
 sg13g2_dfrbp_1 _14581_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net164),
    .D(net2284),
    .Q_N(_05938_),
    .Q(\am_sdr0.cic0.comb2_in_del[11] ));
 sg13g2_dfrbp_1 _14582_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net160),
    .D(net2578),
    .Q_N(_05937_),
    .Q(\am_sdr0.cic0.comb2_in_del[12] ));
 sg13g2_dfrbp_1 _14583_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net156),
    .D(_00970_),
    .Q_N(_05936_),
    .Q(\am_sdr0.cic0.comb2_in_del[13] ));
 sg13g2_dfrbp_1 _14584_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net152),
    .D(net2473),
    .Q_N(_05935_),
    .Q(\am_sdr0.cic0.comb2_in_del[14] ));
 sg13g2_dfrbp_1 _14585_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net148),
    .D(net2744),
    .Q_N(_05934_),
    .Q(\am_sdr0.cic0.comb2_in_del[15] ));
 sg13g2_dfrbp_1 _14586_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net144),
    .D(net2273),
    .Q_N(_05933_),
    .Q(\am_sdr0.cic0.comb2_in_del[16] ));
 sg13g2_dfrbp_1 _14587_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net140),
    .D(net2749),
    .Q_N(_05932_),
    .Q(\am_sdr0.cic0.comb2_in_del[17] ));
 sg13g2_dfrbp_1 _14588_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net136),
    .D(net2590),
    .Q_N(_05931_),
    .Q(\am_sdr0.cic0.comb2_in_del[18] ));
 sg13g2_dfrbp_1 _14589_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net131),
    .D(net2124),
    .Q_N(_05930_),
    .Q(\am_sdr0.cic0.comb2_in_del[19] ));
 sg13g2_dfrbp_1 _14590_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net83),
    .D(_00977_),
    .Q_N(_05929_),
    .Q(\am_sdr0.cic0.comb3[12] ));
 sg13g2_dfrbp_1 _14591_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net75),
    .D(_00978_),
    .Q_N(_05928_),
    .Q(\am_sdr0.cic0.comb3[13] ));
 sg13g2_dfrbp_1 _14592_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net67),
    .D(_00979_),
    .Q_N(_05927_),
    .Q(\am_sdr0.cic0.comb3[14] ));
 sg13g2_dfrbp_1 _14593_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net59),
    .D(_00980_),
    .Q_N(_05926_),
    .Q(\am_sdr0.cic0.comb3[15] ));
 sg13g2_dfrbp_1 _14594_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net51),
    .D(_00981_),
    .Q_N(_05925_),
    .Q(\am_sdr0.cic0.comb3[16] ));
 sg13g2_dfrbp_1 _14595_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net43),
    .D(_00982_),
    .Q_N(_05924_),
    .Q(\am_sdr0.cic0.comb3[17] ));
 sg13g2_dfrbp_1 _14596_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net35),
    .D(_00983_),
    .Q_N(_05923_),
    .Q(\am_sdr0.cic0.comb3[18] ));
 sg13g2_dfrbp_1 _14597_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1157),
    .D(net2135),
    .Q_N(_05922_),
    .Q(\am_sdr0.cic0.comb3[19] ));
 sg13g2_dfrbp_1 _14598_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1125),
    .D(net2171),
    .Q_N(_05921_),
    .Q(\am_sdr0.cic0.comb3_in_del[0] ));
 sg13g2_dfrbp_1 _14599_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1117),
    .D(net2075),
    .Q_N(_05920_),
    .Q(\am_sdr0.cic0.comb3_in_del[1] ));
 sg13g2_dfrbp_1 _14600_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1109),
    .D(net2132),
    .Q_N(_05919_),
    .Q(\am_sdr0.cic0.comb3_in_del[2] ));
 sg13g2_dfrbp_1 _14601_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1100),
    .D(net2080),
    .Q_N(_05918_),
    .Q(\am_sdr0.cic0.comb3_in_del[3] ));
 sg13g2_dfrbp_1 _14602_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1092),
    .D(_00989_),
    .Q_N(_05917_),
    .Q(\am_sdr0.cic0.comb3_in_del[4] ));
 sg13g2_dfrbp_1 _14603_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1084),
    .D(net2276),
    .Q_N(_05916_),
    .Q(\am_sdr0.cic0.comb3_in_del[5] ));
 sg13g2_dfrbp_1 _14604_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1076),
    .D(net2418),
    .Q_N(_05915_),
    .Q(\am_sdr0.cic0.comb3_in_del[6] ));
 sg13g2_dfrbp_1 _14605_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1068),
    .D(net2502),
    .Q_N(_05914_),
    .Q(\am_sdr0.cic0.comb3_in_del[7] ));
 sg13g2_dfrbp_1 _14606_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1023),
    .D(net2320),
    .Q_N(_05913_),
    .Q(\am_sdr0.cic0.comb3_in_del[8] ));
 sg13g2_dfrbp_1 _14607_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1015),
    .D(net2225),
    .Q_N(_05912_),
    .Q(\am_sdr0.cic0.comb3_in_del[9] ));
 sg13g2_dfrbp_1 _14608_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1007),
    .D(_00995_),
    .Q_N(_05911_),
    .Q(\am_sdr0.cic0.comb3_in_del[10] ));
 sg13g2_dfrbp_1 _14609_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net999),
    .D(net2430),
    .Q_N(_05910_),
    .Q(\am_sdr0.cic0.comb3_in_del[11] ));
 sg13g2_dfrbp_1 _14610_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net991),
    .D(_00997_),
    .Q_N(_05909_),
    .Q(\am_sdr0.cic0.comb3_in_del[12] ));
 sg13g2_dfrbp_1 _14611_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net983),
    .D(_00998_),
    .Q_N(_05908_),
    .Q(\am_sdr0.cic0.comb3_in_del[13] ));
 sg13g2_dfrbp_1 _14612_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net975),
    .D(net2266),
    .Q_N(_05907_),
    .Q(\am_sdr0.cic0.comb3_in_del[14] ));
 sg13g2_dfrbp_1 _14613_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net967),
    .D(_01000_),
    .Q_N(_05906_),
    .Q(\am_sdr0.cic0.comb3_in_del[15] ));
 sg13g2_dfrbp_1 _14614_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net959),
    .D(_01001_),
    .Q_N(_05905_),
    .Q(\am_sdr0.cic0.comb3_in_del[16] ));
 sg13g2_dfrbp_1 _14615_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net951),
    .D(net2551),
    .Q_N(_05904_),
    .Q(\am_sdr0.cic0.comb3_in_del[17] ));
 sg13g2_dfrbp_1 _14616_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net943),
    .D(_01003_),
    .Q_N(_05903_),
    .Q(\am_sdr0.cic0.comb3_in_del[18] ));
 sg13g2_dfrbp_1 _14617_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net935),
    .D(_01004_),
    .Q_N(_05902_),
    .Q(\am_sdr0.cic0.comb3_in_del[19] ));
 sg13g2_dfrbp_1 _14618_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net927),
    .D(_01005_),
    .Q_N(_05901_),
    .Q(\am_sdr0.cic0.out_tick ));
 sg13g2_dfrbp_1 _14619_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net923),
    .D(_01006_),
    .Q_N(_00074_),
    .Q(\am_sdr0.cic0.count[0] ));
 sg13g2_dfrbp_1 _14620_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net919),
    .D(_01007_),
    .Q_N(_05900_),
    .Q(\am_sdr0.cic0.count[1] ));
 sg13g2_dfrbp_1 _14621_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net915),
    .D(net1221),
    .Q_N(_05899_),
    .Q(\am_sdr0.cic0.count[2] ));
 sg13g2_dfrbp_1 _14622_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net911),
    .D(_01009_),
    .Q_N(_05898_),
    .Q(\am_sdr0.cic0.count[3] ));
 sg13g2_dfrbp_1 _14623_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net907),
    .D(_01010_),
    .Q_N(_05897_),
    .Q(\am_sdr0.cic0.count[4] ));
 sg13g2_dfrbp_1 _14624_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net903),
    .D(_01011_),
    .Q_N(_05896_),
    .Q(\am_sdr0.cic0.count[5] ));
 sg13g2_dfrbp_1 _14625_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net899),
    .D(net1412),
    .Q_N(_05895_),
    .Q(\am_sdr0.cic0.count[6] ));
 sg13g2_dfrbp_1 _14626_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net895),
    .D(net1253),
    .Q_N(_05894_),
    .Q(\am_sdr0.cic0.count[7] ));
 sg13g2_dfrbp_1 _14627_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net891),
    .D(net2461),
    .Q_N(_05893_),
    .Q(\am_sdr0.cic0.integ1[0] ));
 sg13g2_dfrbp_1 _14628_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net887),
    .D(net3164),
    .Q_N(_05892_),
    .Q(\am_sdr0.cic0.integ1[1] ));
 sg13g2_dfrbp_1 _14629_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net883),
    .D(net3046),
    .Q_N(_05891_),
    .Q(\am_sdr0.cic0.integ1[2] ));
 sg13g2_dfrbp_1 _14630_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net879),
    .D(_01017_),
    .Q_N(_05890_),
    .Q(\am_sdr0.cic0.integ1[3] ));
 sg13g2_dfrbp_1 _14631_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net875),
    .D(_01018_),
    .Q_N(_05889_),
    .Q(\am_sdr0.cic0.integ1[4] ));
 sg13g2_dfrbp_1 _14632_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net871),
    .D(net3104),
    .Q_N(_05888_),
    .Q(\am_sdr0.cic0.integ1[5] ));
 sg13g2_dfrbp_1 _14633_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net867),
    .D(net3136),
    .Q_N(_05887_),
    .Q(\am_sdr0.cic0.integ1[6] ));
 sg13g2_dfrbp_1 _14634_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net863),
    .D(_01021_),
    .Q_N(_05886_),
    .Q(\am_sdr0.cic0.integ1[7] ));
 sg13g2_dfrbp_1 _14635_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net859),
    .D(_01022_),
    .Q_N(_05885_),
    .Q(\am_sdr0.cic0.integ1[8] ));
 sg13g2_dfrbp_1 _14636_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net855),
    .D(_01023_),
    .Q_N(_05884_),
    .Q(\am_sdr0.cic0.integ1[9] ));
 sg13g2_dfrbp_1 _14637_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net851),
    .D(net3214),
    .Q_N(_05883_),
    .Q(\am_sdr0.cic0.integ1[10] ));
 sg13g2_dfrbp_1 _14638_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net847),
    .D(_01025_),
    .Q_N(_05882_),
    .Q(\am_sdr0.cic0.integ1[11] ));
 sg13g2_dfrbp_1 _14639_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net843),
    .D(_01026_),
    .Q_N(_05881_),
    .Q(\am_sdr0.cic0.integ1[12] ));
 sg13g2_dfrbp_1 _14640_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net839),
    .D(net3221),
    .Q_N(_05880_),
    .Q(\am_sdr0.cic0.integ1[13] ));
 sg13g2_dfrbp_1 _14641_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net835),
    .D(net3223),
    .Q_N(_05879_),
    .Q(\am_sdr0.cic0.integ1[14] ));
 sg13g2_dfrbp_1 _14642_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net831),
    .D(_01029_),
    .Q_N(_05878_),
    .Q(\am_sdr0.cic0.integ1[15] ));
 sg13g2_dfrbp_1 _14643_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net827),
    .D(_01030_),
    .Q_N(_05877_),
    .Q(\am_sdr0.cic0.integ1[16] ));
 sg13g2_dfrbp_1 _14644_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net823),
    .D(net3279),
    .Q_N(_05876_),
    .Q(\am_sdr0.cic0.integ1[17] ));
 sg13g2_dfrbp_1 _14645_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net819),
    .D(_01032_),
    .Q_N(_05875_),
    .Q(\am_sdr0.cic0.integ1[18] ));
 sg13g2_dfrbp_1 _14646_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net657),
    .D(_01033_),
    .Q_N(_05874_),
    .Q(\am_sdr0.cic0.integ1[19] ));
 sg13g2_dfrbp_1 _14647_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net653),
    .D(_01034_),
    .Q_N(_05873_),
    .Q(\am_sdr0.cic0.integ1[20] ));
 sg13g2_dfrbp_1 _14648_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net649),
    .D(net3267),
    .Q_N(_05872_),
    .Q(\am_sdr0.cic0.integ1[21] ));
 sg13g2_dfrbp_1 _14649_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net645),
    .D(_01036_),
    .Q_N(_05871_),
    .Q(\am_sdr0.cic0.integ1[22] ));
 sg13g2_dfrbp_1 _14650_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net619),
    .D(_01037_),
    .Q_N(_05870_),
    .Q(\am_sdr0.cic0.integ1[23] ));
 sg13g2_dfrbp_1 _14651_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net615),
    .D(_01038_),
    .Q_N(_05869_),
    .Q(\am_sdr0.cic0.integ1[24] ));
 sg13g2_dfrbp_1 _14652_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net611),
    .D(_01039_),
    .Q_N(_05868_),
    .Q(\am_sdr0.cic0.integ1[25] ));
 sg13g2_dfrbp_1 _14653_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net607),
    .D(net2613),
    .Q_N(_05867_),
    .Q(\am_sdr0.cic0.integ2[0] ));
 sg13g2_dfrbp_1 _14654_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net603),
    .D(net2846),
    .Q_N(_05866_),
    .Q(\am_sdr0.cic0.integ2[1] ));
 sg13g2_dfrbp_1 _14655_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net599),
    .D(_01042_),
    .Q_N(_05865_),
    .Q(\am_sdr0.cic0.integ2[2] ));
 sg13g2_dfrbp_1 _14656_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net595),
    .D(net3204),
    .Q_N(_05864_),
    .Q(\am_sdr0.cic0.integ2[3] ));
 sg13g2_dfrbp_1 _14657_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net591),
    .D(_01044_),
    .Q_N(_05863_),
    .Q(\am_sdr0.cic0.integ2[4] ));
 sg13g2_dfrbp_1 _14658_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net587),
    .D(net3183),
    .Q_N(_05862_),
    .Q(\am_sdr0.cic0.integ2[5] ));
 sg13g2_dfrbp_1 _14659_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net583),
    .D(net3308),
    .Q_N(_05861_),
    .Q(\am_sdr0.cic0.integ2[6] ));
 sg13g2_dfrbp_1 _14660_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net579),
    .D(_01047_),
    .Q_N(_05860_),
    .Q(\am_sdr0.cic0.integ2[7] ));
 sg13g2_dfrbp_1 _14661_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net575),
    .D(_01048_),
    .Q_N(_05859_),
    .Q(\am_sdr0.cic0.integ2[8] ));
 sg13g2_dfrbp_1 _14662_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net571),
    .D(net3233),
    .Q_N(_05858_),
    .Q(\am_sdr0.cic0.integ2[9] ));
 sg13g2_dfrbp_1 _14663_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net567),
    .D(_01050_),
    .Q_N(_05857_),
    .Q(\am_sdr0.cic0.integ2[10] ));
 sg13g2_dfrbp_1 _14664_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net563),
    .D(_01051_),
    .Q_N(_05856_),
    .Q(\am_sdr0.cic0.integ2[11] ));
 sg13g2_dfrbp_1 _14665_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net559),
    .D(_01052_),
    .Q_N(_05855_),
    .Q(\am_sdr0.cic0.integ2[12] ));
 sg13g2_dfrbp_1 _14666_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net555),
    .D(_01053_),
    .Q_N(_05854_),
    .Q(\am_sdr0.cic0.integ2[13] ));
 sg13g2_dfrbp_1 _14667_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net551),
    .D(net3275),
    .Q_N(_05853_),
    .Q(\am_sdr0.cic0.integ2[14] ));
 sg13g2_dfrbp_1 _14668_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net547),
    .D(_01055_),
    .Q_N(_05852_),
    .Q(\am_sdr0.cic0.integ2[15] ));
 sg13g2_dfrbp_1 _14669_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net543),
    .D(_01056_),
    .Q_N(_05851_),
    .Q(\am_sdr0.cic0.integ2[16] ));
 sg13g2_dfrbp_1 _14670_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net539),
    .D(net3201),
    .Q_N(_05850_),
    .Q(\am_sdr0.cic0.integ2[17] ));
 sg13g2_dfrbp_1 _14671_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net535),
    .D(_01058_),
    .Q_N(_05849_),
    .Q(\am_sdr0.cic0.integ2[18] ));
 sg13g2_dfrbp_1 _14672_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net531),
    .D(net3261),
    .Q_N(_05848_),
    .Q(\am_sdr0.cic0.integ2[19] ));
 sg13g2_dfrbp_1 _14673_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net527),
    .D(_01060_),
    .Q_N(_05847_),
    .Q(\am_sdr0.cic0.integ2[20] ));
 sg13g2_dfrbp_1 _14674_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net523),
    .D(net3206),
    .Q_N(_05846_),
    .Q(\am_sdr0.cic0.integ2[21] ));
 sg13g2_dfrbp_1 _14675_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1034),
    .D(_01062_),
    .Q_N(_06819_),
    .Q(\am_sdr0.cic0.integ2[22] ));
 sg13g2_dfrbp_1 _14676_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1035),
    .D(net1168),
    .Q_N(_06820_),
    .Q(\am_sdr0.I_out[0] ));
 sg13g2_dfrbp_1 _14677_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1036),
    .D(_00023_),
    .Q_N(_06821_),
    .Q(\am_sdr0.I_out[1] ));
 sg13g2_dfrbp_1 _14678_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1037),
    .D(net1447),
    .Q_N(_06822_),
    .Q(\am_sdr0.I_out[2] ));
 sg13g2_dfrbp_1 _14679_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1038),
    .D(net1312),
    .Q_N(_06823_),
    .Q(\am_sdr0.I_out[3] ));
 sg13g2_dfrbp_1 _14680_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1039),
    .D(net1268),
    .Q_N(_06824_),
    .Q(\am_sdr0.I_out[4] ));
 sg13g2_dfrbp_1 _14681_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1040),
    .D(net1238),
    .Q_N(_06825_),
    .Q(\am_sdr0.I_out[5] ));
 sg13g2_dfrbp_1 _14682_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1041),
    .D(net2051),
    .Q_N(_06826_),
    .Q(\am_sdr0.I_out[6] ));
 sg13g2_dfrbp_1 _14683_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1042),
    .D(net1216),
    .Q_N(_06827_),
    .Q(\am_sdr0.I_out[7] ));
 sg13g2_dfrbp_1 _14684_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1043),
    .D(net1169),
    .Q_N(_06828_),
    .Q(\am_sdr0.Q_out[0] ));
 sg13g2_dfrbp_1 _14685_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1044),
    .D(_00030_),
    .Q_N(_06829_),
    .Q(\am_sdr0.Q_out[1] ));
 sg13g2_dfrbp_1 _14686_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1045),
    .D(net1461),
    .Q_N(_06830_),
    .Q(\am_sdr0.Q_out[2] ));
 sg13g2_dfrbp_1 _14687_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1046),
    .D(net1251),
    .Q_N(_06831_),
    .Q(\am_sdr0.Q_out[3] ));
 sg13g2_dfrbp_1 _14688_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1047),
    .D(net1327),
    .Q_N(_06832_),
    .Q(\am_sdr0.Q_out[4] ));
 sg13g2_dfrbp_1 _14689_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1048),
    .D(net1199),
    .Q_N(_06833_),
    .Q(\am_sdr0.Q_out[5] ));
 sg13g2_dfrbp_1 _14690_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1161),
    .D(net1207),
    .Q_N(_06834_),
    .Q(\am_sdr0.Q_out[6] ));
 sg13g2_dfrbp_1 _14691_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net519),
    .D(net1197),
    .Q_N(_05845_),
    .Q(\am_sdr0.Q_out[7] ));
 sg13g2_dfrbp_1 _14692_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net515),
    .D(_01063_),
    .Q_N(_05844_),
    .Q(\am_sdr0.cic3.integ_sample[0] ));
 sg13g2_dfrbp_1 _14693_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net511),
    .D(net2350),
    .Q_N(_05843_),
    .Q(\am_sdr0.cic3.integ_sample[1] ));
 sg13g2_dfrbp_1 _14694_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net507),
    .D(net2484),
    .Q_N(_05842_),
    .Q(\am_sdr0.cic3.integ_sample[2] ));
 sg13g2_dfrbp_1 _14695_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net503),
    .D(net2446),
    .Q_N(_05841_),
    .Q(\am_sdr0.cic3.integ_sample[3] ));
 sg13g2_dfrbp_1 _14696_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net499),
    .D(net2514),
    .Q_N(_05840_),
    .Q(\am_sdr0.cic3.integ_sample[4] ));
 sg13g2_dfrbp_1 _14697_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net495),
    .D(net2766),
    .Q_N(_05839_),
    .Q(\am_sdr0.cic3.integ_sample[5] ));
 sg13g2_dfrbp_1 _14698_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net491),
    .D(_01069_),
    .Q_N(_05838_),
    .Q(\am_sdr0.cic3.integ_sample[6] ));
 sg13g2_dfrbp_1 _14699_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net487),
    .D(net2508),
    .Q_N(_05837_),
    .Q(\am_sdr0.cic3.integ_sample[7] ));
 sg13g2_dfrbp_1 _14700_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net483),
    .D(net2505),
    .Q_N(_05836_),
    .Q(\am_sdr0.cic3.integ_sample[8] ));
 sg13g2_dfrbp_1 _14701_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net479),
    .D(net2406),
    .Q_N(_05835_),
    .Q(\am_sdr0.cic3.integ_sample[9] ));
 sg13g2_dfrbp_1 _14702_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net475),
    .D(net2426),
    .Q_N(_05834_),
    .Q(\am_sdr0.cic3.integ_sample[10] ));
 sg13g2_dfrbp_1 _14703_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net471),
    .D(net2303),
    .Q_N(_05833_),
    .Q(\am_sdr0.cic3.integ_sample[11] ));
 sg13g2_dfrbp_1 _14704_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net467),
    .D(net2726),
    .Q_N(_05832_),
    .Q(\am_sdr0.cic3.integ_sample[12] ));
 sg13g2_dfrbp_1 _14705_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net463),
    .D(net2788),
    .Q_N(_05831_),
    .Q(\am_sdr0.cic3.integ_sample[13] ));
 sg13g2_dfrbp_1 _14706_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net459),
    .D(net2280),
    .Q_N(_05830_),
    .Q(\am_sdr0.cic3.integ_sample[14] ));
 sg13g2_dfrbp_1 _14707_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net455),
    .D(net2734),
    .Q_N(_05829_),
    .Q(\am_sdr0.cic3.integ_sample[15] ));
 sg13g2_dfrbp_1 _14708_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net451),
    .D(net2518),
    .Q_N(_05828_),
    .Q(\am_sdr0.cic3.integ_sample[16] ));
 sg13g2_dfrbp_1 _14709_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net447),
    .D(net2792),
    .Q_N(_05827_),
    .Q(\am_sdr0.cic3.integ_sample[17] ));
 sg13g2_dfrbp_1 _14710_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net443),
    .D(net2231),
    .Q_N(_05826_),
    .Q(\am_sdr0.cic3.integ_sample[18] ));
 sg13g2_dfrbp_1 _14711_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net439),
    .D(net2195),
    .Q_N(_05825_),
    .Q(\am_sdr0.cic3.integ_sample[19] ));
 sg13g2_dfrbp_1 _14712_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net435),
    .D(_01083_),
    .Q_N(_05824_),
    .Q(COMP_OUT));
 sg13g2_dfrbp_1 _14713_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net431),
    .D(_01084_),
    .Q_N(_05823_),
    .Q(\am_sdr0.mix0.RF_in_q ));
 sg13g2_dfrbp_1 _14714_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net427),
    .D(_01085_),
    .Q_N(_05822_),
    .Q(\am_sdr0.mix0.RF_in_qq ));
 sg13g2_dfrbp_1 _14715_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net423),
    .D(_01086_),
    .Q_N(_05821_),
    .Q(\am_sdr0.mix0.sin_q[0] ));
 sg13g2_dfrbp_1 _14716_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net419),
    .D(_01087_),
    .Q_N(_05820_),
    .Q(\am_sdr0.mix0.sin_q[1] ));
 sg13g2_dfrbp_1 _14717_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net415),
    .D(_01088_),
    .Q_N(_00040_),
    .Q(\am_sdr0.mix0.sin_q[2] ));
 sg13g2_dfrbp_1 _14718_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net411),
    .D(_01089_),
    .Q_N(_05819_),
    .Q(\am_sdr0.mix0.sin_q[3] ));
 sg13g2_dfrbp_1 _14719_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net407),
    .D(_01090_),
    .Q_N(_00041_),
    .Q(\am_sdr0.mix0.sin_q[4] ));
 sg13g2_dfrbp_1 _14720_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net403),
    .D(_01091_),
    .Q_N(_05818_),
    .Q(\am_sdr0.mix0.sin_q[5] ));
 sg13g2_dfrbp_1 _14721_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net399),
    .D(_01092_),
    .Q_N(_00042_),
    .Q(\am_sdr0.mix0.sin_q[6] ));
 sg13g2_dfrbp_1 _14722_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net395),
    .D(_01093_),
    .Q_N(_05817_),
    .Q(\am_sdr0.mix0.sin_q[7] ));
 sg13g2_dfrbp_1 _14723_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net391),
    .D(_01094_),
    .Q_N(_05816_),
    .Q(\am_sdr0.mix0.cos_q[0] ));
 sg13g2_dfrbp_1 _14724_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net387),
    .D(_01095_),
    .Q_N(_05815_),
    .Q(\am_sdr0.mix0.cos_q[1] ));
 sg13g2_dfrbp_1 _14725_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net383),
    .D(_01096_),
    .Q_N(_00043_),
    .Q(\am_sdr0.mix0.cos_q[2] ));
 sg13g2_dfrbp_1 _14726_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net379),
    .D(_01097_),
    .Q_N(_05814_),
    .Q(\am_sdr0.mix0.cos_q[3] ));
 sg13g2_dfrbp_1 _14727_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net375),
    .D(_01098_),
    .Q_N(_00044_),
    .Q(\am_sdr0.mix0.cos_q[4] ));
 sg13g2_dfrbp_1 _14728_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net371),
    .D(_01099_),
    .Q_N(_05813_),
    .Q(\am_sdr0.mix0.cos_q[5] ));
 sg13g2_dfrbp_1 _14729_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net367),
    .D(_01100_),
    .Q_N(_00045_),
    .Q(\am_sdr0.mix0.cos_q[6] ));
 sg13g2_dfrbp_1 _14730_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net363),
    .D(_01101_),
    .Q_N(_05812_),
    .Q(\am_sdr0.mix0.cos_q[7] ));
 sg13g2_dfrbp_1 _14731_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net359),
    .D(net1176),
    .Q_N(_00073_),
    .Q(\am_sdr0.am0.count[0] ));
 sg13g2_dfrbp_1 _14732_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net351),
    .D(_01103_),
    .Q_N(_05811_),
    .Q(\am_sdr0.am0.count[1] ));
 sg13g2_dfrbp_1 _14733_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net343),
    .D(_01104_),
    .Q_N(_05810_),
    .Q(\am_sdr0.spi0.MOSI_q ));
 sg13g2_dfrbp_1 _14734_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net339),
    .D(_01105_),
    .Q_N(_05809_),
    .Q(\am_sdr0.spi0.SCK_qqq ));
 sg13g2_dfrbp_1 _14735_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net335),
    .D(_01106_),
    .Q_N(_05808_),
    .Q(\am_sdr0.spi0.SCK_qq ));
 sg13g2_dfrbp_1 _14736_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net331),
    .D(_01107_),
    .Q_N(_05807_),
    .Q(\am_sdr0.nco0.phase_inc[0] ));
 sg13g2_dfrbp_1 _14737_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net323),
    .D(_01108_),
    .Q_N(_05806_),
    .Q(\am_sdr0.nco0.phase_inc[1] ));
 sg13g2_dfrbp_1 _14738_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net315),
    .D(net1272),
    .Q_N(_05805_),
    .Q(\am_sdr0.nco0.phase_inc[2] ));
 sg13g2_dfrbp_1 _14739_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net307),
    .D(_01110_),
    .Q_N(_05804_),
    .Q(\am_sdr0.nco0.phase_inc[3] ));
 sg13g2_dfrbp_1 _14740_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net299),
    .D(net1292),
    .Q_N(_05803_),
    .Q(\am_sdr0.nco0.phase_inc[4] ));
 sg13g2_dfrbp_1 _14741_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net291),
    .D(_01112_),
    .Q_N(_05802_),
    .Q(\am_sdr0.nco0.phase_inc[5] ));
 sg13g2_dfrbp_1 _14742_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net283),
    .D(_01113_),
    .Q_N(_05801_),
    .Q(\am_sdr0.nco0.phase_inc[6] ));
 sg13g2_dfrbp_1 _14743_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net275),
    .D(_01114_),
    .Q_N(_05800_),
    .Q(\am_sdr0.nco0.phase_inc[7] ));
 sg13g2_dfrbp_1 _14744_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net267),
    .D(_01115_),
    .Q_N(_05799_),
    .Q(\am_sdr0.nco0.phase_inc[8] ));
 sg13g2_dfrbp_1 _14745_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net259),
    .D(_01116_),
    .Q_N(_05798_),
    .Q(\am_sdr0.nco0.phase_inc[9] ));
 sg13g2_dfrbp_1 _14746_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net251),
    .D(_01117_),
    .Q_N(_05797_),
    .Q(\am_sdr0.nco0.phase_inc[10] ));
 sg13g2_dfrbp_1 _14747_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net243),
    .D(_01118_),
    .Q_N(_05796_),
    .Q(\am_sdr0.nco0.phase_inc[11] ));
 sg13g2_dfrbp_1 _14748_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net235),
    .D(_01119_),
    .Q_N(_05795_),
    .Q(\am_sdr0.nco0.phase_inc[12] ));
 sg13g2_dfrbp_1 _14749_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net186),
    .D(_01120_),
    .Q_N(_05794_),
    .Q(\am_sdr0.nco0.phase_inc[13] ));
 sg13g2_dfrbp_1 _14750_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net178),
    .D(net1346),
    .Q_N(_05793_),
    .Q(\am_sdr0.nco0.phase_inc[14] ));
 sg13g2_dfrbp_1 _14751_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net170),
    .D(net1421),
    .Q_N(_05792_),
    .Q(\am_sdr0.nco0.phase_inc[15] ));
 sg13g2_dfrbp_1 _14752_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net162),
    .D(_01123_),
    .Q_N(_05791_),
    .Q(\am_sdr0.nco0.phase_inc[16] ));
 sg13g2_dfrbp_1 _14753_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net154),
    .D(_01124_),
    .Q_N(_05790_),
    .Q(\am_sdr0.nco0.phase_inc[17] ));
 sg13g2_dfrbp_1 _14754_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net146),
    .D(net2044),
    .Q_N(_05789_),
    .Q(\am_sdr0.nco0.phase_inc[18] ));
 sg13g2_dfrbp_1 _14755_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net138),
    .D(_01126_),
    .Q_N(_05788_),
    .Q(\am_sdr0.nco0.phase_inc[19] ));
 sg13g2_dfrbp_1 _14756_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net127),
    .D(_01127_),
    .Q_N(_05787_),
    .Q(\am_sdr0.nco0.phase_inc[20] ));
 sg13g2_dfrbp_1 _14757_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net71),
    .D(_01128_),
    .Q_N(_05786_),
    .Q(\am_sdr0.nco0.phase_inc[21] ));
 sg13g2_dfrbp_1 _14758_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net55),
    .D(_01129_),
    .Q_N(_05785_),
    .Q(\am_sdr0.nco0.phase_inc[22] ));
 sg13g2_dfrbp_1 _14759_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net39),
    .D(_01130_),
    .Q_N(_05784_),
    .Q(\am_sdr0.nco0.phase_inc[23] ));
 sg13g2_dfrbp_1 _14760_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1153),
    .D(_01131_),
    .Q_N(_05783_),
    .Q(\am_sdr0.nco0.phase_inc[24] ));
 sg13g2_dfrbp_1 _14761_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1113),
    .D(_01132_),
    .Q_N(_05782_),
    .Q(\am_sdr0.nco0.phase_inc[25] ));
 sg13g2_dfrbp_1 _14762_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1096),
    .D(net1405),
    .Q_N(_05781_),
    .Q(\am_sdr0.spi0.state[0] ));
 sg13g2_dfrbp_1 _14763_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1080),
    .D(_01134_),
    .Q_N(_05780_),
    .Q(\am_sdr0.spi0.state[1] ));
 sg13g2_dfrbp_1 _14764_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1027),
    .D(_01135_),
    .Q_N(_05779_),
    .Q(\am_sdr0.gain_spi[0] ));
 sg13g2_dfrbp_1 _14765_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1011),
    .D(_01136_),
    .Q_N(_05778_),
    .Q(\am_sdr0.gain_spi[1] ));
 sg13g2_dfrbp_1 _14766_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net995),
    .D(_01137_),
    .Q_N(_00046_),
    .Q(\am_sdr0.gain_spi[2] ));
 sg13g2_dfrbp_1 _14767_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net979),
    .D(_01138_),
    .Q_N(_05777_),
    .Q(\am_sdr0.nco0.phase[0] ));
 sg13g2_dfrbp_1 _14768_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net971),
    .D(_01139_),
    .Q_N(_05776_),
    .Q(\am_sdr0.nco0.phase[1] ));
 sg13g2_dfrbp_1 _14769_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net963),
    .D(net3067),
    .Q_N(_05775_),
    .Q(\am_sdr0.nco0.phase[2] ));
 sg13g2_dfrbp_1 _14770_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net955),
    .D(_01141_),
    .Q_N(_05774_),
    .Q(\am_sdr0.nco0.phase[3] ));
 sg13g2_dfrbp_1 _14771_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net947),
    .D(_01142_),
    .Q_N(_05773_),
    .Q(\am_sdr0.nco0.phase[4] ));
 sg13g2_dfrbp_1 _14772_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net939),
    .D(net3110),
    .Q_N(_05772_),
    .Q(\am_sdr0.nco0.phase[5] ));
 sg13g2_dfrbp_1 _14773_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net931),
    .D(net3096),
    .Q_N(_05771_),
    .Q(\am_sdr0.nco0.phase[6] ));
 sg13g2_dfrbp_1 _14774_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net355),
    .D(_01145_),
    .Q_N(_05770_),
    .Q(\am_sdr0.nco0.phase[7] ));
 sg13g2_dfrbp_1 _14775_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net347),
    .D(net3083),
    .Q_N(_05769_),
    .Q(\am_sdr0.nco0.phase[8] ));
 sg13g2_dfrbp_1 _14776_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net327),
    .D(_01147_),
    .Q_N(_05768_),
    .Q(\am_sdr0.nco0.phase[9] ));
 sg13g2_dfrbp_1 _14777_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net319),
    .D(_01148_),
    .Q_N(_05767_),
    .Q(\am_sdr0.nco0.phase[10] ));
 sg13g2_dfrbp_1 _14778_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net311),
    .D(_01149_),
    .Q_N(_05766_),
    .Q(\am_sdr0.nco0.phase[11] ));
 sg13g2_dfrbp_1 _14779_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net303),
    .D(_01150_),
    .Q_N(_05765_),
    .Q(\am_sdr0.nco0.phase[12] ));
 sg13g2_dfrbp_1 _14780_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net295),
    .D(net3211),
    .Q_N(_05764_),
    .Q(\am_sdr0.nco0.phase[13] ));
 sg13g2_dfrbp_1 _14781_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net287),
    .D(net3117),
    .Q_N(_05763_),
    .Q(\am_sdr0.nco0.phase[14] ));
 sg13g2_dfrbp_1 _14782_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net279),
    .D(net3194),
    .Q_N(_05762_),
    .Q(\am_sdr0.nco0.phase[15] ));
 sg13g2_dfrbp_1 _14783_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net271),
    .D(_01154_),
    .Q_N(_05761_),
    .Q(\am_sdr0.nco0.phase[16] ));
 sg13g2_dfrbp_1 _14784_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net263),
    .D(_01155_),
    .Q_N(_05760_),
    .Q(\am_sdr0.nco0.phase[17] ));
 sg13g2_dfrbp_1 _14785_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net255),
    .D(net3033),
    .Q_N(_05759_),
    .Q(\am_sdr0.nco0.phase[18] ));
 sg13g2_dfrbp_1 _14786_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net247),
    .D(net3190),
    .Q_N(_05758_),
    .Q(\am_sdr0.nco0.phase[19] ));
 sg13g2_dfrbp_1 _14787_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net239),
    .D(_01158_),
    .Q_N(_05757_),
    .Q(\am_sdr0.nco0.phase[20] ));
 sg13g2_dfrbp_1 _14788_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net190),
    .D(_01159_),
    .Q_N(_05756_),
    .Q(\am_sdr0.nco0.phase[21] ));
 sg13g2_dfrbp_1 _14789_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net182),
    .D(_01160_),
    .Q_N(_00039_),
    .Q(\am_sdr0.nco0.phase[22] ));
 sg13g2_dfrbp_1 _14790_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net174),
    .D(_01161_),
    .Q_N(_00038_),
    .Q(\am_sdr0.nco0.phase[23] ));
 sg13g2_dfrbp_1 _14791_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net166),
    .D(_01162_),
    .Q_N(_00037_),
    .Q(\am_sdr0.nco0.phase[24] ));
 sg13g2_dfrbp_1 _14792_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net158),
    .D(_01163_),
    .Q_N(_05755_),
    .Q(\am_sdr0.nco0.phase[25] ));
 sg13g2_dfrbp_1 _14793_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net150),
    .D(_01164_),
    .Q_N(_05754_),
    .Q(\am_sdr0.spi0.CS_q ));
 sg13g2_dfrbp_1 _14794_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net142),
    .D(_01165_),
    .Q_N(_05753_),
    .Q(\am_sdr0.spi0.CS_qq ));
 sg13g2_dfrbp_1 _14795_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net134),
    .D(_01166_),
    .Q_N(_05752_),
    .Q(\am_sdr0.spi0.CS_qqq ));
 sg13g2_dfrbp_1 _14796_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net79),
    .D(_01167_),
    .Q_N(_05751_),
    .Q(\am_sdr0.spi0.SCK_q ));
 sg13g2_dfrbp_1 _14797_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net63),
    .D(net2482),
    .Q_N(_05750_),
    .Q(PWM_OUT));
 sg13g2_dfrbp_1 _14798_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net47),
    .D(_01169_),
    .Q_N(_05749_),
    .Q(\am_sdr0.am0.demod_out[8] ));
 sg13g2_dfrbp_1 _14799_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1121),
    .D(_01170_),
    .Q_N(_05748_),
    .Q(\am_sdr0.am0.demod_out[9] ));
 sg13g2_dfrbp_1 _14800_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1088),
    .D(_01171_),
    .Q_N(_05747_),
    .Q(\am_sdr0.am0.demod_out[10] ));
 sg13g2_dfrbp_1 _14801_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1019),
    .D(_01172_),
    .Q_N(_05746_),
    .Q(\am_sdr0.am0.demod_out[11] ));
 sg13g2_dfrbp_1 _14802_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net987),
    .D(_01173_),
    .Q_N(_05745_),
    .Q(\am_sdr0.am0.demod_out[12] ));
 sg13g2_dfrbp_1 _14803_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1104),
    .D(_01174_),
    .Q_N(_05744_),
    .Q(\am_sdr0.am0.demod_out[13] ));
 sg13g2_dfrbp_1 _14804_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1003),
    .D(_01175_),
    .Q_N(_05743_),
    .Q(\am_sdr0.am0.demod_out[14] ));
 sg13g2_dfrbp_1 _14805_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1072),
    .D(_01176_),
    .Q_N(_05742_),
    .Q(\am_sdr0.am0.demod_out[15] ));
 sg13g2_tiehi _13676__28 (.L_HI(net28));
 sg13g2_tiehi _13670__29 (.L_HI(net29));
 sg13g2_tiehi _13671__30 (.L_HI(net30));
 sg13g2_tiehi _13672__31 (.L_HI(net31));
 sg13g2_tiehi _13673__32 (.L_HI(net32));
 sg13g2_tiehi _13674__33 (.L_HI(net33));
 sg13g2_tiehi _13731__34 (.L_HI(net34));
 sg13g2_tiehi _14596__35 (.L_HI(net35));
 sg13g2_tiehi _13730__36 (.L_HI(net36));
 sg13g2_tiehi _14322__37 (.L_HI(net37));
 sg13g2_tiehi _13729__38 (.L_HI(net38));
 sg13g2_tiehi _14759__39 (.L_HI(net39));
 sg13g2_tiehi _13728__40 (.L_HI(net40));
 sg13g2_tiehi _14321__41 (.L_HI(net41));
 sg13g2_tiehi _13727__42 (.L_HI(net42));
 sg13g2_tiehi _14595__43 (.L_HI(net43));
 sg13g2_tiehi _13726__44 (.L_HI(net44));
 sg13g2_tiehi _14320__45 (.L_HI(net45));
 sg13g2_tiehi _13725__46 (.L_HI(net46));
 sg13g2_tiehi _14798__47 (.L_HI(net47));
 sg13g2_tiehi _13724__48 (.L_HI(net48));
 sg13g2_tiehi _14319__49 (.L_HI(net49));
 sg13g2_tiehi _13723__50 (.L_HI(net50));
 sg13g2_tiehi _14594__51 (.L_HI(net51));
 sg13g2_tiehi _13722__52 (.L_HI(net52));
 sg13g2_tiehi _14318__53 (.L_HI(net53));
 sg13g2_tiehi _13721__54 (.L_HI(net54));
 sg13g2_tiehi _14758__55 (.L_HI(net55));
 sg13g2_tiehi _13720__56 (.L_HI(net56));
 sg13g2_tiehi _14317__57 (.L_HI(net57));
 sg13g2_tiehi _13719__58 (.L_HI(net58));
 sg13g2_tiehi _14593__59 (.L_HI(net59));
 sg13g2_tiehi _13718__60 (.L_HI(net60));
 sg13g2_tiehi _14316__61 (.L_HI(net61));
 sg13g2_tiehi _13717__62 (.L_HI(net62));
 sg13g2_tiehi _14797__63 (.L_HI(net63));
 sg13g2_tiehi _13716__64 (.L_HI(net64));
 sg13g2_tiehi _14315__65 (.L_HI(net65));
 sg13g2_tiehi _13715__66 (.L_HI(net66));
 sg13g2_tiehi _14592__67 (.L_HI(net67));
 sg13g2_tiehi _13714__68 (.L_HI(net68));
 sg13g2_tiehi _14314__69 (.L_HI(net69));
 sg13g2_tiehi _13713__70 (.L_HI(net70));
 sg13g2_tiehi _14757__71 (.L_HI(net71));
 sg13g2_tiehi _13712__72 (.L_HI(net72));
 sg13g2_tiehi _14313__73 (.L_HI(net73));
 sg13g2_tiehi _13711__74 (.L_HI(net74));
 sg13g2_tiehi _14591__75 (.L_HI(net75));
 sg13g2_tiehi _13710__76 (.L_HI(net76));
 sg13g2_tiehi _14312__77 (.L_HI(net77));
 sg13g2_tiehi _13709__78 (.L_HI(net78));
 sg13g2_tiehi _14796__79 (.L_HI(net79));
 sg13g2_tiehi _13708__80 (.L_HI(net80));
 sg13g2_tiehi _14311__81 (.L_HI(net81));
 sg13g2_tiehi _13707__82 (.L_HI(net82));
 sg13g2_tiehi _14590__83 (.L_HI(net83));
 sg13g2_tiehi _13706__84 (.L_HI(net84));
 sg13g2_tiehi _13705__85 (.L_HI(net85));
 sg13g2_tiehi _13704__86 (.L_HI(net86));
 sg13g2_tiehi _13703__87 (.L_HI(net87));
 sg13g2_tiehi _13702__88 (.L_HI(net88));
 sg13g2_tiehi _13701__89 (.L_HI(net89));
 sg13g2_tiehi _13700__90 (.L_HI(net90));
 sg13g2_tiehi _13699__91 (.L_HI(net91));
 sg13g2_tiehi _13698__92 (.L_HI(net92));
 sg13g2_tiehi _13675__93 (.L_HI(net93));
 sg13g2_tiehi _13735__94 (.L_HI(net94));
 sg13g2_tiehi _13736__95 (.L_HI(net95));
 sg13g2_tiehi _13737__96 (.L_HI(net96));
 sg13g2_tiehi _13738__97 (.L_HI(net97));
 sg13g2_tiehi _13739__98 (.L_HI(net98));
 sg13g2_tiehi _13740__99 (.L_HI(net99));
 sg13g2_tiehi _13697__100 (.L_HI(net100));
 sg13g2_tiehi _13696__101 (.L_HI(net101));
 sg13g2_tiehi _13695__102 (.L_HI(net102));
 sg13g2_tiehi _13694__103 (.L_HI(net103));
 sg13g2_tiehi _13693__104 (.L_HI(net104));
 sg13g2_tiehi _13692__105 (.L_HI(net105));
 sg13g2_tiehi _13691__106 (.L_HI(net106));
 sg13g2_tiehi _13690__107 (.L_HI(net107));
 sg13g2_tiehi _13689__108 (.L_HI(net108));
 sg13g2_tiehi _13688__109 (.L_HI(net109));
 sg13g2_tiehi _13687__110 (.L_HI(net110));
 sg13g2_tiehi _13686__111 (.L_HI(net111));
 sg13g2_tiehi _13685__112 (.L_HI(net112));
 sg13g2_tiehi _13684__113 (.L_HI(net113));
 sg13g2_tiehi _13683__114 (.L_HI(net114));
 sg13g2_tiehi _13682__115 (.L_HI(net115));
 sg13g2_tiehi _13741__116 (.L_HI(net116));
 sg13g2_tiehi _13758__117 (.L_HI(net117));
 sg13g2_tiehi _13759__118 (.L_HI(net118));
 sg13g2_tiehi _13760__119 (.L_HI(net119));
 sg13g2_tiehi _13761__120 (.L_HI(net120));
 sg13g2_tiehi _13762__121 (.L_HI(net121));
 sg13g2_tiehi _13763__122 (.L_HI(net122));
 sg13g2_tiehi _13764__123 (.L_HI(net123));
 sg13g2_tiehi _13681__124 (.L_HI(net124));
 sg13g2_tiehi _14310__125 (.L_HI(net125));
 sg13g2_tiehi _13680__126 (.L_HI(net126));
 sg13g2_tiehi _14756__127 (.L_HI(net127));
 sg13g2_tiehi _13679__128 (.L_HI(net128));
 sg13g2_tiehi _14309__129 (.L_HI(net129));
 sg13g2_tiehi _13678__130 (.L_HI(net130));
 sg13g2_tiehi _14589__131 (.L_HI(net131));
 sg13g2_tiehi _13677__132 (.L_HI(net132));
 sg13g2_tiehi _14308__133 (.L_HI(net133));
 sg13g2_tiehi _14795__134 (.L_HI(net134));
 sg13g2_tiehi _14307__135 (.L_HI(net135));
 sg13g2_tiehi _14588__136 (.L_HI(net136));
 sg13g2_tiehi _14306__137 (.L_HI(net137));
 sg13g2_tiehi _14755__138 (.L_HI(net138));
 sg13g2_tiehi _14305__139 (.L_HI(net139));
 sg13g2_tiehi _14587__140 (.L_HI(net140));
 sg13g2_tiehi _14304__141 (.L_HI(net141));
 sg13g2_tiehi _14794__142 (.L_HI(net142));
 sg13g2_tiehi _14303__143 (.L_HI(net143));
 sg13g2_tiehi _14586__144 (.L_HI(net144));
 sg13g2_tiehi _14302__145 (.L_HI(net145));
 sg13g2_tiehi _14754__146 (.L_HI(net146));
 sg13g2_tiehi _14301__147 (.L_HI(net147));
 sg13g2_tiehi _14585__148 (.L_HI(net148));
 sg13g2_tiehi _14300__149 (.L_HI(net149));
 sg13g2_tiehi _14793__150 (.L_HI(net150));
 sg13g2_tiehi _14299__151 (.L_HI(net151));
 sg13g2_tiehi _14584__152 (.L_HI(net152));
 sg13g2_tiehi _14298__153 (.L_HI(net153));
 sg13g2_tiehi _14753__154 (.L_HI(net154));
 sg13g2_tiehi _14297__155 (.L_HI(net155));
 sg13g2_tiehi _14583__156 (.L_HI(net156));
 sg13g2_tiehi _14296__157 (.L_HI(net157));
 sg13g2_tiehi _14792__158 (.L_HI(net158));
 sg13g2_tiehi _14295__159 (.L_HI(net159));
 sg13g2_tiehi _14582__160 (.L_HI(net160));
 sg13g2_tiehi _14294__161 (.L_HI(net161));
 sg13g2_tiehi _14752__162 (.L_HI(net162));
 sg13g2_tiehi _14293__163 (.L_HI(net163));
 sg13g2_tiehi _14581__164 (.L_HI(net164));
 sg13g2_tiehi _14292__165 (.L_HI(net165));
 sg13g2_tiehi _14791__166 (.L_HI(net166));
 sg13g2_tiehi _14291__167 (.L_HI(net167));
 sg13g2_tiehi _14580__168 (.L_HI(net168));
 sg13g2_tiehi _14290__169 (.L_HI(net169));
 sg13g2_tiehi _14751__170 (.L_HI(net170));
 sg13g2_tiehi _14289__171 (.L_HI(net171));
 sg13g2_tiehi _14579__172 (.L_HI(net172));
 sg13g2_tiehi _14288__173 (.L_HI(net173));
 sg13g2_tiehi _14790__174 (.L_HI(net174));
 sg13g2_tiehi _14287__175 (.L_HI(net175));
 sg13g2_tiehi _14578__176 (.L_HI(net176));
 sg13g2_tiehi _14286__177 (.L_HI(net177));
 sg13g2_tiehi _14750__178 (.L_HI(net178));
 sg13g2_tiehi _14285__179 (.L_HI(net179));
 sg13g2_tiehi _14577__180 (.L_HI(net180));
 sg13g2_tiehi _14284__181 (.L_HI(net181));
 sg13g2_tiehi _14789__182 (.L_HI(net182));
 sg13g2_tiehi _14283__183 (.L_HI(net183));
 sg13g2_tiehi _14576__184 (.L_HI(net184));
 sg13g2_tiehi _14282__185 (.L_HI(net185));
 sg13g2_tiehi _14749__186 (.L_HI(net186));
 sg13g2_tiehi _14281__187 (.L_HI(net187));
 sg13g2_tiehi _14575__188 (.L_HI(net188));
 sg13g2_tiehi _14280__189 (.L_HI(net189));
 sg13g2_tiehi _14788__190 (.L_HI(net190));
 sg13g2_tiehi _14279__191 (.L_HI(net191));
 sg13g2_tiehi _14574__192 (.L_HI(net192));
 sg13g2_tiehi _14278__193 (.L_HI(net193));
 sg13g2_tiehi _14277__194 (.L_HI(net194));
 sg13g2_tiehi _14276__195 (.L_HI(net195));
 sg13g2_tiehi _14275__196 (.L_HI(net196));
 sg13g2_tiehi _14274__197 (.L_HI(net197));
 sg13g2_tiehi _14273__198 (.L_HI(net198));
 sg13g2_tiehi _14272__199 (.L_HI(net199));
 sg13g2_tiehi _14271__200 (.L_HI(net200));
 sg13g2_tiehi _14270__201 (.L_HI(net201));
 sg13g2_tiehi _14269__202 (.L_HI(net202));
 sg13g2_tiehi _14268__203 (.L_HI(net203));
 sg13g2_tiehi _14267__204 (.L_HI(net204));
 sg13g2_tiehi _14266__205 (.L_HI(net205));
 sg13g2_tiehi _14265__206 (.L_HI(net206));
 sg13g2_tiehi _14264__207 (.L_HI(net207));
 sg13g2_tiehi _14263__208 (.L_HI(net208));
 sg13g2_tiehi _14262__209 (.L_HI(net209));
 sg13g2_tiehi _14261__210 (.L_HI(net210));
 sg13g2_tiehi _14260__211 (.L_HI(net211));
 sg13g2_tiehi _14259__212 (.L_HI(net212));
 sg13g2_tiehi _14258__213 (.L_HI(net213));
 sg13g2_tiehi _14257__214 (.L_HI(net214));
 sg13g2_tiehi _14256__215 (.L_HI(net215));
 sg13g2_tiehi _14255__216 (.L_HI(net216));
 sg13g2_tiehi _14254__217 (.L_HI(net217));
 sg13g2_tiehi _14253__218 (.L_HI(net218));
 sg13g2_tiehi _14252__219 (.L_HI(net219));
 sg13g2_tiehi _14251__220 (.L_HI(net220));
 sg13g2_tiehi _14250__221 (.L_HI(net221));
 sg13g2_tiehi _14249__222 (.L_HI(net222));
 sg13g2_tiehi _14248__223 (.L_HI(net223));
 sg13g2_tiehi _14247__224 (.L_HI(net224));
 sg13g2_tiehi _14246__225 (.L_HI(net225));
 sg13g2_tiehi _14245__226 (.L_HI(net226));
 sg13g2_tiehi _14244__227 (.L_HI(net227));
 sg13g2_tiehi _14243__228 (.L_HI(net228));
 sg13g2_tiehi _14242__229 (.L_HI(net229));
 sg13g2_tiehi _14241__230 (.L_HI(net230));
 sg13g2_tiehi _14240__231 (.L_HI(net231));
 sg13g2_tiehi _14239__232 (.L_HI(net232));
 sg13g2_tiehi _14238__233 (.L_HI(net233));
 sg13g2_tiehi _14237__234 (.L_HI(net234));
 sg13g2_tiehi _14748__235 (.L_HI(net235));
 sg13g2_tiehi _14236__236 (.L_HI(net236));
 sg13g2_tiehi _14573__237 (.L_HI(net237));
 sg13g2_tiehi _14235__238 (.L_HI(net238));
 sg13g2_tiehi _14787__239 (.L_HI(net239));
 sg13g2_tiehi _14234__240 (.L_HI(net240));
 sg13g2_tiehi _14572__241 (.L_HI(net241));
 sg13g2_tiehi _14233__242 (.L_HI(net242));
 sg13g2_tiehi _14747__243 (.L_HI(net243));
 sg13g2_tiehi _14232__244 (.L_HI(net244));
 sg13g2_tiehi _14571__245 (.L_HI(net245));
 sg13g2_tiehi _14231__246 (.L_HI(net246));
 sg13g2_tiehi _14786__247 (.L_HI(net247));
 sg13g2_tiehi _14230__248 (.L_HI(net248));
 sg13g2_tiehi _14570__249 (.L_HI(net249));
 sg13g2_tiehi _14229__250 (.L_HI(net250));
 sg13g2_tiehi _14746__251 (.L_HI(net251));
 sg13g2_tiehi _14228__252 (.L_HI(net252));
 sg13g2_tiehi _14569__253 (.L_HI(net253));
 sg13g2_tiehi _14227__254 (.L_HI(net254));
 sg13g2_tiehi _14785__255 (.L_HI(net255));
 sg13g2_tiehi _14226__256 (.L_HI(net256));
 sg13g2_tiehi _14568__257 (.L_HI(net257));
 sg13g2_tiehi _14225__258 (.L_HI(net258));
 sg13g2_tiehi _14745__259 (.L_HI(net259));
 sg13g2_tiehi _14224__260 (.L_HI(net260));
 sg13g2_tiehi _14567__261 (.L_HI(net261));
 sg13g2_tiehi _14223__262 (.L_HI(net262));
 sg13g2_tiehi _14784__263 (.L_HI(net263));
 sg13g2_tiehi _14222__264 (.L_HI(net264));
 sg13g2_tiehi _14566__265 (.L_HI(net265));
 sg13g2_tiehi _14221__266 (.L_HI(net266));
 sg13g2_tiehi _14744__267 (.L_HI(net267));
 sg13g2_tiehi _14220__268 (.L_HI(net268));
 sg13g2_tiehi _14565__269 (.L_HI(net269));
 sg13g2_tiehi _14219__270 (.L_HI(net270));
 sg13g2_tiehi _14783__271 (.L_HI(net271));
 sg13g2_tiehi _14218__272 (.L_HI(net272));
 sg13g2_tiehi _14564__273 (.L_HI(net273));
 sg13g2_tiehi _14217__274 (.L_HI(net274));
 sg13g2_tiehi _14743__275 (.L_HI(net275));
 sg13g2_tiehi _14216__276 (.L_HI(net276));
 sg13g2_tiehi _14563__277 (.L_HI(net277));
 sg13g2_tiehi _14215__278 (.L_HI(net278));
 sg13g2_tiehi _14782__279 (.L_HI(net279));
 sg13g2_tiehi _14214__280 (.L_HI(net280));
 sg13g2_tiehi _14562__281 (.L_HI(net281));
 sg13g2_tiehi _14213__282 (.L_HI(net282));
 sg13g2_tiehi _14742__283 (.L_HI(net283));
 sg13g2_tiehi _14212__284 (.L_HI(net284));
 sg13g2_tiehi _14561__285 (.L_HI(net285));
 sg13g2_tiehi _14211__286 (.L_HI(net286));
 sg13g2_tiehi _14781__287 (.L_HI(net287));
 sg13g2_tiehi _14210__288 (.L_HI(net288));
 sg13g2_tiehi _14560__289 (.L_HI(net289));
 sg13g2_tiehi _14209__290 (.L_HI(net290));
 sg13g2_tiehi _14741__291 (.L_HI(net291));
 sg13g2_tiehi _14208__292 (.L_HI(net292));
 sg13g2_tiehi _14559__293 (.L_HI(net293));
 sg13g2_tiehi _14207__294 (.L_HI(net294));
 sg13g2_tiehi _14780__295 (.L_HI(net295));
 sg13g2_tiehi _14206__296 (.L_HI(net296));
 sg13g2_tiehi _14558__297 (.L_HI(net297));
 sg13g2_tiehi _14205__298 (.L_HI(net298));
 sg13g2_tiehi _14740__299 (.L_HI(net299));
 sg13g2_tiehi _14204__300 (.L_HI(net300));
 sg13g2_tiehi _14557__301 (.L_HI(net301));
 sg13g2_tiehi _14203__302 (.L_HI(net302));
 sg13g2_tiehi _14779__303 (.L_HI(net303));
 sg13g2_tiehi _14202__304 (.L_HI(net304));
 sg13g2_tiehi _14556__305 (.L_HI(net305));
 sg13g2_tiehi _14201__306 (.L_HI(net306));
 sg13g2_tiehi _14739__307 (.L_HI(net307));
 sg13g2_tiehi _14200__308 (.L_HI(net308));
 sg13g2_tiehi _14555__309 (.L_HI(net309));
 sg13g2_tiehi _14199__310 (.L_HI(net310));
 sg13g2_tiehi _14778__311 (.L_HI(net311));
 sg13g2_tiehi _14198__312 (.L_HI(net312));
 sg13g2_tiehi _14554__313 (.L_HI(net313));
 sg13g2_tiehi _14197__314 (.L_HI(net314));
 sg13g2_tiehi _14738__315 (.L_HI(net315));
 sg13g2_tiehi _14196__316 (.L_HI(net316));
 sg13g2_tiehi _14553__317 (.L_HI(net317));
 sg13g2_tiehi _14195__318 (.L_HI(net318));
 sg13g2_tiehi _14777__319 (.L_HI(net319));
 sg13g2_tiehi _14194__320 (.L_HI(net320));
 sg13g2_tiehi _14552__321 (.L_HI(net321));
 sg13g2_tiehi _14193__322 (.L_HI(net322));
 sg13g2_tiehi _14737__323 (.L_HI(net323));
 sg13g2_tiehi _14192__324 (.L_HI(net324));
 sg13g2_tiehi _14551__325 (.L_HI(net325));
 sg13g2_tiehi _14191__326 (.L_HI(net326));
 sg13g2_tiehi _14776__327 (.L_HI(net327));
 sg13g2_tiehi _14190__328 (.L_HI(net328));
 sg13g2_tiehi _14550__329 (.L_HI(net329));
 sg13g2_tiehi _14189__330 (.L_HI(net330));
 sg13g2_tiehi _14736__331 (.L_HI(net331));
 sg13g2_tiehi _14188__332 (.L_HI(net332));
 sg13g2_tiehi _14549__333 (.L_HI(net333));
 sg13g2_tiehi _14187__334 (.L_HI(net334));
 sg13g2_tiehi _14735__335 (.L_HI(net335));
 sg13g2_tiehi _14186__336 (.L_HI(net336));
 sg13g2_tiehi _14548__337 (.L_HI(net337));
 sg13g2_tiehi _14185__338 (.L_HI(net338));
 sg13g2_tiehi _14734__339 (.L_HI(net339));
 sg13g2_tiehi _14184__340 (.L_HI(net340));
 sg13g2_tiehi _14547__341 (.L_HI(net341));
 sg13g2_tiehi _14183__342 (.L_HI(net342));
 sg13g2_tiehi _14733__343 (.L_HI(net343));
 sg13g2_tiehi _14182__344 (.L_HI(net344));
 sg13g2_tiehi _14546__345 (.L_HI(net345));
 sg13g2_tiehi _14181__346 (.L_HI(net346));
 sg13g2_tiehi _14775__347 (.L_HI(net347));
 sg13g2_tiehi _14180__348 (.L_HI(net348));
 sg13g2_tiehi _14545__349 (.L_HI(net349));
 sg13g2_tiehi _14179__350 (.L_HI(net350));
 sg13g2_tiehi _14732__351 (.L_HI(net351));
 sg13g2_tiehi _14178__352 (.L_HI(net352));
 sg13g2_tiehi _14544__353 (.L_HI(net353));
 sg13g2_tiehi _14177__354 (.L_HI(net354));
 sg13g2_tiehi _14774__355 (.L_HI(net355));
 sg13g2_tiehi _14176__356 (.L_HI(net356));
 sg13g2_tiehi _14543__357 (.L_HI(net357));
 sg13g2_tiehi _14175__358 (.L_HI(net358));
 sg13g2_tiehi _14731__359 (.L_HI(net359));
 sg13g2_tiehi _14174__360 (.L_HI(net360));
 sg13g2_tiehi _14542__361 (.L_HI(net361));
 sg13g2_tiehi _14173__362 (.L_HI(net362));
 sg13g2_tiehi _14730__363 (.L_HI(net363));
 sg13g2_tiehi _14172__364 (.L_HI(net364));
 sg13g2_tiehi _14541__365 (.L_HI(net365));
 sg13g2_tiehi _14171__366 (.L_HI(net366));
 sg13g2_tiehi _14729__367 (.L_HI(net367));
 sg13g2_tiehi _14170__368 (.L_HI(net368));
 sg13g2_tiehi _14540__369 (.L_HI(net369));
 sg13g2_tiehi _14169__370 (.L_HI(net370));
 sg13g2_tiehi _14728__371 (.L_HI(net371));
 sg13g2_tiehi _14168__372 (.L_HI(net372));
 sg13g2_tiehi _14539__373 (.L_HI(net373));
 sg13g2_tiehi _14167__374 (.L_HI(net374));
 sg13g2_tiehi _14727__375 (.L_HI(net375));
 sg13g2_tiehi _14166__376 (.L_HI(net376));
 sg13g2_tiehi _14538__377 (.L_HI(net377));
 sg13g2_tiehi _14165__378 (.L_HI(net378));
 sg13g2_tiehi _14726__379 (.L_HI(net379));
 sg13g2_tiehi _14164__380 (.L_HI(net380));
 sg13g2_tiehi _14537__381 (.L_HI(net381));
 sg13g2_tiehi _14163__382 (.L_HI(net382));
 sg13g2_tiehi _14725__383 (.L_HI(net383));
 sg13g2_tiehi _14162__384 (.L_HI(net384));
 sg13g2_tiehi _14536__385 (.L_HI(net385));
 sg13g2_tiehi _14161__386 (.L_HI(net386));
 sg13g2_tiehi _14724__387 (.L_HI(net387));
 sg13g2_tiehi _14160__388 (.L_HI(net388));
 sg13g2_tiehi _14535__389 (.L_HI(net389));
 sg13g2_tiehi _14159__390 (.L_HI(net390));
 sg13g2_tiehi _14723__391 (.L_HI(net391));
 sg13g2_tiehi _14158__392 (.L_HI(net392));
 sg13g2_tiehi _14534__393 (.L_HI(net393));
 sg13g2_tiehi _14157__394 (.L_HI(net394));
 sg13g2_tiehi _14722__395 (.L_HI(net395));
 sg13g2_tiehi _14156__396 (.L_HI(net396));
 sg13g2_tiehi _14533__397 (.L_HI(net397));
 sg13g2_tiehi _14155__398 (.L_HI(net398));
 sg13g2_tiehi _14721__399 (.L_HI(net399));
 sg13g2_tiehi _14154__400 (.L_HI(net400));
 sg13g2_tiehi _14532__401 (.L_HI(net401));
 sg13g2_tiehi _14153__402 (.L_HI(net402));
 sg13g2_tiehi _14720__403 (.L_HI(net403));
 sg13g2_tiehi _14152__404 (.L_HI(net404));
 sg13g2_tiehi _14531__405 (.L_HI(net405));
 sg13g2_tiehi _14151__406 (.L_HI(net406));
 sg13g2_tiehi _14719__407 (.L_HI(net407));
 sg13g2_tiehi _14150__408 (.L_HI(net408));
 sg13g2_tiehi _14530__409 (.L_HI(net409));
 sg13g2_tiehi _14149__410 (.L_HI(net410));
 sg13g2_tiehi _14718__411 (.L_HI(net411));
 sg13g2_tiehi _14148__412 (.L_HI(net412));
 sg13g2_tiehi _14529__413 (.L_HI(net413));
 sg13g2_tiehi _14147__414 (.L_HI(net414));
 sg13g2_tiehi _14717__415 (.L_HI(net415));
 sg13g2_tiehi _14146__416 (.L_HI(net416));
 sg13g2_tiehi _14528__417 (.L_HI(net417));
 sg13g2_tiehi _14145__418 (.L_HI(net418));
 sg13g2_tiehi _14716__419 (.L_HI(net419));
 sg13g2_tiehi _14144__420 (.L_HI(net420));
 sg13g2_tiehi _14527__421 (.L_HI(net421));
 sg13g2_tiehi _14143__422 (.L_HI(net422));
 sg13g2_tiehi _14715__423 (.L_HI(net423));
 sg13g2_tiehi _14142__424 (.L_HI(net424));
 sg13g2_tiehi _14526__425 (.L_HI(net425));
 sg13g2_tiehi _14141__426 (.L_HI(net426));
 sg13g2_tiehi _14714__427 (.L_HI(net427));
 sg13g2_tiehi _14140__428 (.L_HI(net428));
 sg13g2_tiehi _14525__429 (.L_HI(net429));
 sg13g2_tiehi _14139__430 (.L_HI(net430));
 sg13g2_tiehi _14713__431 (.L_HI(net431));
 sg13g2_tiehi _14138__432 (.L_HI(net432));
 sg13g2_tiehi _14524__433 (.L_HI(net433));
 sg13g2_tiehi _14137__434 (.L_HI(net434));
 sg13g2_tiehi _14712__435 (.L_HI(net435));
 sg13g2_tiehi _14136__436 (.L_HI(net436));
 sg13g2_tiehi _14523__437 (.L_HI(net437));
 sg13g2_tiehi _14135__438 (.L_HI(net438));
 sg13g2_tiehi _14711__439 (.L_HI(net439));
 sg13g2_tiehi _14134__440 (.L_HI(net440));
 sg13g2_tiehi _14522__441 (.L_HI(net441));
 sg13g2_tiehi _14133__442 (.L_HI(net442));
 sg13g2_tiehi _14710__443 (.L_HI(net443));
 sg13g2_tiehi _14132__444 (.L_HI(net444));
 sg13g2_tiehi _14521__445 (.L_HI(net445));
 sg13g2_tiehi _14131__446 (.L_HI(net446));
 sg13g2_tiehi _14709__447 (.L_HI(net447));
 sg13g2_tiehi _14130__448 (.L_HI(net448));
 sg13g2_tiehi _14520__449 (.L_HI(net449));
 sg13g2_tiehi _14129__450 (.L_HI(net450));
 sg13g2_tiehi _14708__451 (.L_HI(net451));
 sg13g2_tiehi _14128__452 (.L_HI(net452));
 sg13g2_tiehi _14519__453 (.L_HI(net453));
 sg13g2_tiehi _14127__454 (.L_HI(net454));
 sg13g2_tiehi _14707__455 (.L_HI(net455));
 sg13g2_tiehi _14126__456 (.L_HI(net456));
 sg13g2_tiehi _14518__457 (.L_HI(net457));
 sg13g2_tiehi _14125__458 (.L_HI(net458));
 sg13g2_tiehi _14706__459 (.L_HI(net459));
 sg13g2_tiehi _14124__460 (.L_HI(net460));
 sg13g2_tiehi _14517__461 (.L_HI(net461));
 sg13g2_tiehi _14123__462 (.L_HI(net462));
 sg13g2_tiehi _14705__463 (.L_HI(net463));
 sg13g2_tiehi _14122__464 (.L_HI(net464));
 sg13g2_tiehi _14516__465 (.L_HI(net465));
 sg13g2_tiehi _14121__466 (.L_HI(net466));
 sg13g2_tiehi _14704__467 (.L_HI(net467));
 sg13g2_tiehi _14120__468 (.L_HI(net468));
 sg13g2_tiehi _14515__469 (.L_HI(net469));
 sg13g2_tiehi _14119__470 (.L_HI(net470));
 sg13g2_tiehi _14703__471 (.L_HI(net471));
 sg13g2_tiehi _14118__472 (.L_HI(net472));
 sg13g2_tiehi _14514__473 (.L_HI(net473));
 sg13g2_tiehi _14117__474 (.L_HI(net474));
 sg13g2_tiehi _14702__475 (.L_HI(net475));
 sg13g2_tiehi _14116__476 (.L_HI(net476));
 sg13g2_tiehi _14513__477 (.L_HI(net477));
 sg13g2_tiehi _14115__478 (.L_HI(net478));
 sg13g2_tiehi _14701__479 (.L_HI(net479));
 sg13g2_tiehi _14114__480 (.L_HI(net480));
 sg13g2_tiehi _14512__481 (.L_HI(net481));
 sg13g2_tiehi _14113__482 (.L_HI(net482));
 sg13g2_tiehi _14700__483 (.L_HI(net483));
 sg13g2_tiehi _14112__484 (.L_HI(net484));
 sg13g2_tiehi _14511__485 (.L_HI(net485));
 sg13g2_tiehi _14111__486 (.L_HI(net486));
 sg13g2_tiehi _14699__487 (.L_HI(net487));
 sg13g2_tiehi _14110__488 (.L_HI(net488));
 sg13g2_tiehi _14510__489 (.L_HI(net489));
 sg13g2_tiehi _14109__490 (.L_HI(net490));
 sg13g2_tiehi _14698__491 (.L_HI(net491));
 sg13g2_tiehi _14108__492 (.L_HI(net492));
 sg13g2_tiehi _14509__493 (.L_HI(net493));
 sg13g2_tiehi _14107__494 (.L_HI(net494));
 sg13g2_tiehi _14697__495 (.L_HI(net495));
 sg13g2_tiehi _14106__496 (.L_HI(net496));
 sg13g2_tiehi _14508__497 (.L_HI(net497));
 sg13g2_tiehi _14105__498 (.L_HI(net498));
 sg13g2_tiehi _14696__499 (.L_HI(net499));
 sg13g2_tiehi _14104__500 (.L_HI(net500));
 sg13g2_tiehi _14507__501 (.L_HI(net501));
 sg13g2_tiehi _14103__502 (.L_HI(net502));
 sg13g2_tiehi _14695__503 (.L_HI(net503));
 sg13g2_tiehi _14102__504 (.L_HI(net504));
 sg13g2_tiehi _14506__505 (.L_HI(net505));
 sg13g2_tiehi _14101__506 (.L_HI(net506));
 sg13g2_tiehi _14694__507 (.L_HI(net507));
 sg13g2_tiehi _14100__508 (.L_HI(net508));
 sg13g2_tiehi _14505__509 (.L_HI(net509));
 sg13g2_tiehi _14099__510 (.L_HI(net510));
 sg13g2_tiehi _14693__511 (.L_HI(net511));
 sg13g2_tiehi _14098__512 (.L_HI(net512));
 sg13g2_tiehi _14504__513 (.L_HI(net513));
 sg13g2_tiehi _14097__514 (.L_HI(net514));
 sg13g2_tiehi _14692__515 (.L_HI(net515));
 sg13g2_tiehi _14096__516 (.L_HI(net516));
 sg13g2_tiehi _14503__517 (.L_HI(net517));
 sg13g2_tiehi _14095__518 (.L_HI(net518));
 sg13g2_tiehi _14691__519 (.L_HI(net519));
 sg13g2_tiehi _14094__520 (.L_HI(net520));
 sg13g2_tiehi _14502__521 (.L_HI(net521));
 sg13g2_tiehi _14093__522 (.L_HI(net522));
 sg13g2_tiehi _14674__523 (.L_HI(net523));
 sg13g2_tiehi _14092__524 (.L_HI(net524));
 sg13g2_tiehi _14501__525 (.L_HI(net525));
 sg13g2_tiehi _14091__526 (.L_HI(net526));
 sg13g2_tiehi _14673__527 (.L_HI(net527));
 sg13g2_tiehi _14090__528 (.L_HI(net528));
 sg13g2_tiehi _14500__529 (.L_HI(net529));
 sg13g2_tiehi _14089__530 (.L_HI(net530));
 sg13g2_tiehi _14672__531 (.L_HI(net531));
 sg13g2_tiehi _14088__532 (.L_HI(net532));
 sg13g2_tiehi _14499__533 (.L_HI(net533));
 sg13g2_tiehi _14087__534 (.L_HI(net534));
 sg13g2_tiehi _14671__535 (.L_HI(net535));
 sg13g2_tiehi _14086__536 (.L_HI(net536));
 sg13g2_tiehi _14498__537 (.L_HI(net537));
 sg13g2_tiehi _14085__538 (.L_HI(net538));
 sg13g2_tiehi _14670__539 (.L_HI(net539));
 sg13g2_tiehi _14084__540 (.L_HI(net540));
 sg13g2_tiehi _14497__541 (.L_HI(net541));
 sg13g2_tiehi _14083__542 (.L_HI(net542));
 sg13g2_tiehi _14669__543 (.L_HI(net543));
 sg13g2_tiehi _14082__544 (.L_HI(net544));
 sg13g2_tiehi _14496__545 (.L_HI(net545));
 sg13g2_tiehi _14081__546 (.L_HI(net546));
 sg13g2_tiehi _14668__547 (.L_HI(net547));
 sg13g2_tiehi _14080__548 (.L_HI(net548));
 sg13g2_tiehi _14495__549 (.L_HI(net549));
 sg13g2_tiehi _14079__550 (.L_HI(net550));
 sg13g2_tiehi _14667__551 (.L_HI(net551));
 sg13g2_tiehi _14078__552 (.L_HI(net552));
 sg13g2_tiehi _14494__553 (.L_HI(net553));
 sg13g2_tiehi _14077__554 (.L_HI(net554));
 sg13g2_tiehi _14666__555 (.L_HI(net555));
 sg13g2_tiehi _14076__556 (.L_HI(net556));
 sg13g2_tiehi _14493__557 (.L_HI(net557));
 sg13g2_tiehi _14075__558 (.L_HI(net558));
 sg13g2_tiehi _14665__559 (.L_HI(net559));
 sg13g2_tiehi _14074__560 (.L_HI(net560));
 sg13g2_tiehi _14492__561 (.L_HI(net561));
 sg13g2_tiehi _14073__562 (.L_HI(net562));
 sg13g2_tiehi _14664__563 (.L_HI(net563));
 sg13g2_tiehi _14072__564 (.L_HI(net564));
 sg13g2_tiehi _14491__565 (.L_HI(net565));
 sg13g2_tiehi _14071__566 (.L_HI(net566));
 sg13g2_tiehi _14663__567 (.L_HI(net567));
 sg13g2_tiehi _14070__568 (.L_HI(net568));
 sg13g2_tiehi _14490__569 (.L_HI(net569));
 sg13g2_tiehi _14069__570 (.L_HI(net570));
 sg13g2_tiehi _14662__571 (.L_HI(net571));
 sg13g2_tiehi _14068__572 (.L_HI(net572));
 sg13g2_tiehi _14489__573 (.L_HI(net573));
 sg13g2_tiehi _14067__574 (.L_HI(net574));
 sg13g2_tiehi _14661__575 (.L_HI(net575));
 sg13g2_tiehi _14066__576 (.L_HI(net576));
 sg13g2_tiehi _14488__577 (.L_HI(net577));
 sg13g2_tiehi _14065__578 (.L_HI(net578));
 sg13g2_tiehi _14660__579 (.L_HI(net579));
 sg13g2_tiehi _14064__580 (.L_HI(net580));
 sg13g2_tiehi _14487__581 (.L_HI(net581));
 sg13g2_tiehi _14063__582 (.L_HI(net582));
 sg13g2_tiehi _14659__583 (.L_HI(net583));
 sg13g2_tiehi _14062__584 (.L_HI(net584));
 sg13g2_tiehi _14486__585 (.L_HI(net585));
 sg13g2_tiehi _14061__586 (.L_HI(net586));
 sg13g2_tiehi _14658__587 (.L_HI(net587));
 sg13g2_tiehi _14060__588 (.L_HI(net588));
 sg13g2_tiehi _14485__589 (.L_HI(net589));
 sg13g2_tiehi _14059__590 (.L_HI(net590));
 sg13g2_tiehi _14657__591 (.L_HI(net591));
 sg13g2_tiehi _14058__592 (.L_HI(net592));
 sg13g2_tiehi _14484__593 (.L_HI(net593));
 sg13g2_tiehi _14057__594 (.L_HI(net594));
 sg13g2_tiehi _14656__595 (.L_HI(net595));
 sg13g2_tiehi _14056__596 (.L_HI(net596));
 sg13g2_tiehi _14483__597 (.L_HI(net597));
 sg13g2_tiehi _14055__598 (.L_HI(net598));
 sg13g2_tiehi _14655__599 (.L_HI(net599));
 sg13g2_tiehi _14054__600 (.L_HI(net600));
 sg13g2_tiehi _14482__601 (.L_HI(net601));
 sg13g2_tiehi _14053__602 (.L_HI(net602));
 sg13g2_tiehi _14654__603 (.L_HI(net603));
 sg13g2_tiehi _14052__604 (.L_HI(net604));
 sg13g2_tiehi _14481__605 (.L_HI(net605));
 sg13g2_tiehi _14051__606 (.L_HI(net606));
 sg13g2_tiehi _14653__607 (.L_HI(net607));
 sg13g2_tiehi _14050__608 (.L_HI(net608));
 sg13g2_tiehi _14480__609 (.L_HI(net609));
 sg13g2_tiehi _14049__610 (.L_HI(net610));
 sg13g2_tiehi _14652__611 (.L_HI(net611));
 sg13g2_tiehi _14048__612 (.L_HI(net612));
 sg13g2_tiehi _14479__613 (.L_HI(net613));
 sg13g2_tiehi _14047__614 (.L_HI(net614));
 sg13g2_tiehi _14651__615 (.L_HI(net615));
 sg13g2_tiehi _14046__616 (.L_HI(net616));
 sg13g2_tiehi _14478__617 (.L_HI(net617));
 sg13g2_tiehi _14045__618 (.L_HI(net618));
 sg13g2_tiehi _14650__619 (.L_HI(net619));
 sg13g2_tiehi _14044__620 (.L_HI(net620));
 sg13g2_tiehi _14043__621 (.L_HI(net621));
 sg13g2_tiehi _14042__622 (.L_HI(net622));
 sg13g2_tiehi _14041__623 (.L_HI(net623));
 sg13g2_tiehi _14040__624 (.L_HI(net624));
 sg13g2_tiehi _14039__625 (.L_HI(net625));
 sg13g2_tiehi _14038__626 (.L_HI(net626));
 sg13g2_tiehi _14037__627 (.L_HI(net627));
 sg13g2_tiehi _14036__628 (.L_HI(net628));
 sg13g2_tiehi _14035__629 (.L_HI(net629));
 sg13g2_tiehi _14034__630 (.L_HI(net630));
 sg13g2_tiehi _14033__631 (.L_HI(net631));
 sg13g2_tiehi _14032__632 (.L_HI(net632));
 sg13g2_tiehi _14031__633 (.L_HI(net633));
 sg13g2_tiehi _14030__634 (.L_HI(net634));
 sg13g2_tiehi _14029__635 (.L_HI(net635));
 sg13g2_tiehi _14028__636 (.L_HI(net636));
 sg13g2_tiehi _14027__637 (.L_HI(net637));
 sg13g2_tiehi _14026__638 (.L_HI(net638));
 sg13g2_tiehi _14025__639 (.L_HI(net639));
 sg13g2_tiehi _14024__640 (.L_HI(net640));
 sg13g2_tiehi _14023__641 (.L_HI(net641));
 sg13g2_tiehi _14022__642 (.L_HI(net642));
 sg13g2_tiehi _14477__643 (.L_HI(net643));
 sg13g2_tiehi _14021__644 (.L_HI(net644));
 sg13g2_tiehi _14649__645 (.L_HI(net645));
 sg13g2_tiehi _14020__646 (.L_HI(net646));
 sg13g2_tiehi _14476__647 (.L_HI(net647));
 sg13g2_tiehi _14019__648 (.L_HI(net648));
 sg13g2_tiehi _14648__649 (.L_HI(net649));
 sg13g2_tiehi _14018__650 (.L_HI(net650));
 sg13g2_tiehi _14475__651 (.L_HI(net651));
 sg13g2_tiehi _14017__652 (.L_HI(net652));
 sg13g2_tiehi _14647__653 (.L_HI(net653));
 sg13g2_tiehi _14016__654 (.L_HI(net654));
 sg13g2_tiehi _14474__655 (.L_HI(net655));
 sg13g2_tiehi _14015__656 (.L_HI(net656));
 sg13g2_tiehi _14646__657 (.L_HI(net657));
 sg13g2_tiehi _14014__658 (.L_HI(net658));
 sg13g2_tiehi _14473__659 (.L_HI(net659));
 sg13g2_tiehi _14013__660 (.L_HI(net660));
 sg13g2_tiehi _14472__661 (.L_HI(net661));
 sg13g2_tiehi _14012__662 (.L_HI(net662));
 sg13g2_tiehi _14471__663 (.L_HI(net663));
 sg13g2_tiehi _14011__664 (.L_HI(net664));
 sg13g2_tiehi _14470__665 (.L_HI(net665));
 sg13g2_tiehi _14010__666 (.L_HI(net666));
 sg13g2_tiehi _14469__667 (.L_HI(net667));
 sg13g2_tiehi _14009__668 (.L_HI(net668));
 sg13g2_tiehi _14468__669 (.L_HI(net669));
 sg13g2_tiehi _14008__670 (.L_HI(net670));
 sg13g2_tiehi _14467__671 (.L_HI(net671));
 sg13g2_tiehi _14007__672 (.L_HI(net672));
 sg13g2_tiehi _14466__673 (.L_HI(net673));
 sg13g2_tiehi _14006__674 (.L_HI(net674));
 sg13g2_tiehi _14465__675 (.L_HI(net675));
 sg13g2_tiehi _14005__676 (.L_HI(net676));
 sg13g2_tiehi _14464__677 (.L_HI(net677));
 sg13g2_tiehi _14004__678 (.L_HI(net678));
 sg13g2_tiehi _14463__679 (.L_HI(net679));
 sg13g2_tiehi _14003__680 (.L_HI(net680));
 sg13g2_tiehi _14462__681 (.L_HI(net681));
 sg13g2_tiehi _14002__682 (.L_HI(net682));
 sg13g2_tiehi _14461__683 (.L_HI(net683));
 sg13g2_tiehi _14001__684 (.L_HI(net684));
 sg13g2_tiehi _14460__685 (.L_HI(net685));
 sg13g2_tiehi _14000__686 (.L_HI(net686));
 sg13g2_tiehi _14459__687 (.L_HI(net687));
 sg13g2_tiehi _13999__688 (.L_HI(net688));
 sg13g2_tiehi _14458__689 (.L_HI(net689));
 sg13g2_tiehi _13998__690 (.L_HI(net690));
 sg13g2_tiehi _14457__691 (.L_HI(net691));
 sg13g2_tiehi _13997__692 (.L_HI(net692));
 sg13g2_tiehi _14456__693 (.L_HI(net693));
 sg13g2_tiehi _13996__694 (.L_HI(net694));
 sg13g2_tiehi _14455__695 (.L_HI(net695));
 sg13g2_tiehi _13995__696 (.L_HI(net696));
 sg13g2_tiehi _14454__697 (.L_HI(net697));
 sg13g2_tiehi _13994__698 (.L_HI(net698));
 sg13g2_tiehi _14453__699 (.L_HI(net699));
 sg13g2_tiehi _13993__700 (.L_HI(net700));
 sg13g2_tiehi _14452__701 (.L_HI(net701));
 sg13g2_tiehi _13992__702 (.L_HI(net702));
 sg13g2_tiehi _14451__703 (.L_HI(net703));
 sg13g2_tiehi _13991__704 (.L_HI(net704));
 sg13g2_tiehi _14450__705 (.L_HI(net705));
 sg13g2_tiehi _13990__706 (.L_HI(net706));
 sg13g2_tiehi _14449__707 (.L_HI(net707));
 sg13g2_tiehi _13989__708 (.L_HI(net708));
 sg13g2_tiehi _14448__709 (.L_HI(net709));
 sg13g2_tiehi _13988__710 (.L_HI(net710));
 sg13g2_tiehi _14447__711 (.L_HI(net711));
 sg13g2_tiehi _13987__712 (.L_HI(net712));
 sg13g2_tiehi _14446__713 (.L_HI(net713));
 sg13g2_tiehi _13986__714 (.L_HI(net714));
 sg13g2_tiehi _14445__715 (.L_HI(net715));
 sg13g2_tiehi _13985__716 (.L_HI(net716));
 sg13g2_tiehi _14444__717 (.L_HI(net717));
 sg13g2_tiehi _13984__718 (.L_HI(net718));
 sg13g2_tiehi _14443__719 (.L_HI(net719));
 sg13g2_tiehi _13983__720 (.L_HI(net720));
 sg13g2_tiehi _14442__721 (.L_HI(net721));
 sg13g2_tiehi _13982__722 (.L_HI(net722));
 sg13g2_tiehi _14441__723 (.L_HI(net723));
 sg13g2_tiehi _13981__724 (.L_HI(net724));
 sg13g2_tiehi _14440__725 (.L_HI(net725));
 sg13g2_tiehi _13980__726 (.L_HI(net726));
 sg13g2_tiehi _14439__727 (.L_HI(net727));
 sg13g2_tiehi _13979__728 (.L_HI(net728));
 sg13g2_tiehi _14438__729 (.L_HI(net729));
 sg13g2_tiehi _13978__730 (.L_HI(net730));
 sg13g2_tiehi _14437__731 (.L_HI(net731));
 sg13g2_tiehi _13977__732 (.L_HI(net732));
 sg13g2_tiehi _14436__733 (.L_HI(net733));
 sg13g2_tiehi _13976__734 (.L_HI(net734));
 sg13g2_tiehi _14435__735 (.L_HI(net735));
 sg13g2_tiehi _13975__736 (.L_HI(net736));
 sg13g2_tiehi _14434__737 (.L_HI(net737));
 sg13g2_tiehi _13974__738 (.L_HI(net738));
 sg13g2_tiehi _14433__739 (.L_HI(net739));
 sg13g2_tiehi _13973__740 (.L_HI(net740));
 sg13g2_tiehi _14432__741 (.L_HI(net741));
 sg13g2_tiehi _13972__742 (.L_HI(net742));
 sg13g2_tiehi _14431__743 (.L_HI(net743));
 sg13g2_tiehi _13971__744 (.L_HI(net744));
 sg13g2_tiehi _14430__745 (.L_HI(net745));
 sg13g2_tiehi _13970__746 (.L_HI(net746));
 sg13g2_tiehi _14429__747 (.L_HI(net747));
 sg13g2_tiehi _13969__748 (.L_HI(net748));
 sg13g2_tiehi _14428__749 (.L_HI(net749));
 sg13g2_tiehi _13968__750 (.L_HI(net750));
 sg13g2_tiehi _14427__751 (.L_HI(net751));
 sg13g2_tiehi _13967__752 (.L_HI(net752));
 sg13g2_tiehi _14426__753 (.L_HI(net753));
 sg13g2_tiehi _13966__754 (.L_HI(net754));
 sg13g2_tiehi _14425__755 (.L_HI(net755));
 sg13g2_tiehi _13965__756 (.L_HI(net756));
 sg13g2_tiehi _14424__757 (.L_HI(net757));
 sg13g2_tiehi _13964__758 (.L_HI(net758));
 sg13g2_tiehi _14423__759 (.L_HI(net759));
 sg13g2_tiehi _13963__760 (.L_HI(net760));
 sg13g2_tiehi _14422__761 (.L_HI(net761));
 sg13g2_tiehi _13962__762 (.L_HI(net762));
 sg13g2_tiehi _14421__763 (.L_HI(net763));
 sg13g2_tiehi _13961__764 (.L_HI(net764));
 sg13g2_tiehi _14420__765 (.L_HI(net765));
 sg13g2_tiehi _13960__766 (.L_HI(net766));
 sg13g2_tiehi _14419__767 (.L_HI(net767));
 sg13g2_tiehi _13959__768 (.L_HI(net768));
 sg13g2_tiehi _14418__769 (.L_HI(net769));
 sg13g2_tiehi _13958__770 (.L_HI(net770));
 sg13g2_tiehi _14417__771 (.L_HI(net771));
 sg13g2_tiehi _13957__772 (.L_HI(net772));
 sg13g2_tiehi _14416__773 (.L_HI(net773));
 sg13g2_tiehi _13956__774 (.L_HI(net774));
 sg13g2_tiehi _14415__775 (.L_HI(net775));
 sg13g2_tiehi _13955__776 (.L_HI(net776));
 sg13g2_tiehi _14414__777 (.L_HI(net777));
 sg13g2_tiehi _13954__778 (.L_HI(net778));
 sg13g2_tiehi _14413__779 (.L_HI(net779));
 sg13g2_tiehi _13953__780 (.L_HI(net780));
 sg13g2_tiehi _14412__781 (.L_HI(net781));
 sg13g2_tiehi _13952__782 (.L_HI(net782));
 sg13g2_tiehi _14411__783 (.L_HI(net783));
 sg13g2_tiehi _13951__784 (.L_HI(net784));
 sg13g2_tiehi _14410__785 (.L_HI(net785));
 sg13g2_tiehi _13950__786 (.L_HI(net786));
 sg13g2_tiehi _14409__787 (.L_HI(net787));
 sg13g2_tiehi _13949__788 (.L_HI(net788));
 sg13g2_tiehi _14408__789 (.L_HI(net789));
 sg13g2_tiehi _13948__790 (.L_HI(net790));
 sg13g2_tiehi _14407__791 (.L_HI(net791));
 sg13g2_tiehi _13947__792 (.L_HI(net792));
 sg13g2_tiehi _14406__793 (.L_HI(net793));
 sg13g2_tiehi _13946__794 (.L_HI(net794));
 sg13g2_tiehi _14405__795 (.L_HI(net795));
 sg13g2_tiehi _13945__796 (.L_HI(net796));
 sg13g2_tiehi _14404__797 (.L_HI(net797));
 sg13g2_tiehi _13944__798 (.L_HI(net798));
 sg13g2_tiehi _14403__799 (.L_HI(net799));
 sg13g2_tiehi _13943__800 (.L_HI(net800));
 sg13g2_tiehi _14402__801 (.L_HI(net801));
 sg13g2_tiehi _13942__802 (.L_HI(net802));
 sg13g2_tiehi _14401__803 (.L_HI(net803));
 sg13g2_tiehi _13941__804 (.L_HI(net804));
 sg13g2_tiehi _14400__805 (.L_HI(net805));
 sg13g2_tiehi _13940__806 (.L_HI(net806));
 sg13g2_tiehi _14399__807 (.L_HI(net807));
 sg13g2_tiehi _13939__808 (.L_HI(net808));
 sg13g2_tiehi _14398__809 (.L_HI(net809));
 sg13g2_tiehi _13938__810 (.L_HI(net810));
 sg13g2_tiehi _14397__811 (.L_HI(net811));
 sg13g2_tiehi _13937__812 (.L_HI(net812));
 sg13g2_tiehi _14396__813 (.L_HI(net813));
 sg13g2_tiehi _13936__814 (.L_HI(net814));
 sg13g2_tiehi _14395__815 (.L_HI(net815));
 sg13g2_tiehi _13935__816 (.L_HI(net816));
 sg13g2_tiehi _14394__817 (.L_HI(net817));
 sg13g2_tiehi _13934__818 (.L_HI(net818));
 sg13g2_tiehi _14645__819 (.L_HI(net819));
 sg13g2_tiehi _13933__820 (.L_HI(net820));
 sg13g2_tiehi _14393__821 (.L_HI(net821));
 sg13g2_tiehi _13932__822 (.L_HI(net822));
 sg13g2_tiehi _14644__823 (.L_HI(net823));
 sg13g2_tiehi _13931__824 (.L_HI(net824));
 sg13g2_tiehi _14392__825 (.L_HI(net825));
 sg13g2_tiehi _13930__826 (.L_HI(net826));
 sg13g2_tiehi _14643__827 (.L_HI(net827));
 sg13g2_tiehi _13929__828 (.L_HI(net828));
 sg13g2_tiehi _14391__829 (.L_HI(net829));
 sg13g2_tiehi _13928__830 (.L_HI(net830));
 sg13g2_tiehi _14642__831 (.L_HI(net831));
 sg13g2_tiehi _13927__832 (.L_HI(net832));
 sg13g2_tiehi _14390__833 (.L_HI(net833));
 sg13g2_tiehi _13926__834 (.L_HI(net834));
 sg13g2_tiehi _14641__835 (.L_HI(net835));
 sg13g2_tiehi _13925__836 (.L_HI(net836));
 sg13g2_tiehi _14389__837 (.L_HI(net837));
 sg13g2_tiehi _13924__838 (.L_HI(net838));
 sg13g2_tiehi _14640__839 (.L_HI(net839));
 sg13g2_tiehi _13923__840 (.L_HI(net840));
 sg13g2_tiehi _14388__841 (.L_HI(net841));
 sg13g2_tiehi _13922__842 (.L_HI(net842));
 sg13g2_tiehi _14639__843 (.L_HI(net843));
 sg13g2_tiehi _13921__844 (.L_HI(net844));
 sg13g2_tiehi _14387__845 (.L_HI(net845));
 sg13g2_tiehi _13920__846 (.L_HI(net846));
 sg13g2_tiehi _14638__847 (.L_HI(net847));
 sg13g2_tiehi _13919__848 (.L_HI(net848));
 sg13g2_tiehi _14386__849 (.L_HI(net849));
 sg13g2_tiehi _13918__850 (.L_HI(net850));
 sg13g2_tiehi _14637__851 (.L_HI(net851));
 sg13g2_tiehi _13917__852 (.L_HI(net852));
 sg13g2_tiehi _14385__853 (.L_HI(net853));
 sg13g2_tiehi _13916__854 (.L_HI(net854));
 sg13g2_tiehi _14636__855 (.L_HI(net855));
 sg13g2_tiehi _13915__856 (.L_HI(net856));
 sg13g2_tiehi _14384__857 (.L_HI(net857));
 sg13g2_tiehi _13914__858 (.L_HI(net858));
 sg13g2_tiehi _14635__859 (.L_HI(net859));
 sg13g2_tiehi _13913__860 (.L_HI(net860));
 sg13g2_tiehi _14383__861 (.L_HI(net861));
 sg13g2_tiehi _13912__862 (.L_HI(net862));
 sg13g2_tiehi _14634__863 (.L_HI(net863));
 sg13g2_tiehi _13911__864 (.L_HI(net864));
 sg13g2_tiehi _14382__865 (.L_HI(net865));
 sg13g2_tiehi _13910__866 (.L_HI(net866));
 sg13g2_tiehi _14633__867 (.L_HI(net867));
 sg13g2_tiehi _13909__868 (.L_HI(net868));
 sg13g2_tiehi _14381__869 (.L_HI(net869));
 sg13g2_tiehi _13908__870 (.L_HI(net870));
 sg13g2_tiehi _14632__871 (.L_HI(net871));
 sg13g2_tiehi _13907__872 (.L_HI(net872));
 sg13g2_tiehi _14380__873 (.L_HI(net873));
 sg13g2_tiehi _13906__874 (.L_HI(net874));
 sg13g2_tiehi _14631__875 (.L_HI(net875));
 sg13g2_tiehi _13905__876 (.L_HI(net876));
 sg13g2_tiehi _14379__877 (.L_HI(net877));
 sg13g2_tiehi _13904__878 (.L_HI(net878));
 sg13g2_tiehi _14630__879 (.L_HI(net879));
 sg13g2_tiehi _13903__880 (.L_HI(net880));
 sg13g2_tiehi _14378__881 (.L_HI(net881));
 sg13g2_tiehi _13902__882 (.L_HI(net882));
 sg13g2_tiehi _14629__883 (.L_HI(net883));
 sg13g2_tiehi _13901__884 (.L_HI(net884));
 sg13g2_tiehi _14377__885 (.L_HI(net885));
 sg13g2_tiehi _13900__886 (.L_HI(net886));
 sg13g2_tiehi _14628__887 (.L_HI(net887));
 sg13g2_tiehi _13899__888 (.L_HI(net888));
 sg13g2_tiehi _14376__889 (.L_HI(net889));
 sg13g2_tiehi _13898__890 (.L_HI(net890));
 sg13g2_tiehi _14627__891 (.L_HI(net891));
 sg13g2_tiehi _13897__892 (.L_HI(net892));
 sg13g2_tiehi _14375__893 (.L_HI(net893));
 sg13g2_tiehi _13896__894 (.L_HI(net894));
 sg13g2_tiehi _14626__895 (.L_HI(net895));
 sg13g2_tiehi _13895__896 (.L_HI(net896));
 sg13g2_tiehi _14374__897 (.L_HI(net897));
 sg13g2_tiehi _13894__898 (.L_HI(net898));
 sg13g2_tiehi _14625__899 (.L_HI(net899));
 sg13g2_tiehi _13893__900 (.L_HI(net900));
 sg13g2_tiehi _14373__901 (.L_HI(net901));
 sg13g2_tiehi _13892__902 (.L_HI(net902));
 sg13g2_tiehi _14624__903 (.L_HI(net903));
 sg13g2_tiehi _13891__904 (.L_HI(net904));
 sg13g2_tiehi _14372__905 (.L_HI(net905));
 sg13g2_tiehi _13890__906 (.L_HI(net906));
 sg13g2_tiehi _14623__907 (.L_HI(net907));
 sg13g2_tiehi _13889__908 (.L_HI(net908));
 sg13g2_tiehi _14371__909 (.L_HI(net909));
 sg13g2_tiehi _13888__910 (.L_HI(net910));
 sg13g2_tiehi _14622__911 (.L_HI(net911));
 sg13g2_tiehi _13887__912 (.L_HI(net912));
 sg13g2_tiehi _14370__913 (.L_HI(net913));
 sg13g2_tiehi _13886__914 (.L_HI(net914));
 sg13g2_tiehi _14621__915 (.L_HI(net915));
 sg13g2_tiehi _13885__916 (.L_HI(net916));
 sg13g2_tiehi _14369__917 (.L_HI(net917));
 sg13g2_tiehi _13884__918 (.L_HI(net918));
 sg13g2_tiehi _14620__919 (.L_HI(net919));
 sg13g2_tiehi _13883__920 (.L_HI(net920));
 sg13g2_tiehi _14368__921 (.L_HI(net921));
 sg13g2_tiehi _13882__922 (.L_HI(net922));
 sg13g2_tiehi _14619__923 (.L_HI(net923));
 sg13g2_tiehi _13881__924 (.L_HI(net924));
 sg13g2_tiehi _14367__925 (.L_HI(net925));
 sg13g2_tiehi _13880__926 (.L_HI(net926));
 sg13g2_tiehi _14618__927 (.L_HI(net927));
 sg13g2_tiehi _13879__928 (.L_HI(net928));
 sg13g2_tiehi _14366__929 (.L_HI(net929));
 sg13g2_tiehi _13878__930 (.L_HI(net930));
 sg13g2_tiehi _14773__931 (.L_HI(net931));
 sg13g2_tiehi _13877__932 (.L_HI(net932));
 sg13g2_tiehi _14365__933 (.L_HI(net933));
 sg13g2_tiehi _13876__934 (.L_HI(net934));
 sg13g2_tiehi _14617__935 (.L_HI(net935));
 sg13g2_tiehi _13875__936 (.L_HI(net936));
 sg13g2_tiehi _14364__937 (.L_HI(net937));
 sg13g2_tiehi _13874__938 (.L_HI(net938));
 sg13g2_tiehi _14772__939 (.L_HI(net939));
 sg13g2_tiehi _13873__940 (.L_HI(net940));
 sg13g2_tiehi _14363__941 (.L_HI(net941));
 sg13g2_tiehi _13872__942 (.L_HI(net942));
 sg13g2_tiehi _14616__943 (.L_HI(net943));
 sg13g2_tiehi _13871__944 (.L_HI(net944));
 sg13g2_tiehi _14362__945 (.L_HI(net945));
 sg13g2_tiehi _13870__946 (.L_HI(net946));
 sg13g2_tiehi _14771__947 (.L_HI(net947));
 sg13g2_tiehi _13869__948 (.L_HI(net948));
 sg13g2_tiehi _14361__949 (.L_HI(net949));
 sg13g2_tiehi _13868__950 (.L_HI(net950));
 sg13g2_tiehi _14615__951 (.L_HI(net951));
 sg13g2_tiehi _13867__952 (.L_HI(net952));
 sg13g2_tiehi _14360__953 (.L_HI(net953));
 sg13g2_tiehi _13866__954 (.L_HI(net954));
 sg13g2_tiehi _14770__955 (.L_HI(net955));
 sg13g2_tiehi _13865__956 (.L_HI(net956));
 sg13g2_tiehi _14359__957 (.L_HI(net957));
 sg13g2_tiehi _13864__958 (.L_HI(net958));
 sg13g2_tiehi _14614__959 (.L_HI(net959));
 sg13g2_tiehi _13863__960 (.L_HI(net960));
 sg13g2_tiehi _14358__961 (.L_HI(net961));
 sg13g2_tiehi _13862__962 (.L_HI(net962));
 sg13g2_tiehi _14769__963 (.L_HI(net963));
 sg13g2_tiehi _13861__964 (.L_HI(net964));
 sg13g2_tiehi _14357__965 (.L_HI(net965));
 sg13g2_tiehi _13860__966 (.L_HI(net966));
 sg13g2_tiehi _14613__967 (.L_HI(net967));
 sg13g2_tiehi _13859__968 (.L_HI(net968));
 sg13g2_tiehi _14356__969 (.L_HI(net969));
 sg13g2_tiehi _13858__970 (.L_HI(net970));
 sg13g2_tiehi _14768__971 (.L_HI(net971));
 sg13g2_tiehi _13857__972 (.L_HI(net972));
 sg13g2_tiehi _14355__973 (.L_HI(net973));
 sg13g2_tiehi _13856__974 (.L_HI(net974));
 sg13g2_tiehi _14612__975 (.L_HI(net975));
 sg13g2_tiehi _13855__976 (.L_HI(net976));
 sg13g2_tiehi _14354__977 (.L_HI(net977));
 sg13g2_tiehi _13854__978 (.L_HI(net978));
 sg13g2_tiehi _14767__979 (.L_HI(net979));
 sg13g2_tiehi _13853__980 (.L_HI(net980));
 sg13g2_tiehi _14353__981 (.L_HI(net981));
 sg13g2_tiehi _13852__982 (.L_HI(net982));
 sg13g2_tiehi _14611__983 (.L_HI(net983));
 sg13g2_tiehi _13851__984 (.L_HI(net984));
 sg13g2_tiehi _14352__985 (.L_HI(net985));
 sg13g2_tiehi _13850__986 (.L_HI(net986));
 sg13g2_tiehi _14802__987 (.L_HI(net987));
 sg13g2_tiehi _13849__988 (.L_HI(net988));
 sg13g2_tiehi _14351__989 (.L_HI(net989));
 sg13g2_tiehi _13848__990 (.L_HI(net990));
 sg13g2_tiehi _14610__991 (.L_HI(net991));
 sg13g2_tiehi _13847__992 (.L_HI(net992));
 sg13g2_tiehi _14350__993 (.L_HI(net993));
 sg13g2_tiehi _13846__994 (.L_HI(net994));
 sg13g2_tiehi _14766__995 (.L_HI(net995));
 sg13g2_tiehi _13845__996 (.L_HI(net996));
 sg13g2_tiehi _14349__997 (.L_HI(net997));
 sg13g2_tiehi _13844__998 (.L_HI(net998));
 sg13g2_tiehi _14609__999 (.L_HI(net999));
 sg13g2_tiehi _13843__1000 (.L_HI(net1000));
 sg13g2_tiehi _14348__1001 (.L_HI(net1001));
 sg13g2_tiehi _13842__1002 (.L_HI(net1002));
 sg13g2_tiehi _14804__1003 (.L_HI(net1003));
 sg13g2_tiehi _13841__1004 (.L_HI(net1004));
 sg13g2_tiehi _14347__1005 (.L_HI(net1005));
 sg13g2_tiehi _13840__1006 (.L_HI(net1006));
 sg13g2_tiehi _14608__1007 (.L_HI(net1007));
 sg13g2_tiehi _13839__1008 (.L_HI(net1008));
 sg13g2_tiehi _14346__1009 (.L_HI(net1009));
 sg13g2_tiehi _13838__1010 (.L_HI(net1010));
 sg13g2_tiehi _14765__1011 (.L_HI(net1011));
 sg13g2_tiehi _13837__1012 (.L_HI(net1012));
 sg13g2_tiehi _14345__1013 (.L_HI(net1013));
 sg13g2_tiehi _13836__1014 (.L_HI(net1014));
 sg13g2_tiehi _14607__1015 (.L_HI(net1015));
 sg13g2_tiehi _13835__1016 (.L_HI(net1016));
 sg13g2_tiehi _14344__1017 (.L_HI(net1017));
 sg13g2_tiehi _13834__1018 (.L_HI(net1018));
 sg13g2_tiehi _14801__1019 (.L_HI(net1019));
 sg13g2_tiehi _13833__1020 (.L_HI(net1020));
 sg13g2_tiehi _14343__1021 (.L_HI(net1021));
 sg13g2_tiehi _13832__1022 (.L_HI(net1022));
 sg13g2_tiehi _14606__1023 (.L_HI(net1023));
 sg13g2_tiehi _13831__1024 (.L_HI(net1024));
 sg13g2_tiehi _14342__1025 (.L_HI(net1025));
 sg13g2_tiehi _13830__1026 (.L_HI(net1026));
 sg13g2_tiehi _14764__1027 (.L_HI(net1027));
 sg13g2_tiehi _13829__1028 (.L_HI(net1028));
 sg13g2_tiehi _13828__1029 (.L_HI(net1029));
 sg13g2_tiehi _13827__1030 (.L_HI(net1030));
 sg13g2_tiehi _13826__1031 (.L_HI(net1031));
 sg13g2_tiehi _13825__1032 (.L_HI(net1032));
 sg13g2_tiehi _13765__1033 (.L_HI(net1033));
 sg13g2_tiehi _14675__1034 (.L_HI(net1034));
 sg13g2_tiehi _14676__1035 (.L_HI(net1035));
 sg13g2_tiehi _14677__1036 (.L_HI(net1036));
 sg13g2_tiehi _14678__1037 (.L_HI(net1037));
 sg13g2_tiehi _14679__1038 (.L_HI(net1038));
 sg13g2_tiehi _14680__1039 (.L_HI(net1039));
 sg13g2_tiehi _14681__1040 (.L_HI(net1040));
 sg13g2_tiehi _14682__1041 (.L_HI(net1041));
 sg13g2_tiehi _14683__1042 (.L_HI(net1042));
 sg13g2_tiehi _14684__1043 (.L_HI(net1043));
 sg13g2_tiehi _14685__1044 (.L_HI(net1044));
 sg13g2_tiehi _14686__1045 (.L_HI(net1045));
 sg13g2_tiehi _14687__1046 (.L_HI(net1046));
 sg13g2_tiehi _14688__1047 (.L_HI(net1047));
 sg13g2_tiehi _14689__1048 (.L_HI(net1048));
 sg13g2_tiehi _13824__1049 (.L_HI(net1049));
 sg13g2_tiehi _13823__1050 (.L_HI(net1050));
 sg13g2_tiehi _13822__1051 (.L_HI(net1051));
 sg13g2_tiehi _13821__1052 (.L_HI(net1052));
 sg13g2_tiehi _13820__1053 (.L_HI(net1053));
 sg13g2_tiehi _13819__1054 (.L_HI(net1054));
 sg13g2_tiehi _13818__1055 (.L_HI(net1055));
 sg13g2_tiehi _13817__1056 (.L_HI(net1056));
 sg13g2_tiehi _13816__1057 (.L_HI(net1057));
 sg13g2_tiehi _13815__1058 (.L_HI(net1058));
 sg13g2_tiehi _13814__1059 (.L_HI(net1059));
 sg13g2_tiehi _13813__1060 (.L_HI(net1060));
 sg13g2_tiehi _13812__1061 (.L_HI(net1061));
 sg13g2_tiehi _13811__1062 (.L_HI(net1062));
 sg13g2_tiehi _13810__1063 (.L_HI(net1063));
 sg13g2_tiehi _13809__1064 (.L_HI(net1064));
 sg13g2_tiehi _13808__1065 (.L_HI(net1065));
 sg13g2_tiehi _14341__1066 (.L_HI(net1066));
 sg13g2_tiehi _13807__1067 (.L_HI(net1067));
 sg13g2_tiehi _14605__1068 (.L_HI(net1068));
 sg13g2_tiehi _13806__1069 (.L_HI(net1069));
 sg13g2_tiehi _14340__1070 (.L_HI(net1070));
 sg13g2_tiehi _13805__1071 (.L_HI(net1071));
 sg13g2_tiehi _14805__1072 (.L_HI(net1072));
 sg13g2_tiehi _13804__1073 (.L_HI(net1073));
 sg13g2_tiehi _14339__1074 (.L_HI(net1074));
 sg13g2_tiehi _13803__1075 (.L_HI(net1075));
 sg13g2_tiehi _14604__1076 (.L_HI(net1076));
 sg13g2_tiehi _13802__1077 (.L_HI(net1077));
 sg13g2_tiehi _14338__1078 (.L_HI(net1078));
 sg13g2_tiehi _13801__1079 (.L_HI(net1079));
 sg13g2_tiehi _14763__1080 (.L_HI(net1080));
 sg13g2_tiehi _13800__1081 (.L_HI(net1081));
 sg13g2_tiehi _14337__1082 (.L_HI(net1082));
 sg13g2_tiehi _13799__1083 (.L_HI(net1083));
 sg13g2_tiehi _14603__1084 (.L_HI(net1084));
 sg13g2_tiehi _13798__1085 (.L_HI(net1085));
 sg13g2_tiehi _14336__1086 (.L_HI(net1086));
 sg13g2_tiehi _13797__1087 (.L_HI(net1087));
 sg13g2_tiehi _14800__1088 (.L_HI(net1088));
 sg13g2_tiehi _13796__1089 (.L_HI(net1089));
 sg13g2_tiehi _14335__1090 (.L_HI(net1090));
 sg13g2_tiehi _13795__1091 (.L_HI(net1091));
 sg13g2_tiehi _14602__1092 (.L_HI(net1092));
 sg13g2_tiehi _13794__1093 (.L_HI(net1093));
 sg13g2_tiehi _14334__1094 (.L_HI(net1094));
 sg13g2_tiehi _13793__1095 (.L_HI(net1095));
 sg13g2_tiehi _14762__1096 (.L_HI(net1096));
 sg13g2_tiehi _13792__1097 (.L_HI(net1097));
 sg13g2_tiehi _14333__1098 (.L_HI(net1098));
 sg13g2_tiehi _13791__1099 (.L_HI(net1099));
 sg13g2_tiehi _14601__1100 (.L_HI(net1100));
 sg13g2_tiehi _13790__1101 (.L_HI(net1101));
 sg13g2_tiehi _14332__1102 (.L_HI(net1102));
 sg13g2_tiehi _13789__1103 (.L_HI(net1103));
 sg13g2_tiehi _14803__1104 (.L_HI(net1104));
 sg13g2_tiehi _13788__1105 (.L_HI(net1105));
 sg13g2_tiehi _13787__1106 (.L_HI(net1106));
 sg13g2_tiehi _14331__1107 (.L_HI(net1107));
 sg13g2_tiehi _13786__1108 (.L_HI(net1108));
 sg13g2_tiehi _14600__1109 (.L_HI(net1109));
 sg13g2_tiehi _13785__1110 (.L_HI(net1110));
 sg13g2_tiehi _14330__1111 (.L_HI(net1111));
 sg13g2_tiehi _13784__1112 (.L_HI(net1112));
 sg13g2_tiehi _14761__1113 (.L_HI(net1113));
 sg13g2_tiehi _13783__1114 (.L_HI(net1114));
 sg13g2_tiehi _14329__1115 (.L_HI(net1115));
 sg13g2_tiehi _13782__1116 (.L_HI(net1116));
 sg13g2_tiehi _14599__1117 (.L_HI(net1117));
 sg13g2_tiehi _13781__1118 (.L_HI(net1118));
 sg13g2_tiehi _14328__1119 (.L_HI(net1119));
 sg13g2_tiehi _13780__1120 (.L_HI(net1120));
 sg13g2_tiehi _14799__1121 (.L_HI(net1121));
 sg13g2_tiehi _13779__1122 (.L_HI(net1122));
 sg13g2_tiehi _14327__1123 (.L_HI(net1123));
 sg13g2_tiehi _13778__1124 (.L_HI(net1124));
 sg13g2_tiehi _14598__1125 (.L_HI(net1125));
 sg13g2_tiehi _13777__1126 (.L_HI(net1126));
 sg13g2_tiehi _13776__1127 (.L_HI(net1127));
 sg13g2_tiehi _13775__1128 (.L_HI(net1128));
 sg13g2_tiehi _13774__1129 (.L_HI(net1129));
 sg13g2_tiehi _13773__1130 (.L_HI(net1130));
 sg13g2_tiehi _13772__1131 (.L_HI(net1131));
 sg13g2_tiehi _13771__1132 (.L_HI(net1132));
 sg13g2_tiehi _13770__1133 (.L_HI(net1133));
 sg13g2_tiehi _13769__1134 (.L_HI(net1134));
 sg13g2_tiehi _13768__1135 (.L_HI(net1135));
 sg13g2_tiehi _13767__1136 (.L_HI(net1136));
 sg13g2_tiehi _13766__1137 (.L_HI(net1137));
 sg13g2_tiehi _13757__1138 (.L_HI(net1138));
 sg13g2_tiehi _13756__1139 (.L_HI(net1139));
 sg13g2_tiehi _13755__1140 (.L_HI(net1140));
 sg13g2_tiehi _13754__1141 (.L_HI(net1141));
 sg13g2_tiehi _13753__1142 (.L_HI(net1142));
 sg13g2_tiehi _13752__1143 (.L_HI(net1143));
 sg13g2_tiehi _13751__1144 (.L_HI(net1144));
 sg13g2_tiehi _13750__1145 (.L_HI(net1145));
 sg13g2_tiehi _13749__1146 (.L_HI(net1146));
 sg13g2_tiehi _13748__1147 (.L_HI(net1147));
 sg13g2_tiehi _13747__1148 (.L_HI(net1148));
 sg13g2_tiehi _13746__1149 (.L_HI(net1149));
 sg13g2_tiehi _13745__1150 (.L_HI(net1150));
 sg13g2_tiehi _14326__1151 (.L_HI(net1151));
 sg13g2_tiehi _13744__1152 (.L_HI(net1152));
 sg13g2_tiehi _14760__1153 (.L_HI(net1153));
 sg13g2_tiehi _13743__1154 (.L_HI(net1154));
 sg13g2_tiehi _14325__1155 (.L_HI(net1155));
 sg13g2_tiehi _13742__1156 (.L_HI(net1156));
 sg13g2_tiehi _14597__1157 (.L_HI(net1157));
 sg13g2_tiehi _13734__1158 (.L_HI(net1158));
 sg13g2_tiehi _14324__1159 (.L_HI(net1159));
 sg13g2_tiehi _13733__1160 (.L_HI(net1160));
 sg13g2_tiehi _14690__1161 (.L_HI(net1161));
 sg13g2_tiehi _13732__1162 (.L_HI(net1162));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_6 (.L_LO(net6));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_7 (.L_LO(net7));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_8 (.L_LO(net8));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_9 (.L_LO(net9));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_10 (.L_LO(net10));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_11 (.L_LO(net11));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_12 (.L_LO(net12));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_13 (.L_LO(net13));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_14 (.L_LO(net14));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_15 (.L_LO(net15));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_16 (.L_LO(net16));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_17 (.L_LO(net17));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_18 (.L_LO(net18));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_19 (.L_LO(net19));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_20 (.L_LO(net20));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_21 (.L_LO(net21));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_22 (.L_LO(net22));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_23 (.L_LO(net23));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_24 (.L_LO(net24));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_25 (.L_LO(net25));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_26 (.L_LO(net26));
 sg13g2_tiehi _14323__27 (.L_HI(net27));
 sg13g2_buf_1 _15964_ (.A(COMP_OUT),
    .X(uo_out[0]));
 sg13g2_buf_2 _15965_ (.A(PWM_OUT),
    .X(uo_out[1]));
 sg13g2_buf_2 fanout1530 (.A(net1532),
    .X(net1530));
 sg13g2_buf_1 fanout1531 (.A(net1532),
    .X(net1531));
 sg13g2_buf_2 fanout1532 (.A(net1536),
    .X(net1532));
 sg13g2_buf_2 fanout1533 (.A(net1536),
    .X(net1533));
 sg13g2_buf_2 fanout1534 (.A(net1536),
    .X(net1534));
 sg13g2_buf_2 fanout1535 (.A(net1536),
    .X(net1535));
 sg13g2_buf_2 fanout1536 (.A(_02127_),
    .X(net1536));
 sg13g2_buf_4 fanout1537 (.X(net1537),
    .A(net1539));
 sg13g2_buf_4 fanout1538 (.X(net1538),
    .A(net1539));
 sg13g2_buf_4 fanout1539 (.X(net1539),
    .A(_00409_));
 sg13g2_buf_2 fanout1540 (.A(net1542),
    .X(net1540));
 sg13g2_buf_2 fanout1541 (.A(net1542),
    .X(net1541));
 sg13g2_buf_2 fanout1542 (.A(net1545),
    .X(net1542));
 sg13g2_buf_2 fanout1543 (.A(net1545),
    .X(net1543));
 sg13g2_buf_2 fanout1544 (.A(net1545),
    .X(net1544));
 sg13g2_buf_4 fanout1545 (.X(net1545),
    .A(_00839_));
 sg13g2_buf_2 fanout1546 (.A(net1549),
    .X(net1546));
 sg13g2_buf_2 fanout1547 (.A(net1549),
    .X(net1547));
 sg13g2_buf_2 fanout1548 (.A(net1549),
    .X(net1548));
 sg13g2_buf_1 fanout1549 (.A(net1552),
    .X(net1549));
 sg13g2_buf_2 fanout1550 (.A(net1552),
    .X(net1550));
 sg13g2_buf_2 fanout1551 (.A(net1552),
    .X(net1551));
 sg13g2_buf_2 fanout1552 (.A(_00624_),
    .X(net1552));
 sg13g2_buf_2 fanout1553 (.A(net1554),
    .X(net1553));
 sg13g2_buf_2 fanout1554 (.A(net1555),
    .X(net1554));
 sg13g2_buf_2 fanout1555 (.A(net1560),
    .X(net1555));
 sg13g2_buf_2 fanout1556 (.A(net1557),
    .X(net1556));
 sg13g2_buf_2 fanout1557 (.A(net1560),
    .X(net1557));
 sg13g2_buf_2 fanout1558 (.A(net1560),
    .X(net1558));
 sg13g2_buf_1 fanout1559 (.A(net1560),
    .X(net1559));
 sg13g2_buf_2 fanout1560 (.A(_04752_),
    .X(net1560));
 sg13g2_buf_2 fanout1561 (.A(_04752_),
    .X(net1561));
 sg13g2_buf_1 fanout1562 (.A(_04752_),
    .X(net1562));
 sg13g2_buf_2 fanout1563 (.A(_01935_),
    .X(net1563));
 sg13g2_buf_2 fanout1564 (.A(_01739_),
    .X(net1564));
 sg13g2_buf_2 fanout1565 (.A(_01739_),
    .X(net1565));
 sg13g2_buf_4 fanout1566 (.X(net1566),
    .A(_01737_));
 sg13g2_buf_2 fanout1567 (.A(net1568),
    .X(net1567));
 sg13g2_buf_2 fanout1568 (.A(_01709_),
    .X(net1568));
 sg13g2_buf_4 fanout1569 (.X(net1569),
    .A(net1571));
 sg13g2_buf_4 fanout1570 (.X(net1570),
    .A(net1571));
 sg13g2_buf_2 fanout1571 (.A(_02101_),
    .X(net1571));
 sg13g2_buf_2 fanout1572 (.A(_02030_),
    .X(net1572));
 sg13g2_buf_1 fanout1573 (.A(_02030_),
    .X(net1573));
 sg13g2_buf_2 fanout1574 (.A(net1576),
    .X(net1574));
 sg13g2_buf_1 fanout1575 (.A(net1576),
    .X(net1575));
 sg13g2_buf_2 fanout1576 (.A(_02030_),
    .X(net1576));
 sg13g2_buf_4 fanout1577 (.X(net1577),
    .A(net1578));
 sg13g2_buf_2 fanout1578 (.A(_02029_),
    .X(net1578));
 sg13g2_buf_4 fanout1579 (.X(net1579),
    .A(_02029_));
 sg13g2_buf_2 fanout1580 (.A(_01937_),
    .X(net1580));
 sg13g2_buf_2 fanout1581 (.A(net1583),
    .X(net1581));
 sg13g2_buf_2 fanout1582 (.A(net1583),
    .X(net1582));
 sg13g2_buf_2 fanout1583 (.A(_01924_),
    .X(net1583));
 sg13g2_buf_2 fanout1584 (.A(_01736_),
    .X(net1584));
 sg13g2_buf_2 fanout1585 (.A(net1586),
    .X(net1585));
 sg13g2_buf_1 fanout1586 (.A(net1587),
    .X(net1586));
 sg13g2_buf_2 fanout1587 (.A(net1588),
    .X(net1587));
 sg13g2_buf_2 fanout1588 (.A(net1590),
    .X(net1588));
 sg13g2_buf_2 fanout1589 (.A(net1590),
    .X(net1589));
 sg13g2_buf_2 fanout1590 (.A(_01671_),
    .X(net1590));
 sg13g2_buf_2 fanout1591 (.A(net1592),
    .X(net1591));
 sg13g2_buf_2 fanout1592 (.A(net1593),
    .X(net1592));
 sg13g2_buf_2 fanout1593 (.A(net1596),
    .X(net1593));
 sg13g2_buf_2 fanout1594 (.A(net1595),
    .X(net1594));
 sg13g2_buf_2 fanout1595 (.A(net1596),
    .X(net1595));
 sg13g2_buf_2 fanout1596 (.A(net1599),
    .X(net1596));
 sg13g2_buf_2 fanout1597 (.A(net1599),
    .X(net1597));
 sg13g2_buf_2 fanout1598 (.A(net1599),
    .X(net1598));
 sg13g2_buf_4 fanout1599 (.X(net1599),
    .A(_05495_));
 sg13g2_buf_2 fanout1600 (.A(net1602),
    .X(net1600));
 sg13g2_buf_2 fanout1601 (.A(net1602),
    .X(net1601));
 sg13g2_buf_2 fanout1602 (.A(_01918_),
    .X(net1602));
 sg13g2_buf_2 fanout1603 (.A(_01918_),
    .X(net1603));
 sg13g2_buf_2 fanout1604 (.A(net1605),
    .X(net1604));
 sg13g2_buf_2 fanout1605 (.A(net1607),
    .X(net1605));
 sg13g2_buf_2 fanout1606 (.A(net1607),
    .X(net1606));
 sg13g2_buf_2 fanout1607 (.A(_01673_),
    .X(net1607));
 sg13g2_buf_4 fanout1608 (.X(net1608),
    .A(_01599_));
 sg13g2_buf_2 fanout1609 (.A(net1611),
    .X(net1609));
 sg13g2_buf_2 fanout1610 (.A(_01598_),
    .X(net1610));
 sg13g2_buf_2 fanout1611 (.A(_01598_),
    .X(net1611));
 sg13g2_buf_2 fanout1612 (.A(net1613),
    .X(net1612));
 sg13g2_buf_2 fanout1613 (.A(net1614),
    .X(net1613));
 sg13g2_buf_4 fanout1614 (.X(net1614),
    .A(_04748_));
 sg13g2_buf_2 fanout1615 (.A(_04748_),
    .X(net1615));
 sg13g2_buf_4 fanout1616 (.X(net1616),
    .A(_02099_));
 sg13g2_buf_2 fanout1617 (.A(_01920_),
    .X(net1617));
 sg13g2_buf_2 fanout1618 (.A(net1619),
    .X(net1618));
 sg13g2_buf_2 fanout1619 (.A(_01919_),
    .X(net1619));
 sg13g2_buf_2 fanout1620 (.A(_01669_),
    .X(net1620));
 sg13g2_buf_2 fanout1621 (.A(_01582_),
    .X(net1621));
 sg13g2_buf_2 fanout1622 (.A(net1623),
    .X(net1622));
 sg13g2_buf_4 fanout1623 (.X(net1623),
    .A(net1624));
 sg13g2_buf_4 fanout1624 (.X(net1624),
    .A(_01481_));
 sg13g2_buf_1 fanout1625 (.A(_01481_),
    .X(net1625));
 sg13g2_buf_4 fanout1626 (.X(net1626),
    .A(net1627));
 sg13g2_buf_4 fanout1627 (.X(net1627),
    .A(_01470_));
 sg13g2_buf_4 fanout1628 (.X(net1628),
    .A(_01395_));
 sg13g2_buf_2 fanout1629 (.A(_01395_),
    .X(net1629));
 sg13g2_buf_2 fanout1630 (.A(net1632),
    .X(net1630));
 sg13g2_buf_1 fanout1631 (.A(net1632),
    .X(net1631));
 sg13g2_buf_1 fanout1632 (.A(net1634),
    .X(net1632));
 sg13g2_buf_2 fanout1633 (.A(net1634),
    .X(net1633));
 sg13g2_buf_2 fanout1634 (.A(_01395_),
    .X(net1634));
 sg13g2_buf_4 fanout1635 (.X(net1635),
    .A(_01384_));
 sg13g2_buf_4 fanout1636 (.X(net1636),
    .A(_01384_));
 sg13g2_buf_4 fanout1637 (.X(net1637),
    .A(net1638));
 sg13g2_buf_4 fanout1638 (.X(net1638),
    .A(net1641));
 sg13g2_buf_4 fanout1639 (.X(net1639),
    .A(net1640));
 sg13g2_buf_4 fanout1640 (.X(net1640),
    .A(net1641));
 sg13g2_buf_2 fanout1641 (.A(_01306_),
    .X(net1641));
 sg13g2_buf_4 fanout1642 (.X(net1642),
    .A(net1646));
 sg13g2_buf_2 fanout1643 (.A(net1645),
    .X(net1643));
 sg13g2_buf_2 fanout1644 (.A(net1645),
    .X(net1644));
 sg13g2_buf_2 fanout1645 (.A(net1646),
    .X(net1645));
 sg13g2_buf_4 fanout1646 (.X(net1646),
    .A(_01223_));
 sg13g2_buf_2 fanout1647 (.A(\am_sdr0.am0.demod_out[9] ),
    .X(net1647));
 sg13g2_buf_2 fanout1648 (.A(net1650),
    .X(net1648));
 sg13g2_buf_2 fanout1649 (.A(net1650),
    .X(net1649));
 sg13g2_buf_2 fanout1650 (.A(net2956),
    .X(net1650));
 sg13g2_buf_2 fanout1651 (.A(net1652),
    .X(net1651));
 sg13g2_buf_2 fanout1652 (.A(net2130),
    .X(net1652));
 sg13g2_buf_2 fanout1653 (.A(net2947),
    .X(net1653));
 sg13g2_buf_2 fanout1654 (.A(net3018),
    .X(net1654));
 sg13g2_buf_2 fanout1655 (.A(\am_sdr0.mix0.RF_in_qq ),
    .X(net1655));
 sg13g2_buf_2 fanout1656 (.A(\am_sdr0.mix0.RF_in_qq ),
    .X(net1656));
 sg13g2_buf_2 fanout1657 (.A(net1659),
    .X(net1657));
 sg13g2_buf_2 fanout1658 (.A(net1659),
    .X(net1658));
 sg13g2_buf_2 fanout1659 (.A(\am_sdr0.Q_out[7] ),
    .X(net1659));
 sg13g2_buf_4 fanout1660 (.X(net1660),
    .A(net1662));
 sg13g2_buf_2 fanout1661 (.A(\am_sdr0.Q_out[7] ),
    .X(net1661));
 sg13g2_buf_1 fanout1662 (.A(\am_sdr0.Q_out[7] ),
    .X(net1662));
 sg13g2_buf_2 fanout1663 (.A(net1664),
    .X(net1663));
 sg13g2_buf_2 fanout1664 (.A(\am_sdr0.I_out[7] ),
    .X(net1664));
 sg13g2_buf_1 fanout1665 (.A(\am_sdr0.I_out[7] ),
    .X(net1665));
 sg13g2_buf_2 fanout1666 (.A(net1667),
    .X(net1666));
 sg13g2_buf_1 fanout1667 (.A(net1668),
    .X(net1667));
 sg13g2_buf_2 fanout1668 (.A(net1669),
    .X(net1668));
 sg13g2_buf_2 fanout1669 (.A(\am_sdr0.I_out[7] ),
    .X(net1669));
 sg13g2_buf_2 fanout1670 (.A(net1671),
    .X(net1670));
 sg13g2_buf_2 fanout1671 (.A(net1682),
    .X(net1671));
 sg13g2_buf_1 fanout1672 (.A(net1682),
    .X(net1672));
 sg13g2_buf_2 fanout1673 (.A(net1674),
    .X(net1673));
 sg13g2_buf_2 fanout1674 (.A(net1676),
    .X(net1674));
 sg13g2_buf_2 fanout1675 (.A(net1676),
    .X(net1675));
 sg13g2_buf_2 fanout1676 (.A(net1682),
    .X(net1676));
 sg13g2_buf_2 fanout1677 (.A(net1678),
    .X(net1677));
 sg13g2_buf_2 fanout1678 (.A(net1681),
    .X(net1678));
 sg13g2_buf_2 fanout1679 (.A(net1681),
    .X(net1679));
 sg13g2_buf_1 fanout1680 (.A(net1681),
    .X(net1680));
 sg13g2_buf_2 fanout1681 (.A(net1682),
    .X(net1681));
 sg13g2_buf_2 fanout1682 (.A(\am_sdr0.cic0.out_tick ),
    .X(net1682));
 sg13g2_buf_2 fanout1683 (.A(net1688),
    .X(net1683));
 sg13g2_buf_1 fanout1684 (.A(net1688),
    .X(net1684));
 sg13g2_buf_2 fanout1685 (.A(net1687),
    .X(net1685));
 sg13g2_buf_2 fanout1686 (.A(net1688),
    .X(net1686));
 sg13g2_buf_1 fanout1687 (.A(net1688),
    .X(net1687));
 sg13g2_buf_1 fanout1688 (.A(\am_sdr0.cic0.out_tick ),
    .X(net1688));
 sg13g2_buf_2 fanout1689 (.A(net1692),
    .X(net1689));
 sg13g2_buf_2 fanout1690 (.A(net1691),
    .X(net1690));
 sg13g2_buf_2 fanout1691 (.A(net1692),
    .X(net1691));
 sg13g2_buf_1 fanout1692 (.A(\am_sdr0.cic0.out_tick ),
    .X(net1692));
 sg13g2_buf_2 fanout1693 (.A(net1696),
    .X(net1693));
 sg13g2_buf_4 fanout1694 (.X(net1694),
    .A(net1696));
 sg13g2_buf_2 fanout1695 (.A(net1696),
    .X(net1695));
 sg13g2_buf_2 fanout1696 (.A(\am_sdr0.cic0.x_out[15] ),
    .X(net1696));
 sg13g2_buf_4 fanout1697 (.X(net1697),
    .A(net1698));
 sg13g2_buf_2 fanout1698 (.A(\am_sdr0.cic0.x_out[15] ),
    .X(net1698));
 sg13g2_buf_2 fanout1699 (.A(net1702),
    .X(net1699));
 sg13g2_buf_2 fanout1700 (.A(net1702),
    .X(net1700));
 sg13g2_buf_2 fanout1701 (.A(net1702),
    .X(net1701));
 sg13g2_buf_2 fanout1702 (.A(net1706),
    .X(net1702));
 sg13g2_buf_2 fanout1703 (.A(net1704),
    .X(net1703));
 sg13g2_buf_2 fanout1704 (.A(net1706),
    .X(net1704));
 sg13g2_buf_2 fanout1705 (.A(net1706),
    .X(net1705));
 sg13g2_buf_2 fanout1706 (.A(\am_sdr0.cic0.sample ),
    .X(net1706));
 sg13g2_buf_2 fanout1707 (.A(net1708),
    .X(net1707));
 sg13g2_buf_2 fanout1708 (.A(net1709),
    .X(net1708));
 sg13g2_buf_2 fanout1709 (.A(net1715),
    .X(net1709));
 sg13g2_buf_2 fanout1710 (.A(net1714),
    .X(net1710));
 sg13g2_buf_2 fanout1711 (.A(net1714),
    .X(net1711));
 sg13g2_buf_2 fanout1712 (.A(net1714),
    .X(net1712));
 sg13g2_buf_1 fanout1713 (.A(net1714),
    .X(net1713));
 sg13g2_buf_1 fanout1714 (.A(net1715),
    .X(net1714));
 sg13g2_buf_2 fanout1715 (.A(\am_sdr0.cic0.sample ),
    .X(net1715));
 sg13g2_buf_2 fanout1716 (.A(net1720),
    .X(net1716));
 sg13g2_buf_2 fanout1717 (.A(net1719),
    .X(net1717));
 sg13g2_buf_2 fanout1718 (.A(net1719),
    .X(net1718));
 sg13g2_buf_2 fanout1719 (.A(net1720),
    .X(net1719));
 sg13g2_buf_1 fanout1720 (.A(net1734),
    .X(net1720));
 sg13g2_buf_2 fanout1721 (.A(net1726),
    .X(net1721));
 sg13g2_buf_2 fanout1722 (.A(net1725),
    .X(net1722));
 sg13g2_buf_2 fanout1723 (.A(net1725),
    .X(net1723));
 sg13g2_buf_1 fanout1724 (.A(net1725),
    .X(net1724));
 sg13g2_buf_1 fanout1725 (.A(net1726),
    .X(net1725));
 sg13g2_buf_1 fanout1726 (.A(net1734),
    .X(net1726));
 sg13g2_buf_2 fanout1727 (.A(net1730),
    .X(net1727));
 sg13g2_buf_2 fanout1728 (.A(net1730),
    .X(net1728));
 sg13g2_buf_1 fanout1729 (.A(net1730),
    .X(net1729));
 sg13g2_buf_2 fanout1730 (.A(net1734),
    .X(net1730));
 sg13g2_buf_2 fanout1731 (.A(net1732),
    .X(net1731));
 sg13g2_buf_2 fanout1732 (.A(net1733),
    .X(net1732));
 sg13g2_buf_2 fanout1733 (.A(net1734),
    .X(net1733));
 sg13g2_buf_2 fanout1734 (.A(\am_sdr0.cic0.sample ),
    .X(net1734));
 sg13g2_buf_2 fanout1735 (.A(net1737),
    .X(net1735));
 sg13g2_buf_2 fanout1736 (.A(net1737),
    .X(net1736));
 sg13g2_buf_2 fanout1737 (.A(net1739),
    .X(net1737));
 sg13g2_buf_2 fanout1738 (.A(net1739),
    .X(net1738));
 sg13g2_buf_2 fanout1739 (.A(\am_sdr0.cic1.out_tick ),
    .X(net1739));
 sg13g2_buf_2 fanout1740 (.A(net1741),
    .X(net1740));
 sg13g2_buf_2 fanout1741 (.A(net1748),
    .X(net1741));
 sg13g2_buf_2 fanout1742 (.A(net1743),
    .X(net1742));
 sg13g2_buf_2 fanout1743 (.A(net1748),
    .X(net1743));
 sg13g2_buf_2 fanout1744 (.A(net1748),
    .X(net1744));
 sg13g2_buf_1 fanout1745 (.A(net1748),
    .X(net1745));
 sg13g2_buf_2 fanout1746 (.A(net1747),
    .X(net1746));
 sg13g2_buf_2 fanout1747 (.A(net1748),
    .X(net1747));
 sg13g2_buf_2 fanout1748 (.A(\am_sdr0.cic1.out_tick ),
    .X(net1748));
 sg13g2_buf_2 fanout1749 (.A(net1750),
    .X(net1749));
 sg13g2_buf_2 fanout1750 (.A(net1755),
    .X(net1750));
 sg13g2_buf_2 fanout1751 (.A(net1755),
    .X(net1751));
 sg13g2_buf_2 fanout1752 (.A(net1755),
    .X(net1752));
 sg13g2_buf_2 fanout1753 (.A(net1754),
    .X(net1753));
 sg13g2_buf_2 fanout1754 (.A(net1755),
    .X(net1754));
 sg13g2_buf_2 fanout1755 (.A(\am_sdr0.cic1.out_tick ),
    .X(net1755));
 sg13g2_buf_4 fanout1756 (.X(net1756),
    .A(net1758));
 sg13g2_buf_2 fanout1757 (.A(net1758),
    .X(net1757));
 sg13g2_buf_1 fanout1758 (.A(\am_sdr0.cic1.x_out[15] ),
    .X(net1758));
 sg13g2_buf_2 fanout1759 (.A(net1761),
    .X(net1759));
 sg13g2_buf_2 fanout1760 (.A(net1761),
    .X(net1760));
 sg13g2_buf_2 fanout1761 (.A(\am_sdr0.cic1.x_out[15] ),
    .X(net1761));
 sg13g2_buf_2 fanout1762 (.A(net1765),
    .X(net1762));
 sg13g2_buf_1 fanout1763 (.A(net1765),
    .X(net1763));
 sg13g2_buf_2 fanout1764 (.A(net1765),
    .X(net1764));
 sg13g2_buf_1 fanout1765 (.A(net1783),
    .X(net1765));
 sg13g2_buf_2 fanout1766 (.A(net1767),
    .X(net1766));
 sg13g2_buf_2 fanout1767 (.A(net1771),
    .X(net1767));
 sg13g2_buf_2 fanout1768 (.A(net1771),
    .X(net1768));
 sg13g2_buf_2 fanout1769 (.A(net1770),
    .X(net1769));
 sg13g2_buf_2 fanout1770 (.A(net1771),
    .X(net1770));
 sg13g2_buf_2 fanout1771 (.A(net1783),
    .X(net1771));
 sg13g2_buf_2 fanout1772 (.A(net1777),
    .X(net1772));
 sg13g2_buf_2 fanout1773 (.A(net1777),
    .X(net1773));
 sg13g2_buf_2 fanout1774 (.A(net1776),
    .X(net1774));
 sg13g2_buf_2 fanout1775 (.A(net1777),
    .X(net1775));
 sg13g2_buf_1 fanout1776 (.A(net1777),
    .X(net1776));
 sg13g2_buf_1 fanout1777 (.A(net1783),
    .X(net1777));
 sg13g2_buf_2 fanout1778 (.A(net1779),
    .X(net1778));
 sg13g2_buf_2 fanout1779 (.A(net1783),
    .X(net1779));
 sg13g2_buf_2 fanout1780 (.A(net1782),
    .X(net1780));
 sg13g2_buf_2 fanout1781 (.A(net1782),
    .X(net1781));
 sg13g2_buf_2 fanout1782 (.A(net1783),
    .X(net1782));
 sg13g2_buf_2 fanout1783 (.A(\am_sdr0.cic1.sample ),
    .X(net1783));
 sg13g2_buf_2 fanout1784 (.A(net1785),
    .X(net1784));
 sg13g2_buf_2 fanout1785 (.A(net1788),
    .X(net1785));
 sg13g2_buf_2 fanout1786 (.A(net1787),
    .X(net1786));
 sg13g2_buf_2 fanout1787 (.A(net1788),
    .X(net1787));
 sg13g2_buf_2 fanout1788 (.A(net1793),
    .X(net1788));
 sg13g2_buf_2 fanout1789 (.A(net1790),
    .X(net1789));
 sg13g2_buf_2 fanout1790 (.A(net1793),
    .X(net1790));
 sg13g2_buf_2 fanout1791 (.A(net1793),
    .X(net1791));
 sg13g2_buf_1 fanout1792 (.A(net1793),
    .X(net1792));
 sg13g2_buf_1 fanout1793 (.A(\am_sdr0.cic1.sample ),
    .X(net1793));
 sg13g2_buf_2 fanout1794 (.A(net1795),
    .X(net1794));
 sg13g2_buf_1 fanout1795 (.A(net1796),
    .X(net1795));
 sg13g2_buf_1 fanout1796 (.A(\am_sdr0.cic1.sample ),
    .X(net1796));
 sg13g2_buf_2 fanout1797 (.A(net1799),
    .X(net1797));
 sg13g2_buf_2 fanout1798 (.A(net1799),
    .X(net1798));
 sg13g2_buf_2 fanout1799 (.A(net1800),
    .X(net1799));
 sg13g2_buf_2 fanout1800 (.A(net1803),
    .X(net1800));
 sg13g2_buf_2 fanout1801 (.A(net1802),
    .X(net1801));
 sg13g2_buf_2 fanout1802 (.A(net1803),
    .X(net1802));
 sg13g2_buf_1 fanout1803 (.A(\am_sdr0.cic2.sample ),
    .X(net1803));
 sg13g2_buf_2 fanout1804 (.A(net1806),
    .X(net1804));
 sg13g2_buf_2 fanout1805 (.A(net1806),
    .X(net1805));
 sg13g2_buf_1 fanout1806 (.A(net3009),
    .X(net1806));
 sg13g2_buf_2 fanout1807 (.A(net1811),
    .X(net1807));
 sg13g2_buf_1 fanout1808 (.A(net1811),
    .X(net1808));
 sg13g2_buf_2 fanout1809 (.A(net1811),
    .X(net1809));
 sg13g2_buf_1 fanout1810 (.A(net1811),
    .X(net1810));
 sg13g2_buf_1 fanout1811 (.A(net1812),
    .X(net1811));
 sg13g2_buf_2 fanout1812 (.A(net1830),
    .X(net1812));
 sg13g2_buf_2 fanout1813 (.A(net1815),
    .X(net1813));
 sg13g2_buf_2 fanout1814 (.A(net1815),
    .X(net1814));
 sg13g2_buf_2 fanout1815 (.A(net1830),
    .X(net1815));
 sg13g2_buf_2 fanout1816 (.A(net1818),
    .X(net1816));
 sg13g2_buf_2 fanout1817 (.A(net1818),
    .X(net1817));
 sg13g2_buf_2 fanout1818 (.A(net1830),
    .X(net1818));
 sg13g2_buf_2 fanout1819 (.A(net1821),
    .X(net1819));
 sg13g2_buf_1 fanout1820 (.A(net1821),
    .X(net1820));
 sg13g2_buf_2 fanout1821 (.A(net1826),
    .X(net1821));
 sg13g2_buf_2 fanout1822 (.A(net1826),
    .X(net1822));
 sg13g2_buf_2 fanout1823 (.A(net1824),
    .X(net1823));
 sg13g2_buf_1 fanout1824 (.A(net1825),
    .X(net1824));
 sg13g2_buf_1 fanout1825 (.A(net1826),
    .X(net1825));
 sg13g2_buf_2 fanout1826 (.A(net1830),
    .X(net1826));
 sg13g2_buf_2 fanout1827 (.A(net1828),
    .X(net1827));
 sg13g2_buf_2 fanout1828 (.A(net1829),
    .X(net1828));
 sg13g2_buf_2 fanout1829 (.A(net1830),
    .X(net1829));
 sg13g2_buf_2 fanout1830 (.A(\am_sdr0.cic2.sample ),
    .X(net1830));
 sg13g2_buf_2 fanout1831 (.A(net1835),
    .X(net1831));
 sg13g2_buf_1 fanout1832 (.A(net1835),
    .X(net1832));
 sg13g2_buf_2 fanout1833 (.A(net1835),
    .X(net1833));
 sg13g2_buf_1 fanout1834 (.A(net1835),
    .X(net1834));
 sg13g2_buf_2 fanout1835 (.A(net1869),
    .X(net1835));
 sg13g2_buf_2 fanout1836 (.A(net1838),
    .X(net1836));
 sg13g2_buf_1 fanout1837 (.A(net1838),
    .X(net1837));
 sg13g2_buf_2 fanout1838 (.A(net1842),
    .X(net1838));
 sg13g2_buf_2 fanout1839 (.A(net1841),
    .X(net1839));
 sg13g2_buf_2 fanout1840 (.A(net1841),
    .X(net1840));
 sg13g2_buf_2 fanout1841 (.A(net1842),
    .X(net1841));
 sg13g2_buf_1 fanout1842 (.A(net1869),
    .X(net1842));
 sg13g2_buf_2 fanout1843 (.A(net1849),
    .X(net1843));
 sg13g2_buf_1 fanout1844 (.A(net1849),
    .X(net1844));
 sg13g2_buf_2 fanout1845 (.A(net1849),
    .X(net1845));
 sg13g2_buf_2 fanout1846 (.A(net1847),
    .X(net1846));
 sg13g2_buf_1 fanout1847 (.A(net1848),
    .X(net1847));
 sg13g2_buf_2 fanout1848 (.A(net1849),
    .X(net1848));
 sg13g2_buf_1 fanout1849 (.A(net1869),
    .X(net1849));
 sg13g2_buf_2 fanout1850 (.A(net1852),
    .X(net1850));
 sg13g2_buf_1 fanout1851 (.A(net1852),
    .X(net1851));
 sg13g2_buf_2 fanout1852 (.A(net1868),
    .X(net1852));
 sg13g2_buf_2 fanout1853 (.A(net1855),
    .X(net1853));
 sg13g2_buf_1 fanout1854 (.A(net1855),
    .X(net1854));
 sg13g2_buf_1 fanout1855 (.A(net1868),
    .X(net1855));
 sg13g2_buf_2 fanout1856 (.A(net1859),
    .X(net1856));
 sg13g2_buf_2 fanout1857 (.A(net1859),
    .X(net1857));
 sg13g2_buf_1 fanout1858 (.A(net1859),
    .X(net1858));
 sg13g2_buf_2 fanout1859 (.A(net1868),
    .X(net1859));
 sg13g2_buf_2 fanout1860 (.A(net1863),
    .X(net1860));
 sg13g2_buf_2 fanout1861 (.A(net1863),
    .X(net1861));
 sg13g2_buf_2 fanout1862 (.A(net1863),
    .X(net1862));
 sg13g2_buf_1 fanout1863 (.A(net1868),
    .X(net1863));
 sg13g2_buf_2 fanout1864 (.A(net1865),
    .X(net1864));
 sg13g2_buf_2 fanout1865 (.A(net1867),
    .X(net1865));
 sg13g2_buf_2 fanout1866 (.A(net1867),
    .X(net1866));
 sg13g2_buf_2 fanout1867 (.A(net1868),
    .X(net1867));
 sg13g2_buf_2 fanout1868 (.A(net1869),
    .X(net1868));
 sg13g2_buf_2 fanout1869 (.A(\am_sdr0.cic3.sample ),
    .X(net1869));
 sg13g2_buf_2 fanout1870 (.A(net3225),
    .X(net1870));
 sg13g2_buf_2 fanout1871 (.A(net1872),
    .X(net1871));
 sg13g2_buf_2 fanout1872 (.A(\am_sdr0.am0.r[9] ),
    .X(net1872));
 sg13g2_buf_2 fanout1873 (.A(net2897),
    .X(net1873));
 sg13g2_buf_4 fanout1874 (.X(net1874),
    .A(net1875));
 sg13g2_buf_2 fanout1875 (.A(net1878),
    .X(net1875));
 sg13g2_buf_4 fanout1876 (.X(net1876),
    .A(net1877));
 sg13g2_buf_2 fanout1877 (.A(net1878),
    .X(net1877));
 sg13g2_buf_8 fanout1878 (.A(net1895),
    .X(net1878));
 sg13g2_buf_4 fanout1879 (.X(net1879),
    .A(net1880));
 sg13g2_buf_2 fanout1880 (.A(net1887),
    .X(net1880));
 sg13g2_buf_4 fanout1881 (.X(net1881),
    .A(net1883));
 sg13g2_buf_4 fanout1882 (.X(net1882),
    .A(net1887));
 sg13g2_buf_2 fanout1883 (.A(net1887),
    .X(net1883));
 sg13g2_buf_4 fanout1884 (.X(net1884),
    .A(net1886));
 sg13g2_buf_1 fanout1885 (.A(net1886),
    .X(net1885));
 sg13g2_buf_4 fanout1886 (.X(net1886),
    .A(net1887));
 sg13g2_buf_2 fanout1887 (.A(net1895),
    .X(net1887));
 sg13g2_buf_4 fanout1888 (.X(net1888),
    .A(net1889));
 sg13g2_buf_4 fanout1889 (.X(net1889),
    .A(net1890));
 sg13g2_buf_4 fanout1890 (.X(net1890),
    .A(net1895));
 sg13g2_buf_4 fanout1891 (.X(net1891),
    .A(net1894));
 sg13g2_buf_2 fanout1892 (.A(net1893),
    .X(net1892));
 sg13g2_buf_4 fanout1893 (.X(net1893),
    .A(net1894));
 sg13g2_buf_1 fanout1894 (.A(net1895),
    .X(net1894));
 sg13g2_buf_8 fanout1895 (.A(_01565_),
    .X(net1895));
 sg13g2_buf_2 fanout1896 (.A(net1900),
    .X(net1896));
 sg13g2_buf_2 fanout1897 (.A(net1900),
    .X(net1897));
 sg13g2_buf_4 fanout1898 (.X(net1898),
    .A(net1900));
 sg13g2_buf_1 fanout1899 (.A(net1900),
    .X(net1899));
 sg13g2_buf_1 fanout1900 (.A(net1906),
    .X(net1900));
 sg13g2_buf_2 fanout1901 (.A(net1905),
    .X(net1901));
 sg13g2_buf_2 fanout1902 (.A(net1903),
    .X(net1902));
 sg13g2_buf_2 fanout1903 (.A(net1905),
    .X(net1903));
 sg13g2_buf_2 fanout1904 (.A(net1905),
    .X(net1904));
 sg13g2_buf_2 fanout1905 (.A(net1906),
    .X(net1905));
 sg13g2_buf_2 fanout1906 (.A(net1960),
    .X(net1906));
 sg13g2_buf_2 fanout1907 (.A(net1908),
    .X(net1907));
 sg13g2_buf_2 fanout1908 (.A(net1916),
    .X(net1908));
 sg13g2_buf_2 fanout1909 (.A(net1910),
    .X(net1909));
 sg13g2_buf_2 fanout1910 (.A(net1916),
    .X(net1910));
 sg13g2_buf_2 fanout1911 (.A(net1912),
    .X(net1911));
 sg13g2_buf_2 fanout1912 (.A(net1915),
    .X(net1912));
 sg13g2_buf_2 fanout1913 (.A(net1915),
    .X(net1913));
 sg13g2_buf_2 fanout1914 (.A(net1915),
    .X(net1914));
 sg13g2_buf_2 fanout1915 (.A(net1916),
    .X(net1915));
 sg13g2_buf_2 fanout1916 (.A(net1926),
    .X(net1916));
 sg13g2_buf_2 fanout1917 (.A(net1918),
    .X(net1917));
 sg13g2_buf_2 fanout1918 (.A(net1926),
    .X(net1918));
 sg13g2_buf_4 fanout1919 (.X(net1919),
    .A(net1920));
 sg13g2_buf_4 fanout1920 (.X(net1920),
    .A(net1926));
 sg13g2_buf_2 fanout1921 (.A(net1922),
    .X(net1921));
 sg13g2_buf_2 fanout1922 (.A(net1925),
    .X(net1922));
 sg13g2_buf_2 fanout1923 (.A(net1924),
    .X(net1923));
 sg13g2_buf_4 fanout1924 (.X(net1924),
    .A(net1925));
 sg13g2_buf_2 fanout1925 (.A(net1926),
    .X(net1925));
 sg13g2_buf_2 fanout1926 (.A(net1960),
    .X(net1926));
 sg13g2_buf_2 fanout1927 (.A(net1933),
    .X(net1927));
 sg13g2_buf_2 fanout1928 (.A(net1929),
    .X(net1928));
 sg13g2_buf_2 fanout1929 (.A(net1933),
    .X(net1929));
 sg13g2_buf_2 fanout1930 (.A(net1931),
    .X(net1930));
 sg13g2_buf_4 fanout1931 (.X(net1931),
    .A(net1933));
 sg13g2_buf_1 fanout1932 (.A(net1933),
    .X(net1932));
 sg13g2_buf_2 fanout1933 (.A(net1960),
    .X(net1933));
 sg13g2_buf_2 fanout1934 (.A(net1935),
    .X(net1934));
 sg13g2_buf_2 fanout1935 (.A(net1939),
    .X(net1935));
 sg13g2_buf_2 fanout1936 (.A(net1938),
    .X(net1936));
 sg13g2_buf_4 fanout1937 (.X(net1937),
    .A(net1938));
 sg13g2_buf_2 fanout1938 (.A(net1939),
    .X(net1938));
 sg13g2_buf_2 fanout1939 (.A(net1960),
    .X(net1939));
 sg13g2_buf_4 fanout1940 (.X(net1940),
    .A(net1943));
 sg13g2_buf_2 fanout1941 (.A(net1942),
    .X(net1941));
 sg13g2_buf_2 fanout1942 (.A(net1943),
    .X(net1942));
 sg13g2_buf_2 fanout1943 (.A(net1959),
    .X(net1943));
 sg13g2_buf_2 fanout1944 (.A(net1945),
    .X(net1944));
 sg13g2_buf_2 fanout1945 (.A(net1949),
    .X(net1945));
 sg13g2_buf_2 fanout1946 (.A(net1949),
    .X(net1946));
 sg13g2_buf_2 fanout1947 (.A(net1949),
    .X(net1947));
 sg13g2_buf_2 fanout1948 (.A(net1949),
    .X(net1948));
 sg13g2_buf_2 fanout1949 (.A(net1959),
    .X(net1949));
 sg13g2_buf_2 fanout1950 (.A(net1953),
    .X(net1950));
 sg13g2_buf_2 fanout1951 (.A(net1952),
    .X(net1951));
 sg13g2_buf_2 fanout1952 (.A(net1953),
    .X(net1952));
 sg13g2_buf_2 fanout1953 (.A(net1959),
    .X(net1953));
 sg13g2_buf_2 fanout1954 (.A(net1955),
    .X(net1954));
 sg13g2_buf_2 fanout1955 (.A(net1958),
    .X(net1955));
 sg13g2_buf_2 fanout1956 (.A(net1957),
    .X(net1956));
 sg13g2_buf_2 fanout1957 (.A(net1958),
    .X(net1957));
 sg13g2_buf_2 fanout1958 (.A(net1959),
    .X(net1958));
 sg13g2_buf_2 fanout1959 (.A(net1960),
    .X(net1959));
 sg13g2_buf_8 fanout1960 (.A(net2026),
    .X(net1960));
 sg13g2_buf_2 fanout1961 (.A(net1962),
    .X(net1961));
 sg13g2_buf_2 fanout1962 (.A(net1965),
    .X(net1962));
 sg13g2_buf_2 fanout1963 (.A(net1964),
    .X(net1963));
 sg13g2_buf_2 fanout1964 (.A(net1965),
    .X(net1964));
 sg13g2_buf_1 fanout1965 (.A(net1980),
    .X(net1965));
 sg13g2_buf_4 fanout1966 (.X(net1966),
    .A(net1967));
 sg13g2_buf_4 fanout1967 (.X(net1967),
    .A(net1969));
 sg13g2_buf_4 fanout1968 (.X(net1968),
    .A(net1969));
 sg13g2_buf_2 fanout1969 (.A(net1980),
    .X(net1969));
 sg13g2_buf_4 fanout1970 (.X(net1970),
    .A(net1974));
 sg13g2_buf_1 fanout1971 (.A(net1974),
    .X(net1971));
 sg13g2_buf_4 fanout1972 (.X(net1972),
    .A(net1974));
 sg13g2_buf_2 fanout1973 (.A(net1974),
    .X(net1973));
 sg13g2_buf_2 fanout1974 (.A(net1980),
    .X(net1974));
 sg13g2_buf_2 fanout1975 (.A(net1976),
    .X(net1975));
 sg13g2_buf_2 fanout1976 (.A(net1979),
    .X(net1976));
 sg13g2_buf_2 fanout1977 (.A(net1978),
    .X(net1977));
 sg13g2_buf_4 fanout1978 (.X(net1978),
    .A(net1979));
 sg13g2_buf_2 fanout1979 (.A(net1980),
    .X(net1979));
 sg13g2_buf_2 fanout1980 (.A(net2002),
    .X(net1980));
 sg13g2_buf_4 fanout1981 (.X(net1981),
    .A(net1982));
 sg13g2_buf_2 fanout1982 (.A(net1992),
    .X(net1982));
 sg13g2_buf_2 fanout1983 (.A(net1992),
    .X(net1983));
 sg13g2_buf_2 fanout1984 (.A(net1992),
    .X(net1984));
 sg13g2_buf_2 fanout1985 (.A(net1988),
    .X(net1985));
 sg13g2_buf_2 fanout1986 (.A(net1988),
    .X(net1986));
 sg13g2_buf_2 fanout1987 (.A(net1988),
    .X(net1987));
 sg13g2_buf_2 fanout1988 (.A(net1992),
    .X(net1988));
 sg13g2_buf_2 fanout1989 (.A(net1991),
    .X(net1989));
 sg13g2_buf_2 fanout1990 (.A(net1991),
    .X(net1990));
 sg13g2_buf_2 fanout1991 (.A(net1992),
    .X(net1991));
 sg13g2_buf_2 fanout1992 (.A(net2002),
    .X(net1992));
 sg13g2_buf_4 fanout1993 (.X(net1993),
    .A(net1996));
 sg13g2_buf_4 fanout1994 (.X(net1994),
    .A(net1996));
 sg13g2_buf_2 fanout1995 (.A(net1996),
    .X(net1995));
 sg13g2_buf_2 fanout1996 (.A(net2002),
    .X(net1996));
 sg13g2_buf_2 fanout1997 (.A(net2001),
    .X(net1997));
 sg13g2_buf_2 fanout1998 (.A(net2001),
    .X(net1998));
 sg13g2_buf_2 fanout1999 (.A(net2000),
    .X(net1999));
 sg13g2_buf_2 fanout2000 (.A(net2001),
    .X(net2000));
 sg13g2_buf_2 fanout2001 (.A(net2002),
    .X(net2001));
 sg13g2_buf_2 fanout2002 (.A(net2026),
    .X(net2002));
 sg13g2_buf_4 fanout2003 (.X(net2003),
    .A(net2007));
 sg13g2_buf_2 fanout2004 (.A(net2007),
    .X(net2004));
 sg13g2_buf_4 fanout2005 (.X(net2005),
    .A(net2007));
 sg13g2_buf_2 fanout2006 (.A(net2007),
    .X(net2006));
 sg13g2_buf_2 fanout2007 (.A(net2016),
    .X(net2007));
 sg13g2_buf_4 fanout2008 (.X(net2008),
    .A(net2009));
 sg13g2_buf_2 fanout2009 (.A(net2012),
    .X(net2009));
 sg13g2_buf_2 fanout2010 (.A(net2012),
    .X(net2010));
 sg13g2_buf_4 fanout2011 (.X(net2011),
    .A(net2012));
 sg13g2_buf_2 fanout2012 (.A(net2016),
    .X(net2012));
 sg13g2_buf_2 fanout2013 (.A(net2014),
    .X(net2013));
 sg13g2_buf_2 fanout2014 (.A(net2015),
    .X(net2014));
 sg13g2_buf_4 fanout2015 (.X(net2015),
    .A(net2016));
 sg13g2_buf_2 fanout2016 (.A(net2026),
    .X(net2016));
 sg13g2_buf_2 fanout2017 (.A(net2021),
    .X(net2017));
 sg13g2_buf_1 fanout2018 (.A(net2019),
    .X(net2018));
 sg13g2_buf_2 fanout2019 (.A(net2021),
    .X(net2019));
 sg13g2_buf_2 fanout2020 (.A(net2021),
    .X(net2020));
 sg13g2_buf_2 fanout2021 (.A(net2025),
    .X(net2021));
 sg13g2_buf_2 fanout2022 (.A(net2023),
    .X(net2022));
 sg13g2_buf_2 fanout2023 (.A(net2024),
    .X(net2023));
 sg13g2_buf_1 fanout2024 (.A(net2025),
    .X(net2024));
 sg13g2_buf_2 fanout2025 (.A(net2026),
    .X(net2025));
 sg13g2_buf_4 fanout2026 (.X(net2026),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_tielo tt_um_jamesrosssharp_1bitam_5 (.L_LO(net5));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_leaf_82_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_2 clkbuf_leaf_83_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_2 clkbuf_leaf_84_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_2 clkbuf_leaf_85_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_2 clkbuf_leaf_86_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_2 clkbuf_leaf_87_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_2 clkbuf_leaf_88_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_2 clkbuf_leaf_89_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_2 clkbuf_leaf_90_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_2 clkbuf_leaf_91_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_2 clkbuf_leaf_92_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_2 clkbuf_leaf_93_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_2 clkbuf_leaf_94_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_2 clkbuf_leaf_95_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_2 clkbuf_leaf_96_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_2 clkbuf_leaf_97_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_2 clkbuf_leaf_98_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_2 clkbuf_leaf_99_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_2 clkbuf_leaf_100_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_2 clkbuf_leaf_101_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_2 clkbuf_leaf_102_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_2 clkbuf_leaf_103_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_2 clkbuf_leaf_104_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_2 clkbuf_leaf_105_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_2 clkbuf_leaf_106_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_2 clkbuf_leaf_107_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_2 clkbuf_leaf_108_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_2 clkbuf_leaf_109_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_2 clkbuf_leaf_110_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_2 clkbuf_leaf_111_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_2 clkbuf_leaf_112_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_2 clkbuf_leaf_113_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_2 clkbuf_leaf_114_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_2 clkbuf_leaf_115_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_2 clkbuf_leaf_116_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_2 clkbuf_leaf_117_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_2 clkbuf_leaf_118_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_2 clkbuf_leaf_119_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_2 clkbuf_leaf_120_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_2 clkbuf_leaf_121_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_2 clkbuf_leaf_122_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_2 clkbuf_leaf_123_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_2 clkbuf_leaf_124_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_2 clkbuf_leaf_125_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_2 clkbuf_leaf_126_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_2 clkbuf_leaf_127_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_2 clkbuf_leaf_128_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_2 clkbuf_leaf_129_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_2 clkbuf_leaf_130_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_2 clkbuf_leaf_131_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_2 clkbuf_leaf_132_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_2 clkbuf_leaf_133_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_2 clkbuf_leaf_134_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_2 clkbuf_leaf_135_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_2 clkbuf_leaf_136_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_2 clkbuf_leaf_137_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_2 clkbuf_leaf_138_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_2 clkbuf_leaf_139_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_2 clkbuf_leaf_140_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_2 clkbuf_leaf_141_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_2 clkbuf_leaf_142_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_2 clkbuf_leaf_143_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_2 clkbuf_leaf_145_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkload7 (.A(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkload9 (.A(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkload10 (.A(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkload11 (.A(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkload12 (.A(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkload13 (.A(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkload14 (.A(clknet_5_31__leaf_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_145_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_141_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_127_clk));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_25_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_33_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_116_clk));
 sg13g2_inv_2 clkload21 (.A(clknet_leaf_91_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_125_clk));
 sg13g2_inv_2 clkload23 (.A(clknet_leaf_100_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_62_clk));
 sg13g2_inv_2 clkload25 (.A(clknet_leaf_63_clk));
 sg13g2_inv_2 clkload26 (.A(clknet_leaf_67_clk));
 sg13g2_inv_1 clkload27 (.A(clknet_leaf_75_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_00074_),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold2 (.A(_00075_),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold3 (.A(_00076_),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold4 (.A(_00078_),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold5 (.A(_01674_),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold6 (.A(\am_sdr0.mix0.cos_q[0] ),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold7 (.A(\am_sdr0.mix0.sin_q[0] ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold8 (.A(_00077_),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold9 (.A(_00125_),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold10 (.A(_00022_),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold11 (.A(_00164_),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold12 (.A(_00073_),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold13 (.A(_05494_),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold14 (.A(_01102_),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold15 (.A(\am_sdr0.cos[5] ),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold16 (.A(\am_sdr0.mix0.sin_in[4] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold17 (.A(\am_sdr0.spi0.MOSI_q ),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold18 (.A(\am_sdr0.cos[1] ),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold19 (.A(\am_sdr0.spi0.CS_q ),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold20 (.A(\am_sdr0.mix0.sin_in[7] ),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold21 (.A(\am_sdr0.spi0.SCK_q ),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold22 (.A(\am_sdr0.mix0.sin_in[1] ),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold23 (.A(\am_sdr0.mix0.sin_in[6] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold24 (.A(\am_sdr0.cos[0] ),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold25 (.A(\am_sdr0.mix0.sin_in[5] ),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold26 (.A(\am_sdr0.mix0.sin_in[2] ),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold27 (.A(\am_sdr0.mix0.sin_in[0] ),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold28 (.A(\am_sdr0.mix0.sin_in[3] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold29 (.A(\am_sdr0.cos[6] ),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold30 (.A(\am_sdr0.cos[7] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold31 (.A(\am_sdr0.cos[2] ),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold32 (.A(\am_sdr0.cos[3] ),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold33 (.A(\am_sdr0.spi0.SCK_qq ),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold34 (.A(\am_sdr0.mix0.sin_q[7] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold35 (.A(_00036_),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold36 (.A(\am_sdr0.mix0.sin_q[5] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold37 (.A(_00034_),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold38 (.A(\am_sdr0.am0.r[6] ),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold39 (.A(_02110_),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold40 (.A(\am_sdr0.cic1.count[2] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold41 (.A(_04364_),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold42 (.A(_00784_),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold43 (.A(\am_sdr0.mix0.RF_in_q ),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold44 (.A(\am_sdr0.mix0.sin_q[6] ),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold45 (.A(_00035_),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold46 (.A(\am_sdr0.cic1.count[7] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold47 (.A(_00789_),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold48 (.A(\am_sdr0.am0.r[2] ),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold49 (.A(_02106_),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold50 (.A(\am_sdr0.am0.r[0] ),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold51 (.A(_02104_),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold52 (.A(\am_sdr0.cos[4] ),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold53 (.A(\am_sdr0.mix0.cos_q[7] ),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold54 (.A(_00029_),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold55 (.A(\am_sdr0.am0.r[1] ),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold56 (.A(_02105_),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold57 (.A(\am_sdr0.cic0.count[2] ),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold58 (.A(_05198_),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold59 (.A(_01008_),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold60 (.A(\am_sdr0.am0.r[3] ),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold61 (.A(_02107_),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold62 (.A(\am_sdr0.am0.r[4] ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold63 (.A(_02108_),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold64 (.A(\am_sdr0.cic1.comb3[15] ),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold65 (.A(_00668_),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold66 (.A(\am_sdr0.cic2.count[1] ),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold67 (.A(_03391_),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold68 (.A(_00548_),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold69 (.A(\am_sdr0.cic2.comb3[12] ),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold70 (.A(_00431_),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold71 (.A(\am_sdr0.am0.left[0] ),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold72 (.A(_01939_),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold73 (.A(\am_sdr0.spi0.shift_reg[28] ),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold74 (.A(_00888_),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold75 (.A(\am_sdr0.mix0.cos_q[5] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold76 (.A(_00027_),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold77 (.A(\am_sdr0.am0.a[1] ),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold78 (.A(_02032_),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold79 (.A(\am_sdr0.cic1.comb3[14] ),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold80 (.A(_00667_),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold81 (.A(\am_sdr0.cic3.count[1] ),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold82 (.A(_02520_),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold83 (.A(_00333_),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold84 (.A(\am_sdr0.cic2.comb3[18] ),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold85 (.A(_00437_),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold86 (.A(\am_sdr0.am0.a[0] ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold87 (.A(_02031_),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold88 (.A(\am_sdr0.mix0.sin_q[3] ),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold89 (.A(_00032_),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold90 (.A(\am_sdr0.cic0.count[7] ),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold91 (.A(_01013_),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold92 (.A(\am_sdr0.am0.count2[2] ),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold93 (.A(_00127_),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold94 (.A(\am_sdr0.am0.count[1] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold95 (.A(_01934_),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold96 (.A(\am_sdr0.am0.state[6] ),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold97 (.A(_00018_),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold98 (.A(\am_sdr0.am0.state[3] ),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold99 (.A(_01601_),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold100 (.A(\am_sdr0.cic2.comb3[16] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold101 (.A(_00435_),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold102 (.A(\am_sdr0.cic1.comb3[18] ),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold103 (.A(_00671_),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold104 (.A(\am_sdr0.mix0.cos_q[4] ),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold105 (.A(_01653_),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold106 (.A(_00026_),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold107 (.A(\am_sdr0.cic0.comb3[16] ),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold108 (.A(_00893_),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold109 (.A(\am_sdr0.spi0.shift_reg[2] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold110 (.A(_01109_),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold111 (.A(\am_sdr0.am0.state[0] ),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold112 (.A(_00016_),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold113 (.A(\am_sdr0.am0.state[4] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold114 (.A(_01600_),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold115 (.A(\am_sdr0.cic3.integ1[0] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold116 (.A(_02529_),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold117 (.A(_00340_),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold118 (.A(\am_sdr0.cic2.integ1[0] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold119 (.A(_03400_),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold120 (.A(_00555_),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold121 (.A(\am_sdr0.cic1.comb3[12] ),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold122 (.A(_00665_),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold123 (.A(\am_sdr0.cic2.comb3[17] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold124 (.A(_00436_),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold125 (.A(\am_sdr0.cic2.comb3[19] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold126 (.A(_00438_),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold127 (.A(\am_sdr0.spi0.shift_reg[19] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold128 (.A(_00879_),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold129 (.A(\am_sdr0.spi0.shift_reg[4] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold130 (.A(_01111_),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold131 (.A(\am_sdr0.cic0.comb3[18] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold132 (.A(_00895_),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold133 (.A(\am_sdr0.cic2.comb3[14] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold134 (.A(_00433_),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold135 (.A(\am_sdr0.cic3.integ1[25] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold136 (.A(\am_sdr0.spi0.shift_reg[13] ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold137 (.A(_00873_),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold138 (.A(\am_sdr0.cic2.integ2[0] ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold139 (.A(_03560_),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold140 (.A(\am_sdr0.spi0.MOSI_qq ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold141 (.A(_00860_),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold142 (.A(\am_sdr0.am0.a[15] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold143 (.A(_02103_),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold144 (.A(\am_sdr0.cic0.comb3[17] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold145 (.A(_00894_),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold146 (.A(\am_sdr0.am0.a[14] ),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold147 (.A(\am_sdr0.cic0.integ3[19] ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold148 (.A(_00664_),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold149 (.A(\am_sdr0.mix0.cos_q[3] ),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold150 (.A(_00025_),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold151 (.A(\am_sdr0.am0.r[5] ),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold152 (.A(_02109_),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold153 (.A(\am_sdr0.spi0.shift_reg[10] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold154 (.A(_00870_),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold155 (.A(\am_sdr0.am0.a[10] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold156 (.A(_00148_),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold157 (.A(\am_sdr0.cic3.comb3[16] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold158 (.A(_00220_),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold159 (.A(\am_sdr0.cic3.integ2[0] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold160 (.A(_02688_),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold161 (.A(\am_sdr0.am0.q[7] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold162 (.A(_02120_),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold163 (.A(\am_sdr0.spi0.shift_reg[3] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold164 (.A(\am_sdr0.mix0.sin_q[4] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold165 (.A(_00033_),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold166 (.A(\am_sdr0.cic2.count[7] ),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold167 (.A(_00554_),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold168 (.A(\am_sdr0.spi0.shift_reg[5] ),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold169 (.A(_00865_),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold170 (.A(\am_sdr0.cic3.comb3[19] ),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold171 (.A(_00223_),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold172 (.A(\am_sdr0.cic1.integ3[6] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold173 (.A(_00417_),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold174 (.A(_00051_),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold175 (.A(\am_sdr0.cic1.comb3[13] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold176 (.A(_00666_),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold177 (.A(\am_sdr0.cic0.comb3[13] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold178 (.A(_00890_),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold179 (.A(\am_sdr0.spi0.state[1] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold180 (.A(_04748_),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold181 (.A(\am_sdr0.spi0.shift_reg[24] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold182 (.A(_00884_),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold183 (.A(\am_sdr0.spi0.shift_reg[14] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold184 (.A(_01121_),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold185 (.A(\am_sdr0.cic1.comb3[17] ),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold186 (.A(_00670_),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold187 (.A(\am_sdr0.cic3.comb3[17] ),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold188 (.A(_00221_),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold189 (.A(\am_sdr0.cic2.integ1[25] ),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold190 (.A(\am_sdr0.am0.r[7] ),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold191 (.A(_02111_),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold192 (.A(\am_sdr0.nco0.phase_inc[13] ),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold193 (.A(\am_sdr0.cic3.comb3[18] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold194 (.A(_00222_),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold195 (.A(\am_sdr0.spi0.state[0] ),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold196 (.A(\am_sdr0.am0.a[12] ),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold197 (.A(_00150_),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold198 (.A(\am_sdr0.spi0.shift_reg[17] ),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold199 (.A(_00877_),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold200 (.A(\am_sdr0.spi0.shift_reg[12] ),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold201 (.A(_00872_),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold202 (.A(\am_sdr0.am0.right[6] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold203 (.A(_02117_),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold204 (.A(\am_sdr0.cic1.comb3[16] ),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold205 (.A(_00669_),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold206 (.A(\am_sdr0.cic0.comb3[19] ),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold207 (.A(\am_sdr0.cic2.comb3[13] ),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold208 (.A(_00432_),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold209 (.A(\am_sdr0.am0.demod_out[15] ),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold210 (.A(\am_sdr0.cic1.count[6] ),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold211 (.A(_04368_),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold212 (.A(_00788_),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold213 (.A(\am_sdr0.cic3.count[7] ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold214 (.A(_00339_),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold215 (.A(\am_sdr0.am0.a[13] ),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold216 (.A(_02073_),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold217 (.A(\am_sdr0.cic1.integ3[19] ),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold218 (.A(_00430_),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold219 (.A(\am_sdr0.spi0.shift_reg[20] ),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold220 (.A(\am_sdr0.spi0.shift_reg[9] ),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold221 (.A(_00869_),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold222 (.A(\am_sdr0.cic2.integ_sample[14] ),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold223 (.A(_00210_),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold224 (.A(\am_sdr0.am0.a[2] ),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold225 (.A(_00140_),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold226 (.A(\am_sdr0.spi0.shift_reg[1] ),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold227 (.A(\am_sdr0.cic1.integ3[1] ),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold228 (.A(_00412_),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold229 (.A(\am_sdr0.nco0.phase_inc[10] ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold230 (.A(\am_sdr0.am0.left[6] ),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold231 (.A(\am_sdr0.spi0.shift_reg[16] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold232 (.A(_00876_),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold233 (.A(\am_sdr0.am0.right[4] ),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold234 (.A(_02115_),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold235 (.A(\am_sdr0.cic2.count[0] ),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold236 (.A(\am_sdr0.cic1.integ3[13] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold237 (.A(_00424_),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold238 (.A(\am_sdr0.cic0.integ3[6] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold239 (.A(_00651_),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold240 (.A(\am_sdr0.am0.demod_out[9] ),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold241 (.A(_05735_),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold242 (.A(\am_sdr0.spi0.CS_qq ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold243 (.A(_01133_),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold244 (.A(\am_sdr0.cic1.integ3[18] ),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold245 (.A(_00429_),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold246 (.A(\am_sdr0.spi0.shift_reg[6] ),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold247 (.A(\am_sdr0.spi0.shift_reg[11] ),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold248 (.A(\am_sdr0.cic0.count[6] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold249 (.A(_05202_),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold250 (.A(_01012_),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold251 (.A(\am_sdr0.am0.a[8] ),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold252 (.A(_00146_),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold253 (.A(\am_sdr0.spi0.shift_reg[23] ),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold254 (.A(_00883_),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold255 (.A(\am_sdr0.nco0.phase_inc[23] ),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold256 (.A(\am_sdr0.spi0.shift_reg[7] ),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold257 (.A(\am_sdr0.spi0.shift_reg[21] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold258 (.A(\am_sdr0.spi0.shift_reg[15] ),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold259 (.A(_01122_),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold260 (.A(\am_sdr0.spi0.shift_reg[8] ),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold261 (.A(\am_sdr0.cic1.integ3[9] ),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold262 (.A(_00420_),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold263 (.A(\am_sdr0.cic0.count[4] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold264 (.A(_05200_),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold265 (.A(\am_sdr0.am0.multB[7] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold266 (.A(_00089_),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold267 (.A(\am_sdr0.cic1.count[4] ),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold268 (.A(_04366_),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold269 (.A(\am_sdr0.am0.sum[0] ),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold270 (.A(_00108_),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold271 (.A(\am_sdr0.cic0.integ3[3] ),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold272 (.A(_00648_),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold273 (.A(\am_sdr0.am0.q[6] ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold274 (.A(_02119_),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold275 (.A(\am_sdr0.cic0.integ3[8] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold276 (.A(_00653_),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold277 (.A(\am_sdr0.cic1.count[3] ),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold278 (.A(_04365_),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold279 (.A(\am_sdr0.cic1.integ3[7] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold280 (.A(_00418_),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold281 (.A(\am_sdr0.cic0.integ3[9] ),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold282 (.A(_00654_),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold283 (.A(\am_sdr0.mix0.cos_q[2] ),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold284 (.A(_01648_),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold285 (.A(_00024_),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold286 (.A(\am_sdr0.am0.a[9] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold287 (.A(_00147_),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold288 (.A(\am_sdr0.cic2.comb3[15] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold289 (.A(_00434_),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold290 (.A(\am_sdr0.cic3.comb3[14] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold291 (.A(_00218_),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold292 (.A(\am_sdr0.nco0.phase_inc[21] ),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold293 (.A(\am_sdr0.spi0.shift_reg[22] ),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold294 (.A(\am_sdr0.am0.a[5] ),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold295 (.A(_00143_),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold296 (.A(\am_sdr0.am0.a[3] ),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold297 (.A(_00141_),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold298 (.A(\am_sdr0.mix0.sin_q[2] ),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold299 (.A(_00031_),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold300 (.A(\am_sdr0.cic3.comb3[15] ),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold301 (.A(_00219_),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold302 (.A(\am_sdr0.cic2.integ3[0] ),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold303 (.A(_03711_),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold304 (.A(\am_sdr0.cic2.comb2[0] ),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold305 (.A(_00527_),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold306 (.A(\am_sdr0.am0.a[11] ),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold307 (.A(_02067_),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold308 (.A(\am_sdr0.spi0.shift_reg[0] ),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold309 (.A(\am_sdr0.am0.sqrt_done ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold310 (.A(_02100_),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold311 (.A(_00174_),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold312 (.A(\am_sdr0.am0.right[2] ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold313 (.A(_02113_),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold314 (.A(\am_sdr0.cic1.integ3[8] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold315 (.A(_00419_),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold316 (.A(\am_sdr0.cic0.comb3[14] ),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold317 (.A(_00891_),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold318 (.A(\am_sdr0.am0.sum[12] ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold319 (.A(\am_sdr0.nco0.phase_inc[19] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold320 (.A(\am_sdr0.spi0.shift_reg[27] ),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold321 (.A(_00887_),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold322 (.A(\am_sdr0.cic1.comb3[19] ),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold323 (.A(_00672_),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold324 (.A(\am_sdr0.cic2.integ_sample[19] ),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold325 (.A(_00478_),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold326 (.A(\am_sdr0.am0.q[5] ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold327 (.A(_02118_),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold328 (.A(\am_sdr0.cic3.count[0] ),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold329 (.A(\am_sdr0.am0.a[7] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold330 (.A(_00145_),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold331 (.A(\am_sdr0.am0.multB[3] ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold332 (.A(_00085_),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold333 (.A(\am_sdr0.cic0.comb3[15] ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold334 (.A(_00892_),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold335 (.A(\am_sdr0.cic1.integ3[10] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold336 (.A(_00421_),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold337 (.A(\am_sdr0.cic0.integ3[2] ),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold338 (.A(_00647_),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold339 (.A(\am_sdr0.cic0.integ3[4] ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold340 (.A(_00649_),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold341 (.A(\am_sdr0.cic0.comb3[12] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold342 (.A(_00889_),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold343 (.A(\am_sdr0.mix0.sin_q[1] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold344 (.A(\am_sdr0.nco0.phase_inc[8] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold345 (.A(\am_sdr0.nco0.phase_inc[11] ),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold346 (.A(\am_sdr0.am0.a[6] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold347 (.A(_00144_),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold348 (.A(\am_sdr0.am0.multB[5] ),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold349 (.A(_00087_),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold350 (.A(\am_sdr0.cic0.integ3[10] ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold351 (.A(_00655_),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold352 (.A(\am_sdr0.cic0.integ3[18] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold353 (.A(_00663_),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold354 (.A(\am_sdr0.cic3.comb3[12] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold355 (.A(_00216_),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold356 (.A(\am_sdr0.cic0.integ3[16] ),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold357 (.A(_00661_),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold358 (.A(\am_sdr0.am0.multB[4] ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold359 (.A(_00086_),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold360 (.A(\am_sdr0.am0.q[3] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold361 (.A(_05737_),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold362 (.A(\am_sdr0.am0.right[5] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold363 (.A(_00037_),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold364 (.A(_01608_),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold365 (.A(_00007_),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold366 (.A(\am_sdr0.cic3.comb2[0] ),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold367 (.A(_00312_),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold368 (.A(\am_sdr0.am0.a[4] ),
    .X(net2027));
 sg13g2_dlygate4sd3_1 hold369 (.A(_00142_),
    .X(net2028));
 sg13g2_dlygate4sd3_1 hold370 (.A(\am_sdr0.cic1.comb3_in_del[17] ),
    .X(net2029));
 sg13g2_dlygate4sd3_1 hold371 (.A(_04330_),
    .X(net2030));
 sg13g2_dlygate4sd3_1 hold372 (.A(_00758_),
    .X(net2031));
 sg13g2_dlygate4sd3_1 hold373 (.A(\am_sdr0.am0.sum[15] ),
    .X(net2032));
 sg13g2_dlygate4sd3_1 hold374 (.A(\am_sdr0.cic0.count[3] ),
    .X(net2033));
 sg13g2_dlygate4sd3_1 hold375 (.A(_05199_),
    .X(net2034));
 sg13g2_dlygate4sd3_1 hold376 (.A(\am_sdr0.cic1.comb1_in_del[0] ),
    .X(net2035));
 sg13g2_dlygate4sd3_1 hold377 (.A(_00693_),
    .X(net2036));
 sg13g2_dlygate4sd3_1 hold378 (.A(\am_sdr0.am0.multB[6] ),
    .X(net2037));
 sg13g2_dlygate4sd3_1 hold379 (.A(_00088_),
    .X(net2038));
 sg13g2_dlygate4sd3_1 hold380 (.A(\am_sdr0.cic2.comb2[17] ),
    .X(net2039));
 sg13g2_dlygate4sd3_1 hold381 (.A(_03357_),
    .X(net2040));
 sg13g2_dlygate4sd3_1 hold382 (.A(_03359_),
    .X(net2041));
 sg13g2_dlygate4sd3_1 hold383 (.A(_00524_),
    .X(net2042));
 sg13g2_dlygate4sd3_1 hold384 (.A(\am_sdr0.spi0.shift_reg[18] ),
    .X(net2043));
 sg13g2_dlygate4sd3_1 hold385 (.A(_01125_),
    .X(net2044));
 sg13g2_dlygate4sd3_1 hold386 (.A(\am_sdr0.cic3.comb2[1] ),
    .X(net2045));
 sg13g2_dlygate4sd3_1 hold387 (.A(_00313_),
    .X(net2046));
 sg13g2_dlygate4sd3_1 hold388 (.A(\am_sdr0.am0.demod_out[14] ),
    .X(net2047));
 sg13g2_dlygate4sd3_1 hold389 (.A(\am_sdr0.am0.multB[2] ),
    .X(net2048));
 sg13g2_dlygate4sd3_1 hold390 (.A(_00084_),
    .X(net2049));
 sg13g2_dlygate4sd3_1 hold391 (.A(\am_sdr0.mix0.cos_q[6] ),
    .X(net2050));
 sg13g2_dlygate4sd3_1 hold392 (.A(_00028_),
    .X(net2051));
 sg13g2_dlygate4sd3_1 hold393 (.A(\am_sdr0.cic0.integ3[5] ),
    .X(net2052));
 sg13g2_dlygate4sd3_1 hold394 (.A(_00650_),
    .X(net2053));
 sg13g2_dlygate4sd3_1 hold395 (.A(\am_sdr0.nco0.phase_inc[0] ),
    .X(net2054));
 sg13g2_dlygate4sd3_1 hold396 (.A(\am_sdr0.cic0.integ3[7] ),
    .X(net2055));
 sg13g2_dlygate4sd3_1 hold397 (.A(_00652_),
    .X(net2056));
 sg13g2_dlygate4sd3_1 hold398 (.A(\am_sdr0.cic2.comb2[19] ),
    .X(net2057));
 sg13g2_dlygate4sd3_1 hold399 (.A(_03367_),
    .X(net2058));
 sg13g2_dlygate4sd3_1 hold400 (.A(_03368_),
    .X(net2059));
 sg13g2_dlygate4sd3_1 hold401 (.A(_00526_),
    .X(net2060));
 sg13g2_dlygate4sd3_1 hold402 (.A(\am_sdr0.cic1.comb2[19] ),
    .X(net2061));
 sg13g2_dlygate4sd3_1 hold403 (.A(_00780_),
    .X(net2062));
 sg13g2_dlygate4sd3_1 hold404 (.A(\am_sdr0.cic2.count[6] ),
    .X(net2063));
 sg13g2_dlygate4sd3_1 hold405 (.A(_03397_),
    .X(net2064));
 sg13g2_dlygate4sd3_1 hold406 (.A(_00553_),
    .X(net2065));
 sg13g2_dlygate4sd3_1 hold407 (.A(\am_sdr0.cic2.integ_sample[11] ),
    .X(net2066));
 sg13g2_dlygate4sd3_1 hold408 (.A(_00470_),
    .X(net2067));
 sg13g2_dlygate4sd3_1 hold409 (.A(\am_sdr0.cic2.comb1_in_del[0] ),
    .X(net2068));
 sg13g2_dlygate4sd3_1 hold410 (.A(_00459_),
    .X(net2069));
 sg13g2_dlygate4sd3_1 hold411 (.A(\am_sdr0.cic1.integ3[3] ),
    .X(net2070));
 sg13g2_dlygate4sd3_1 hold412 (.A(_00414_),
    .X(net2071));
 sg13g2_dlygate4sd3_1 hold413 (.A(\am_sdr0.cic1.integ1[21] ),
    .X(net2072));
 sg13g2_dlygate4sd3_1 hold414 (.A(_04606_),
    .X(net2073));
 sg13g2_dlygate4sd3_1 hold415 (.A(\am_sdr0.cic0.comb2[1] ),
    .X(net2074));
 sg13g2_dlygate4sd3_1 hold416 (.A(_00986_),
    .X(net2075));
 sg13g2_dlygate4sd3_1 hold417 (.A(\am_sdr0.nco0.phase_inc[9] ),
    .X(net2076));
 sg13g2_dlygate4sd3_1 hold418 (.A(\am_sdr0.cic2.integ_sample[10] ),
    .X(net2077));
 sg13g2_dlygate4sd3_1 hold419 (.A(_00469_),
    .X(net2078));
 sg13g2_dlygate4sd3_1 hold420 (.A(\am_sdr0.cic0.comb3_in_del[3] ),
    .X(net2079));
 sg13g2_dlygate4sd3_1 hold421 (.A(_00988_),
    .X(net2080));
 sg13g2_dlygate4sd3_1 hold422 (.A(\am_sdr0.cic1.integ3[2] ),
    .X(net2081));
 sg13g2_dlygate4sd3_1 hold423 (.A(_00413_),
    .X(net2082));
 sg13g2_dlygate4sd3_1 hold424 (.A(\am_sdr0.cic2.comb2[1] ),
    .X(net2083));
 sg13g2_dlygate4sd3_1 hold425 (.A(_00528_),
    .X(net2084));
 sg13g2_dlygate4sd3_1 hold426 (.A(\am_sdr0.cic1.integ3[5] ),
    .X(net2085));
 sg13g2_dlygate4sd3_1 hold427 (.A(_00416_),
    .X(net2086));
 sg13g2_dlygate4sd3_1 hold428 (.A(\am_sdr0.cic1.comb3_in_del[10] ),
    .X(net2087));
 sg13g2_dlygate4sd3_1 hold429 (.A(_00771_),
    .X(net2088));
 sg13g2_dlygate4sd3_1 hold430 (.A(\am_sdr0.cic3.comb3_in_del[2] ),
    .X(net2089));
 sg13g2_dlygate4sd3_1 hold431 (.A(_00314_),
    .X(net2090));
 sg13g2_dlygate4sd3_1 hold432 (.A(\am_sdr0.nco0.phase_inc[7] ),
    .X(net2091));
 sg13g2_dlygate4sd3_1 hold433 (.A(\am_sdr0.cic0.comb2[13] ),
    .X(net2092));
 sg13g2_dlygate4sd3_1 hold434 (.A(\am_sdr0.nco0.phase_inc[17] ),
    .X(net2093));
 sg13g2_dlygate4sd3_1 hold435 (.A(\am_sdr0.cic3.count[6] ),
    .X(net2094));
 sg13g2_dlygate4sd3_1 hold436 (.A(_02526_),
    .X(net2095));
 sg13g2_dlygate4sd3_1 hold437 (.A(_00338_),
    .X(net2096));
 sg13g2_dlygate4sd3_1 hold438 (.A(\am_sdr0.am0.count2[3] ),
    .X(net2097));
 sg13g2_dlygate4sd3_1 hold439 (.A(_00128_),
    .X(net2098));
 sg13g2_dlygate4sd3_1 hold440 (.A(\am_sdr0.am0.sum[4] ),
    .X(net2099));
 sg13g2_dlygate4sd3_1 hold441 (.A(_01778_),
    .X(net2100));
 sg13g2_dlygate4sd3_1 hold442 (.A(\am_sdr0.am0.demod_out[13] ),
    .X(net2101));
 sg13g2_dlygate4sd3_1 hold443 (.A(\am_sdr0.cic1.comb3_in_del[5] ),
    .X(net2102));
 sg13g2_dlygate4sd3_1 hold444 (.A(_00766_),
    .X(net2103));
 sg13g2_dlygate4sd3_1 hold445 (.A(\am_sdr0.cic2.comb2[15] ),
    .X(net2104));
 sg13g2_dlygate4sd3_1 hold446 (.A(_03339_),
    .X(net2105));
 sg13g2_dlygate4sd3_1 hold447 (.A(_03343_),
    .X(net2106));
 sg13g2_dlygate4sd3_1 hold448 (.A(\am_sdr0.cic0.comb1[7] ),
    .X(net2107));
 sg13g2_dlygate4sd3_1 hold449 (.A(_00964_),
    .X(net2108));
 sg13g2_dlygate4sd3_1 hold450 (.A(\am_sdr0.cic0.integ3[14] ),
    .X(net2109));
 sg13g2_dlygate4sd3_1 hold451 (.A(_00659_),
    .X(net2110));
 sg13g2_dlygate4sd3_1 hold452 (.A(\am_sdr0.cic2.comb3_in_del[2] ),
    .X(net2111));
 sg13g2_dlygate4sd3_1 hold453 (.A(_00529_),
    .X(net2112));
 sg13g2_dlygate4sd3_1 hold454 (.A(\am_sdr0.spi0.CS_qqq ),
    .X(net2113));
 sg13g2_dlygate4sd3_1 hold455 (.A(\am_sdr0.cic1.integ3[11] ),
    .X(net2114));
 sg13g2_dlygate4sd3_1 hold456 (.A(_00422_),
    .X(net2115));
 sg13g2_dlygate4sd3_1 hold457 (.A(\am_sdr0.cic3.integ3[0] ),
    .X(net2116));
 sg13g2_dlygate4sd3_1 hold458 (.A(_02846_),
    .X(net2117));
 sg13g2_dlygate4sd3_1 hold459 (.A(\am_sdr0.am0.sqrt_state[0] ),
    .X(net2118));
 sg13g2_dlygate4sd3_1 hold460 (.A(\am_sdr0.cic1.comb1[19] ),
    .X(net2119));
 sg13g2_dlygate4sd3_1 hold461 (.A(_00752_),
    .X(net2120));
 sg13g2_dlygate4sd3_1 hold462 (.A(\am_sdr0.cic0.comb1_in_del[0] ),
    .X(net2121));
 sg13g2_dlygate4sd3_1 hold463 (.A(_00917_),
    .X(net2122));
 sg13g2_dlygate4sd3_1 hold464 (.A(\am_sdr0.cic0.comb1[19] ),
    .X(net2123));
 sg13g2_dlygate4sd3_1 hold465 (.A(_00976_),
    .X(net2124));
 sg13g2_dlygate4sd3_1 hold466 (.A(\am_sdr0.cic2.comb3_in_del[3] ),
    .X(net2125));
 sg13g2_dlygate4sd3_1 hold467 (.A(_00530_),
    .X(net2126));
 sg13g2_dlygate4sd3_1 hold468 (.A(\am_sdr0.am0.q[2] ),
    .X(net2127));
 sg13g2_dlygate4sd3_1 hold469 (.A(_05736_),
    .X(net2128));
 sg13g2_dlygate4sd3_1 hold470 (.A(\am_sdr0.nco0.phase_inc[22] ),
    .X(net2129));
 sg13g2_dlygate4sd3_1 hold471 (.A(\am_sdr0.nco0.phase[24] ),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold472 (.A(\am_sdr0.cic0.comb3_in_del[2] ),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold473 (.A(_00987_),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold474 (.A(\am_sdr0.cic0.comb2[19] ),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold475 (.A(_05173_),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold476 (.A(_00984_),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold477 (.A(\am_sdr0.nco0.phase[0] ),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold478 (.A(\am_sdr0.cic2.integ_sample[3] ),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold479 (.A(_00199_),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold480 (.A(\am_sdr0.am0.q[1] ),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold481 (.A(_02114_),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold482 (.A(\am_sdr0.cic1.integ_sample[19] ),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold483 (.A(_00712_),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold484 (.A(\am_sdr0.cic0.comb3_in_del[15] ),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold485 (.A(_05149_),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold486 (.A(\am_sdr0.cic1.comb2[18] ),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold487 (.A(_00779_),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold488 (.A(\am_sdr0.cic1.comb2[16] ),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold489 (.A(_00777_),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold490 (.A(\am_sdr0.cic3.comb3[13] ),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold491 (.A(_00217_),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold492 (.A(\am_sdr0.cic2.integ_sample[8] ),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold493 (.A(_00467_),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold494 (.A(\am_sdr0.cic0.comb3_in_del[15] ),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold495 (.A(_05158_),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold496 (.A(\am_sdr0.cic3.comb3_in_del[7] ),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold497 (.A(_00319_),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold498 (.A(\am_sdr0.cic1.integ3[16] ),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold499 (.A(_00427_),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold500 (.A(\am_sdr0.cic1.integ3[4] ),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold501 (.A(_00415_),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold502 (.A(\am_sdr0.spi0.shift_reg[25] ),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold503 (.A(\am_sdr0.am0.m_count[1] ),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold504 (.A(_01675_),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold505 (.A(_00080_),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold506 (.A(\am_sdr0.cic0.comb3_in_del[19] ),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold507 (.A(\am_sdr0.cic1.comb2[0] ),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold508 (.A(_00761_),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold509 (.A(\am_sdr0.am0.q[4] ),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold510 (.A(_05738_),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold511 (.A(\am_sdr0.cic0.comb2[0] ),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold512 (.A(_00985_),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold513 (.A(\am_sdr0.cic2.comb2[9] ),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold514 (.A(_00536_),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold515 (.A(\am_sdr0.cic1.count[1] ),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold516 (.A(_04363_),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold517 (.A(\am_sdr0.cic1.integ3[15] ),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold518 (.A(_00426_),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold519 (.A(\am_sdr0.cic1.comb3_in_del[19] ),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold520 (.A(_04341_),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold521 (.A(_00760_),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold522 (.A(\am_sdr0.cic3.comb3_in_del[9] ),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold523 (.A(_00321_),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold524 (.A(\am_sdr0.cic1.comb3_in_del[3] ),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold525 (.A(_00764_),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold526 (.A(\am_sdr0.cic1.integ1[0] ),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold527 (.A(_04372_),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold528 (.A(_00790_),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold529 (.A(\am_sdr0.cic3.comb2[3] ),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold530 (.A(\am_sdr0.cic1.comb3_in_del[2] ),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold531 (.A(_00763_),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold532 (.A(\am_sdr0.cic3.comb2[19] ),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold533 (.A(_00331_),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold534 (.A(\am_sdr0.nco0.phase_inc[5] ),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold535 (.A(\am_sdr0.cic3.integ_sample[19] ),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold536 (.A(_01082_),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold537 (.A(\am_sdr0.cic1.integ2[0] ),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold538 (.A(_04511_),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold539 (.A(\am_sdr0.cic3.comb1_in_del[19] ),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold540 (.A(\am_sdr0.cic3.comb3_in_del[6] ),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold541 (.A(_00318_),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold542 (.A(\am_sdr0.cic0.comb2[18] ),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold543 (.A(_05168_),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold544 (.A(\am_sdr0.cic3.comb2[17] ),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold545 (.A(_00329_),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold546 (.A(\am_sdr0.cic0.integ3[13] ),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold547 (.A(_00658_),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold548 (.A(\am_sdr0.cic1.comb3_in_del[9] ),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold549 (.A(_00770_),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold550 (.A(\am_sdr0.am0.sum[16] ),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold551 (.A(\am_sdr0.cic3.comb3_in_del[8] ),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold552 (.A(_00320_),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold553 (.A(\am_sdr0.cic0.comb2[10] ),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold554 (.A(\am_sdr0.cic3.comb2[11] ),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold555 (.A(_00323_),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold556 (.A(\am_sdr0.cic3.comb3_in_del[3] ),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold557 (.A(\am_sdr0.cic0.comb1_in_del[13] ),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold558 (.A(_00930_),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold559 (.A(\am_sdr0.cic0.comb3_in_del[16] ),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold560 (.A(_05165_),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold561 (.A(\am_sdr0.nco0.phase_inc[24] ),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold562 (.A(\am_sdr0.cic0.comb1[3] ),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold563 (.A(\am_sdr0.cic2.comb1[4] ),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold564 (.A(_00503_),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold565 (.A(\am_sdr0.cic0.comb3_in_del[9] ),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold566 (.A(_00994_),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold567 (.A(\am_sdr0.cic2.integ_sample[15] ),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold568 (.A(_00211_),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold569 (.A(\am_sdr0.cic3.comb2[4] ),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold570 (.A(_00316_),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold571 (.A(\am_sdr0.cic3.integ3[18] ),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold572 (.A(_01081_),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold573 (.A(\am_sdr0.cic3.comb2[5] ),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold574 (.A(_00317_),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold575 (.A(\am_sdr0.cic2.integ_sample[17] ),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold576 (.A(_00213_),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold577 (.A(\am_sdr0.cic3.comb1[11] ),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold578 (.A(_00295_),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold579 (.A(\am_sdr0.cic3.comb1[2] ),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold580 (.A(_00286_),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold581 (.A(\am_sdr0.cic0.integ3[11] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold582 (.A(_00656_),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold583 (.A(\am_sdr0.cic1.comb2_in_del[11] ),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold584 (.A(_00744_),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold585 (.A(\am_sdr0.nco0.phase_inc[6] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold586 (.A(\am_sdr0.cic2.comb1[18] ),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold587 (.A(_00517_),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold588 (.A(\am_sdr0.am0.sum[8] ),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold589 (.A(_00116_),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold590 (.A(\am_sdr0.cic2.comb3_in_del[6] ),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold591 (.A(_00533_),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold592 (.A(\am_sdr0.cic2.comb1[11] ),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold593 (.A(_00510_),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold594 (.A(\am_sdr0.cic0.count[1] ),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold595 (.A(_05197_),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold596 (.A(\am_sdr0.mix0.cos_q[1] ),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold597 (.A(\am_sdr0.cic1.comb2[17] ),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold598 (.A(_04329_),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold599 (.A(_04334_),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold600 (.A(_04336_),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold601 (.A(\am_sdr0.cic3.comb1[0] ),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold602 (.A(_00284_),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold603 (.A(\am_sdr0.cic3.integ_sample[0] ),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold604 (.A(\am_sdr0.cic1.comb1[3] ),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold605 (.A(\am_sdr0.cic3.comb2[7] ),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold606 (.A(\am_sdr0.cic0.comb2[14] ),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold607 (.A(_00999_),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold608 (.A(\am_sdr0.cic0.integ3[12] ),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold609 (.A(_00657_),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold610 (.A(\am_sdr0.cic1.comb3_in_del[16] ),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold611 (.A(\am_sdr0.cic3.comb2[12] ),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold612 (.A(_00324_),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold613 (.A(\am_sdr0.cic0.comb1[16] ),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold614 (.A(_00973_),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold615 (.A(\am_sdr0.cic2.integ3[11] ),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold616 (.A(\am_sdr0.cic0.comb3_in_del[5] ),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold617 (.A(_00990_),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold618 (.A(\am_sdr0.am0.sum[2] ),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold619 (.A(_00110_),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold620 (.A(\am_sdr0.cic3.integ3[14] ),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold621 (.A(_01077_),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold622 (.A(\am_sdr0.cic2.comb1[9] ),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold623 (.A(_00508_),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold624 (.A(\am_sdr0.cic0.comb2_in_del[11] ),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold625 (.A(_00968_),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold626 (.A(\am_sdr0.cic3.comb3_in_del[15] ),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold627 (.A(_00327_),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold628 (.A(\am_sdr0.cic0.integ_sample[19] ),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold629 (.A(_00936_),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold630 (.A(\am_sdr0.cic0.comb3_in_del[12] ),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold631 (.A(\am_sdr0.cic0.integ3[1] ),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold632 (.A(_00646_),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold633 (.A(\am_sdr0.cic0.integ_sample[11] ),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold634 (.A(_00928_),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold635 (.A(\am_sdr0.cic3.comb3_in_del[10] ),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold636 (.A(_00322_),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold637 (.A(\am_sdr0.cic2.integ_sample[16] ),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold638 (.A(_00212_),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold639 (.A(\am_sdr0.cic1.integ_sample[11] ),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold640 (.A(_00704_),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold641 (.A(\am_sdr0.cic3.comb2[14] ),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold642 (.A(\am_sdr0.am0.q[0] ),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold643 (.A(\am_sdr0.cic3.integ_sample[11] ),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold644 (.A(_01074_),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold645 (.A(\am_sdr0.cic2.comb1_in_del[14] ),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold646 (.A(\am_sdr0.cic2.integ3[19] ),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold647 (.A(\am_sdr0.cic3.comb1_in_del[11] ),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold648 (.A(\am_sdr0.cic1.comb2[1] ),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold649 (.A(_00762_),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold650 (.A(\am_sdr0.cic1.comb2_in_del[19] ),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold651 (.A(_04248_),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold652 (.A(_00732_),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold653 (.A(\am_sdr0.cic2.comb1[1] ),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold654 (.A(_00500_),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold655 (.A(\am_sdr0.cic2.comb2[14] ),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold656 (.A(\am_sdr0.cic2.comb1[19] ),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold657 (.A(_00518_),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold658 (.A(\am_sdr0.am0.right[1] ),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold659 (.A(_02112_),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold660 (.A(\am_sdr0.cic0.comb2[8] ),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold661 (.A(_00993_),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold662 (.A(\am_sdr0.cic3.comb1[14] ),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold663 (.A(_00298_),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold664 (.A(\am_sdr0.cic1.comb3_in_del[14] ),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold665 (.A(_04305_),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold666 (.A(\am_sdr0.cic2.comb2[8] ),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold667 (.A(_00535_),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold668 (.A(\am_sdr0.cic1.comb1[13] ),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold669 (.A(_00746_),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold670 (.A(\am_sdr0.cic1.comb1[10] ),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold671 (.A(_00743_),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold672 (.A(\am_sdr0.cic0.comb1[6] ),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold673 (.A(_00963_),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold674 (.A(\am_sdr0.cic2.comb2[10] ),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold675 (.A(_00537_),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold676 (.A(\am_sdr0.cic1.comb2[13] ),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold677 (.A(_04299_),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold678 (.A(_04302_),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold679 (.A(\am_sdr0.cic2.integ3[8] ),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold680 (.A(\am_sdr0.cic2.comb2[18] ),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold681 (.A(_03362_),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold682 (.A(_03364_),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold683 (.A(\am_sdr0.cic2.integ_sample[18] ),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold684 (.A(_00214_),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold685 (.A(\am_sdr0.cic2.comb2[16] ),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold686 (.A(_03346_),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold687 (.A(_03352_),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold688 (.A(\am_sdr0.cic3.comb1[1] ),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold689 (.A(_00285_),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold690 (.A(\am_sdr0.cic3.integ_sample[1] ),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold691 (.A(_01064_),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold692 (.A(\am_sdr0.cic1.integ_sample[17] ),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold693 (.A(_00428_),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold694 (.A(\am_sdr0.cic3.comb2[17] ),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold695 (.A(\am_sdr0.cic1.integ3[14] ),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold696 (.A(_00425_),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold697 (.A(\am_sdr0.cic2.integ_sample[12] ),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold698 (.A(_00208_),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold699 (.A(\am_sdr0.cic3.comb2_in_del[0] ),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold700 (.A(\am_sdr0.cic1.integ_sample[1] ),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold701 (.A(_00694_),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold702 (.A(\am_sdr0.cic2.integ_sample[9] ),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold703 (.A(_00468_),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold704 (.A(\am_sdr0.cic3.comb1[18] ),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold705 (.A(_00302_),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold706 (.A(\am_sdr0.cic3.comb1[16] ),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold707 (.A(_00300_),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold708 (.A(\am_sdr0.cic1.comb3_in_del[12] ),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold709 (.A(\am_sdr0.cic2.comb3_in_del[12] ),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold710 (.A(\am_sdr0.cic2.comb2_in_del[8] ),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold711 (.A(\am_sdr0.cic1.comb2[4] ),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold712 (.A(_00765_),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold713 (.A(\am_sdr0.cic3.comb1_in_del[1] ),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold714 (.A(_00245_),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold715 (.A(\am_sdr0.cic2.integ_sample[6] ),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold716 (.A(_00465_),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold717 (.A(\am_sdr0.cic1.comb2[15] ),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold718 (.A(\am_sdr0.cic0.comb2_in_del[0] ),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold719 (.A(_00957_),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold720 (.A(\am_sdr0.cic3.comb1[10] ),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold721 (.A(_00294_),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold722 (.A(\am_sdr0.cic2.comb2[5] ),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold723 (.A(_00532_),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold724 (.A(\am_sdr0.cic2.comb1[0] ),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold725 (.A(_03147_),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold726 (.A(_00479_),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold727 (.A(\am_sdr0.cic2.comb1[5] ),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold728 (.A(_00504_),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold729 (.A(\am_sdr0.cic1.comb1[0] ),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold730 (.A(_00733_),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold731 (.A(\am_sdr0.cic0.comb2[14] ),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold732 (.A(\am_sdr0.cic2.comb3_in_del[19] ),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold733 (.A(\am_sdr0.cic1.comb2[6] ),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold734 (.A(_00767_),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold735 (.A(\am_sdr0.cic2.comb1[6] ),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold736 (.A(_00505_),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold737 (.A(\am_sdr0.cic2.integ_sample[7] ),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold738 (.A(_00466_),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold739 (.A(\am_sdr0.cic1.comb1[14] ),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold740 (.A(\am_sdr0.cic0.comb2[4] ),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold741 (.A(_00941_),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold742 (.A(\am_sdr0.cic0.comb1[10] ),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold743 (.A(_00967_),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold744 (.A(\am_sdr0.cic1.comb2[8] ),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold745 (.A(_00769_),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold746 (.A(\am_sdr0.cic3.integ3[9] ),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold747 (.A(_01072_),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold748 (.A(\am_sdr0.cic1.integ3[0] ),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold749 (.A(_00411_),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold750 (.A(_00039_),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold751 (.A(_00003_),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold752 (.A(\am_sdr0.cic1.comb1_in_del[15] ),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold753 (.A(_00708_),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold754 (.A(\am_sdr0.cic3.comb1_in_del[0] ),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold755 (.A(\am_sdr0.cic1.comb3_in_del[15] ),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold756 (.A(\am_sdr0.spi0.shift_reg[26] ),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold757 (.A(\am_sdr0.cic2.comb2_in_del[0] ),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold758 (.A(\am_sdr0.cic0.comb3_in_del[6] ),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold759 (.A(_00991_),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold760 (.A(\am_sdr0.cic0.comb3_in_del[18] ),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold761 (.A(\am_sdr0.cic2.comb1[2] ),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold762 (.A(_00501_),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold763 (.A(\am_sdr0.cic2.integ_sample[0] ),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold764 (.A(\am_sdr0.cic3.comb2[18] ),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold765 (.A(_02493_),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold766 (.A(\am_sdr0.cic3.integ_sample[10] ),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold767 (.A(_01073_),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold768 (.A(\am_sdr0.cic1.comb3_in_del[11] ),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold769 (.A(_00772_),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold770 (.A(\am_sdr0.cic0.comb3_in_del[11] ),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold771 (.A(_00996_),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold772 (.A(\am_sdr0.cic0.comb1[5] ),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold773 (.A(_00962_),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold774 (.A(\am_sdr0.count[0] ),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold775 (.A(_00157_),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold776 (.A(\am_sdr0.cic3.comb2_in_del[19] ),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold777 (.A(_00303_),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold778 (.A(\am_sdr0.cic2.comb3_in_del[14] ),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold779 (.A(\am_sdr0.cic3.comb3_in_del[14] ),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold780 (.A(\am_sdr0.nco0.phase_inc[12] ),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold781 (.A(\am_sdr0.cic0.comb1[8] ),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold782 (.A(_05004_),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold783 (.A(\am_sdr0.cic1.comb1[7] ),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold784 (.A(_00740_),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold785 (.A(\am_sdr0.cic0.comb2[6] ),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold786 (.A(\am_sdr0.cic3.integ_sample[3] ),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold787 (.A(_01066_),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold788 (.A(\am_sdr0.cic2.integ_sample[4] ),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold789 (.A(_00200_),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold790 (.A(\am_sdr0.cic3.comb1[5] ),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold791 (.A(_02311_),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold792 (.A(\am_sdr0.am0.multA[15] ),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold793 (.A(_01735_),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold794 (.A(\am_sdr0.cic2.integ_sample[1] ),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold795 (.A(_00460_),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold796 (.A(\am_sdr0.am0.count[0] ),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold797 (.A(_00172_),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold798 (.A(\am_sdr0.cic0.comb3_in_del[4] ),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold799 (.A(\am_sdr0.cic1.comb2_in_del[0] ),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold800 (.A(\am_sdr0.cic0.integ1[0] ),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold801 (.A(_05206_),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold802 (.A(_01014_),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold803 (.A(\am_sdr0.cic0.comb1_in_del[14] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold804 (.A(_00931_),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold805 (.A(\am_sdr0.cic0.integ_sample[3] ),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold806 (.A(_00920_),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold807 (.A(\am_sdr0.cic2.comb1_in_del[12] ),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold808 (.A(\am_sdr0.cic3.integ3[3] ),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold809 (.A(\am_sdr0.cic1.comb1[1] ),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold810 (.A(_00734_),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold811 (.A(\am_sdr0.am0.sum[11] ),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold812 (.A(_00119_),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold813 (.A(\am_sdr0.cic0.comb1[14] ),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold814 (.A(_00971_),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold815 (.A(\am_sdr0.cic3.comb3_in_del[19] ),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold816 (.A(_02497_),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold817 (.A(\am_sdr0.cic3.integ_sample[18] ),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold818 (.A(_00262_),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold819 (.A(\am_sdr0.cic3.integ3[6] ),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold820 (.A(\am_sdr0.cic2.comb1[8] ),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold821 (.A(_00046_),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold822 (.A(_05720_),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold823 (.A(_01168_),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold824 (.A(\am_sdr0.cic3.integ_sample[2] ),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold825 (.A(_01065_),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold826 (.A(\am_sdr0.cic1.comb1[8] ),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold827 (.A(_00741_),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold828 (.A(\am_sdr0.cic0.comb2_in_del[19] ),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold829 (.A(_05077_),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold830 (.A(_00956_),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold831 (.A(\am_sdr0.cic3.comb2[16] ),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold832 (.A(_00328_),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold833 (.A(\am_sdr0.cic1.comb1[2] ),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold834 (.A(_00735_),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold835 (.A(\am_sdr0.cic1.comb2[7] ),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold836 (.A(_00768_),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold837 (.A(\am_sdr0.cic2.comb1[10] ),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold838 (.A(_00509_),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold839 (.A(\am_sdr0.nco0.phase_inc[16] ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold840 (.A(\am_sdr0.cic2.comb1_in_del[18] ),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold841 (.A(\am_sdr0.cic1.comb2[14] ),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold842 (.A(\am_sdr0.cic0.comb3_in_del[7] ),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold843 (.A(_00992_),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold844 (.A(\am_sdr0.am0.sum[1] ),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold845 (.A(\am_sdr0.cic3.integ_sample[8] ),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold846 (.A(_01071_),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold847 (.A(\am_sdr0.cic3.comb1_in_del[3] ),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold848 (.A(\am_sdr0.cic3.integ_sample[7] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold849 (.A(_01070_),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold850 (.A(\am_sdr0.cic2.comb2[13] ),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold851 (.A(_03324_),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold852 (.A(\am_sdr0.cic2.comb3_in_del[11] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold853 (.A(_00538_),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold854 (.A(\am_sdr0.cic3.integ_sample[4] ),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold855 (.A(_01067_),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold856 (.A(\am_sdr0.cic2.comb2_in_del[3] ),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold857 (.A(_00502_),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold858 (.A(\am_sdr0.cic3.integ3[16] ),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold859 (.A(_01079_),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold860 (.A(\am_sdr0.cic2.integ3[10] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold861 (.A(\am_sdr0.cic2.comb1[7] ),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold862 (.A(_00506_),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold863 (.A(\am_sdr0.cic3.comb1[12] ),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold864 (.A(\am_sdr0.cic0.integ3[0] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold865 (.A(_00645_),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold866 (.A(\am_sdr0.cic2.comb1_in_del[16] ),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold867 (.A(\am_sdr0.count[2] ),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold868 (.A(_02076_),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold869 (.A(_00158_),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold870 (.A(\am_sdr0.cic2.comb2[4] ),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold871 (.A(_00531_),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold872 (.A(\am_sdr0.cic2.comb3_in_del[16] ),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold873 (.A(\am_sdr0.cic2.comb3_in_del[18] ),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold874 (.A(\am_sdr0.cic3.comb2_in_del[3] ),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold875 (.A(_00287_),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold876 (.A(\am_sdr0.cic2.comb1_in_del[3] ),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold877 (.A(\am_sdr0.cic3.comb2[16] ),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold878 (.A(\am_sdr0.nco0.phase_inc[25] ),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold879 (.A(\am_sdr0.cic2.comb1[13] ),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold880 (.A(_03227_),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold881 (.A(\am_sdr0.cic3.comb2_in_del[13] ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold882 (.A(_00297_),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold883 (.A(\am_sdr0.cic3.comb2[13] ),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold884 (.A(_02460_),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold885 (.A(\am_sdr0.cic0.comb3_in_del[10] ),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold886 (.A(\am_sdr0.cic0.comb1[2] ),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold887 (.A(_00959_),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold888 (.A(\am_sdr0.cic0.comb1[0] ),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold889 (.A(\am_sdr0.cic2.count[3] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold890 (.A(_03394_),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold891 (.A(\am_sdr0.cic0.comb2[17] ),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold892 (.A(_01002_),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold893 (.A(\am_sdr0.cic3.comb1_in_del[7] ),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold894 (.A(\am_sdr0.cic3.comb1[3] ),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold895 (.A(\am_sdr0.nco0.phase_inc[1] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold896 (.A(\am_sdr0.cic0.comb1_in_del[16] ),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold897 (.A(_00933_),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold898 (.A(\am_sdr0.nco0.phase_inc[20] ),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold899 (.A(\am_sdr0.cic3.comb1[10] ),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold900 (.A(_02338_),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold901 (.A(\am_sdr0.cic0.comb2[16] ),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold902 (.A(\am_sdr0.cic1.integ_sample[2] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold903 (.A(_00695_),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold904 (.A(\am_sdr0.cic1.comb2_in_del[14] ),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold905 (.A(\am_sdr0.cic2.comb1_in_del[4] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold906 (.A(_00463_),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold907 (.A(\am_sdr0.cic1.comb2_in_del[3] ),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold908 (.A(\am_sdr0.cic2.comb1[14] ),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold909 (.A(_00513_),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold910 (.A(\am_sdr0.cic1.integ_sample[7] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold911 (.A(_00700_),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold912 (.A(\am_sdr0.cic1.comb2[11] ),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold913 (.A(\am_sdr0.cic0.comb2_in_del[3] ),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold914 (.A(\am_sdr0.cic0.comb1_in_del[12] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold915 (.A(_00929_),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold916 (.A(\am_sdr0.cic3.comb1[7] ),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold917 (.A(_00291_),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold918 (.A(\am_sdr0.cic0.comb2_in_del[12] ),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold919 (.A(_00969_),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold920 (.A(\am_sdr0.cic1.integ_sample[14] ),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold921 (.A(_00707_),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold922 (.A(\am_sdr0.cic2.comb1[3] ),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold923 (.A(\am_sdr0.am0.demod_out[8] ),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold924 (.A(\am_sdr0.cic1.comb2_in_del[5] ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold925 (.A(_00738_),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold926 (.A(\am_sdr0.cic2.comb3_in_del[7] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold927 (.A(_00534_),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold928 (.A(\am_sdr0.cic3.integ_sample[6] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold929 (.A(\am_sdr0.cic1.integ2[3] ),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold930 (.A(\am_sdr0.cic0.comb1[18] ),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold931 (.A(_00975_),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold932 (.A(\am_sdr0.cic3.count[3] ),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold933 (.A(_02523_),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold934 (.A(\am_sdr0.cic1.integ_sample[3] ),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold935 (.A(_00696_),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold936 (.A(\am_sdr0.cic3.comb1[4] ),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold937 (.A(_02306_),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold938 (.A(\am_sdr0.cic0.integ_sample[17] ),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold939 (.A(_00662_),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold940 (.A(\am_sdr0.cic2.integ_sample[2] ),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold941 (.A(_00461_),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold942 (.A(\am_sdr0.cic3.count[4] ),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold943 (.A(\am_sdr0.cic3.comb1_in_del[2] ),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold944 (.A(_00038_),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold945 (.A(\am_sdr0.cic2.integ3[2] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold946 (.A(\am_sdr0.cic1.comb2_in_del[3] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold947 (.A(\am_sdr0.cic1.comb2_in_del[15] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold948 (.A(_00748_),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold949 (.A(\am_sdr0.cic1.comb2_in_del[6] ),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold950 (.A(\am_sdr0.cic1.comb2_in_del[18] ),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold951 (.A(_04239_),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold952 (.A(\am_sdr0.cic0.integ2[0] ),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold953 (.A(_05346_),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold954 (.A(_01040_),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold955 (.A(\am_sdr0.cic0.integ_sample[0] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold956 (.A(\am_sdr0.cic2.comb2_in_del[19] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold957 (.A(\am_sdr0.cic2.comb1_in_del[13] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold958 (.A(_00472_),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold959 (.A(\am_sdr0.am0.sum[13] ),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold960 (.A(\am_sdr0.cic2.count[4] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold961 (.A(\am_sdr0.cic2.integ3[7] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold962 (.A(\am_sdr0.cic3.integ_sample[16] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold963 (.A(_00260_),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold964 (.A(\am_sdr0.cic3.comb3_in_del[18] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold965 (.A(\am_sdr0.cic0.comb1_in_del[7] ),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold966 (.A(_00924_),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold967 (.A(\am_sdr0.cic0.integ_sample[5] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold968 (.A(_04842_),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold969 (.A(_04844_),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold970 (.A(\am_sdr0.cic2.integ3[1] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold971 (.A(\am_sdr0.cic1.integ_sample[0] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold972 (.A(\am_sdr0.cic2.comb1[16] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold973 (.A(_00515_),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold974 (.A(\am_sdr0.cic0.comb2[15] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold975 (.A(\am_sdr0.cic2.integ3[3] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold976 (.A(\am_sdr0.cic3.comb1_in_del[6] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold977 (.A(\am_sdr0.cic0.integ_sample[10] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold978 (.A(_00927_),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold979 (.A(\am_sdr0.cic0.comb1_in_del[17] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold980 (.A(\am_sdr0.cic2.comb2_in_del[1] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold981 (.A(\am_sdr0.gain_spi[1] ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold982 (.A(\am_sdr0.cic0.comb2[7] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold983 (.A(\am_sdr0.cic0.comb1[16] ),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold984 (.A(_05053_),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold985 (.A(\am_sdr0.gain_spi[2] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold986 (.A(\am_sdr0.cic1.integ3[12] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold987 (.A(_00423_),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold988 (.A(\am_sdr0.cic2.comb3_in_del[17] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold989 (.A(\am_sdr0.cic1.comb2_in_del[12] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold990 (.A(_00745_),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold991 (.A(\am_sdr0.cic3.comb2[9] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold992 (.A(_00273_),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold993 (.A(\am_sdr0.cic3.integ2[2] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold994 (.A(_00368_),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold995 (.A(\am_sdr0.cic2.comb1_in_del[5] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold996 (.A(_00464_),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold997 (.A(\am_sdr0.cic1.comb1_in_del[10] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold998 (.A(_00703_),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold999 (.A(\am_sdr0.cic2.integ3[9] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\am_sdr0.cic2.comb1[17] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold1001 (.A(_00456_),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\am_sdr0.cic0.integ_sample[18] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold1003 (.A(_04928_),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\am_sdr0.cic1.comb1_in_del[18] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold1005 (.A(_00711_),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\am_sdr0.cic3.comb2_in_del[8] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold1007 (.A(_00292_),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\am_sdr0.cic0.comb1_in_del[1] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold1009 (.A(_00918_),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\am_sdr0.cic2.comb1_in_del[19] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\am_sdr0.cic1.comb1[4] ),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold1012 (.A(_00737_),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\am_sdr0.cic0.comb2_in_del[1] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold1014 (.A(_00958_),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\am_sdr0.cic2.comb2[12] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\am_sdr0.cic2.comb2_in_del[12] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold1017 (.A(_03229_),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold1018 (.A(_03231_),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\am_sdr0.am0.multA[7] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold1020 (.A(_00098_),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\am_sdr0.cic3.integ_sample[14] ),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold1022 (.A(_00258_),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\am_sdr0.cic0.comb1_in_del[19] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold1024 (.A(_04937_),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\am_sdr0.cic0.comb2[12] ),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\am_sdr0.cic0.comb1_in_del[6] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold1027 (.A(_00923_),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\am_sdr0.am0.sum[3] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\am_sdr0.cic0.comb1_in_del[18] ),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\am_sdr0.cic1.comb2_in_del[16] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\am_sdr0.cic1.comb1_in_del[19] ),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold1032 (.A(_04103_),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\am_sdr0.cic1.comb1_in_del[4] ),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold1034 (.A(_00697_),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\am_sdr0.cic0.comb1[13] ),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold1036 (.A(_00910_),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\am_sdr0.cic3.comb1_in_del[10] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\am_sdr0.am0.multA[13] ),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold1039 (.A(_00105_),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\am_sdr0.cic3.integ1[2] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\am_sdr0.cic1.comb1_in_del[8] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold1042 (.A(_00701_),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\am_sdr0.am0.sum[12] ),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\am_sdr0.cic0.integ_sample[8] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\am_sdr0.cic2.integ3[6] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\am_sdr0.cic0.integ_sample[2] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold1047 (.A(_00919_),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\am_sdr0.cic2.comb3_in_del[15] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\am_sdr0.cic3.comb2_in_del[4] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\am_sdr0.cic0.comb1_in_del[15] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold1051 (.A(_00932_),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\am_sdr0.cic0.comb2[5] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold1053 (.A(_00942_),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\am_sdr0.cic1.comb1_in_del[12] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold1055 (.A(_00705_),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\am_sdr0.cic2.integ2[2] ),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold1057 (.A(_00583_),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\am_sdr0.cic0.comb2_in_del[8] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\am_sdr0.cic1.comb2[12] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\am_sdr0.cic3.comb2_in_del[6] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold1061 (.A(_00290_),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\am_sdr0.cic0.comb2_in_del[18] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\am_sdr0.cic0.comb1[1] ),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold1064 (.A(_04962_),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\am_sdr0.cic3.comb1[6] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\am_sdr0.cic3.integ_sample[12] ),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold1067 (.A(_01075_),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\am_sdr0.cic3.comb1[8] ),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\am_sdr0.cic3.comb1_in_del[8] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\am_sdr0.am0.sum[5] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\am_sdr0.am0.multA[8] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\am_sdr0.cic0.comb1[14] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\am_sdr0.cic1.comb1[6] ),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\am_sdr0.cic3.integ3[15] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold1075 (.A(_01078_),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\am_sdr0.cic3.comb1_in_del[4] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\am_sdr0.cic3.comb1[17] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold1078 (.A(_00241_),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\am_sdr0.cic0.integ_sample[4] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold1080 (.A(_00921_),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\am_sdr0.am0.sum[6] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\am_sdr0.cic3.integ2[1] ),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\am_sdr0.cic3.comb2_in_del[12] ),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\am_sdr0.cic0.comb1[15] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold1085 (.A(_00972_),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\am_sdr0.nco0.phase_inc[3] ),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\am_sdr0.cic0.comb1[13] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold1088 (.A(_05039_),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\am_sdr0.cic0.comb1[17] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold1090 (.A(_00974_),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\am_sdr0.cic2.comb2_in_del[5] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\am_sdr0.cic1.integ_sample[6] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold1093 (.A(_00699_),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\am_sdr0.cic1.comb1_in_del[16] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold1095 (.A(_00709_),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\am_sdr0.cic3.integ3[9] ),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\am_sdr0.cic0.integ2[3] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\am_sdr0.cic3.comb2[10] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\am_sdr0.cic3.comb1[15] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold1100 (.A(_00299_),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\am_sdr0.cic1.comb1[18] ),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\am_sdr0.cic2.comb1_in_del[15] ),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\am_sdr0.cic3.integ_sample[14] ),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\am_sdr0.cic1.comb2_in_del[1] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\am_sdr0.cic3.comb1[16] ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\am_sdr0.cic3.integ3[5] ),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold1107 (.A(_01068_),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\am_sdr0.am0.sum[14] ),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\am_sdr0.cic2.integ_sample[10] ),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\am_sdr0.cic3.comb1_in_del[12] ),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\am_sdr0.cic3.comb2[6] ),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold1112 (.A(_00270_),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\am_sdr0.cic3.comb2_in_del[1] ),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\am_sdr0.cic1.comb1[16] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\am_sdr0.cic1.comb1_in_del[4] ),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold1116 (.A(_03999_),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\am_sdr0.cic3.comb1[9] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold1118 (.A(_00293_),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\am_sdr0.am0.m_count[2] ),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold1120 (.A(_01679_),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\am_sdr0.cic1.comb2[10] ),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\am_sdr0.am0.multA[14] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\am_sdr0.cic0.comb1_in_del[8] ),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\am_sdr0.cic2.comb2_in_del[13] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\am_sdr0.cic3.comb2[8] ),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\am_sdr0.cic2.comb2[7] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold1127 (.A(_00486_),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\am_sdr0.cic3.integ3[13] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold1129 (.A(_01076_),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\am_sdr0.cic2.comb1[18] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold1131 (.A(_03263_),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\am_sdr0.cic3.integ3[17] ),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold1133 (.A(_01080_),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\am_sdr0.cic0.comb2[3] ),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\am_sdr0.cic2.comb1[12] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\am_sdr0.cic2.comb1_in_del[17] ),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\am_sdr0.cic3.integ_sample[16] ),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\am_sdr0.cic2.comb3_in_del[13] ),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\am_sdr0.cic3.comb1[19] ),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\am_sdr0.cic2.comb2[11] ),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\am_sdr0.mix0.RF_in_qq ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\am_sdr0.am0.state[2] ),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\am_sdr0.cic2.integ1[2] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold1144 (.A(_00557_),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\am_sdr0.cic1.integ_sample[13] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\am_sdr0.cic3.integ1[1] ),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold1147 (.A(_00341_),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\am_sdr0.cic1.integ_sample[8] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold1149 (.A(_04027_),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\am_sdr0.cic2.integ2[22] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\am_sdr0.cic0.count[5] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\am_sdr0.cic2.integ3[5] ),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold1153 (.A(_00201_),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\am_sdr0.cic3.comb1_in_del[15] ),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold1155 (.A(_00259_),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\am_sdr0.cic2.integ2[1] ),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\am_sdr0.cic1.comb1[17] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold1158 (.A(_00690_),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\am_sdr0.cic2.integ3[4] ),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\am_sdr0.am0.multA[9] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold1161 (.A(_01727_),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\am_sdr0.am0.multB[1] ),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold1163 (.A(_01683_),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\am_sdr0.cic0.comb1[4] ),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold1165 (.A(_00901_),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\am_sdr0.cic1.comb3_in_del[13] ),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\am_sdr0.cic3.comb1[18] ),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\am_sdr0.am0.state[1] ),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\am_sdr0.cic0.comb2_in_del[4] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\am_sdr0.am0.multA[2] ),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold1171 (.A(_00094_),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\am_sdr0.am0.multA[5] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold1173 (.A(_00097_),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\am_sdr0.cic3.comb1_in_del[3] ),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\am_sdr0.cic2.integ2[6] ),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\am_sdr0.am0.sum[7] ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\am_sdr0.cic1.comb2[9] ),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\am_sdr0.cic3.comb3_in_del[13] ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\am_sdr0.cic0.comb2[11] ),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\am_sdr0.cic2.comb2[3] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\am_sdr0.cic2.integ1[1] ),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold1182 (.A(_00556_),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\am_sdr0.cic1.comb2[3] ),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\am_sdr0.cic0.comb1_in_del[9] ),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold1185 (.A(_00926_),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\am_sdr0.cic0.integ1[3] ),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold1187 (.A(_01041_),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\am_sdr0.cic1.comb2_in_del[9] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold1189 (.A(_00742_),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\am_sdr0.cic2.integ_sample[13] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold1191 (.A(_00209_),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\am_sdr0.cic2.count[5] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\am_sdr0.cic0.integ_sample[16] ),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\am_sdr0.cic3.comb1_in_del[18] ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold1195 (.A(_02262_),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\am_sdr0.cic2.comb1[15] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold1197 (.A(_00514_),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\am_sdr0.cic1.count[5] ),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\am_sdr0.cic0.integ_sample[6] ),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\am_sdr0.cic3.comb2[2] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold1201 (.A(_00266_),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\am_sdr0.cic3.count[5] ),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\am_sdr0.cic3.comb1[17] ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\am_sdr0.cic1.comb1[11] ),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\am_sdr0.cic1.comb2[5] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold1206 (.A(_00718_),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\am_sdr0.cic2.comb1[16] ),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\am_sdr0.cic0.integ_sample[15] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold1209 (.A(_00660_),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\am_sdr0.cic2.integ_sample[6] ),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\am_sdr0.cic2.comb1_in_del[1] ),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\am_sdr0.cic2.comb2[2] ),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold1213 (.A(_00481_),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\am_sdr0.cic0.comb2_in_del[13] ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\am_sdr0.cic3.integ3[19] ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold1216 (.A(_00408_),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\am_sdr0.cic2.comb2[6] ),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\am_sdr0.cic1.integ_sample[5] ),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold1219 (.A(_00698_),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\am_sdr0.cic3.integ2[3] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\am_sdr0.cic0.comb2[9] ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold1222 (.A(_00946_),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\am_sdr0.cic1.comb2_in_del[6] ),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold1224 (.A(_04153_),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\am_sdr0.cic2.comb1_in_del[14] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\am_sdr0.cic3.comb2[15] ),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold1227 (.A(_00279_),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\am_sdr0.cic3.comb1_in_del[17] ),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold1229 (.A(_00261_),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\am_sdr0.cic3.comb1_in_del[9] ),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold1231 (.A(_02191_),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\am_sdr0.cic3.integ_sample[5] ),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold1233 (.A(_02170_),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold1234 (.A(_00229_),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\am_sdr0.cic0.comb1[9] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold1236 (.A(_00966_),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\am_sdr0.cic3.integ2[22] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\am_sdr0.am0.state[5] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\am_sdr0.cic2.integ1[20] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\am_sdr0.cic3.integ3[14] ),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold1241 (.A(_02932_),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\am_sdr0.cic1.comb2[2] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold1243 (.A(_00715_),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\am_sdr0.cic1.integ_sample[9] ),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold1245 (.A(_00702_),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\am_sdr0.am0.multA[4] ),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold1247 (.A(_00096_),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\am_sdr0.cic2.comb2_in_del[17] ),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\am_sdr0.cic2.integ3[16] ),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\am_sdr0.am0.multA[3] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold1251 (.A(_00095_),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\am_sdr0.cic0.comb1[11] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\am_sdr0.cic2.integ3[14] ),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\am_sdr0.cic0.comb2[2] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold1255 (.A(_00939_),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\am_sdr0.cic2.integ2[3] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\am_sdr0.cic0.comb1_in_del[14] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold1258 (.A(_04910_),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\am_sdr0.cic2.count[2] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\am_sdr0.cic2.integ1[21] ),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\am_sdr0.cic1.comb1_in_del[10] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\am_sdr0.cic3.integ_sample[9] ),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\am_sdr0.cic0.integ_sample[1] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\am_sdr0.cic2.integ2[21] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\am_sdr0.cic0.comb3_in_del[13] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\am_sdr0.am0.multA[1] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold1267 (.A(_00093_),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\am_sdr0.cic1.comb1_in_del[17] ),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\am_sdr0.cic0.integ_sample[2] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\am_sdr0.cic1.comb2_in_del[17] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\am_sdr0.cic1.comb1_in_del[13] ),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\am_sdr0.cic1.comb1_in_del[1] ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold1273 (.A(_03990_),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\am_sdr0.cic3.comb2_in_del[17] ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\am_sdr0.cic2.integ_sample[8] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\am_sdr0.cic3.integ1[6] ),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\am_sdr0.cic0.integ_sample[17] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold1278 (.A(_04925_),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\am_sdr0.am0.sum[10] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\am_sdr0.cic3.comb1_in_del[13] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold1281 (.A(_00257_),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\am_sdr0.cic1.integ2[1] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold1283 (.A(_04513_),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold1284 (.A(_00817_),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\am_sdr0.cic0.comb1[17] ),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\am_sdr0.cic3.comb2_in_del[5] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\am_sdr0.cic3.integ1[20] ),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\am_sdr0.nco0.phase[23] ),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\am_sdr0.am0.multA[12] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\am_sdr0.cic2.integ3[8] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\am_sdr0.cic1.comb1[9] ),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold1292 (.A(_00682_),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\am_sdr0.cic2.comb2_in_del[14] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold1294 (.A(_03243_),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\am_sdr0.cic3.integ3[16] ),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\am_sdr0.am0.sum[9] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\am_sdr0.nco0.phase[25] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\am_sdr0.cic3.comb1_in_del[5] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\am_sdr0.cic2.integ3[18] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\am_sdr0.cic3.integ3[11] ),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold1301 (.A(_00400_),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\am_sdr0.cic2.integ1[3] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold1303 (.A(_00558_),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\am_sdr0.cic3.count[2] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\am_sdr0.cic1.comb1[12] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold1306 (.A(\am_sdr0.cic1.integ_sample[6] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\am_sdr0.cic3.integ1[5] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\am_sdr0.cic3.integ3[8] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\am_sdr0.cic2.integ2[9] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\am_sdr0.cic2.integ3[17] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold1311 (.A(_00621_),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\am_sdr0.cic0.integ_sample[9] ),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold1313 (.A(_04865_),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\am_sdr0.cic1.comb1[15] ),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\am_sdr0.cic3.integ3[2] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold1316 (.A(_00391_),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\am_sdr0.cic1.integ2[4] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\am_sdr0.cic3.integ3[7] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\am_sdr0.cic2.integ1[5] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold1320 (.A(_00560_),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\am_sdr0.cic3.integ3[5] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold1322 (.A(_02873_),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\am_sdr0.cic1.integ2[22] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold1324 (.A(_00644_),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\am_sdr0.cic3.integ3[12] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\am_sdr0.am0.multA[10] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold1327 (.A(_00102_),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\am_sdr0.cic2.integ3[13] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold1329 (.A(_00617_),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\am_sdr0.cic3.integ2[17] ),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\am_sdr0.cic0.integ2[4] ),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\am_sdr0.cic2.integ3[6] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\am_sdr0.cic2.comb1_in_del[2] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\am_sdr0.cic2.integ1[6] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\am_sdr0.cic0.comb1_in_del[5] ),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\am_sdr0.cic3.integ3[10] ),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\am_sdr0.cic2.integ3[12] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\am_sdr0.cic1.integ3[17] ),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold1339 (.A(_03943_),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold1340 (.A(_00643_),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\am_sdr0.cic3.integ1[23] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\am_sdr0.cic2.integ1[13] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\am_sdr0.cic2.integ1[7] ),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold1344 (.A(_00562_),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\am_sdr0.am0.count2[1] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold1346 (.A(_01928_),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold1347 (.A(_00126_),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\am_sdr0.cic3.integ3[4] ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\am_sdr0.cic2.integ3[10] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\am_sdr0.cic2.sample ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\am_sdr0.cic2.integ1[9] ),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\am_sdr0.am0.multA[11] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold1353 (.A(\am_sdr0.cic1.comb1[5] ),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold1354 (.A(_00678_),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\am_sdr0.cic2.integ1[12] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\am_sdr0.cic3.integ3[1] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\am_sdr0.cic3.integ2[9] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\am_sdr0.cic3.integ_sample[15] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\am_sdr0.nco0.phase[22] ),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\am_sdr0.cic0.integ2[22] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold1361 (.A(_00859_),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\am_sdr0.cic2.integ3[15] ),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold1363 (.A(_00619_),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\am_sdr0.cic2.integ1[11] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\am_sdr0.cic3.integ2[21] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\am_sdr0.cic0.integ3[17] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold1367 (.A(_04741_),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold1368 (.A(_00858_),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\am_sdr0.cic2.integ2[17] ),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\am_sdr0.am0.right[0] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\am_sdr0.cic3.comb1[13] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\am_sdr0.nco0.phase[18] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold1373 (.A(_05632_),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold1374 (.A(_01156_),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\am_sdr0.cic1.integ1[24] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\am_sdr0.cic3.integ1[3] ),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold1377 (.A(_00343_),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\am_sdr0.cic2.integ1[19] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\am_sdr0.cic3.integ2[11] ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\am_sdr0.cic3.integ1[19] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\am_sdr0.cic3.integ3[12] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\am_sdr0.cic3.integ2[20] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\am_sdr0.cic1.integ1[25] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold1384 (.A(_00838_),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\am_sdr0.I_out[1] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold1386 (.A(_05214_),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold1387 (.A(_01016_),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\am_sdr0.cic0.comb1[12] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold1389 (.A(_00909_),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\am_sdr0.cic3.integ2[7] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\am_sdr0.cic3.integ1[17] ),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\am_sdr0.gain_spi[0] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\am_sdr0.cic3.integ1[21] ),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\am_sdr0.cic3.integ1[12] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\am_sdr0.cic3.integ1[9] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\am_sdr0.cic3.integ1[16] ),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\am_sdr0.cic2.integ1[23] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\am_sdr0.Q_out[4] ),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold1399 (.A(_04396_),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold1400 (.A(_00795_),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\am_sdr0.cic2.integ2[10] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\am_sdr0.cic3.integ2[13] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\am_sdr0.cic3.integ1[10] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\am_sdr0.cic2.integ1[4] ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\am_sdr0.cic2.integ1[17] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\am_sdr0.cic2.integ1[8] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold1407 (.A(\am_sdr0.nco0.phase[1] ),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold1408 (.A(_01140_),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold1409 (.A(\am_sdr0.cic2.integ2[19] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\am_sdr0.cic3.integ2[14] ),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\am_sdr0.cic2.integ2[16] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\am_sdr0.cic1.comb2_in_del[12] ),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\am_sdr0.cic0.integ1[25] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\am_sdr0.nco0.phase[10] ),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold1415 (.A(\am_sdr0.count[5] ),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold1416 (.A(_02084_),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\am_sdr0.cic3.integ2[6] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\am_sdr0.cic3.integ2[12] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\am_sdr0.cic3.integ1[11] ),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\am_sdr0.cic2.integ2[18] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\am_sdr0.cic2.integ2[14] ),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\am_sdr0.cic1.integ2[15] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\am_sdr0.nco0.phase[8] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold1424 (.A(_01146_),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\am_sdr0.Q_out[2] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold1426 (.A(_04378_),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold1427 (.A(_00792_),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\am_sdr0.cic1.integ2[19] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold1429 (.A(_00641_),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\am_sdr0.cic3.integ1[8] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\am_sdr0.nco0.phase[20] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\am_sdr0.cic3.integ1[13] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\am_sdr0.count[4] ),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\am_sdr0.cic0.integ2[19] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold1435 (.A(_00856_),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\am_sdr0.nco0.phase[6] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold1437 (.A(_01144_),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\am_sdr0.cic3.integ2[10] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\am_sdr0.cic3.integ2[19] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\am_sdr0.cic0.integ2[8] ),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold1441 (.A(_00845_),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\am_sdr0.cic2.integ2[20] ),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\am_sdr0.I_out[4] ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold1444 (.A(_05230_),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold1445 (.A(_01019_),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold1446 (.A(\am_sdr0.cic1.integ2[8] ),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold1447 (.A(_00630_),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\am_sdr0.cic2.integ2[5] ),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\am_sdr0.nco0.phase[4] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold1450 (.A(_05550_),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold1451 (.A(_01143_),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\am_sdr0.cic3.integ1[7] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold1453 (.A(_00347_),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\am_sdr0.am0.multA[0] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold1455 (.A(_00092_),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\am_sdr0.nco0.phase[14] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold1457 (.A(_05604_),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold1458 (.A(_01152_),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\am_sdr0.cic1.integ1[23] ),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold1460 (.A(_04500_),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\am_sdr0.cic2.integ2[8] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\am_sdr0.cic2.integ1[14] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\am_sdr0.Q_out[0] ),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold1464 (.A(_04375_),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold1465 (.A(_00791_),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\am_sdr0.cic2.integ1[10] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\am_sdr0.cic0.integ2[13] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\am_sdr0.cic3.integ1[15] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\am_sdr0.cic3.integ2[16] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\am_sdr0.cic3.integ2[4] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\am_sdr0.cic1.integ2[6] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold1472 (.A(_00628_),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\am_sdr0.cic3.integ1[4] ),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\am_sdr0.cic1.integ2[13] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\am_sdr0.I_out[6] ),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold1476 (.A(_05233_),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold1477 (.A(_01020_),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\am_sdr0.cic3.integ2[18] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\am_sdr0.cic3.integ1[24] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\am_sdr0.cic2.integ2[12] ),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold1481 (.A(\am_sdr0.cic3.integ2[5] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\am_sdr0.cic2.integ2[13] ),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\am_sdr0.cic0.integ2[6] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold1484 (.A(_00843_),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\am_sdr0.cic0.integ2[20] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold1486 (.A(\am_sdr0.cic3.integ2[8] ),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\am_sdr0.cic2.integ1[15] ),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\am_sdr0.cic3.integ2[15] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\am_sdr0.cic0.integ1[24] ),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold1490 (.A(\am_sdr0.Q_out[6] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold1491 (.A(_04399_),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold1492 (.A(_00796_),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\am_sdr0.cic3.integ1[14] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\am_sdr0.cic1.integ2[20] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\am_sdr0.cic3.integ1[18] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\am_sdr0.cic2.integ2[7] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\am_sdr0.cic2.integ1[16] ),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\am_sdr0.count[3] ),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\am_sdr0.cic2.integ1[24] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\am_sdr0.am0.I_in[0] ),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold1501 (.A(_01681_),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\am_sdr0.cic2.integ1[22] ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\am_sdr0.I_out[0] ),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold1504 (.A(_05209_),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold1505 (.A(_01015_),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\am_sdr0.cic1.integ1[19] ),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold1507 (.A(_04604_),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold1508 (.A(_00833_),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\am_sdr0.nco0.phase_inc[1] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\am_sdr0.cic1.integ2[5] ),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold1511 (.A(_04531_),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold1512 (.A(_00821_),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\am_sdr0.cic2.integ2[4] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold1514 (.A(_00585_),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\am_sdr0.nco0.phase[21] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\am_sdr0.cic1.integ2[2] ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold1517 (.A(_04515_),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold1518 (.A(_00819_),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\am_sdr0.am0.m_count[3] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\am_sdr0.cic0.integ2[15] ),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold1521 (.A(_00853_),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\am_sdr0.cic0.integ2[5] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold1523 (.A(_05366_),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold1524 (.A(_01045_),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\am_sdr0.nco0.phase[9] ),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\am_sdr0.cic2.integ2[15] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\am_sdr0.cic2.integ2[11] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\am_sdr0.cic2.integ1[18] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\am_sdr0.nco0.phase[19] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold1530 (.A(_05641_),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold1531 (.A(_01157_),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\am_sdr0.nco0.phase[15] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold1533 (.A(_05611_),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold1534 (.A(_05613_),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold1535 (.A(_01153_),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\am_sdr0.cic3.integ1[22] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\am_sdr0.nco0.phase[11] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\am_sdr0.cic1.integ1[7] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold1539 (.A(_00798_),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\am_sdr0.cic0.integ1[19] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold1541 (.A(_05439_),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold1542 (.A(_01057_),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\am_sdr0.cic0.integ2[2] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold1544 (.A(_05350_),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold1545 (.A(_01043_),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\am_sdr0.cic0.integ2[21] ),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold1547 (.A(_01061_),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\am_sdr0.cic0.integ2[12] ),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold1549 (.A(_04681_),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold1550 (.A(_00849_),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\am_sdr0.nco0.phase[12] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold1552 (.A(_01151_),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\am_sdr0.cic1.integ2[14] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\am_sdr0.cic0.integ1[10] ),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold1555 (.A(_01024_),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\am_sdr0.cic0.integ2[14] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\am_sdr0.cic1.integ1[5] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\am_sdr0.cic0.integ1[22] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\am_sdr0.cic1.integ1[12] ),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold1560 (.A(_00803_),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\am_sdr0.cic0.integ1[12] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold1562 (.A(_01027_),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\am_sdr0.cic0.integ1[13] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold1564 (.A(_01028_),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\am_sdr0.cic0.integ1[23] ),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\am_sdr0.count[6] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\am_sdr0.count[0] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\am_sdr0.cic1.integ2[11] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold1569 (.A(_00634_),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\am_sdr0.nco0.phase[16] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\am_sdr0.Q_out[3] ),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\am_sdr0.cic0.integ2[9] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold1573 (.A(_05387_),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold1574 (.A(_01049_),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\am_sdr0.cic1.integ2[12] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold1576 (.A(_04566_),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold1577 (.A(_04581_),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\am_sdr0.cic1.integ1[11] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\am_sdr0.cic1.integ1[22] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\am_sdr0.cic0.integ1[15] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold1581 (.A(_05416_),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\am_sdr0.cic0.integ2[1] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold1583 (.A(_05353_),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\am_sdr0.cic1.integ2[9] ),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold1585 (.A(_04552_),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\am_sdr0.cic1.integ2[21] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\am_sdr0.cic0.integ1[11] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\am_sdr0.nco0.phase[3] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\am_sdr0.cic1.integ1[14] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\am_sdr0.I_out[3] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\am_sdr0.cic1.integ2[10] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\am_sdr0.cic1.integ2[11] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\am_sdr0.cic1.integ3[5] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold1594 (.A(_03864_),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold1595 (.A(_00631_),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\am_sdr0.cic0.integ2[10] ),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold1597 (.A(_04669_),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\am_sdr0.cic1.integ1[13] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold1599 (.A(_00827_),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\am_sdr0.cic0.integ1[22] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold1601 (.A(_05453_),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold1602 (.A(_01059_),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\am_sdr0.cic0.integ2[11] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold1604 (.A(_04675_),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold1605 (.A(\am_sdr0.cic1.integ1[17] ),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold1606 (.A(_00807_),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\am_sdr0.cic0.integ1[20] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold1608 (.A(_01035_),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\am_sdr0.cic0.integ3[5] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\am_sdr0.cic0.integ1[8] ),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold1611 (.A(_00056_),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold1612 (.A(_02026_),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\am_sdr0.cic0.integ1[14] ),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\am_sdr0.cic1.integ2[15] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\am_sdr0.cic0.integ2[13] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold1616 (.A(_01054_),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\am_sdr0.cic0.integ1[18] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold1618 (.A(_05304_),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\am_sdr0.cic0.integ1[17] ),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold1620 (.A(_01031_),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\am_sdr0.cic1.integ2[13] ),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\am_sdr0.nco0.phase_inc[3] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\am_sdr0.cic1.integ1[2] ),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\am_sdr0.cic1.integ1[9] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold1625 (.A(_04541_),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\am_sdr0.cic1.integ1[8] ),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\am_sdr0.I_out[2] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\am_sdr0.cic0.integ1[18] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold1629 (.A(\am_sdr0.cic0.integ1[10] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold1630 (.A(_05375_),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\am_sdr0.cic1.integ2[8] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\am_sdr0.cic0.integ1[21] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold1633 (.A(\am_sdr0.cic1.integ2[5] ),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\am_sdr0.cic0.integ1[24] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold1635 (.A(_05339_),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\am_sdr0.cic1.integ2[19] ),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\am_sdr0.cic2.comb2[12] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold1638 (.A(\am_sdr0.cic1.comb1[4] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\am_sdr0.cic0.comb2[12] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\am_sdr0.cic3.integ1[1] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\am_sdr0.cic0.comb2[15] ),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\am_sdr0.cic1.integ_sample[2] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\am_sdr0.cic2.integ3[18] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\am_sdr0.cic0.comb2[17] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\am_sdr0.cic0.integ1[11] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold1646 (.A(_05381_),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold1647 (.A(\am_sdr0.cic0.integ3[7] ),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\am_sdr0.cic0.integ2[6] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold1649 (.A(_01046_),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\am_sdr0.cic1.integ3[14] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\am_sdr0.cic2.comb1[8] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\am_sdr0.cic1.comb1[6] ),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\am_sdr0.cic0.integ1[19] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\am_sdr0.cic1.integ2[6] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold1655 (.A(_03847_),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\am_sdr0.cic3.comb1[18] ),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\am_sdr0.cic0.integ3[14] ),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\am_sdr0.cic2.integ1[12] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\am_sdr0.cic2.comb3_in_del[14] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\am_sdr0.cic2.comb3_in_del[15] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\am_sdr0.cic2.comb1[14] ),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\am_sdr0.cic1.comb2_in_del[9] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\am_sdr0.cic3.comb2_in_del[4] ),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\am_sdr0.cic0.comb1[10] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\am_sdr0.cic0.comb1_in_del[5] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\am_sdr0.cic1.integ1[12] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold1667 (.A(\am_sdr0.cic1.comb2[12] ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\am_sdr0.cic0.integ1[24] ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\am_sdr0.cic0.comb1[10] ),
    .X(net3328));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(rst_n));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(rst_n));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_antennanp ANTENNA_6 (.A(rst_n));
 sg13g2_antennanp ANTENNA_7 (.A(rst_n));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_fill_2 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_188 ();
 sg13g2_decap_4 FILLER_0_195 ();
 sg13g2_fill_1 FILLER_0_208 ();
 sg13g2_decap_4 FILLER_0_221 ();
 sg13g2_fill_2 FILLER_0_225 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_fill_2 FILLER_0_238 ();
 sg13g2_fill_2 FILLER_0_253 ();
 sg13g2_fill_2 FILLER_0_291 ();
 sg13g2_fill_1 FILLER_0_293 ();
 sg13g2_fill_2 FILLER_0_342 ();
 sg13g2_fill_2 FILLER_0_389 ();
 sg13g2_fill_1 FILLER_0_426 ();
 sg13g2_decap_4 FILLER_0_432 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_4 FILLER_0_469 ();
 sg13g2_fill_2 FILLER_0_473 ();
 sg13g2_fill_2 FILLER_0_501 ();
 sg13g2_fill_2 FILLER_0_516 ();
 sg13g2_fill_2 FILLER_0_531 ();
 sg13g2_fill_2 FILLER_0_563 ();
 sg13g2_fill_1 FILLER_0_599 ();
 sg13g2_fill_1 FILLER_0_608 ();
 sg13g2_decap_8 FILLER_0_617 ();
 sg13g2_fill_2 FILLER_0_624 ();
 sg13g2_fill_1 FILLER_0_626 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_fill_2 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_678 ();
 sg13g2_decap_8 FILLER_0_685 ();
 sg13g2_decap_8 FILLER_0_692 ();
 sg13g2_decap_8 FILLER_0_699 ();
 sg13g2_decap_8 FILLER_0_706 ();
 sg13g2_decap_8 FILLER_0_713 ();
 sg13g2_decap_8 FILLER_0_720 ();
 sg13g2_decap_8 FILLER_0_727 ();
 sg13g2_decap_8 FILLER_0_734 ();
 sg13g2_decap_8 FILLER_0_741 ();
 sg13g2_decap_8 FILLER_0_748 ();
 sg13g2_decap_8 FILLER_0_755 ();
 sg13g2_decap_8 FILLER_0_762 ();
 sg13g2_decap_8 FILLER_0_769 ();
 sg13g2_decap_8 FILLER_0_776 ();
 sg13g2_decap_8 FILLER_0_783 ();
 sg13g2_decap_8 FILLER_0_790 ();
 sg13g2_decap_8 FILLER_0_797 ();
 sg13g2_decap_8 FILLER_0_804 ();
 sg13g2_decap_8 FILLER_0_811 ();
 sg13g2_decap_8 FILLER_0_822 ();
 sg13g2_fill_2 FILLER_0_829 ();
 sg13g2_fill_2 FILLER_0_883 ();
 sg13g2_fill_1 FILLER_0_885 ();
 sg13g2_decap_4 FILLER_0_912 ();
 sg13g2_fill_1 FILLER_0_916 ();
 sg13g2_fill_2 FILLER_0_944 ();
 sg13g2_fill_1 FILLER_0_946 ();
 sg13g2_decap_4 FILLER_0_961 ();
 sg13g2_fill_2 FILLER_0_975 ();
 sg13g2_fill_1 FILLER_0_977 ();
 sg13g2_decap_8 FILLER_0_1017 ();
 sg13g2_decap_4 FILLER_0_1024 ();
 sg13g2_fill_1 FILLER_0_1028 ();
 sg13g2_fill_1 FILLER_0_1109 ();
 sg13g2_fill_2 FILLER_0_1136 ();
 sg13g2_fill_1 FILLER_0_1217 ();
 sg13g2_decap_8 FILLER_0_1246 ();
 sg13g2_decap_8 FILLER_0_1253 ();
 sg13g2_decap_8 FILLER_0_1260 ();
 sg13g2_decap_8 FILLER_0_1267 ();
 sg13g2_decap_8 FILLER_0_1274 ();
 sg13g2_decap_8 FILLER_0_1281 ();
 sg13g2_decap_8 FILLER_0_1288 ();
 sg13g2_decap_8 FILLER_0_1295 ();
 sg13g2_decap_8 FILLER_0_1302 ();
 sg13g2_decap_4 FILLER_0_1309 ();
 sg13g2_fill_2 FILLER_0_1313 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_4 FILLER_1_168 ();
 sg13g2_fill_2 FILLER_1_172 ();
 sg13g2_fill_2 FILLER_1_242 ();
 sg13g2_fill_1 FILLER_1_244 ();
 sg13g2_fill_2 FILLER_1_253 ();
 sg13g2_fill_1 FILLER_1_255 ();
 sg13g2_fill_1 FILLER_1_264 ();
 sg13g2_fill_1 FILLER_1_314 ();
 sg13g2_fill_1 FILLER_1_328 ();
 sg13g2_fill_2 FILLER_1_360 ();
 sg13g2_fill_2 FILLER_1_376 ();
 sg13g2_fill_1 FILLER_1_413 ();
 sg13g2_fill_2 FILLER_1_449 ();
 sg13g2_fill_1 FILLER_1_451 ();
 sg13g2_fill_1 FILLER_1_461 ();
 sg13g2_fill_2 FILLER_1_475 ();
 sg13g2_fill_2 FILLER_1_496 ();
 sg13g2_fill_1 FILLER_1_568 ();
 sg13g2_fill_2 FILLER_1_597 ();
 sg13g2_fill_1 FILLER_1_657 ();
 sg13g2_decap_8 FILLER_1_689 ();
 sg13g2_decap_8 FILLER_1_696 ();
 sg13g2_decap_4 FILLER_1_703 ();
 sg13g2_fill_2 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_4 FILLER_1_777 ();
 sg13g2_fill_1 FILLER_1_781 ();
 sg13g2_decap_8 FILLER_1_786 ();
 sg13g2_decap_8 FILLER_1_793 ();
 sg13g2_decap_8 FILLER_1_800 ();
 sg13g2_fill_2 FILLER_1_833 ();
 sg13g2_fill_2 FILLER_1_844 ();
 sg13g2_decap_4 FILLER_1_860 ();
 sg13g2_decap_8 FILLER_1_883 ();
 sg13g2_decap_8 FILLER_1_890 ();
 sg13g2_fill_2 FILLER_1_901 ();
 sg13g2_fill_1 FILLER_1_912 ();
 sg13g2_fill_1 FILLER_1_944 ();
 sg13g2_fill_1 FILLER_1_987 ();
 sg13g2_fill_1 FILLER_1_1002 ();
 sg13g2_fill_2 FILLER_1_1042 ();
 sg13g2_fill_1 FILLER_1_1044 ();
 sg13g2_fill_2 FILLER_1_1053 ();
 sg13g2_fill_1 FILLER_1_1105 ();
 sg13g2_fill_2 FILLER_1_1119 ();
 sg13g2_fill_2 FILLER_1_1125 ();
 sg13g2_fill_1 FILLER_1_1127 ();
 sg13g2_fill_1 FILLER_1_1150 ();
 sg13g2_decap_8 FILLER_1_1243 ();
 sg13g2_decap_8 FILLER_1_1250 ();
 sg13g2_decap_8 FILLER_1_1257 ();
 sg13g2_decap_8 FILLER_1_1264 ();
 sg13g2_decap_8 FILLER_1_1271 ();
 sg13g2_decap_8 FILLER_1_1278 ();
 sg13g2_decap_8 FILLER_1_1285 ();
 sg13g2_decap_8 FILLER_1_1292 ();
 sg13g2_decap_8 FILLER_1_1299 ();
 sg13g2_decap_8 FILLER_1_1306 ();
 sg13g2_fill_2 FILLER_1_1313 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_fill_2 FILLER_2_182 ();
 sg13g2_fill_1 FILLER_2_198 ();
 sg13g2_decap_4 FILLER_2_221 ();
 sg13g2_fill_1 FILLER_2_284 ();
 sg13g2_decap_4 FILLER_2_289 ();
 sg13g2_fill_1 FILLER_2_314 ();
 sg13g2_fill_1 FILLER_2_460 ();
 sg13g2_fill_2 FILLER_2_469 ();
 sg13g2_fill_2 FILLER_2_485 ();
 sg13g2_fill_2 FILLER_2_518 ();
 sg13g2_fill_1 FILLER_2_536 ();
 sg13g2_fill_2 FILLER_2_554 ();
 sg13g2_fill_1 FILLER_2_653 ();
 sg13g2_fill_1 FILLER_2_697 ();
 sg13g2_decap_8 FILLER_2_731 ();
 sg13g2_decap_4 FILLER_2_738 ();
 sg13g2_fill_2 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_4 FILLER_2_756 ();
 sg13g2_fill_1 FILLER_2_760 ();
 sg13g2_fill_1 FILLER_2_821 ();
 sg13g2_fill_1 FILLER_2_848 ();
 sg13g2_fill_2 FILLER_2_921 ();
 sg13g2_fill_2 FILLER_2_927 ();
 sg13g2_decap_8 FILLER_2_933 ();
 sg13g2_fill_2 FILLER_2_940 ();
 sg13g2_decap_4 FILLER_2_950 ();
 sg13g2_fill_2 FILLER_2_971 ();
 sg13g2_fill_2 FILLER_2_978 ();
 sg13g2_fill_1 FILLER_2_980 ();
 sg13g2_fill_2 FILLER_2_997 ();
 sg13g2_fill_1 FILLER_2_1018 ();
 sg13g2_fill_1 FILLER_2_1033 ();
 sg13g2_fill_1 FILLER_2_1060 ();
 sg13g2_fill_2 FILLER_2_1101 ();
 sg13g2_decap_4 FILLER_2_1108 ();
 sg13g2_fill_1 FILLER_2_1112 ();
 sg13g2_fill_1 FILLER_2_1175 ();
 sg13g2_fill_2 FILLER_2_1188 ();
 sg13g2_fill_1 FILLER_2_1190 ();
 sg13g2_fill_1 FILLER_2_1217 ();
 sg13g2_decap_8 FILLER_2_1250 ();
 sg13g2_decap_8 FILLER_2_1257 ();
 sg13g2_decap_8 FILLER_2_1264 ();
 sg13g2_decap_8 FILLER_2_1271 ();
 sg13g2_decap_8 FILLER_2_1278 ();
 sg13g2_decap_8 FILLER_2_1285 ();
 sg13g2_decap_8 FILLER_2_1292 ();
 sg13g2_decap_8 FILLER_2_1299 ();
 sg13g2_decap_8 FILLER_2_1306 ();
 sg13g2_fill_2 FILLER_2_1313 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_4 FILLER_3_168 ();
 sg13g2_fill_1 FILLER_3_172 ();
 sg13g2_fill_1 FILLER_3_238 ();
 sg13g2_fill_1 FILLER_3_247 ();
 sg13g2_fill_2 FILLER_3_369 ();
 sg13g2_fill_1 FILLER_3_371 ();
 sg13g2_fill_1 FILLER_3_402 ();
 sg13g2_decap_4 FILLER_3_463 ();
 sg13g2_decap_8 FILLER_3_500 ();
 sg13g2_fill_2 FILLER_3_507 ();
 sg13g2_fill_2 FILLER_3_543 ();
 sg13g2_fill_2 FILLER_3_586 ();
 sg13g2_fill_1 FILLER_3_597 ();
 sg13g2_fill_2 FILLER_3_608 ();
 sg13g2_fill_1 FILLER_3_615 ();
 sg13g2_fill_2 FILLER_3_621 ();
 sg13g2_fill_1 FILLER_3_627 ();
 sg13g2_fill_1 FILLER_3_637 ();
 sg13g2_fill_1 FILLER_3_642 ();
 sg13g2_decap_4 FILLER_3_659 ();
 sg13g2_fill_1 FILLER_3_672 ();
 sg13g2_fill_1 FILLER_3_727 ();
 sg13g2_fill_2 FILLER_3_767 ();
 sg13g2_fill_1 FILLER_3_769 ();
 sg13g2_fill_1 FILLER_3_784 ();
 sg13g2_fill_1 FILLER_3_799 ();
 sg13g2_decap_8 FILLER_3_813 ();
 sg13g2_fill_2 FILLER_3_820 ();
 sg13g2_fill_1 FILLER_3_822 ();
 sg13g2_decap_4 FILLER_3_839 ();
 sg13g2_fill_1 FILLER_3_843 ();
 sg13g2_fill_2 FILLER_3_849 ();
 sg13g2_fill_1 FILLER_3_851 ();
 sg13g2_fill_2 FILLER_3_856 ();
 sg13g2_decap_4 FILLER_3_867 ();
 sg13g2_fill_1 FILLER_3_880 ();
 sg13g2_fill_2 FILLER_3_884 ();
 sg13g2_fill_1 FILLER_3_886 ();
 sg13g2_fill_2 FILLER_3_907 ();
 sg13g2_fill_1 FILLER_3_909 ();
 sg13g2_fill_2 FILLER_3_944 ();
 sg13g2_fill_2 FILLER_3_950 ();
 sg13g2_fill_1 FILLER_3_952 ();
 sg13g2_fill_2 FILLER_3_975 ();
 sg13g2_fill_1 FILLER_3_977 ();
 sg13g2_fill_2 FILLER_3_991 ();
 sg13g2_fill_1 FILLER_3_993 ();
 sg13g2_fill_2 FILLER_3_1050 ();
 sg13g2_fill_1 FILLER_3_1052 ();
 sg13g2_fill_1 FILLER_3_1056 ();
 sg13g2_fill_1 FILLER_3_1074 ();
 sg13g2_fill_2 FILLER_3_1088 ();
 sg13g2_fill_1 FILLER_3_1090 ();
 sg13g2_fill_1 FILLER_3_1123 ();
 sg13g2_decap_8 FILLER_3_1133 ();
 sg13g2_decap_4 FILLER_3_1140 ();
 sg13g2_fill_1 FILLER_3_1144 ();
 sg13g2_decap_8 FILLER_3_1188 ();
 sg13g2_fill_1 FILLER_3_1195 ();
 sg13g2_fill_1 FILLER_3_1201 ();
 sg13g2_decap_8 FILLER_3_1206 ();
 sg13g2_decap_8 FILLER_3_1254 ();
 sg13g2_decap_8 FILLER_3_1261 ();
 sg13g2_decap_8 FILLER_3_1268 ();
 sg13g2_decap_8 FILLER_3_1275 ();
 sg13g2_decap_8 FILLER_3_1282 ();
 sg13g2_decap_8 FILLER_3_1289 ();
 sg13g2_decap_8 FILLER_3_1296 ();
 sg13g2_decap_8 FILLER_3_1303 ();
 sg13g2_decap_4 FILLER_3_1310 ();
 sg13g2_fill_1 FILLER_3_1314 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_fill_2 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_188 ();
 sg13g2_fill_2 FILLER_4_195 ();
 sg13g2_fill_1 FILLER_4_209 ();
 sg13g2_decap_8 FILLER_4_242 ();
 sg13g2_fill_2 FILLER_4_258 ();
 sg13g2_decap_8 FILLER_4_264 ();
 sg13g2_fill_2 FILLER_4_271 ();
 sg13g2_decap_8 FILLER_4_277 ();
 sg13g2_fill_2 FILLER_4_355 ();
 sg13g2_fill_2 FILLER_4_366 ();
 sg13g2_fill_1 FILLER_4_368 ();
 sg13g2_fill_1 FILLER_4_382 ();
 sg13g2_fill_2 FILLER_4_399 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_fill_1 FILLER_4_439 ();
 sg13g2_fill_1 FILLER_4_448 ();
 sg13g2_fill_1 FILLER_4_465 ();
 sg13g2_fill_2 FILLER_4_536 ();
 sg13g2_fill_2 FILLER_4_585 ();
 sg13g2_decap_4 FILLER_4_613 ();
 sg13g2_fill_2 FILLER_4_617 ();
 sg13g2_fill_2 FILLER_4_648 ();
 sg13g2_fill_1 FILLER_4_650 ();
 sg13g2_fill_1 FILLER_4_746 ();
 sg13g2_fill_2 FILLER_4_777 ();
 sg13g2_fill_1 FILLER_4_779 ();
 sg13g2_decap_4 FILLER_4_801 ();
 sg13g2_fill_2 FILLER_4_805 ();
 sg13g2_decap_4 FILLER_4_833 ();
 sg13g2_fill_2 FILLER_4_837 ();
 sg13g2_decap_4 FILLER_4_843 ();
 sg13g2_fill_2 FILLER_4_857 ();
 sg13g2_fill_1 FILLER_4_864 ();
 sg13g2_fill_2 FILLER_4_873 ();
 sg13g2_fill_1 FILLER_4_898 ();
 sg13g2_fill_1 FILLER_4_925 ();
 sg13g2_fill_1 FILLER_4_944 ();
 sg13g2_decap_4 FILLER_4_971 ();
 sg13g2_fill_1 FILLER_4_975 ();
 sg13g2_fill_2 FILLER_4_1030 ();
 sg13g2_fill_1 FILLER_4_1032 ();
 sg13g2_decap_8 FILLER_4_1108 ();
 sg13g2_fill_2 FILLER_4_1115 ();
 sg13g2_fill_2 FILLER_4_1148 ();
 sg13g2_fill_1 FILLER_4_1150 ();
 sg13g2_fill_2 FILLER_4_1156 ();
 sg13g2_decap_8 FILLER_4_1210 ();
 sg13g2_decap_8 FILLER_4_1251 ();
 sg13g2_decap_8 FILLER_4_1258 ();
 sg13g2_decap_8 FILLER_4_1265 ();
 sg13g2_decap_8 FILLER_4_1272 ();
 sg13g2_decap_8 FILLER_4_1279 ();
 sg13g2_decap_8 FILLER_4_1286 ();
 sg13g2_decap_8 FILLER_4_1293 ();
 sg13g2_decap_8 FILLER_4_1300 ();
 sg13g2_decap_8 FILLER_4_1307 ();
 sg13g2_fill_1 FILLER_4_1314 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_fill_1 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_180 ();
 sg13g2_decap_4 FILLER_5_205 ();
 sg13g2_fill_2 FILLER_5_239 ();
 sg13g2_fill_2 FILLER_5_275 ();
 sg13g2_fill_2 FILLER_5_303 ();
 sg13g2_fill_1 FILLER_5_305 ();
 sg13g2_fill_1 FILLER_5_311 ();
 sg13g2_fill_1 FILLER_5_384 ();
 sg13g2_fill_2 FILLER_5_421 ();
 sg13g2_fill_1 FILLER_5_423 ();
 sg13g2_decap_4 FILLER_5_434 ();
 sg13g2_fill_1 FILLER_5_438 ();
 sg13g2_decap_4 FILLER_5_442 ();
 sg13g2_decap_8 FILLER_5_463 ();
 sg13g2_fill_1 FILLER_5_470 ();
 sg13g2_decap_4 FILLER_5_476 ();
 sg13g2_fill_2 FILLER_5_480 ();
 sg13g2_decap_8 FILLER_5_486 ();
 sg13g2_fill_2 FILLER_5_501 ();
 sg13g2_decap_4 FILLER_5_507 ();
 sg13g2_fill_1 FILLER_5_525 ();
 sg13g2_fill_1 FILLER_5_538 ();
 sg13g2_fill_2 FILLER_5_573 ();
 sg13g2_decap_8 FILLER_5_587 ();
 sg13g2_fill_2 FILLER_5_594 ();
 sg13g2_fill_1 FILLER_5_596 ();
 sg13g2_fill_1 FILLER_5_606 ();
 sg13g2_decap_4 FILLER_5_612 ();
 sg13g2_fill_2 FILLER_5_616 ();
 sg13g2_fill_2 FILLER_5_747 ();
 sg13g2_fill_2 FILLER_5_759 ();
 sg13g2_fill_1 FILLER_5_770 ();
 sg13g2_fill_2 FILLER_5_776 ();
 sg13g2_fill_1 FILLER_5_778 ();
 sg13g2_fill_2 FILLER_5_884 ();
 sg13g2_decap_4 FILLER_5_904 ();
 sg13g2_fill_2 FILLER_5_908 ();
 sg13g2_decap_4 FILLER_5_923 ();
 sg13g2_fill_1 FILLER_5_927 ();
 sg13g2_fill_2 FILLER_5_935 ();
 sg13g2_fill_1 FILLER_5_944 ();
 sg13g2_fill_2 FILLER_5_960 ();
 sg13g2_decap_4 FILLER_5_976 ();
 sg13g2_fill_1 FILLER_5_980 ();
 sg13g2_fill_2 FILLER_5_1001 ();
 sg13g2_fill_1 FILLER_5_1003 ();
 sg13g2_fill_1 FILLER_5_1021 ();
 sg13g2_fill_2 FILLER_5_1062 ();
 sg13g2_decap_4 FILLER_5_1078 ();
 sg13g2_fill_1 FILLER_5_1087 ();
 sg13g2_fill_2 FILLER_5_1098 ();
 sg13g2_fill_1 FILLER_5_1100 ();
 sg13g2_decap_8 FILLER_5_1124 ();
 sg13g2_fill_1 FILLER_5_1131 ();
 sg13g2_fill_2 FILLER_5_1149 ();
 sg13g2_fill_2 FILLER_5_1221 ();
 sg13g2_fill_1 FILLER_5_1223 ();
 sg13g2_decap_8 FILLER_5_1263 ();
 sg13g2_decap_8 FILLER_5_1270 ();
 sg13g2_decap_8 FILLER_5_1277 ();
 sg13g2_decap_8 FILLER_5_1284 ();
 sg13g2_decap_8 FILLER_5_1291 ();
 sg13g2_decap_8 FILLER_5_1298 ();
 sg13g2_decap_8 FILLER_5_1305 ();
 sg13g2_fill_2 FILLER_5_1312 ();
 sg13g2_fill_1 FILLER_5_1314 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_4 FILLER_6_161 ();
 sg13g2_fill_1 FILLER_6_165 ();
 sg13g2_fill_2 FILLER_6_200 ();
 sg13g2_fill_1 FILLER_6_202 ();
 sg13g2_fill_1 FILLER_6_221 ();
 sg13g2_fill_1 FILLER_6_280 ();
 sg13g2_fill_2 FILLER_6_311 ();
 sg13g2_fill_1 FILLER_6_313 ();
 sg13g2_fill_2 FILLER_6_354 ();
 sg13g2_fill_1 FILLER_6_365 ();
 sg13g2_decap_8 FILLER_6_404 ();
 sg13g2_fill_1 FILLER_6_416 ();
 sg13g2_fill_2 FILLER_6_426 ();
 sg13g2_fill_1 FILLER_6_428 ();
 sg13g2_fill_1 FILLER_6_439 ();
 sg13g2_decap_8 FILLER_6_456 ();
 sg13g2_fill_1 FILLER_6_507 ();
 sg13g2_fill_2 FILLER_6_548 ();
 sg13g2_fill_1 FILLER_6_563 ();
 sg13g2_decap_4 FILLER_6_580 ();
 sg13g2_fill_2 FILLER_6_584 ();
 sg13g2_decap_4 FILLER_6_591 ();
 sg13g2_decap_4 FILLER_6_599 ();
 sg13g2_fill_1 FILLER_6_603 ();
 sg13g2_fill_2 FILLER_6_635 ();
 sg13g2_fill_1 FILLER_6_651 ();
 sg13g2_fill_2 FILLER_6_689 ();
 sg13g2_fill_1 FILLER_6_760 ();
 sg13g2_fill_2 FILLER_6_801 ();
 sg13g2_decap_8 FILLER_6_855 ();
 sg13g2_decap_4 FILLER_6_862 ();
 sg13g2_fill_2 FILLER_6_872 ();
 sg13g2_fill_2 FILLER_6_895 ();
 sg13g2_fill_2 FILLER_6_907 ();
 sg13g2_fill_2 FILLER_6_927 ();
 sg13g2_decap_4 FILLER_6_948 ();
 sg13g2_fill_1 FILLER_6_982 ();
 sg13g2_fill_1 FILLER_6_999 ();
 sg13g2_fill_2 FILLER_6_1026 ();
 sg13g2_fill_1 FILLER_6_1162 ();
 sg13g2_fill_2 FILLER_6_1172 ();
 sg13g2_fill_1 FILLER_6_1174 ();
 sg13g2_fill_2 FILLER_6_1258 ();
 sg13g2_fill_1 FILLER_6_1260 ();
 sg13g2_decap_8 FILLER_6_1270 ();
 sg13g2_decap_8 FILLER_6_1277 ();
 sg13g2_decap_8 FILLER_6_1284 ();
 sg13g2_decap_8 FILLER_6_1291 ();
 sg13g2_decap_8 FILLER_6_1298 ();
 sg13g2_decap_8 FILLER_6_1305 ();
 sg13g2_fill_2 FILLER_6_1312 ();
 sg13g2_fill_1 FILLER_6_1314 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_4 FILLER_7_184 ();
 sg13g2_fill_2 FILLER_7_188 ();
 sg13g2_fill_2 FILLER_7_214 ();
 sg13g2_decap_8 FILLER_7_251 ();
 sg13g2_decap_8 FILLER_7_258 ();
 sg13g2_decap_8 FILLER_7_269 ();
 sg13g2_fill_2 FILLER_7_276 ();
 sg13g2_fill_2 FILLER_7_283 ();
 sg13g2_fill_2 FILLER_7_301 ();
 sg13g2_fill_1 FILLER_7_303 ();
 sg13g2_fill_2 FILLER_7_312 ();
 sg13g2_fill_1 FILLER_7_314 ();
 sg13g2_fill_1 FILLER_7_349 ();
 sg13g2_fill_1 FILLER_7_374 ();
 sg13g2_fill_1 FILLER_7_383 ();
 sg13g2_fill_1 FILLER_7_432 ();
 sg13g2_decap_4 FILLER_7_458 ();
 sg13g2_fill_1 FILLER_7_462 ();
 sg13g2_fill_1 FILLER_7_476 ();
 sg13g2_fill_1 FILLER_7_518 ();
 sg13g2_fill_2 FILLER_7_555 ();
 sg13g2_fill_1 FILLER_7_557 ();
 sg13g2_fill_2 FILLER_7_570 ();
 sg13g2_decap_4 FILLER_7_580 ();
 sg13g2_fill_1 FILLER_7_615 ();
 sg13g2_fill_2 FILLER_7_621 ();
 sg13g2_fill_2 FILLER_7_667 ();
 sg13g2_fill_1 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_739 ();
 sg13g2_decap_8 FILLER_7_746 ();
 sg13g2_decap_4 FILLER_7_753 ();
 sg13g2_decap_8 FILLER_7_766 ();
 sg13g2_decap_8 FILLER_7_773 ();
 sg13g2_fill_2 FILLER_7_824 ();
 sg13g2_fill_2 FILLER_7_867 ();
 sg13g2_fill_2 FILLER_7_882 ();
 sg13g2_decap_8 FILLER_7_889 ();
 sg13g2_decap_4 FILLER_7_896 ();
 sg13g2_fill_1 FILLER_7_900 ();
 sg13g2_decap_4 FILLER_7_927 ();
 sg13g2_fill_1 FILLER_7_931 ();
 sg13g2_decap_8 FILLER_7_947 ();
 sg13g2_decap_8 FILLER_7_968 ();
 sg13g2_decap_4 FILLER_7_975 ();
 sg13g2_fill_1 FILLER_7_979 ();
 sg13g2_fill_1 FILLER_7_1015 ();
 sg13g2_fill_2 FILLER_7_1090 ();
 sg13g2_fill_1 FILLER_7_1092 ();
 sg13g2_fill_1 FILLER_7_1102 ();
 sg13g2_fill_2 FILLER_7_1127 ();
 sg13g2_decap_8 FILLER_7_1133 ();
 sg13g2_fill_2 FILLER_7_1140 ();
 sg13g2_fill_1 FILLER_7_1142 ();
 sg13g2_fill_1 FILLER_7_1186 ();
 sg13g2_decap_8 FILLER_7_1192 ();
 sg13g2_fill_2 FILLER_7_1199 ();
 sg13g2_fill_1 FILLER_7_1217 ();
 sg13g2_decap_8 FILLER_7_1261 ();
 sg13g2_decap_8 FILLER_7_1268 ();
 sg13g2_decap_8 FILLER_7_1275 ();
 sg13g2_decap_8 FILLER_7_1282 ();
 sg13g2_decap_8 FILLER_7_1289 ();
 sg13g2_decap_8 FILLER_7_1296 ();
 sg13g2_decap_8 FILLER_7_1303 ();
 sg13g2_decap_4 FILLER_7_1310 ();
 sg13g2_fill_1 FILLER_7_1314 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_4 FILLER_8_161 ();
 sg13g2_fill_1 FILLER_8_165 ();
 sg13g2_fill_1 FILLER_8_170 ();
 sg13g2_fill_2 FILLER_8_200 ();
 sg13g2_fill_1 FILLER_8_216 ();
 sg13g2_fill_1 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_275 ();
 sg13g2_decap_8 FILLER_8_282 ();
 sg13g2_fill_1 FILLER_8_289 ();
 sg13g2_fill_2 FILLER_8_316 ();
 sg13g2_fill_2 FILLER_8_332 ();
 sg13g2_fill_1 FILLER_8_342 ();
 sg13g2_fill_2 FILLER_8_386 ();
 sg13g2_fill_2 FILLER_8_402 ();
 sg13g2_fill_2 FILLER_8_415 ();
 sg13g2_fill_2 FILLER_8_422 ();
 sg13g2_fill_2 FILLER_8_455 ();
 sg13g2_decap_4 FILLER_8_462 ();
 sg13g2_fill_1 FILLER_8_494 ();
 sg13g2_fill_1 FILLER_8_527 ();
 sg13g2_fill_1 FILLER_8_542 ();
 sg13g2_fill_1 FILLER_8_561 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_fill_2 FILLER_8_581 ();
 sg13g2_fill_1 FILLER_8_583 ();
 sg13g2_decap_8 FILLER_8_589 ();
 sg13g2_fill_2 FILLER_8_596 ();
 sg13g2_decap_8 FILLER_8_603 ();
 sg13g2_fill_2 FILLER_8_652 ();
 sg13g2_fill_1 FILLER_8_654 ();
 sg13g2_fill_2 FILLER_8_698 ();
 sg13g2_fill_1 FILLER_8_712 ();
 sg13g2_fill_2 FILLER_8_799 ();
 sg13g2_fill_1 FILLER_8_801 ();
 sg13g2_decap_8 FILLER_8_815 ();
 sg13g2_fill_1 FILLER_8_822 ();
 sg13g2_decap_4 FILLER_8_854 ();
 sg13g2_decap_8 FILLER_8_866 ();
 sg13g2_fill_2 FILLER_8_873 ();
 sg13g2_decap_4 FILLER_8_884 ();
 sg13g2_fill_1 FILLER_8_888 ();
 sg13g2_fill_1 FILLER_8_907 ();
 sg13g2_decap_8 FILLER_8_921 ();
 sg13g2_fill_1 FILLER_8_928 ();
 sg13g2_fill_2 FILLER_8_951 ();
 sg13g2_fill_1 FILLER_8_953 ();
 sg13g2_fill_2 FILLER_8_1026 ();
 sg13g2_fill_2 FILLER_8_1056 ();
 sg13g2_fill_2 FILLER_8_1116 ();
 sg13g2_fill_1 FILLER_8_1118 ();
 sg13g2_fill_2 FILLER_8_1145 ();
 sg13g2_fill_1 FILLER_8_1147 ();
 sg13g2_fill_2 FILLER_8_1242 ();
 sg13g2_decap_8 FILLER_8_1251 ();
 sg13g2_decap_8 FILLER_8_1258 ();
 sg13g2_decap_8 FILLER_8_1265 ();
 sg13g2_decap_8 FILLER_8_1272 ();
 sg13g2_decap_8 FILLER_8_1279 ();
 sg13g2_decap_8 FILLER_8_1286 ();
 sg13g2_decap_8 FILLER_8_1293 ();
 sg13g2_decap_8 FILLER_8_1300 ();
 sg13g2_decap_8 FILLER_8_1307 ();
 sg13g2_fill_1 FILLER_8_1314 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_fill_1 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_185 ();
 sg13g2_fill_1 FILLER_9_192 ();
 sg13g2_decap_8 FILLER_9_197 ();
 sg13g2_decap_8 FILLER_9_218 ();
 sg13g2_fill_2 FILLER_9_225 ();
 sg13g2_fill_1 FILLER_9_288 ();
 sg13g2_fill_1 FILLER_9_297 ();
 sg13g2_decap_4 FILLER_9_307 ();
 sg13g2_fill_1 FILLER_9_315 ();
 sg13g2_fill_2 FILLER_9_331 ();
 sg13g2_fill_1 FILLER_9_359 ();
 sg13g2_fill_2 FILLER_9_369 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_443 ();
 sg13g2_fill_1 FILLER_9_449 ();
 sg13g2_fill_2 FILLER_9_541 ();
 sg13g2_fill_1 FILLER_9_553 ();
 sg13g2_fill_2 FILLER_9_565 ();
 sg13g2_fill_2 FILLER_9_619 ();
 sg13g2_fill_2 FILLER_9_631 ();
 sg13g2_fill_2 FILLER_9_689 ();
 sg13g2_fill_2 FILLER_9_753 ();
 sg13g2_fill_1 FILLER_9_760 ();
 sg13g2_decap_8 FILLER_9_766 ();
 sg13g2_fill_1 FILLER_9_773 ();
 sg13g2_decap_4 FILLER_9_782 ();
 sg13g2_fill_1 FILLER_9_786 ();
 sg13g2_decap_4 FILLER_9_805 ();
 sg13g2_fill_2 FILLER_9_809 ();
 sg13g2_fill_1 FILLER_9_824 ();
 sg13g2_fill_1 FILLER_9_843 ();
 sg13g2_decap_4 FILLER_9_848 ();
 sg13g2_fill_1 FILLER_9_852 ();
 sg13g2_fill_2 FILLER_9_858 ();
 sg13g2_fill_1 FILLER_9_860 ();
 sg13g2_fill_2 FILLER_9_874 ();
 sg13g2_fill_1 FILLER_9_876 ();
 sg13g2_fill_1 FILLER_9_926 ();
 sg13g2_decap_8 FILLER_9_950 ();
 sg13g2_fill_2 FILLER_9_957 ();
 sg13g2_fill_1 FILLER_9_959 ();
 sg13g2_decap_4 FILLER_9_969 ();
 sg13g2_fill_2 FILLER_9_982 ();
 sg13g2_decap_4 FILLER_9_995 ();
 sg13g2_fill_1 FILLER_9_999 ();
 sg13g2_fill_2 FILLER_9_1015 ();
 sg13g2_fill_1 FILLER_9_1017 ();
 sg13g2_fill_2 FILLER_9_1036 ();
 sg13g2_fill_2 FILLER_9_1064 ();
 sg13g2_fill_2 FILLER_9_1091 ();
 sg13g2_fill_2 FILLER_9_1121 ();
 sg13g2_fill_1 FILLER_9_1123 ();
 sg13g2_fill_2 FILLER_9_1143 ();
 sg13g2_fill_2 FILLER_9_1150 ();
 sg13g2_fill_1 FILLER_9_1220 ();
 sg13g2_fill_2 FILLER_9_1233 ();
 sg13g2_decap_8 FILLER_9_1261 ();
 sg13g2_decap_8 FILLER_9_1268 ();
 sg13g2_decap_8 FILLER_9_1275 ();
 sg13g2_decap_8 FILLER_9_1282 ();
 sg13g2_decap_8 FILLER_9_1289 ();
 sg13g2_decap_8 FILLER_9_1296 ();
 sg13g2_decap_8 FILLER_9_1303 ();
 sg13g2_decap_4 FILLER_9_1310 ();
 sg13g2_fill_1 FILLER_9_1314 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_fill_2 FILLER_10_168 ();
 sg13g2_fill_1 FILLER_10_170 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_fill_2 FILLER_10_182 ();
 sg13g2_fill_2 FILLER_10_189 ();
 sg13g2_fill_1 FILLER_10_191 ();
 sg13g2_fill_1 FILLER_10_197 ();
 sg13g2_decap_8 FILLER_10_216 ();
 sg13g2_decap_8 FILLER_10_223 ();
 sg13g2_fill_2 FILLER_10_253 ();
 sg13g2_fill_1 FILLER_10_255 ();
 sg13g2_fill_2 FILLER_10_260 ();
 sg13g2_fill_1 FILLER_10_262 ();
 sg13g2_fill_1 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_decap_4 FILLER_10_289 ();
 sg13g2_fill_1 FILLER_10_293 ();
 sg13g2_fill_2 FILLER_10_315 ();
 sg13g2_fill_1 FILLER_10_317 ();
 sg13g2_decap_4 FILLER_10_339 ();
 sg13g2_fill_2 FILLER_10_343 ();
 sg13g2_fill_2 FILLER_10_349 ();
 sg13g2_fill_1 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_412 ();
 sg13g2_fill_1 FILLER_10_440 ();
 sg13g2_fill_2 FILLER_10_451 ();
 sg13g2_decap_4 FILLER_10_501 ();
 sg13g2_fill_2 FILLER_10_514 ();
 sg13g2_fill_1 FILLER_10_516 ();
 sg13g2_fill_2 FILLER_10_534 ();
 sg13g2_fill_1 FILLER_10_536 ();
 sg13g2_fill_1 FILLER_10_551 ();
 sg13g2_decap_4 FILLER_10_590 ();
 sg13g2_decap_8 FILLER_10_598 ();
 sg13g2_fill_2 FILLER_10_605 ();
 sg13g2_fill_1 FILLER_10_607 ();
 sg13g2_fill_2 FILLER_10_649 ();
 sg13g2_fill_2 FILLER_10_669 ();
 sg13g2_fill_2 FILLER_10_685 ();
 sg13g2_fill_2 FILLER_10_695 ();
 sg13g2_decap_4 FILLER_10_737 ();
 sg13g2_fill_2 FILLER_10_745 ();
 sg13g2_decap_4 FILLER_10_752 ();
 sg13g2_fill_1 FILLER_10_756 ();
 sg13g2_decap_4 FILLER_10_765 ();
 sg13g2_fill_1 FILLER_10_769 ();
 sg13g2_fill_2 FILLER_10_832 ();
 sg13g2_fill_2 FILLER_10_893 ();
 sg13g2_fill_1 FILLER_10_895 ();
 sg13g2_decap_4 FILLER_10_909 ();
 sg13g2_fill_2 FILLER_10_913 ();
 sg13g2_decap_8 FILLER_10_919 ();
 sg13g2_fill_2 FILLER_10_926 ();
 sg13g2_fill_1 FILLER_10_928 ();
 sg13g2_fill_1 FILLER_10_945 ();
 sg13g2_fill_2 FILLER_10_954 ();
 sg13g2_fill_1 FILLER_10_956 ();
 sg13g2_fill_2 FILLER_10_988 ();
 sg13g2_fill_1 FILLER_10_990 ();
 sg13g2_fill_2 FILLER_10_1012 ();
 sg13g2_fill_1 FILLER_10_1014 ();
 sg13g2_fill_1 FILLER_10_1019 ();
 sg13g2_fill_2 FILLER_10_1030 ();
 sg13g2_fill_1 FILLER_10_1032 ();
 sg13g2_decap_4 FILLER_10_1059 ();
 sg13g2_fill_2 FILLER_10_1063 ();
 sg13g2_fill_2 FILLER_10_1070 ();
 sg13g2_fill_1 FILLER_10_1085 ();
 sg13g2_fill_2 FILLER_10_1095 ();
 sg13g2_fill_2 FILLER_10_1119 ();
 sg13g2_fill_2 FILLER_10_1143 ();
 sg13g2_fill_1 FILLER_10_1145 ();
 sg13g2_fill_2 FILLER_10_1197 ();
 sg13g2_fill_1 FILLER_10_1234 ();
 sg13g2_decap_8 FILLER_10_1258 ();
 sg13g2_decap_8 FILLER_10_1265 ();
 sg13g2_decap_8 FILLER_10_1272 ();
 sg13g2_decap_8 FILLER_10_1279 ();
 sg13g2_decap_8 FILLER_10_1286 ();
 sg13g2_decap_8 FILLER_10_1293 ();
 sg13g2_decap_8 FILLER_10_1300 ();
 sg13g2_decap_8 FILLER_10_1307 ();
 sg13g2_fill_1 FILLER_10_1314 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_4 FILLER_11_154 ();
 sg13g2_fill_2 FILLER_11_158 ();
 sg13g2_fill_2 FILLER_11_194 ();
 sg13g2_fill_1 FILLER_11_315 ();
 sg13g2_fill_2 FILLER_11_442 ();
 sg13g2_fill_2 FILLER_11_448 ();
 sg13g2_decap_4 FILLER_11_458 ();
 sg13g2_fill_1 FILLER_11_493 ();
 sg13g2_fill_2 FILLER_11_520 ();
 sg13g2_decap_4 FILLER_11_582 ();
 sg13g2_fill_2 FILLER_11_617 ();
 sg13g2_fill_1 FILLER_11_619 ();
 sg13g2_fill_1 FILLER_11_655 ();
 sg13g2_fill_2 FILLER_11_673 ();
 sg13g2_fill_1 FILLER_11_675 ();
 sg13g2_fill_1 FILLER_11_702 ();
 sg13g2_fill_1 FILLER_11_773 ();
 sg13g2_fill_2 FILLER_11_793 ();
 sg13g2_fill_2 FILLER_11_800 ();
 sg13g2_fill_1 FILLER_11_811 ();
 sg13g2_fill_2 FILLER_11_826 ();
 sg13g2_fill_1 FILLER_11_833 ();
 sg13g2_fill_1 FILLER_11_843 ();
 sg13g2_fill_2 FILLER_11_857 ();
 sg13g2_fill_1 FILLER_11_859 ();
 sg13g2_fill_2 FILLER_11_868 ();
 sg13g2_fill_2 FILLER_11_888 ();
 sg13g2_fill_1 FILLER_11_898 ();
 sg13g2_fill_2 FILLER_11_944 ();
 sg13g2_fill_1 FILLER_11_946 ();
 sg13g2_decap_8 FILLER_11_977 ();
 sg13g2_decap_4 FILLER_11_984 ();
 sg13g2_fill_2 FILLER_11_996 ();
 sg13g2_fill_1 FILLER_11_998 ();
 sg13g2_fill_1 FILLER_11_1042 ();
 sg13g2_fill_2 FILLER_11_1051 ();
 sg13g2_decap_4 FILLER_11_1057 ();
 sg13g2_fill_1 FILLER_11_1061 ();
 sg13g2_decap_4 FILLER_11_1113 ();
 sg13g2_fill_2 FILLER_11_1117 ();
 sg13g2_fill_1 FILLER_11_1164 ();
 sg13g2_fill_2 FILLER_11_1195 ();
 sg13g2_fill_1 FILLER_11_1197 ();
 sg13g2_fill_1 FILLER_11_1224 ();
 sg13g2_decap_8 FILLER_11_1256 ();
 sg13g2_decap_8 FILLER_11_1263 ();
 sg13g2_decap_8 FILLER_11_1270 ();
 sg13g2_decap_8 FILLER_11_1277 ();
 sg13g2_decap_8 FILLER_11_1284 ();
 sg13g2_decap_8 FILLER_11_1291 ();
 sg13g2_decap_8 FILLER_11_1298 ();
 sg13g2_decap_8 FILLER_11_1305 ();
 sg13g2_fill_2 FILLER_11_1312 ();
 sg13g2_fill_1 FILLER_11_1314 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_fill_2 FILLER_12_175 ();
 sg13g2_fill_1 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_206 ();
 sg13g2_decap_8 FILLER_12_216 ();
 sg13g2_fill_1 FILLER_12_236 ();
 sg13g2_fill_2 FILLER_12_254 ();
 sg13g2_fill_2 FILLER_12_260 ();
 sg13g2_fill_1 FILLER_12_262 ();
 sg13g2_fill_1 FILLER_12_297 ();
 sg13g2_fill_1 FILLER_12_307 ();
 sg13g2_fill_2 FILLER_12_321 ();
 sg13g2_fill_2 FILLER_12_327 ();
 sg13g2_fill_2 FILLER_12_390 ();
 sg13g2_fill_1 FILLER_12_436 ();
 sg13g2_fill_1 FILLER_12_448 ();
 sg13g2_fill_1 FILLER_12_475 ();
 sg13g2_fill_1 FILLER_12_504 ();
 sg13g2_fill_2 FILLER_12_536 ();
 sg13g2_fill_2 FILLER_12_546 ();
 sg13g2_fill_2 FILLER_12_608 ();
 sg13g2_fill_1 FILLER_12_610 ();
 sg13g2_fill_2 FILLER_12_616 ();
 sg13g2_fill_1 FILLER_12_618 ();
 sg13g2_fill_2 FILLER_12_660 ();
 sg13g2_fill_1 FILLER_12_662 ();
 sg13g2_fill_1 FILLER_12_673 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_fill_2 FILLER_12_690 ();
 sg13g2_fill_1 FILLER_12_692 ();
 sg13g2_fill_1 FILLER_12_706 ();
 sg13g2_fill_1 FILLER_12_715 ();
 sg13g2_fill_2 FILLER_12_757 ();
 sg13g2_fill_1 FILLER_12_778 ();
 sg13g2_fill_2 FILLER_12_805 ();
 sg13g2_fill_2 FILLER_12_872 ();
 sg13g2_decap_4 FILLER_12_911 ();
 sg13g2_fill_2 FILLER_12_929 ();
 sg13g2_fill_2 FILLER_12_943 ();
 sg13g2_fill_1 FILLER_12_945 ();
 sg13g2_decap_8 FILLER_12_982 ();
 sg13g2_fill_2 FILLER_12_989 ();
 sg13g2_decap_4 FILLER_12_995 ();
 sg13g2_fill_1 FILLER_12_999 ();
 sg13g2_fill_2 FILLER_12_1005 ();
 sg13g2_fill_2 FILLER_12_1012 ();
 sg13g2_fill_2 FILLER_12_1058 ();
 sg13g2_decap_4 FILLER_12_1065 ();
 sg13g2_fill_1 FILLER_12_1082 ();
 sg13g2_decap_4 FILLER_12_1092 ();
 sg13g2_fill_2 FILLER_12_1096 ();
 sg13g2_fill_1 FILLER_12_1142 ();
 sg13g2_fill_1 FILLER_12_1175 ();
 sg13g2_fill_1 FILLER_12_1224 ();
 sg13g2_fill_2 FILLER_12_1239 ();
 sg13g2_decap_8 FILLER_12_1245 ();
 sg13g2_decap_8 FILLER_12_1252 ();
 sg13g2_decap_8 FILLER_12_1259 ();
 sg13g2_decap_8 FILLER_12_1266 ();
 sg13g2_decap_8 FILLER_12_1273 ();
 sg13g2_decap_8 FILLER_12_1280 ();
 sg13g2_decap_8 FILLER_12_1287 ();
 sg13g2_decap_8 FILLER_12_1294 ();
 sg13g2_decap_8 FILLER_12_1301 ();
 sg13g2_decap_8 FILLER_12_1308 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_4 FILLER_13_154 ();
 sg13g2_fill_2 FILLER_13_158 ();
 sg13g2_fill_2 FILLER_13_194 ();
 sg13g2_fill_1 FILLER_13_196 ();
 sg13g2_fill_2 FILLER_13_215 ();
 sg13g2_decap_8 FILLER_13_225 ();
 sg13g2_fill_2 FILLER_13_232 ();
 sg13g2_fill_2 FILLER_13_263 ();
 sg13g2_fill_2 FILLER_13_291 ();
 sg13g2_fill_1 FILLER_13_327 ();
 sg13g2_fill_2 FILLER_13_354 ();
 sg13g2_fill_1 FILLER_13_387 ();
 sg13g2_fill_2 FILLER_13_449 ();
 sg13g2_fill_1 FILLER_13_451 ();
 sg13g2_fill_2 FILLER_13_457 ();
 sg13g2_fill_1 FILLER_13_459 ();
 sg13g2_decap_4 FILLER_13_464 ();
 sg13g2_fill_2 FILLER_13_468 ();
 sg13g2_fill_2 FILLER_13_475 ();
 sg13g2_fill_1 FILLER_13_482 ();
 sg13g2_fill_2 FILLER_13_497 ();
 sg13g2_fill_1 FILLER_13_509 ();
 sg13g2_fill_2 FILLER_13_529 ();
 sg13g2_fill_1 FILLER_13_531 ();
 sg13g2_decap_8 FILLER_13_545 ();
 sg13g2_decap_4 FILLER_13_556 ();
 sg13g2_fill_2 FILLER_13_560 ();
 sg13g2_fill_2 FILLER_13_619 ();
 sg13g2_fill_1 FILLER_13_630 ();
 sg13g2_fill_1 FILLER_13_674 ();
 sg13g2_fill_1 FILLER_13_701 ();
 sg13g2_fill_2 FILLER_13_742 ();
 sg13g2_fill_2 FILLER_13_787 ();
 sg13g2_fill_2 FILLER_13_807 ();
 sg13g2_fill_1 FILLER_13_809 ();
 sg13g2_fill_1 FILLER_13_823 ();
 sg13g2_fill_2 FILLER_13_833 ();
 sg13g2_fill_1 FILLER_13_835 ();
 sg13g2_fill_1 FILLER_13_846 ();
 sg13g2_fill_2 FILLER_13_856 ();
 sg13g2_fill_1 FILLER_13_858 ();
 sg13g2_fill_1 FILLER_13_864 ();
 sg13g2_decap_8 FILLER_13_909 ();
 sg13g2_fill_1 FILLER_13_916 ();
 sg13g2_decap_8 FILLER_13_922 ();
 sg13g2_decap_8 FILLER_13_944 ();
 sg13g2_decap_4 FILLER_13_964 ();
 sg13g2_fill_2 FILLER_13_977 ();
 sg13g2_fill_1 FILLER_13_1010 ();
 sg13g2_fill_2 FILLER_13_1068 ();
 sg13g2_decap_4 FILLER_13_1104 ();
 sg13g2_fill_2 FILLER_13_1108 ();
 sg13g2_fill_2 FILLER_13_1192 ();
 sg13g2_fill_1 FILLER_13_1194 ();
 sg13g2_fill_2 FILLER_13_1217 ();
 sg13g2_fill_1 FILLER_13_1219 ();
 sg13g2_fill_1 FILLER_13_1225 ();
 sg13g2_decap_8 FILLER_13_1235 ();
 sg13g2_decap_8 FILLER_13_1242 ();
 sg13g2_fill_2 FILLER_13_1249 ();
 sg13g2_decap_8 FILLER_13_1254 ();
 sg13g2_decap_8 FILLER_13_1261 ();
 sg13g2_decap_8 FILLER_13_1268 ();
 sg13g2_decap_8 FILLER_13_1275 ();
 sg13g2_decap_8 FILLER_13_1282 ();
 sg13g2_decap_8 FILLER_13_1289 ();
 sg13g2_decap_8 FILLER_13_1296 ();
 sg13g2_decap_8 FILLER_13_1303 ();
 sg13g2_decap_4 FILLER_13_1310 ();
 sg13g2_fill_1 FILLER_13_1314 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_fill_2 FILLER_14_168 ();
 sg13g2_fill_1 FILLER_14_170 ();
 sg13g2_decap_4 FILLER_14_175 ();
 sg13g2_fill_2 FILLER_14_215 ();
 sg13g2_decap_4 FILLER_14_221 ();
 sg13g2_fill_2 FILLER_14_225 ();
 sg13g2_fill_2 FILLER_14_235 ();
 sg13g2_fill_1 FILLER_14_237 ();
 sg13g2_fill_2 FILLER_14_251 ();
 sg13g2_fill_1 FILLER_14_253 ();
 sg13g2_fill_2 FILLER_14_280 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_1 FILLER_14_308 ();
 sg13g2_fill_2 FILLER_14_313 ();
 sg13g2_fill_1 FILLER_14_315 ();
 sg13g2_fill_2 FILLER_14_408 ();
 sg13g2_decap_4 FILLER_14_429 ();
 sg13g2_fill_2 FILLER_14_519 ();
 sg13g2_fill_1 FILLER_14_521 ();
 sg13g2_fill_2 FILLER_14_529 ();
 sg13g2_fill_2 FILLER_14_539 ();
 sg13g2_fill_2 FILLER_14_581 ();
 sg13g2_decap_4 FILLER_14_611 ();
 sg13g2_fill_1 FILLER_14_615 ();
 sg13g2_fill_1 FILLER_14_715 ();
 sg13g2_fill_2 FILLER_14_742 ();
 sg13g2_fill_1 FILLER_14_788 ();
 sg13g2_fill_1 FILLER_14_797 ();
 sg13g2_fill_2 FILLER_14_816 ();
 sg13g2_fill_1 FILLER_14_826 ();
 sg13g2_fill_2 FILLER_14_832 ();
 sg13g2_decap_8 FILLER_14_880 ();
 sg13g2_decap_8 FILLER_14_905 ();
 sg13g2_decap_4 FILLER_14_937 ();
 sg13g2_decap_4 FILLER_14_967 ();
 sg13g2_fill_1 FILLER_14_971 ();
 sg13g2_decap_4 FILLER_14_976 ();
 sg13g2_fill_1 FILLER_14_989 ();
 sg13g2_decap_8 FILLER_14_1000 ();
 sg13g2_decap_4 FILLER_14_1012 ();
 sg13g2_fill_2 FILLER_14_1028 ();
 sg13g2_fill_1 FILLER_14_1030 ();
 sg13g2_fill_2 FILLER_14_1035 ();
 sg13g2_fill_1 FILLER_14_1041 ();
 sg13g2_fill_2 FILLER_14_1055 ();
 sg13g2_fill_1 FILLER_14_1057 ();
 sg13g2_decap_4 FILLER_14_1117 ();
 sg13g2_fill_1 FILLER_14_1121 ();
 sg13g2_decap_4 FILLER_14_1127 ();
 sg13g2_fill_1 FILLER_14_1131 ();
 sg13g2_decap_4 FILLER_14_1136 ();
 sg13g2_fill_2 FILLER_14_1140 ();
 sg13g2_fill_1 FILLER_14_1164 ();
 sg13g2_fill_1 FILLER_14_1251 ();
 sg13g2_decap_8 FILLER_14_1261 ();
 sg13g2_decap_8 FILLER_14_1268 ();
 sg13g2_decap_8 FILLER_14_1275 ();
 sg13g2_decap_8 FILLER_14_1282 ();
 sg13g2_decap_8 FILLER_14_1289 ();
 sg13g2_decap_8 FILLER_14_1296 ();
 sg13g2_decap_8 FILLER_14_1303 ();
 sg13g2_decap_4 FILLER_14_1310 ();
 sg13g2_fill_1 FILLER_14_1314 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_fill_2 FILLER_15_175 ();
 sg13g2_fill_2 FILLER_15_289 ();
 sg13g2_fill_1 FILLER_15_291 ();
 sg13g2_fill_2 FILLER_15_315 ();
 sg13g2_fill_1 FILLER_15_317 ();
 sg13g2_fill_2 FILLER_15_322 ();
 sg13g2_fill_1 FILLER_15_324 ();
 sg13g2_fill_2 FILLER_15_337 ();
 sg13g2_fill_1 FILLER_15_339 ();
 sg13g2_fill_2 FILLER_15_359 ();
 sg13g2_fill_1 FILLER_15_361 ();
 sg13g2_fill_1 FILLER_15_388 ();
 sg13g2_fill_1 FILLER_15_415 ();
 sg13g2_fill_2 FILLER_15_429 ();
 sg13g2_fill_2 FILLER_15_438 ();
 sg13g2_decap_8 FILLER_15_454 ();
 sg13g2_decap_4 FILLER_15_465 ();
 sg13g2_fill_2 FILLER_15_469 ();
 sg13g2_fill_1 FILLER_15_488 ();
 sg13g2_fill_2 FILLER_15_514 ();
 sg13g2_fill_1 FILLER_15_516 ();
 sg13g2_fill_2 FILLER_15_525 ();
 sg13g2_fill_1 FILLER_15_527 ();
 sg13g2_decap_4 FILLER_15_542 ();
 sg13g2_fill_2 FILLER_15_546 ();
 sg13g2_fill_1 FILLER_15_585 ();
 sg13g2_fill_1 FILLER_15_690 ();
 sg13g2_fill_1 FILLER_15_696 ();
 sg13g2_fill_2 FILLER_15_702 ();
 sg13g2_fill_2 FILLER_15_713 ();
 sg13g2_fill_2 FILLER_15_732 ();
 sg13g2_fill_2 FILLER_15_752 ();
 sg13g2_fill_1 FILLER_15_772 ();
 sg13g2_fill_1 FILLER_15_808 ();
 sg13g2_fill_2 FILLER_15_866 ();
 sg13g2_fill_1 FILLER_15_868 ();
 sg13g2_fill_2 FILLER_15_881 ();
 sg13g2_fill_1 FILLER_15_921 ();
 sg13g2_fill_2 FILLER_15_948 ();
 sg13g2_fill_2 FILLER_15_955 ();
 sg13g2_fill_1 FILLER_15_957 ();
 sg13g2_fill_2 FILLER_15_976 ();
 sg13g2_fill_1 FILLER_15_983 ();
 sg13g2_fill_1 FILLER_15_991 ();
 sg13g2_fill_2 FILLER_15_1046 ();
 sg13g2_fill_2 FILLER_15_1074 ();
 sg13g2_fill_2 FILLER_15_1119 ();
 sg13g2_fill_2 FILLER_15_1181 ();
 sg13g2_fill_1 FILLER_15_1183 ();
 sg13g2_fill_2 FILLER_15_1194 ();
 sg13g2_decap_4 FILLER_15_1217 ();
 sg13g2_fill_2 FILLER_15_1221 ();
 sg13g2_decap_8 FILLER_15_1242 ();
 sg13g2_decap_8 FILLER_15_1249 ();
 sg13g2_decap_8 FILLER_15_1256 ();
 sg13g2_decap_8 FILLER_15_1263 ();
 sg13g2_decap_8 FILLER_15_1270 ();
 sg13g2_decap_8 FILLER_15_1277 ();
 sg13g2_decap_8 FILLER_15_1284 ();
 sg13g2_decap_8 FILLER_15_1291 ();
 sg13g2_decap_8 FILLER_15_1298 ();
 sg13g2_decap_8 FILLER_15_1305 ();
 sg13g2_fill_2 FILLER_15_1312 ();
 sg13g2_fill_1 FILLER_15_1314 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_4 FILLER_16_175 ();
 sg13g2_fill_1 FILLER_16_179 ();
 sg13g2_fill_2 FILLER_16_199 ();
 sg13g2_fill_2 FILLER_16_217 ();
 sg13g2_fill_1 FILLER_16_219 ();
 sg13g2_fill_2 FILLER_16_250 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_fill_1 FILLER_16_388 ();
 sg13g2_fill_2 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_451 ();
 sg13g2_decap_8 FILLER_16_547 ();
 sg13g2_decap_4 FILLER_16_554 ();
 sg13g2_fill_1 FILLER_16_558 ();
 sg13g2_fill_2 FILLER_16_572 ();
 sg13g2_fill_1 FILLER_16_583 ();
 sg13g2_fill_2 FILLER_16_617 ();
 sg13g2_fill_2 FILLER_16_633 ();
 sg13g2_fill_1 FILLER_16_635 ();
 sg13g2_fill_1 FILLER_16_640 ();
 sg13g2_decap_8 FILLER_16_645 ();
 sg13g2_fill_2 FILLER_16_652 ();
 sg13g2_fill_1 FILLER_16_657 ();
 sg13g2_fill_1 FILLER_16_731 ();
 sg13g2_fill_1 FILLER_16_736 ();
 sg13g2_fill_1 FILLER_16_820 ();
 sg13g2_decap_8 FILLER_16_871 ();
 sg13g2_decap_4 FILLER_16_878 ();
 sg13g2_fill_2 FILLER_16_882 ();
 sg13g2_fill_1 FILLER_16_901 ();
 sg13g2_fill_1 FILLER_16_934 ();
 sg13g2_fill_2 FILLER_16_943 ();
 sg13g2_fill_1 FILLER_16_945 ();
 sg13g2_fill_2 FILLER_16_977 ();
 sg13g2_fill_1 FILLER_16_983 ();
 sg13g2_fill_1 FILLER_16_1007 ();
 sg13g2_fill_2 FILLER_16_1017 ();
 sg13g2_fill_1 FILLER_16_1028 ();
 sg13g2_fill_1 FILLER_16_1069 ();
 sg13g2_fill_2 FILLER_16_1075 ();
 sg13g2_fill_2 FILLER_16_1086 ();
 sg13g2_fill_1 FILLER_16_1088 ();
 sg13g2_decap_8 FILLER_16_1118 ();
 sg13g2_fill_1 FILLER_16_1130 ();
 sg13g2_fill_1 FILLER_16_1176 ();
 sg13g2_decap_8 FILLER_16_1235 ();
 sg13g2_decap_8 FILLER_16_1242 ();
 sg13g2_decap_8 FILLER_16_1249 ();
 sg13g2_decap_8 FILLER_16_1256 ();
 sg13g2_decap_8 FILLER_16_1263 ();
 sg13g2_decap_8 FILLER_16_1270 ();
 sg13g2_decap_8 FILLER_16_1277 ();
 sg13g2_decap_8 FILLER_16_1284 ();
 sg13g2_decap_8 FILLER_16_1291 ();
 sg13g2_decap_8 FILLER_16_1298 ();
 sg13g2_decap_8 FILLER_16_1305 ();
 sg13g2_fill_2 FILLER_16_1312 ();
 sg13g2_fill_1 FILLER_16_1314 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_175 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_decap_4 FILLER_17_191 ();
 sg13g2_fill_1 FILLER_17_200 ();
 sg13g2_fill_2 FILLER_17_216 ();
 sg13g2_fill_1 FILLER_17_261 ();
 sg13g2_fill_1 FILLER_17_356 ();
 sg13g2_fill_1 FILLER_17_392 ();
 sg13g2_fill_2 FILLER_17_400 ();
 sg13g2_fill_1 FILLER_17_402 ();
 sg13g2_fill_2 FILLER_17_416 ();
 sg13g2_fill_1 FILLER_17_418 ();
 sg13g2_fill_2 FILLER_17_486 ();
 sg13g2_fill_1 FILLER_17_488 ();
 sg13g2_decap_4 FILLER_17_507 ();
 sg13g2_fill_1 FILLER_17_511 ();
 sg13g2_fill_2 FILLER_17_533 ();
 sg13g2_fill_1 FILLER_17_543 ();
 sg13g2_decap_4 FILLER_17_570 ();
 sg13g2_fill_1 FILLER_17_579 ();
 sg13g2_decap_8 FILLER_17_648 ();
 sg13g2_fill_2 FILLER_17_655 ();
 sg13g2_fill_1 FILLER_17_661 ();
 sg13g2_fill_1 FILLER_17_671 ();
 sg13g2_fill_1 FILLER_17_676 ();
 sg13g2_fill_2 FILLER_17_715 ();
 sg13g2_decap_8 FILLER_17_743 ();
 sg13g2_fill_1 FILLER_17_750 ();
 sg13g2_fill_1 FILLER_17_774 ();
 sg13g2_fill_2 FILLER_17_801 ();
 sg13g2_fill_2 FILLER_17_843 ();
 sg13g2_fill_2 FILLER_17_909 ();
 sg13g2_decap_8 FILLER_17_919 ();
 sg13g2_fill_2 FILLER_17_926 ();
 sg13g2_fill_1 FILLER_17_933 ();
 sg13g2_decap_8 FILLER_17_957 ();
 sg13g2_fill_2 FILLER_17_964 ();
 sg13g2_fill_1 FILLER_17_966 ();
 sg13g2_fill_2 FILLER_17_976 ();
 sg13g2_fill_1 FILLER_17_978 ();
 sg13g2_fill_1 FILLER_17_991 ();
 sg13g2_decap_4 FILLER_17_1005 ();
 sg13g2_fill_2 FILLER_17_1040 ();
 sg13g2_fill_1 FILLER_17_1080 ();
 sg13g2_fill_2 FILLER_17_1160 ();
 sg13g2_fill_2 FILLER_17_1188 ();
 sg13g2_fill_1 FILLER_17_1190 ();
 sg13g2_fill_2 FILLER_17_1201 ();
 sg13g2_fill_1 FILLER_17_1203 ();
 sg13g2_decap_4 FILLER_17_1230 ();
 sg13g2_fill_2 FILLER_17_1234 ();
 sg13g2_decap_8 FILLER_17_1240 ();
 sg13g2_decap_8 FILLER_17_1247 ();
 sg13g2_decap_8 FILLER_17_1254 ();
 sg13g2_decap_8 FILLER_17_1261 ();
 sg13g2_decap_8 FILLER_17_1268 ();
 sg13g2_decap_8 FILLER_17_1275 ();
 sg13g2_decap_8 FILLER_17_1282 ();
 sg13g2_decap_8 FILLER_17_1289 ();
 sg13g2_decap_8 FILLER_17_1296 ();
 sg13g2_decap_8 FILLER_17_1303 ();
 sg13g2_decap_4 FILLER_17_1310 ();
 sg13g2_fill_1 FILLER_17_1314 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_4 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_132 ();
 sg13g2_decap_4 FILLER_18_139 ();
 sg13g2_decap_4 FILLER_18_147 ();
 sg13g2_fill_2 FILLER_18_151 ();
 sg13g2_fill_2 FILLER_18_164 ();
 sg13g2_fill_2 FILLER_18_200 ();
 sg13g2_fill_1 FILLER_18_202 ();
 sg13g2_fill_2 FILLER_18_208 ();
 sg13g2_fill_2 FILLER_18_220 ();
 sg13g2_fill_2 FILLER_18_243 ();
 sg13g2_fill_1 FILLER_18_245 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_fill_2 FILLER_18_321 ();
 sg13g2_fill_2 FILLER_18_335 ();
 sg13g2_fill_2 FILLER_18_443 ();
 sg13g2_fill_2 FILLER_18_463 ();
 sg13g2_fill_1 FILLER_18_493 ();
 sg13g2_fill_2 FILLER_18_499 ();
 sg13g2_fill_2 FILLER_18_514 ();
 sg13g2_fill_1 FILLER_18_529 ();
 sg13g2_fill_2 FILLER_18_544 ();
 sg13g2_fill_1 FILLER_18_546 ();
 sg13g2_fill_2 FILLER_18_586 ();
 sg13g2_fill_1 FILLER_18_701 ();
 sg13g2_fill_1 FILLER_18_715 ();
 sg13g2_fill_2 FILLER_18_779 ();
 sg13g2_fill_1 FILLER_18_799 ();
 sg13g2_fill_2 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_853 ();
 sg13g2_decap_8 FILLER_18_860 ();
 sg13g2_fill_2 FILLER_18_872 ();
 sg13g2_fill_2 FILLER_18_884 ();
 sg13g2_fill_1 FILLER_18_886 ();
 sg13g2_decap_8 FILLER_18_905 ();
 sg13g2_fill_2 FILLER_18_912 ();
 sg13g2_fill_1 FILLER_18_914 ();
 sg13g2_decap_4 FILLER_18_920 ();
 sg13g2_decap_4 FILLER_18_942 ();
 sg13g2_fill_2 FILLER_18_946 ();
 sg13g2_fill_2 FILLER_18_1008 ();
 sg13g2_fill_2 FILLER_18_1037 ();
 sg13g2_fill_2 FILLER_18_1095 ();
 sg13g2_fill_1 FILLER_18_1097 ();
 sg13g2_decap_8 FILLER_18_1124 ();
 sg13g2_decap_8 FILLER_18_1131 ();
 sg13g2_fill_1 FILLER_18_1138 ();
 sg13g2_decap_4 FILLER_18_1148 ();
 sg13g2_fill_1 FILLER_18_1152 ();
 sg13g2_fill_2 FILLER_18_1173 ();
 sg13g2_fill_2 FILLER_18_1180 ();
 sg13g2_fill_1 FILLER_18_1182 ();
 sg13g2_fill_1 FILLER_18_1209 ();
 sg13g2_fill_1 FILLER_18_1219 ();
 sg13g2_decap_8 FILLER_18_1251 ();
 sg13g2_decap_8 FILLER_18_1258 ();
 sg13g2_decap_8 FILLER_18_1265 ();
 sg13g2_decap_8 FILLER_18_1272 ();
 sg13g2_decap_8 FILLER_18_1279 ();
 sg13g2_decap_8 FILLER_18_1286 ();
 sg13g2_decap_8 FILLER_18_1293 ();
 sg13g2_decap_8 FILLER_18_1300 ();
 sg13g2_decap_8 FILLER_18_1307 ();
 sg13g2_fill_1 FILLER_18_1314 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_4 FILLER_19_112 ();
 sg13g2_fill_2 FILLER_19_125 ();
 sg13g2_fill_1 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_155 ();
 sg13g2_decap_8 FILLER_19_162 ();
 sg13g2_decap_8 FILLER_19_169 ();
 sg13g2_decap_8 FILLER_19_176 ();
 sg13g2_decap_8 FILLER_19_183 ();
 sg13g2_decap_4 FILLER_19_209 ();
 sg13g2_fill_2 FILLER_19_213 ();
 sg13g2_fill_1 FILLER_19_232 ();
 sg13g2_fill_2 FILLER_19_260 ();
 sg13g2_fill_2 FILLER_19_272 ();
 sg13g2_fill_1 FILLER_19_274 ();
 sg13g2_fill_2 FILLER_19_301 ();
 sg13g2_fill_2 FILLER_19_368 ();
 sg13g2_fill_2 FILLER_19_396 ();
 sg13g2_fill_2 FILLER_19_422 ();
 sg13g2_fill_1 FILLER_19_424 ();
 sg13g2_fill_2 FILLER_19_468 ();
 sg13g2_fill_2 FILLER_19_541 ();
 sg13g2_fill_1 FILLER_19_543 ();
 sg13g2_fill_1 FILLER_19_580 ();
 sg13g2_decap_8 FILLER_19_646 ();
 sg13g2_fill_2 FILLER_19_670 ();
 sg13g2_fill_1 FILLER_19_672 ();
 sg13g2_fill_2 FILLER_19_710 ();
 sg13g2_decap_8 FILLER_19_743 ();
 sg13g2_fill_1 FILLER_19_750 ();
 sg13g2_decap_4 FILLER_19_774 ();
 sg13g2_fill_2 FILLER_19_778 ();
 sg13g2_fill_2 FILLER_19_811 ();
 sg13g2_decap_4 FILLER_19_856 ();
 sg13g2_fill_2 FILLER_19_878 ();
 sg13g2_fill_1 FILLER_19_880 ();
 sg13g2_fill_2 FILLER_19_897 ();
 sg13g2_fill_2 FILLER_19_914 ();
 sg13g2_fill_1 FILLER_19_916 ();
 sg13g2_fill_1 FILLER_19_935 ();
 sg13g2_decap_8 FILLER_19_967 ();
 sg13g2_decap_4 FILLER_19_974 ();
 sg13g2_fill_1 FILLER_19_978 ();
 sg13g2_fill_2 FILLER_19_986 ();
 sg13g2_fill_1 FILLER_19_988 ();
 sg13g2_decap_8 FILLER_19_993 ();
 sg13g2_fill_2 FILLER_19_1000 ();
 sg13g2_fill_2 FILLER_19_1077 ();
 sg13g2_fill_1 FILLER_19_1097 ();
 sg13g2_decap_8 FILLER_19_1133 ();
 sg13g2_fill_2 FILLER_19_1163 ();
 sg13g2_fill_2 FILLER_19_1188 ();
 sg13g2_fill_1 FILLER_19_1190 ();
 sg13g2_decap_8 FILLER_19_1257 ();
 sg13g2_decap_8 FILLER_19_1264 ();
 sg13g2_decap_8 FILLER_19_1271 ();
 sg13g2_decap_8 FILLER_19_1278 ();
 sg13g2_decap_8 FILLER_19_1285 ();
 sg13g2_decap_8 FILLER_19_1292 ();
 sg13g2_decap_8 FILLER_19_1299 ();
 sg13g2_decap_8 FILLER_19_1306 ();
 sg13g2_fill_2 FILLER_19_1313 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_4 FILLER_20_98 ();
 sg13g2_fill_1 FILLER_20_128 ();
 sg13g2_decap_8 FILLER_20_164 ();
 sg13g2_decap_4 FILLER_20_171 ();
 sg13g2_fill_1 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_fill_2 FILLER_20_205 ();
 sg13g2_fill_1 FILLER_20_212 ();
 sg13g2_fill_1 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_264 ();
 sg13g2_fill_2 FILLER_20_274 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_fill_2 FILLER_20_317 ();
 sg13g2_fill_1 FILLER_20_319 ();
 sg13g2_fill_2 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_428 ();
 sg13g2_fill_1 FILLER_20_435 ();
 sg13g2_fill_1 FILLER_20_450 ();
 sg13g2_fill_1 FILLER_20_460 ();
 sg13g2_fill_2 FILLER_20_466 ();
 sg13g2_fill_2 FILLER_20_473 ();
 sg13g2_fill_1 FILLER_20_518 ();
 sg13g2_fill_2 FILLER_20_528 ();
 sg13g2_fill_1 FILLER_20_530 ();
 sg13g2_fill_1 FILLER_20_535 ();
 sg13g2_fill_1 FILLER_20_540 ();
 sg13g2_fill_2 FILLER_20_572 ();
 sg13g2_fill_2 FILLER_20_588 ();
 sg13g2_decap_4 FILLER_20_598 ();
 sg13g2_decap_4 FILLER_20_606 ();
 sg13g2_fill_1 FILLER_20_610 ();
 sg13g2_decap_4 FILLER_20_677 ();
 sg13g2_fill_2 FILLER_20_681 ();
 sg13g2_fill_1 FILLER_20_687 ();
 sg13g2_fill_2 FILLER_20_697 ();
 sg13g2_fill_2 FILLER_20_839 ();
 sg13g2_fill_1 FILLER_20_841 ();
 sg13g2_decap_4 FILLER_20_876 ();
 sg13g2_fill_1 FILLER_20_880 ();
 sg13g2_fill_1 FILLER_20_886 ();
 sg13g2_decap_8 FILLER_20_908 ();
 sg13g2_decap_4 FILLER_20_915 ();
 sg13g2_fill_2 FILLER_20_919 ();
 sg13g2_decap_4 FILLER_20_926 ();
 sg13g2_fill_1 FILLER_20_930 ();
 sg13g2_fill_1 FILLER_20_941 ();
 sg13g2_decap_4 FILLER_20_968 ();
 sg13g2_decap_8 FILLER_20_976 ();
 sg13g2_decap_8 FILLER_20_983 ();
 sg13g2_fill_1 FILLER_20_993 ();
 sg13g2_decap_4 FILLER_20_999 ();
 sg13g2_fill_2 FILLER_20_1023 ();
 sg13g2_fill_1 FILLER_20_1025 ();
 sg13g2_decap_4 FILLER_20_1035 ();
 sg13g2_fill_1 FILLER_20_1057 ();
 sg13g2_fill_1 FILLER_20_1063 ();
 sg13g2_fill_1 FILLER_20_1077 ();
 sg13g2_fill_2 FILLER_20_1110 ();
 sg13g2_fill_1 FILLER_20_1207 ();
 sg13g2_decap_8 FILLER_20_1256 ();
 sg13g2_decap_8 FILLER_20_1263 ();
 sg13g2_decap_8 FILLER_20_1270 ();
 sg13g2_decap_8 FILLER_20_1277 ();
 sg13g2_decap_8 FILLER_20_1284 ();
 sg13g2_decap_8 FILLER_20_1291 ();
 sg13g2_decap_8 FILLER_20_1298 ();
 sg13g2_decap_8 FILLER_20_1305 ();
 sg13g2_fill_2 FILLER_20_1312 ();
 sg13g2_fill_1 FILLER_20_1314 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_fill_2 FILLER_21_164 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_decap_8 FILLER_21_225 ();
 sg13g2_decap_4 FILLER_21_232 ();
 sg13g2_fill_1 FILLER_21_273 ();
 sg13g2_fill_1 FILLER_21_300 ();
 sg13g2_fill_2 FILLER_21_390 ();
 sg13g2_fill_1 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_419 ();
 sg13g2_fill_1 FILLER_21_451 ();
 sg13g2_fill_1 FILLER_21_492 ();
 sg13g2_fill_2 FILLER_21_502 ();
 sg13g2_fill_2 FILLER_21_549 ();
 sg13g2_decap_4 FILLER_21_603 ();
 sg13g2_fill_2 FILLER_21_607 ();
 sg13g2_fill_1 FILLER_21_613 ();
 sg13g2_decap_4 FILLER_21_640 ();
 sg13g2_fill_2 FILLER_21_644 ();
 sg13g2_fill_2 FILLER_21_650 ();
 sg13g2_fill_1 FILLER_21_652 ();
 sg13g2_decap_4 FILLER_21_657 ();
 sg13g2_fill_2 FILLER_21_661 ();
 sg13g2_fill_2 FILLER_21_711 ();
 sg13g2_fill_1 FILLER_21_713 ();
 sg13g2_fill_2 FILLER_21_719 ();
 sg13g2_fill_2 FILLER_21_731 ();
 sg13g2_fill_1 FILLER_21_733 ();
 sg13g2_fill_2 FILLER_21_751 ();
 sg13g2_decap_8 FILLER_21_776 ();
 sg13g2_decap_4 FILLER_21_783 ();
 sg13g2_fill_2 FILLER_21_808 ();
 sg13g2_decap_8 FILLER_21_855 ();
 sg13g2_decap_8 FILLER_21_866 ();
 sg13g2_fill_2 FILLER_21_878 ();
 sg13g2_decap_8 FILLER_21_885 ();
 sg13g2_fill_2 FILLER_21_892 ();
 sg13g2_fill_2 FILLER_21_904 ();
 sg13g2_decap_4 FILLER_21_932 ();
 sg13g2_fill_2 FILLER_21_936 ();
 sg13g2_fill_2 FILLER_21_954 ();
 sg13g2_fill_1 FILLER_21_987 ();
 sg13g2_fill_2 FILLER_21_1009 ();
 sg13g2_fill_1 FILLER_21_1011 ();
 sg13g2_fill_2 FILLER_21_1097 ();
 sg13g2_fill_2 FILLER_21_1115 ();
 sg13g2_decap_8 FILLER_21_1122 ();
 sg13g2_fill_1 FILLER_21_1129 ();
 sg13g2_fill_1 FILLER_21_1134 ();
 sg13g2_decap_4 FILLER_21_1139 ();
 sg13g2_fill_2 FILLER_21_1143 ();
 sg13g2_fill_2 FILLER_21_1169 ();
 sg13g2_fill_1 FILLER_21_1184 ();
 sg13g2_fill_1 FILLER_21_1190 ();
 sg13g2_fill_2 FILLER_21_1226 ();
 sg13g2_decap_8 FILLER_21_1257 ();
 sg13g2_decap_8 FILLER_21_1264 ();
 sg13g2_decap_8 FILLER_21_1271 ();
 sg13g2_decap_8 FILLER_21_1278 ();
 sg13g2_decap_8 FILLER_21_1285 ();
 sg13g2_decap_8 FILLER_21_1292 ();
 sg13g2_decap_8 FILLER_21_1299 ();
 sg13g2_decap_8 FILLER_21_1306 ();
 sg13g2_fill_2 FILLER_21_1313 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_fill_1 FILLER_22_131 ();
 sg13g2_decap_4 FILLER_22_172 ();
 sg13g2_fill_2 FILLER_22_176 ();
 sg13g2_fill_2 FILLER_22_182 ();
 sg13g2_fill_1 FILLER_22_184 ();
 sg13g2_decap_8 FILLER_22_199 ();
 sg13g2_decap_4 FILLER_22_206 ();
 sg13g2_decap_4 FILLER_22_232 ();
 sg13g2_fill_1 FILLER_22_236 ();
 sg13g2_decap_4 FILLER_22_241 ();
 sg13g2_fill_1 FILLER_22_257 ();
 sg13g2_fill_1 FILLER_22_273 ();
 sg13g2_fill_2 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_302 ();
 sg13g2_fill_2 FILLER_22_321 ();
 sg13g2_fill_1 FILLER_22_323 ();
 sg13g2_fill_2 FILLER_22_337 ();
 sg13g2_fill_1 FILLER_22_344 ();
 sg13g2_fill_1 FILLER_22_354 ();
 sg13g2_fill_2 FILLER_22_368 ();
 sg13g2_fill_1 FILLER_22_401 ();
 sg13g2_fill_2 FILLER_22_415 ();
 sg13g2_decap_4 FILLER_22_427 ();
 sg13g2_fill_2 FILLER_22_431 ();
 sg13g2_decap_4 FILLER_22_437 ();
 sg13g2_fill_2 FILLER_22_441 ();
 sg13g2_fill_2 FILLER_22_454 ();
 sg13g2_fill_2 FILLER_22_544 ();
 sg13g2_fill_2 FILLER_22_551 ();
 sg13g2_fill_1 FILLER_22_568 ();
 sg13g2_fill_1 FILLER_22_597 ();
 sg13g2_fill_1 FILLER_22_624 ();
 sg13g2_fill_1 FILLER_22_629 ();
 sg13g2_fill_1 FILLER_22_733 ();
 sg13g2_fill_1 FILLER_22_747 ();
 sg13g2_fill_2 FILLER_22_826 ();
 sg13g2_fill_1 FILLER_22_828 ();
 sg13g2_fill_1 FILLER_22_844 ();
 sg13g2_fill_2 FILLER_22_850 ();
 sg13g2_decap_8 FILLER_22_923 ();
 sg13g2_decap_4 FILLER_22_930 ();
 sg13g2_fill_2 FILLER_22_934 ();
 sg13g2_fill_2 FILLER_22_955 ();
 sg13g2_fill_1 FILLER_22_957 ();
 sg13g2_fill_2 FILLER_22_968 ();
 sg13g2_fill_1 FILLER_22_970 ();
 sg13g2_fill_2 FILLER_22_1009 ();
 sg13g2_fill_1 FILLER_22_1011 ();
 sg13g2_fill_1 FILLER_22_1021 ();
 sg13g2_fill_2 FILLER_22_1036 ();
 sg13g2_fill_1 FILLER_22_1038 ();
 sg13g2_fill_1 FILLER_22_1061 ();
 sg13g2_fill_2 FILLER_22_1103 ();
 sg13g2_fill_1 FILLER_22_1105 ();
 sg13g2_fill_2 FILLER_22_1111 ();
 sg13g2_fill_1 FILLER_22_1113 ();
 sg13g2_fill_2 FILLER_22_1145 ();
 sg13g2_fill_2 FILLER_22_1160 ();
 sg13g2_decap_8 FILLER_22_1238 ();
 sg13g2_decap_8 FILLER_22_1245 ();
 sg13g2_decap_8 FILLER_22_1252 ();
 sg13g2_decap_8 FILLER_22_1259 ();
 sg13g2_decap_8 FILLER_22_1266 ();
 sg13g2_decap_8 FILLER_22_1273 ();
 sg13g2_decap_8 FILLER_22_1280 ();
 sg13g2_decap_8 FILLER_22_1287 ();
 sg13g2_decap_8 FILLER_22_1294 ();
 sg13g2_decap_8 FILLER_22_1301 ();
 sg13g2_decap_8 FILLER_22_1308 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_4 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_125 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_fill_2 FILLER_23_210 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_fill_1 FILLER_23_319 ();
 sg13g2_fill_2 FILLER_23_346 ();
 sg13g2_fill_2 FILLER_23_374 ();
 sg13g2_fill_1 FILLER_23_393 ();
 sg13g2_fill_2 FILLER_23_415 ();
 sg13g2_decap_4 FILLER_23_519 ();
 sg13g2_fill_1 FILLER_23_523 ();
 sg13g2_fill_1 FILLER_23_528 ();
 sg13g2_fill_2 FILLER_23_577 ();
 sg13g2_decap_4 FILLER_23_597 ();
 sg13g2_fill_2 FILLER_23_615 ();
 sg13g2_fill_1 FILLER_23_617 ();
 sg13g2_fill_1 FILLER_23_641 ();
 sg13g2_decap_8 FILLER_23_664 ();
 sg13g2_decap_4 FILLER_23_671 ();
 sg13g2_fill_1 FILLER_23_675 ();
 sg13g2_decap_4 FILLER_23_680 ();
 sg13g2_decap_4 FILLER_23_700 ();
 sg13g2_fill_2 FILLER_23_704 ();
 sg13g2_decap_8 FILLER_23_711 ();
 sg13g2_fill_1 FILLER_23_735 ();
 sg13g2_fill_1 FILLER_23_750 ();
 sg13g2_fill_2 FILLER_23_769 ();
 sg13g2_fill_1 FILLER_23_771 ();
 sg13g2_fill_2 FILLER_23_781 ();
 sg13g2_fill_1 FILLER_23_783 ();
 sg13g2_decap_8 FILLER_23_788 ();
 sg13g2_decap_4 FILLER_23_795 ();
 sg13g2_fill_1 FILLER_23_827 ();
 sg13g2_fill_2 FILLER_23_838 ();
 sg13g2_decap_8 FILLER_23_866 ();
 sg13g2_fill_1 FILLER_23_873 ();
 sg13g2_decap_4 FILLER_23_891 ();
 sg13g2_decap_4 FILLER_23_908 ();
 sg13g2_fill_2 FILLER_23_985 ();
 sg13g2_fill_1 FILLER_23_1041 ();
 sg13g2_fill_2 FILLER_23_1102 ();
 sg13g2_decap_4 FILLER_23_1130 ();
 sg13g2_fill_1 FILLER_23_1134 ();
 sg13g2_fill_2 FILLER_23_1170 ();
 sg13g2_fill_2 FILLER_23_1189 ();
 sg13g2_decap_8 FILLER_23_1240 ();
 sg13g2_decap_8 FILLER_23_1247 ();
 sg13g2_decap_8 FILLER_23_1254 ();
 sg13g2_decap_8 FILLER_23_1261 ();
 sg13g2_decap_8 FILLER_23_1268 ();
 sg13g2_decap_8 FILLER_23_1275 ();
 sg13g2_decap_8 FILLER_23_1282 ();
 sg13g2_decap_8 FILLER_23_1289 ();
 sg13g2_decap_8 FILLER_23_1296 ();
 sg13g2_decap_8 FILLER_23_1303 ();
 sg13g2_decap_4 FILLER_23_1310 ();
 sg13g2_fill_1 FILLER_23_1314 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_4 FILLER_24_98 ();
 sg13g2_fill_2 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_139 ();
 sg13g2_decap_4 FILLER_24_180 ();
 sg13g2_fill_1 FILLER_24_193 ();
 sg13g2_fill_2 FILLER_24_206 ();
 sg13g2_fill_1 FILLER_24_233 ();
 sg13g2_decap_4 FILLER_24_243 ();
 sg13g2_fill_2 FILLER_24_247 ();
 sg13g2_fill_2 FILLER_24_267 ();
 sg13g2_fill_2 FILLER_24_317 ();
 sg13g2_fill_1 FILLER_24_319 ();
 sg13g2_fill_1 FILLER_24_398 ();
 sg13g2_fill_1 FILLER_24_435 ();
 sg13g2_fill_1 FILLER_24_464 ();
 sg13g2_fill_1 FILLER_24_475 ();
 sg13g2_fill_2 FILLER_24_494 ();
 sg13g2_fill_2 FILLER_24_527 ();
 sg13g2_fill_2 FILLER_24_551 ();
 sg13g2_fill_1 FILLER_24_559 ();
 sg13g2_fill_1 FILLER_24_586 ();
 sg13g2_fill_1 FILLER_24_596 ();
 sg13g2_fill_2 FILLER_24_610 ();
 sg13g2_fill_1 FILLER_24_612 ();
 sg13g2_fill_2 FILLER_24_625 ();
 sg13g2_fill_1 FILLER_24_627 ();
 sg13g2_fill_2 FILLER_24_669 ();
 sg13g2_fill_1 FILLER_24_671 ();
 sg13g2_fill_1 FILLER_24_687 ();
 sg13g2_fill_1 FILLER_24_702 ();
 sg13g2_fill_2 FILLER_24_733 ();
 sg13g2_fill_2 FILLER_24_741 ();
 sg13g2_fill_1 FILLER_24_756 ();
 sg13g2_fill_1 FILLER_24_793 ();
 sg13g2_fill_2 FILLER_24_799 ();
 sg13g2_fill_2 FILLER_24_826 ();
 sg13g2_fill_2 FILLER_24_850 ();
 sg13g2_fill_1 FILLER_24_881 ();
 sg13g2_fill_2 FILLER_24_909 ();
 sg13g2_fill_1 FILLER_24_916 ();
 sg13g2_decap_8 FILLER_24_930 ();
 sg13g2_fill_2 FILLER_24_937 ();
 sg13g2_fill_1 FILLER_24_949 ();
 sg13g2_decap_4 FILLER_24_954 ();
 sg13g2_fill_2 FILLER_24_958 ();
 sg13g2_decap_8 FILLER_24_970 ();
 sg13g2_decap_8 FILLER_24_977 ();
 sg13g2_decap_4 FILLER_24_984 ();
 sg13g2_fill_2 FILLER_24_988 ();
 sg13g2_fill_2 FILLER_24_1009 ();
 sg13g2_decap_8 FILLER_24_1016 ();
 sg13g2_fill_2 FILLER_24_1023 ();
 sg13g2_fill_1 FILLER_24_1025 ();
 sg13g2_fill_2 FILLER_24_1034 ();
 sg13g2_fill_2 FILLER_24_1073 ();
 sg13g2_fill_1 FILLER_24_1075 ();
 sg13g2_fill_1 FILLER_24_1080 ();
 sg13g2_decap_4 FILLER_24_1102 ();
 sg13g2_decap_8 FILLER_24_1119 ();
 sg13g2_fill_1 FILLER_24_1126 ();
 sg13g2_fill_1 FILLER_24_1191 ();
 sg13g2_fill_1 FILLER_24_1201 ();
 sg13g2_fill_1 FILLER_24_1206 ();
 sg13g2_fill_2 FILLER_24_1212 ();
 sg13g2_decap_8 FILLER_24_1255 ();
 sg13g2_decap_8 FILLER_24_1262 ();
 sg13g2_decap_8 FILLER_24_1269 ();
 sg13g2_decap_8 FILLER_24_1276 ();
 sg13g2_decap_8 FILLER_24_1283 ();
 sg13g2_decap_8 FILLER_24_1290 ();
 sg13g2_decap_8 FILLER_24_1297 ();
 sg13g2_decap_8 FILLER_24_1304 ();
 sg13g2_decap_4 FILLER_24_1311 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_fill_2 FILLER_25_124 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_fill_1 FILLER_25_173 ();
 sg13g2_decap_4 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_183 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_fill_2 FILLER_25_310 ();
 sg13g2_fill_1 FILLER_25_399 ();
 sg13g2_fill_1 FILLER_25_413 ();
 sg13g2_fill_1 FILLER_25_478 ();
 sg13g2_fill_2 FILLER_25_495 ();
 sg13g2_fill_1 FILLER_25_497 ();
 sg13g2_fill_2 FILLER_25_503 ();
 sg13g2_fill_1 FILLER_25_529 ();
 sg13g2_fill_1 FILLER_25_562 ();
 sg13g2_decap_4 FILLER_25_566 ();
 sg13g2_fill_1 FILLER_25_582 ();
 sg13g2_fill_2 FILLER_25_614 ();
 sg13g2_fill_1 FILLER_25_616 ();
 sg13g2_fill_1 FILLER_25_623 ();
 sg13g2_decap_8 FILLER_25_643 ();
 sg13g2_decap_4 FILLER_25_650 ();
 sg13g2_decap_8 FILLER_25_658 ();
 sg13g2_decap_8 FILLER_25_668 ();
 sg13g2_fill_2 FILLER_25_675 ();
 sg13g2_fill_2 FILLER_25_682 ();
 sg13g2_fill_2 FILLER_25_691 ();
 sg13g2_fill_1 FILLER_25_706 ();
 sg13g2_fill_2 FILLER_25_727 ();
 sg13g2_fill_1 FILLER_25_729 ();
 sg13g2_fill_1 FILLER_25_789 ();
 sg13g2_fill_2 FILLER_25_830 ();
 sg13g2_fill_1 FILLER_25_832 ();
 sg13g2_decap_8 FILLER_25_868 ();
 sg13g2_fill_2 FILLER_25_899 ();
 sg13g2_decap_4 FILLER_25_924 ();
 sg13g2_fill_2 FILLER_25_936 ();
 sg13g2_fill_2 FILLER_25_948 ();
 sg13g2_fill_2 FILLER_25_958 ();
 sg13g2_fill_1 FILLER_25_960 ();
 sg13g2_fill_1 FILLER_25_987 ();
 sg13g2_fill_2 FILLER_25_1031 ();
 sg13g2_fill_2 FILLER_25_1090 ();
 sg13g2_fill_1 FILLER_25_1092 ();
 sg13g2_decap_4 FILLER_25_1116 ();
 sg13g2_fill_2 FILLER_25_1120 ();
 sg13g2_decap_8 FILLER_25_1127 ();
 sg13g2_decap_8 FILLER_25_1134 ();
 sg13g2_fill_2 FILLER_25_1150 ();
 sg13g2_fill_1 FILLER_25_1152 ();
 sg13g2_decap_8 FILLER_25_1196 ();
 sg13g2_fill_1 FILLER_25_1223 ();
 sg13g2_decap_8 FILLER_25_1249 ();
 sg13g2_decap_8 FILLER_25_1256 ();
 sg13g2_decap_8 FILLER_25_1263 ();
 sg13g2_decap_8 FILLER_25_1270 ();
 sg13g2_decap_8 FILLER_25_1277 ();
 sg13g2_decap_8 FILLER_25_1284 ();
 sg13g2_decap_8 FILLER_25_1291 ();
 sg13g2_decap_8 FILLER_25_1298 ();
 sg13g2_decap_8 FILLER_25_1305 ();
 sg13g2_fill_2 FILLER_25_1312 ();
 sg13g2_fill_1 FILLER_25_1314 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_fill_2 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_126 ();
 sg13g2_fill_2 FILLER_26_146 ();
 sg13g2_fill_1 FILLER_26_152 ();
 sg13g2_fill_2 FILLER_26_161 ();
 sg13g2_fill_2 FILLER_26_202 ();
 sg13g2_fill_1 FILLER_26_227 ();
 sg13g2_fill_2 FILLER_26_246 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_fill_2 FILLER_26_412 ();
 sg13g2_fill_2 FILLER_26_466 ();
 sg13g2_fill_1 FILLER_26_481 ();
 sg13g2_decap_8 FILLER_26_490 ();
 sg13g2_fill_2 FILLER_26_497 ();
 sg13g2_fill_1 FILLER_26_525 ();
 sg13g2_decap_4 FILLER_26_564 ();
 sg13g2_fill_1 FILLER_26_568 ();
 sg13g2_fill_2 FILLER_26_573 ();
 sg13g2_fill_2 FILLER_26_596 ();
 sg13g2_fill_2 FILLER_26_611 ();
 sg13g2_fill_1 FILLER_26_621 ();
 sg13g2_fill_2 FILLER_26_627 ();
 sg13g2_decap_4 FILLER_26_637 ();
 sg13g2_fill_2 FILLER_26_641 ();
 sg13g2_fill_1 FILLER_26_681 ();
 sg13g2_decap_4 FILLER_26_714 ();
 sg13g2_fill_2 FILLER_26_728 ();
 sg13g2_fill_1 FILLER_26_730 ();
 sg13g2_fill_1 FILLER_26_756 ();
 sg13g2_decap_8 FILLER_26_761 ();
 sg13g2_fill_2 FILLER_26_768 ();
 sg13g2_fill_1 FILLER_26_796 ();
 sg13g2_decap_4 FILLER_26_806 ();
 sg13g2_fill_1 FILLER_26_845 ();
 sg13g2_fill_2 FILLER_26_856 ();
 sg13g2_fill_1 FILLER_26_884 ();
 sg13g2_decap_8 FILLER_26_890 ();
 sg13g2_decap_8 FILLER_26_897 ();
 sg13g2_fill_2 FILLER_26_904 ();
 sg13g2_fill_1 FILLER_26_906 ();
 sg13g2_fill_2 FILLER_26_915 ();
 sg13g2_decap_4 FILLER_26_922 ();
 sg13g2_fill_2 FILLER_26_935 ();
 sg13g2_fill_1 FILLER_26_937 ();
 sg13g2_fill_2 FILLER_26_958 ();
 sg13g2_fill_1 FILLER_26_960 ();
 sg13g2_fill_2 FILLER_26_999 ();
 sg13g2_fill_1 FILLER_26_1014 ();
 sg13g2_fill_2 FILLER_26_1041 ();
 sg13g2_fill_1 FILLER_26_1043 ();
 sg13g2_fill_2 FILLER_26_1053 ();
 sg13g2_fill_2 FILLER_26_1064 ();
 sg13g2_fill_1 FILLER_26_1095 ();
 sg13g2_fill_1 FILLER_26_1119 ();
 sg13g2_fill_2 FILLER_26_1181 ();
 sg13g2_fill_1 FILLER_26_1191 ();
 sg13g2_fill_1 FILLER_26_1218 ();
 sg13g2_decap_8 FILLER_26_1245 ();
 sg13g2_decap_8 FILLER_26_1252 ();
 sg13g2_decap_8 FILLER_26_1259 ();
 sg13g2_decap_8 FILLER_26_1266 ();
 sg13g2_decap_8 FILLER_26_1273 ();
 sg13g2_decap_8 FILLER_26_1280 ();
 sg13g2_decap_8 FILLER_26_1287 ();
 sg13g2_decap_8 FILLER_26_1294 ();
 sg13g2_decap_8 FILLER_26_1301 ();
 sg13g2_decap_8 FILLER_26_1308 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_4 FILLER_27_98 ();
 sg13g2_fill_2 FILLER_27_102 ();
 sg13g2_fill_2 FILLER_27_118 ();
 sg13g2_fill_1 FILLER_27_125 ();
 sg13g2_fill_1 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_163 ();
 sg13g2_fill_2 FILLER_27_194 ();
 sg13g2_fill_2 FILLER_27_249 ();
 sg13g2_fill_1 FILLER_27_251 ();
 sg13g2_fill_1 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_289 ();
 sg13g2_fill_2 FILLER_27_333 ();
 sg13g2_fill_2 FILLER_27_416 ();
 sg13g2_fill_1 FILLER_27_418 ();
 sg13g2_fill_2 FILLER_27_445 ();
 sg13g2_fill_2 FILLER_27_478 ();
 sg13g2_fill_1 FILLER_27_524 ();
 sg13g2_decap_4 FILLER_27_554 ();
 sg13g2_fill_1 FILLER_27_558 ();
 sg13g2_fill_1 FILLER_27_585 ();
 sg13g2_fill_1 FILLER_27_595 ();
 sg13g2_fill_2 FILLER_27_609 ();
 sg13g2_fill_1 FILLER_27_611 ();
 sg13g2_fill_2 FILLER_27_621 ();
 sg13g2_fill_1 FILLER_27_623 ();
 sg13g2_fill_1 FILLER_27_628 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_4 FILLER_27_657 ();
 sg13g2_fill_1 FILLER_27_661 ();
 sg13g2_fill_2 FILLER_27_669 ();
 sg13g2_fill_2 FILLER_27_720 ();
 sg13g2_decap_8 FILLER_27_748 ();
 sg13g2_decap_4 FILLER_27_755 ();
 sg13g2_decap_8 FILLER_27_767 ();
 sg13g2_decap_8 FILLER_27_774 ();
 sg13g2_decap_4 FILLER_27_781 ();
 sg13g2_fill_2 FILLER_27_785 ();
 sg13g2_fill_1 FILLER_27_846 ();
 sg13g2_fill_2 FILLER_27_872 ();
 sg13g2_decap_8 FILLER_27_893 ();
 sg13g2_fill_2 FILLER_27_900 ();
 sg13g2_fill_1 FILLER_27_902 ();
 sg13g2_fill_1 FILLER_27_908 ();
 sg13g2_fill_2 FILLER_27_935 ();
 sg13g2_fill_1 FILLER_27_937 ();
 sg13g2_fill_1 FILLER_27_946 ();
 sg13g2_decap_4 FILLER_27_955 ();
 sg13g2_decap_4 FILLER_27_985 ();
 sg13g2_fill_2 FILLER_27_1034 ();
 sg13g2_fill_1 FILLER_27_1036 ();
 sg13g2_fill_1 FILLER_27_1097 ();
 sg13g2_fill_2 FILLER_27_1122 ();
 sg13g2_fill_1 FILLER_27_1124 ();
 sg13g2_fill_1 FILLER_27_1130 ();
 sg13g2_fill_2 FILLER_27_1135 ();
 sg13g2_decap_4 FILLER_27_1146 ();
 sg13g2_fill_2 FILLER_27_1150 ();
 sg13g2_fill_2 FILLER_27_1156 ();
 sg13g2_decap_8 FILLER_27_1200 ();
 sg13g2_decap_8 FILLER_27_1207 ();
 sg13g2_fill_1 FILLER_27_1214 ();
 sg13g2_fill_1 FILLER_27_1229 ();
 sg13g2_decap_8 FILLER_27_1234 ();
 sg13g2_decap_8 FILLER_27_1241 ();
 sg13g2_decap_8 FILLER_27_1248 ();
 sg13g2_decap_8 FILLER_27_1255 ();
 sg13g2_decap_8 FILLER_27_1262 ();
 sg13g2_decap_8 FILLER_27_1269 ();
 sg13g2_decap_8 FILLER_27_1276 ();
 sg13g2_decap_8 FILLER_27_1283 ();
 sg13g2_decap_8 FILLER_27_1290 ();
 sg13g2_decap_8 FILLER_27_1297 ();
 sg13g2_decap_8 FILLER_27_1304 ();
 sg13g2_decap_4 FILLER_27_1311 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_137 ();
 sg13g2_fill_2 FILLER_28_181 ();
 sg13g2_fill_2 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_194 ();
 sg13g2_fill_2 FILLER_28_200 ();
 sg13g2_fill_2 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_216 ();
 sg13g2_fill_2 FILLER_28_303 ();
 sg13g2_fill_2 FILLER_28_319 ();
 sg13g2_fill_1 FILLER_28_365 ();
 sg13g2_fill_2 FILLER_28_389 ();
 sg13g2_fill_1 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_430 ();
 sg13g2_fill_2 FILLER_28_468 ();
 sg13g2_fill_2 FILLER_28_488 ();
 sg13g2_fill_2 FILLER_28_495 ();
 sg13g2_fill_1 FILLER_28_497 ();
 sg13g2_fill_1 FILLER_28_508 ();
 sg13g2_decap_4 FILLER_28_513 ();
 sg13g2_fill_2 FILLER_28_517 ();
 sg13g2_decap_8 FILLER_28_565 ();
 sg13g2_fill_2 FILLER_28_572 ();
 sg13g2_fill_1 FILLER_28_592 ();
 sg13g2_fill_1 FILLER_28_603 ();
 sg13g2_fill_1 FILLER_28_627 ();
 sg13g2_fill_2 FILLER_28_664 ();
 sg13g2_fill_1 FILLER_28_666 ();
 sg13g2_fill_1 FILLER_28_682 ();
 sg13g2_fill_1 FILLER_28_687 ();
 sg13g2_fill_2 FILLER_28_718 ();
 sg13g2_fill_1 FILLER_28_729 ();
 sg13g2_fill_2 FILLER_28_739 ();
 sg13g2_fill_1 FILLER_28_741 ();
 sg13g2_fill_1 FILLER_28_818 ();
 sg13g2_fill_1 FILLER_28_845 ();
 sg13g2_fill_1 FILLER_28_882 ();
 sg13g2_decap_4 FILLER_28_914 ();
 sg13g2_fill_1 FILLER_28_918 ();
 sg13g2_fill_2 FILLER_28_937 ();
 sg13g2_fill_1 FILLER_28_939 ();
 sg13g2_decap_4 FILLER_28_953 ();
 sg13g2_fill_1 FILLER_28_957 ();
 sg13g2_fill_1 FILLER_28_1081 ();
 sg13g2_fill_1 FILLER_28_1115 ();
 sg13g2_decap_4 FILLER_28_1147 ();
 sg13g2_fill_1 FILLER_28_1151 ();
 sg13g2_decap_8 FILLER_28_1193 ();
 sg13g2_decap_8 FILLER_28_1200 ();
 sg13g2_decap_8 FILLER_28_1207 ();
 sg13g2_decap_8 FILLER_28_1214 ();
 sg13g2_decap_8 FILLER_28_1221 ();
 sg13g2_decap_8 FILLER_28_1228 ();
 sg13g2_decap_8 FILLER_28_1235 ();
 sg13g2_decap_8 FILLER_28_1242 ();
 sg13g2_decap_8 FILLER_28_1249 ();
 sg13g2_decap_8 FILLER_28_1256 ();
 sg13g2_decap_8 FILLER_28_1263 ();
 sg13g2_decap_8 FILLER_28_1270 ();
 sg13g2_decap_8 FILLER_28_1277 ();
 sg13g2_decap_8 FILLER_28_1284 ();
 sg13g2_decap_8 FILLER_28_1291 ();
 sg13g2_decap_8 FILLER_28_1298 ();
 sg13g2_decap_8 FILLER_28_1305 ();
 sg13g2_fill_2 FILLER_28_1312 ();
 sg13g2_fill_1 FILLER_28_1314 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_91 ();
 sg13g2_fill_1 FILLER_29_93 ();
 sg13g2_fill_1 FILLER_29_98 ();
 sg13g2_fill_1 FILLER_29_122 ();
 sg13g2_fill_1 FILLER_29_156 ();
 sg13g2_fill_2 FILLER_29_178 ();
 sg13g2_fill_1 FILLER_29_180 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_fill_2 FILLER_29_263 ();
 sg13g2_fill_2 FILLER_29_270 ();
 sg13g2_fill_1 FILLER_29_272 ();
 sg13g2_fill_1 FILLER_29_309 ();
 sg13g2_fill_2 FILLER_29_336 ();
 sg13g2_fill_2 FILLER_29_356 ();
 sg13g2_fill_2 FILLER_29_389 ();
 sg13g2_fill_1 FILLER_29_446 ();
 sg13g2_fill_1 FILLER_29_481 ();
 sg13g2_fill_1 FILLER_29_493 ();
 sg13g2_fill_1 FILLER_29_548 ();
 sg13g2_fill_1 FILLER_29_556 ();
 sg13g2_fill_2 FILLER_29_616 ();
 sg13g2_fill_1 FILLER_29_618 ();
 sg13g2_fill_2 FILLER_29_631 ();
 sg13g2_fill_1 FILLER_29_633 ();
 sg13g2_decap_8 FILLER_29_639 ();
 sg13g2_decap_4 FILLER_29_646 ();
 sg13g2_fill_2 FILLER_29_650 ();
 sg13g2_fill_2 FILLER_29_660 ();
 sg13g2_fill_1 FILLER_29_662 ();
 sg13g2_fill_2 FILLER_29_698 ();
 sg13g2_fill_2 FILLER_29_714 ();
 sg13g2_fill_1 FILLER_29_747 ();
 sg13g2_fill_2 FILLER_29_767 ();
 sg13g2_fill_1 FILLER_29_769 ();
 sg13g2_fill_1 FILLER_29_818 ();
 sg13g2_fill_1 FILLER_29_824 ();
 sg13g2_fill_2 FILLER_29_882 ();
 sg13g2_decap_4 FILLER_29_943 ();
 sg13g2_fill_1 FILLER_29_955 ();
 sg13g2_fill_2 FILLER_29_970 ();
 sg13g2_fill_1 FILLER_29_972 ();
 sg13g2_fill_2 FILLER_29_982 ();
 sg13g2_fill_2 FILLER_29_997 ();
 sg13g2_fill_1 FILLER_29_999 ();
 sg13g2_fill_2 FILLER_29_1014 ();
 sg13g2_fill_1 FILLER_29_1016 ();
 sg13g2_fill_2 FILLER_29_1095 ();
 sg13g2_fill_1 FILLER_29_1097 ();
 sg13g2_fill_1 FILLER_29_1152 ();
 sg13g2_fill_2 FILLER_29_1177 ();
 sg13g2_fill_2 FILLER_29_1184 ();
 sg13g2_fill_1 FILLER_29_1186 ();
 sg13g2_decap_8 FILLER_29_1213 ();
 sg13g2_decap_8 FILLER_29_1220 ();
 sg13g2_decap_8 FILLER_29_1227 ();
 sg13g2_decap_8 FILLER_29_1234 ();
 sg13g2_decap_8 FILLER_29_1241 ();
 sg13g2_decap_8 FILLER_29_1248 ();
 sg13g2_decap_8 FILLER_29_1255 ();
 sg13g2_decap_8 FILLER_29_1262 ();
 sg13g2_decap_8 FILLER_29_1269 ();
 sg13g2_decap_8 FILLER_29_1276 ();
 sg13g2_decap_8 FILLER_29_1283 ();
 sg13g2_decap_8 FILLER_29_1290 ();
 sg13g2_decap_8 FILLER_29_1297 ();
 sg13g2_decap_8 FILLER_29_1304 ();
 sg13g2_decap_4 FILLER_29_1311 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_4 FILLER_30_77 ();
 sg13g2_fill_1 FILLER_30_81 ();
 sg13g2_fill_2 FILLER_30_108 ();
 sg13g2_fill_2 FILLER_30_205 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_213 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_decap_4 FILLER_30_242 ();
 sg13g2_fill_1 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_277 ();
 sg13g2_fill_2 FILLER_30_309 ();
 sg13g2_fill_1 FILLER_30_311 ();
 sg13g2_fill_1 FILLER_30_387 ();
 sg13g2_fill_2 FILLER_30_438 ();
 sg13g2_fill_1 FILLER_30_457 ();
 sg13g2_fill_2 FILLER_30_462 ();
 sg13g2_fill_2 FILLER_30_490 ();
 sg13g2_fill_2 FILLER_30_497 ();
 sg13g2_decap_4 FILLER_30_517 ();
 sg13g2_fill_1 FILLER_30_521 ();
 sg13g2_decap_4 FILLER_30_527 ();
 sg13g2_fill_2 FILLER_30_553 ();
 sg13g2_fill_2 FILLER_30_574 ();
 sg13g2_fill_1 FILLER_30_576 ();
 sg13g2_decap_8 FILLER_30_586 ();
 sg13g2_fill_2 FILLER_30_593 ();
 sg13g2_fill_1 FILLER_30_595 ();
 sg13g2_fill_1 FILLER_30_606 ();
 sg13g2_fill_2 FILLER_30_631 ();
 sg13g2_decap_4 FILLER_30_674 ();
 sg13g2_fill_1 FILLER_30_678 ();
 sg13g2_decap_8 FILLER_30_684 ();
 sg13g2_fill_1 FILLER_30_691 ();
 sg13g2_decap_4 FILLER_30_697 ();
 sg13g2_fill_2 FILLER_30_701 ();
 sg13g2_fill_1 FILLER_30_752 ();
 sg13g2_fill_1 FILLER_30_808 ();
 sg13g2_fill_2 FILLER_30_835 ();
 sg13g2_fill_2 FILLER_30_916 ();
 sg13g2_fill_1 FILLER_30_918 ();
 sg13g2_decap_4 FILLER_30_928 ();
 sg13g2_fill_1 FILLER_30_932 ();
 sg13g2_fill_1 FILLER_30_955 ();
 sg13g2_fill_2 FILLER_30_1016 ();
 sg13g2_fill_1 FILLER_30_1109 ();
 sg13g2_decap_8 FILLER_30_1127 ();
 sg13g2_fill_2 FILLER_30_1138 ();
 sg13g2_decap_4 FILLER_30_1143 ();
 sg13g2_fill_2 FILLER_30_1147 ();
 sg13g2_fill_1 FILLER_30_1165 ();
 sg13g2_decap_8 FILLER_30_1208 ();
 sg13g2_decap_8 FILLER_30_1215 ();
 sg13g2_decap_8 FILLER_30_1222 ();
 sg13g2_decap_8 FILLER_30_1229 ();
 sg13g2_decap_8 FILLER_30_1236 ();
 sg13g2_decap_8 FILLER_30_1243 ();
 sg13g2_decap_8 FILLER_30_1250 ();
 sg13g2_decap_8 FILLER_30_1257 ();
 sg13g2_decap_8 FILLER_30_1264 ();
 sg13g2_decap_8 FILLER_30_1271 ();
 sg13g2_decap_8 FILLER_30_1278 ();
 sg13g2_decap_8 FILLER_30_1285 ();
 sg13g2_decap_8 FILLER_30_1292 ();
 sg13g2_decap_8 FILLER_30_1299 ();
 sg13g2_decap_8 FILLER_30_1306 ();
 sg13g2_fill_2 FILLER_30_1313 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_111 ();
 sg13g2_fill_1 FILLER_31_113 ();
 sg13g2_fill_2 FILLER_31_159 ();
 sg13g2_fill_2 FILLER_31_255 ();
 sg13g2_fill_1 FILLER_31_288 ();
 sg13g2_fill_2 FILLER_31_346 ();
 sg13g2_fill_2 FILLER_31_353 ();
 sg13g2_fill_2 FILLER_31_395 ();
 sg13g2_fill_1 FILLER_31_444 ();
 sg13g2_fill_1 FILLER_31_457 ();
 sg13g2_fill_1 FILLER_31_523 ();
 sg13g2_fill_2 FILLER_31_532 ();
 sg13g2_decap_4 FILLER_31_560 ();
 sg13g2_fill_2 FILLER_31_595 ();
 sg13g2_fill_1 FILLER_31_597 ();
 sg13g2_fill_2 FILLER_31_606 ();
 sg13g2_fill_1 FILLER_31_616 ();
 sg13g2_fill_2 FILLER_31_625 ();
 sg13g2_fill_1 FILLER_31_627 ();
 sg13g2_fill_2 FILLER_31_666 ();
 sg13g2_decap_8 FILLER_31_742 ();
 sg13g2_decap_8 FILLER_31_749 ();
 sg13g2_fill_2 FILLER_31_756 ();
 sg13g2_fill_1 FILLER_31_758 ();
 sg13g2_fill_2 FILLER_31_771 ();
 sg13g2_fill_2 FILLER_31_781 ();
 sg13g2_decap_4 FILLER_31_815 ();
 sg13g2_fill_1 FILLER_31_819 ();
 sg13g2_decap_8 FILLER_31_824 ();
 sg13g2_fill_2 FILLER_31_831 ();
 sg13g2_fill_1 FILLER_31_833 ();
 sg13g2_fill_1 FILLER_31_860 ();
 sg13g2_fill_2 FILLER_31_887 ();
 sg13g2_fill_2 FILLER_31_933 ();
 sg13g2_fill_2 FILLER_31_943 ();
 sg13g2_decap_8 FILLER_31_953 ();
 sg13g2_decap_8 FILLER_31_960 ();
 sg13g2_decap_8 FILLER_31_967 ();
 sg13g2_decap_4 FILLER_31_1003 ();
 sg13g2_fill_2 FILLER_31_1007 ();
 sg13g2_fill_2 FILLER_31_1017 ();
 sg13g2_fill_2 FILLER_31_1071 ();
 sg13g2_fill_2 FILLER_31_1174 ();
 sg13g2_fill_1 FILLER_31_1176 ();
 sg13g2_decap_8 FILLER_31_1213 ();
 sg13g2_decap_8 FILLER_31_1220 ();
 sg13g2_decap_8 FILLER_31_1227 ();
 sg13g2_decap_8 FILLER_31_1234 ();
 sg13g2_decap_8 FILLER_31_1241 ();
 sg13g2_decap_8 FILLER_31_1248 ();
 sg13g2_decap_8 FILLER_31_1255 ();
 sg13g2_decap_8 FILLER_31_1262 ();
 sg13g2_decap_8 FILLER_31_1269 ();
 sg13g2_decap_8 FILLER_31_1276 ();
 sg13g2_decap_8 FILLER_31_1283 ();
 sg13g2_decap_8 FILLER_31_1290 ();
 sg13g2_decap_8 FILLER_31_1297 ();
 sg13g2_decap_8 FILLER_31_1304 ();
 sg13g2_decap_4 FILLER_31_1311 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_4 FILLER_32_70 ();
 sg13g2_fill_1 FILLER_32_74 ();
 sg13g2_fill_2 FILLER_32_101 ();
 sg13g2_fill_1 FILLER_32_103 ();
 sg13g2_fill_2 FILLER_32_130 ();
 sg13g2_fill_1 FILLER_32_132 ();
 sg13g2_fill_2 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_174 ();
 sg13g2_fill_1 FILLER_32_189 ();
 sg13g2_fill_2 FILLER_32_204 ();
 sg13g2_fill_2 FILLER_32_211 ();
 sg13g2_fill_2 FILLER_32_239 ();
 sg13g2_fill_1 FILLER_32_241 ();
 sg13g2_decap_4 FILLER_32_250 ();
 sg13g2_fill_1 FILLER_32_268 ();
 sg13g2_fill_2 FILLER_32_320 ();
 sg13g2_fill_2 FILLER_32_353 ();
 sg13g2_fill_1 FILLER_32_461 ();
 sg13g2_fill_2 FILLER_32_471 ();
 sg13g2_fill_1 FILLER_32_511 ();
 sg13g2_decap_4 FILLER_32_527 ();
 sg13g2_fill_1 FILLER_32_544 ();
 sg13g2_fill_1 FILLER_32_552 ();
 sg13g2_fill_2 FILLER_32_577 ();
 sg13g2_fill_1 FILLER_32_579 ();
 sg13g2_fill_2 FILLER_32_589 ();
 sg13g2_fill_1 FILLER_32_591 ();
 sg13g2_decap_8 FILLER_32_601 ();
 sg13g2_fill_2 FILLER_32_608 ();
 sg13g2_fill_1 FILLER_32_610 ();
 sg13g2_fill_1 FILLER_32_623 ();
 sg13g2_fill_2 FILLER_32_633 ();
 sg13g2_fill_1 FILLER_32_635 ();
 sg13g2_decap_8 FILLER_32_649 ();
 sg13g2_fill_2 FILLER_32_671 ();
 sg13g2_decap_4 FILLER_32_680 ();
 sg13g2_fill_2 FILLER_32_690 ();
 sg13g2_fill_1 FILLER_32_718 ();
 sg13g2_decap_8 FILLER_32_743 ();
 sg13g2_fill_2 FILLER_32_750 ();
 sg13g2_fill_2 FILLER_32_794 ();
 sg13g2_fill_2 FILLER_32_803 ();
 sg13g2_fill_2 FILLER_32_817 ();
 sg13g2_fill_1 FILLER_32_819 ();
 sg13g2_fill_2 FILLER_32_825 ();
 sg13g2_fill_1 FILLER_32_827 ();
 sg13g2_decap_8 FILLER_32_832 ();
 sg13g2_fill_2 FILLER_32_839 ();
 sg13g2_fill_2 FILLER_32_868 ();
 sg13g2_fill_1 FILLER_32_870 ();
 sg13g2_fill_2 FILLER_32_880 ();
 sg13g2_decap_8 FILLER_32_892 ();
 sg13g2_fill_2 FILLER_32_899 ();
 sg13g2_fill_2 FILLER_32_909 ();
 sg13g2_fill_2 FILLER_32_966 ();
 sg13g2_fill_2 FILLER_32_981 ();
 sg13g2_fill_1 FILLER_32_983 ();
 sg13g2_fill_2 FILLER_32_997 ();
 sg13g2_fill_1 FILLER_32_999 ();
 sg13g2_fill_1 FILLER_32_1047 ();
 sg13g2_fill_2 FILLER_32_1060 ();
 sg13g2_fill_2 FILLER_32_1094 ();
 sg13g2_fill_2 FILLER_32_1101 ();
 sg13g2_fill_1 FILLER_32_1103 ();
 sg13g2_decap_4 FILLER_32_1121 ();
 sg13g2_fill_2 FILLER_32_1125 ();
 sg13g2_fill_2 FILLER_32_1140 ();
 sg13g2_fill_2 FILLER_32_1188 ();
 sg13g2_decap_8 FILLER_32_1220 ();
 sg13g2_decap_8 FILLER_32_1227 ();
 sg13g2_decap_8 FILLER_32_1234 ();
 sg13g2_decap_8 FILLER_32_1241 ();
 sg13g2_decap_8 FILLER_32_1248 ();
 sg13g2_decap_8 FILLER_32_1255 ();
 sg13g2_decap_8 FILLER_32_1262 ();
 sg13g2_decap_8 FILLER_32_1269 ();
 sg13g2_decap_8 FILLER_32_1276 ();
 sg13g2_decap_8 FILLER_32_1283 ();
 sg13g2_decap_8 FILLER_32_1290 ();
 sg13g2_decap_8 FILLER_32_1297 ();
 sg13g2_decap_8 FILLER_32_1304 ();
 sg13g2_decap_4 FILLER_32_1311 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_4 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_81 ();
 sg13g2_fill_2 FILLER_33_108 ();
 sg13g2_fill_2 FILLER_33_174 ();
 sg13g2_fill_1 FILLER_33_190 ();
 sg13g2_fill_2 FILLER_33_243 ();
 sg13g2_fill_1 FILLER_33_245 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_290 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_374 ();
 sg13g2_fill_2 FILLER_33_384 ();
 sg13g2_fill_2 FILLER_33_411 ();
 sg13g2_fill_1 FILLER_33_501 ();
 sg13g2_fill_1 FILLER_33_515 ();
 sg13g2_fill_2 FILLER_33_568 ();
 sg13g2_fill_1 FILLER_33_570 ();
 sg13g2_decap_4 FILLER_33_579 ();
 sg13g2_decap_8 FILLER_33_621 ();
 sg13g2_fill_1 FILLER_33_658 ();
 sg13g2_decap_8 FILLER_33_673 ();
 sg13g2_fill_2 FILLER_33_680 ();
 sg13g2_decap_8 FILLER_33_687 ();
 sg13g2_fill_1 FILLER_33_735 ();
 sg13g2_fill_2 FILLER_33_767 ();
 sg13g2_fill_1 FILLER_33_769 ();
 sg13g2_fill_1 FILLER_33_843 ();
 sg13g2_fill_1 FILLER_33_859 ();
 sg13g2_fill_1 FILLER_33_881 ();
 sg13g2_fill_2 FILLER_33_986 ();
 sg13g2_fill_1 FILLER_33_988 ();
 sg13g2_fill_2 FILLER_33_1020 ();
 sg13g2_fill_2 FILLER_33_1045 ();
 sg13g2_fill_2 FILLER_33_1064 ();
 sg13g2_decap_4 FILLER_33_1160 ();
 sg13g2_fill_2 FILLER_33_1164 ();
 sg13g2_decap_8 FILLER_33_1170 ();
 sg13g2_decap_4 FILLER_33_1177 ();
 sg13g2_fill_1 FILLER_33_1181 ();
 sg13g2_fill_1 FILLER_33_1198 ();
 sg13g2_decap_8 FILLER_33_1225 ();
 sg13g2_decap_8 FILLER_33_1232 ();
 sg13g2_decap_8 FILLER_33_1239 ();
 sg13g2_decap_8 FILLER_33_1246 ();
 sg13g2_decap_8 FILLER_33_1253 ();
 sg13g2_decap_8 FILLER_33_1260 ();
 sg13g2_decap_8 FILLER_33_1267 ();
 sg13g2_decap_8 FILLER_33_1274 ();
 sg13g2_decap_8 FILLER_33_1281 ();
 sg13g2_decap_8 FILLER_33_1288 ();
 sg13g2_decap_8 FILLER_33_1295 ();
 sg13g2_decap_8 FILLER_33_1302 ();
 sg13g2_decap_4 FILLER_33_1309 ();
 sg13g2_fill_2 FILLER_33_1313 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_fill_2 FILLER_34_124 ();
 sg13g2_fill_1 FILLER_34_126 ();
 sg13g2_fill_1 FILLER_34_161 ();
 sg13g2_fill_1 FILLER_34_167 ();
 sg13g2_fill_2 FILLER_34_172 ();
 sg13g2_fill_1 FILLER_34_174 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_212 ();
 sg13g2_fill_1 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_decap_4 FILLER_34_252 ();
 sg13g2_fill_1 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_261 ();
 sg13g2_fill_2 FILLER_34_271 ();
 sg13g2_fill_1 FILLER_34_286 ();
 sg13g2_fill_1 FILLER_34_348 ();
 sg13g2_fill_2 FILLER_34_358 ();
 sg13g2_fill_1 FILLER_34_386 ();
 sg13g2_fill_2 FILLER_34_396 ();
 sg13g2_fill_1 FILLER_34_418 ();
 sg13g2_fill_2 FILLER_34_424 ();
 sg13g2_fill_1 FILLER_34_454 ();
 sg13g2_fill_2 FILLER_34_534 ();
 sg13g2_fill_1 FILLER_34_546 ();
 sg13g2_fill_1 FILLER_34_561 ();
 sg13g2_fill_2 FILLER_34_577 ();
 sg13g2_fill_2 FILLER_34_594 ();
 sg13g2_fill_1 FILLER_34_622 ();
 sg13g2_fill_2 FILLER_34_649 ();
 sg13g2_fill_1 FILLER_34_651 ();
 sg13g2_fill_2 FILLER_34_661 ();
 sg13g2_decap_4 FILLER_34_671 ();
 sg13g2_fill_2 FILLER_34_688 ();
 sg13g2_fill_1 FILLER_34_690 ();
 sg13g2_fill_2 FILLER_34_699 ();
 sg13g2_fill_2 FILLER_34_718 ();
 sg13g2_fill_2 FILLER_34_727 ();
 sg13g2_fill_1 FILLER_34_729 ();
 sg13g2_fill_1 FILLER_34_751 ();
 sg13g2_fill_1 FILLER_34_761 ();
 sg13g2_fill_1 FILLER_34_771 ();
 sg13g2_fill_2 FILLER_34_818 ();
 sg13g2_fill_1 FILLER_34_820 ();
 sg13g2_fill_2 FILLER_34_862 ();
 sg13g2_fill_1 FILLER_34_864 ();
 sg13g2_fill_2 FILLER_34_906 ();
 sg13g2_fill_1 FILLER_34_908 ();
 sg13g2_fill_2 FILLER_34_919 ();
 sg13g2_fill_1 FILLER_34_956 ();
 sg13g2_decap_4 FILLER_34_961 ();
 sg13g2_fill_1 FILLER_34_975 ();
 sg13g2_fill_2 FILLER_34_995 ();
 sg13g2_fill_1 FILLER_34_997 ();
 sg13g2_fill_2 FILLER_34_1007 ();
 sg13g2_fill_1 FILLER_34_1078 ();
 sg13g2_fill_2 FILLER_34_1088 ();
 sg13g2_fill_2 FILLER_34_1099 ();
 sg13g2_fill_1 FILLER_34_1101 ();
 sg13g2_fill_2 FILLER_34_1138 ();
 sg13g2_fill_1 FILLER_34_1153 ();
 sg13g2_fill_1 FILLER_34_1211 ();
 sg13g2_decap_8 FILLER_34_1229 ();
 sg13g2_decap_8 FILLER_34_1236 ();
 sg13g2_decap_8 FILLER_34_1243 ();
 sg13g2_decap_8 FILLER_34_1250 ();
 sg13g2_decap_8 FILLER_34_1257 ();
 sg13g2_decap_8 FILLER_34_1264 ();
 sg13g2_decap_8 FILLER_34_1271 ();
 sg13g2_decap_8 FILLER_34_1278 ();
 sg13g2_decap_8 FILLER_34_1285 ();
 sg13g2_decap_8 FILLER_34_1292 ();
 sg13g2_decap_8 FILLER_34_1299 ();
 sg13g2_decap_8 FILLER_34_1306 ();
 sg13g2_fill_2 FILLER_34_1313 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_4 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_85 ();
 sg13g2_fill_1 FILLER_35_87 ();
 sg13g2_fill_2 FILLER_35_111 ();
 sg13g2_fill_2 FILLER_35_139 ();
 sg13g2_fill_2 FILLER_35_150 ();
 sg13g2_fill_2 FILLER_35_178 ();
 sg13g2_fill_1 FILLER_35_180 ();
 sg13g2_decap_4 FILLER_35_234 ();
 sg13g2_fill_2 FILLER_35_277 ();
 sg13g2_fill_2 FILLER_35_322 ();
 sg13g2_fill_1 FILLER_35_385 ();
 sg13g2_fill_1 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_496 ();
 sg13g2_fill_2 FILLER_35_619 ();
 sg13g2_fill_2 FILLER_35_626 ();
 sg13g2_decap_8 FILLER_35_632 ();
 sg13g2_fill_2 FILLER_35_639 ();
 sg13g2_fill_1 FILLER_35_641 ();
 sg13g2_fill_2 FILLER_35_655 ();
 sg13g2_fill_1 FILLER_35_657 ();
 sg13g2_decap_4 FILLER_35_665 ();
 sg13g2_fill_2 FILLER_35_669 ();
 sg13g2_fill_2 FILLER_35_676 ();
 sg13g2_fill_1 FILLER_35_678 ();
 sg13g2_fill_2 FILLER_35_693 ();
 sg13g2_fill_1 FILLER_35_695 ();
 sg13g2_fill_1 FILLER_35_701 ();
 sg13g2_decap_8 FILLER_35_720 ();
 sg13g2_fill_1 FILLER_35_727 ();
 sg13g2_fill_2 FILLER_35_747 ();
 sg13g2_fill_2 FILLER_35_783 ();
 sg13g2_fill_1 FILLER_35_798 ();
 sg13g2_fill_1 FILLER_35_851 ();
 sg13g2_decap_8 FILLER_35_872 ();
 sg13g2_decap_8 FILLER_35_879 ();
 sg13g2_decap_4 FILLER_35_886 ();
 sg13g2_fill_1 FILLER_35_890 ();
 sg13g2_decap_8 FILLER_35_895 ();
 sg13g2_fill_1 FILLER_35_912 ();
 sg13g2_fill_2 FILLER_35_922 ();
 sg13g2_fill_2 FILLER_35_933 ();
 sg13g2_fill_1 FILLER_35_964 ();
 sg13g2_fill_2 FILLER_35_1026 ();
 sg13g2_fill_1 FILLER_35_1028 ();
 sg13g2_fill_1 FILLER_35_1038 ();
 sg13g2_fill_2 FILLER_35_1044 ();
 sg13g2_fill_1 FILLER_35_1059 ();
 sg13g2_fill_2 FILLER_35_1070 ();
 sg13g2_fill_1 FILLER_35_1103 ();
 sg13g2_fill_1 FILLER_35_1145 ();
 sg13g2_fill_1 FILLER_35_1162 ();
 sg13g2_fill_1 FILLER_35_1203 ();
 sg13g2_decap_8 FILLER_35_1230 ();
 sg13g2_decap_8 FILLER_35_1237 ();
 sg13g2_decap_8 FILLER_35_1244 ();
 sg13g2_decap_8 FILLER_35_1251 ();
 sg13g2_decap_8 FILLER_35_1258 ();
 sg13g2_decap_8 FILLER_35_1265 ();
 sg13g2_decap_8 FILLER_35_1272 ();
 sg13g2_decap_8 FILLER_35_1279 ();
 sg13g2_decap_8 FILLER_35_1286 ();
 sg13g2_decap_8 FILLER_35_1293 ();
 sg13g2_decap_8 FILLER_35_1300 ();
 sg13g2_decap_8 FILLER_35_1307 ();
 sg13g2_fill_1 FILLER_35_1314 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_4 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_74 ();
 sg13g2_fill_2 FILLER_36_102 ();
 sg13g2_fill_1 FILLER_36_104 ();
 sg13g2_fill_2 FILLER_36_166 ();
 sg13g2_fill_1 FILLER_36_168 ();
 sg13g2_fill_1 FILLER_36_196 ();
 sg13g2_fill_1 FILLER_36_206 ();
 sg13g2_decap_8 FILLER_36_215 ();
 sg13g2_decap_4 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_fill_2 FILLER_36_257 ();
 sg13g2_fill_1 FILLER_36_276 ();
 sg13g2_fill_1 FILLER_36_320 ();
 sg13g2_fill_1 FILLER_36_334 ();
 sg13g2_fill_1 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_419 ();
 sg13g2_fill_1 FILLER_36_421 ();
 sg13g2_fill_2 FILLER_36_432 ();
 sg13g2_fill_1 FILLER_36_447 ();
 sg13g2_fill_2 FILLER_36_544 ();
 sg13g2_fill_1 FILLER_36_546 ();
 sg13g2_decap_8 FILLER_36_569 ();
 sg13g2_decap_4 FILLER_36_576 ();
 sg13g2_fill_2 FILLER_36_580 ();
 sg13g2_decap_8 FILLER_36_600 ();
 sg13g2_fill_2 FILLER_36_624 ();
 sg13g2_fill_1 FILLER_36_670 ();
 sg13g2_fill_1 FILLER_36_697 ();
 sg13g2_fill_1 FILLER_36_724 ();
 sg13g2_fill_1 FILLER_36_797 ();
 sg13g2_decap_4 FILLER_36_841 ();
 sg13g2_decap_4 FILLER_36_850 ();
 sg13g2_decap_4 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_863 ();
 sg13g2_fill_2 FILLER_36_899 ();
 sg13g2_fill_1 FILLER_36_901 ();
 sg13g2_fill_1 FILLER_36_923 ();
 sg13g2_fill_1 FILLER_36_950 ();
 sg13g2_fill_1 FILLER_36_984 ();
 sg13g2_fill_2 FILLER_36_1029 ();
 sg13g2_fill_1 FILLER_36_1031 ();
 sg13g2_fill_1 FILLER_36_1124 ();
 sg13g2_fill_1 FILLER_36_1151 ();
 sg13g2_fill_1 FILLER_36_1189 ();
 sg13g2_decap_8 FILLER_36_1215 ();
 sg13g2_decap_8 FILLER_36_1222 ();
 sg13g2_decap_8 FILLER_36_1229 ();
 sg13g2_decap_8 FILLER_36_1236 ();
 sg13g2_decap_8 FILLER_36_1243 ();
 sg13g2_decap_8 FILLER_36_1250 ();
 sg13g2_decap_8 FILLER_36_1257 ();
 sg13g2_decap_8 FILLER_36_1264 ();
 sg13g2_decap_8 FILLER_36_1271 ();
 sg13g2_decap_8 FILLER_36_1278 ();
 sg13g2_decap_8 FILLER_36_1285 ();
 sg13g2_decap_8 FILLER_36_1292 ();
 sg13g2_decap_8 FILLER_36_1299 ();
 sg13g2_decap_8 FILLER_36_1306 ();
 sg13g2_fill_2 FILLER_36_1313 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_4 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_fill_2 FILLER_37_85 ();
 sg13g2_decap_4 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_95 ();
 sg13g2_decap_4 FILLER_37_100 ();
 sg13g2_fill_2 FILLER_37_144 ();
 sg13g2_fill_1 FILLER_37_146 ();
 sg13g2_fill_2 FILLER_37_243 ();
 sg13g2_fill_1 FILLER_37_370 ();
 sg13g2_fill_1 FILLER_37_480 ();
 sg13g2_fill_2 FILLER_37_496 ();
 sg13g2_decap_4 FILLER_37_578 ();
 sg13g2_fill_1 FILLER_37_582 ();
 sg13g2_decap_8 FILLER_37_588 ();
 sg13g2_fill_2 FILLER_37_595 ();
 sg13g2_decap_8 FILLER_37_620 ();
 sg13g2_fill_2 FILLER_37_627 ();
 sg13g2_fill_1 FILLER_37_629 ();
 sg13g2_decap_8 FILLER_37_640 ();
 sg13g2_decap_8 FILLER_37_647 ();
 sg13g2_decap_4 FILLER_37_654 ();
 sg13g2_fill_2 FILLER_37_662 ();
 sg13g2_decap_4 FILLER_37_668 ();
 sg13g2_fill_1 FILLER_37_677 ();
 sg13g2_decap_8 FILLER_37_687 ();
 sg13g2_decap_4 FILLER_37_699 ();
 sg13g2_fill_1 FILLER_37_703 ();
 sg13g2_fill_2 FILLER_37_717 ();
 sg13g2_fill_1 FILLER_37_719 ();
 sg13g2_fill_2 FILLER_37_728 ();
 sg13g2_fill_1 FILLER_37_730 ();
 sg13g2_fill_1 FILLER_37_736 ();
 sg13g2_fill_2 FILLER_37_742 ();
 sg13g2_fill_1 FILLER_37_744 ();
 sg13g2_fill_2 FILLER_37_790 ();
 sg13g2_decap_4 FILLER_37_839 ();
 sg13g2_decap_4 FILLER_37_850 ();
 sg13g2_fill_1 FILLER_37_885 ();
 sg13g2_fill_1 FILLER_37_895 ();
 sg13g2_fill_1 FILLER_37_908 ();
 sg13g2_fill_1 FILLER_37_915 ();
 sg13g2_fill_2 FILLER_37_931 ();
 sg13g2_fill_1 FILLER_37_933 ();
 sg13g2_decap_4 FILLER_37_951 ();
 sg13g2_fill_1 FILLER_37_981 ();
 sg13g2_decap_4 FILLER_37_1008 ();
 sg13g2_fill_2 FILLER_37_1012 ();
 sg13g2_fill_2 FILLER_37_1062 ();
 sg13g2_fill_2 FILLER_37_1095 ();
 sg13g2_fill_2 FILLER_37_1106 ();
 sg13g2_fill_2 FILLER_37_1135 ();
 sg13g2_fill_2 FILLER_37_1154 ();
 sg13g2_fill_2 FILLER_37_1190 ();
 sg13g2_fill_2 FILLER_37_1220 ();
 sg13g2_fill_1 FILLER_37_1222 ();
 sg13g2_decap_8 FILLER_37_1226 ();
 sg13g2_decap_8 FILLER_37_1233 ();
 sg13g2_decap_8 FILLER_37_1240 ();
 sg13g2_decap_8 FILLER_37_1247 ();
 sg13g2_decap_8 FILLER_37_1254 ();
 sg13g2_decap_8 FILLER_37_1261 ();
 sg13g2_decap_8 FILLER_37_1268 ();
 sg13g2_decap_8 FILLER_37_1275 ();
 sg13g2_decap_8 FILLER_37_1282 ();
 sg13g2_decap_8 FILLER_37_1289 ();
 sg13g2_decap_8 FILLER_37_1296 ();
 sg13g2_decap_8 FILLER_37_1303 ();
 sg13g2_decap_4 FILLER_37_1310 ();
 sg13g2_fill_1 FILLER_37_1314 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_56 ();
 sg13g2_fill_2 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_74 ();
 sg13g2_fill_2 FILLER_38_129 ();
 sg13g2_fill_2 FILLER_38_136 ();
 sg13g2_fill_1 FILLER_38_138 ();
 sg13g2_fill_1 FILLER_38_153 ();
 sg13g2_fill_1 FILLER_38_167 ();
 sg13g2_fill_1 FILLER_38_193 ();
 sg13g2_fill_1 FILLER_38_217 ();
 sg13g2_fill_2 FILLER_38_258 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_fill_2 FILLER_38_281 ();
 sg13g2_fill_1 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_298 ();
 sg13g2_fill_2 FILLER_38_324 ();
 sg13g2_fill_2 FILLER_38_340 ();
 sg13g2_fill_1 FILLER_38_403 ();
 sg13g2_fill_1 FILLER_38_425 ();
 sg13g2_fill_1 FILLER_38_473 ();
 sg13g2_fill_1 FILLER_38_487 ();
 sg13g2_decap_4 FILLER_38_500 ();
 sg13g2_fill_2 FILLER_38_504 ();
 sg13g2_fill_2 FILLER_38_569 ();
 sg13g2_fill_1 FILLER_38_571 ();
 sg13g2_fill_1 FILLER_38_604 ();
 sg13g2_fill_1 FILLER_38_664 ();
 sg13g2_decap_4 FILLER_38_670 ();
 sg13g2_fill_1 FILLER_38_674 ();
 sg13g2_decap_4 FILLER_38_682 ();
 sg13g2_fill_2 FILLER_38_686 ();
 sg13g2_fill_2 FILLER_38_719 ();
 sg13g2_fill_1 FILLER_38_743 ();
 sg13g2_fill_2 FILLER_38_774 ();
 sg13g2_fill_2 FILLER_38_828 ();
 sg13g2_fill_1 FILLER_38_830 ();
 sg13g2_fill_2 FILLER_38_841 ();
 sg13g2_decap_8 FILLER_38_857 ();
 sg13g2_decap_4 FILLER_38_868 ();
 sg13g2_fill_1 FILLER_38_908 ();
 sg13g2_decap_8 FILLER_38_950 ();
 sg13g2_fill_1 FILLER_38_957 ();
 sg13g2_decap_4 FILLER_38_962 ();
 sg13g2_decap_8 FILLER_38_970 ();
 sg13g2_decap_8 FILLER_38_977 ();
 sg13g2_decap_4 FILLER_38_988 ();
 sg13g2_fill_1 FILLER_38_992 ();
 sg13g2_fill_2 FILLER_38_1001 ();
 sg13g2_fill_1 FILLER_38_1003 ();
 sg13g2_decap_4 FILLER_38_1047 ();
 sg13g2_fill_1 FILLER_38_1073 ();
 sg13g2_decap_8 FILLER_38_1159 ();
 sg13g2_decap_4 FILLER_38_1170 ();
 sg13g2_decap_8 FILLER_38_1177 ();
 sg13g2_decap_4 FILLER_38_1184 ();
 sg13g2_fill_1 FILLER_38_1188 ();
 sg13g2_fill_1 FILLER_38_1223 ();
 sg13g2_decap_8 FILLER_38_1233 ();
 sg13g2_decap_8 FILLER_38_1240 ();
 sg13g2_decap_8 FILLER_38_1247 ();
 sg13g2_decap_8 FILLER_38_1254 ();
 sg13g2_decap_8 FILLER_38_1261 ();
 sg13g2_decap_8 FILLER_38_1268 ();
 sg13g2_decap_8 FILLER_38_1275 ();
 sg13g2_decap_8 FILLER_38_1282 ();
 sg13g2_decap_8 FILLER_38_1289 ();
 sg13g2_decap_8 FILLER_38_1296 ();
 sg13g2_decap_8 FILLER_38_1303 ();
 sg13g2_decap_4 FILLER_38_1310 ();
 sg13g2_fill_1 FILLER_38_1314 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_fill_2 FILLER_39_70 ();
 sg13g2_fill_1 FILLER_39_72 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_fill_1 FILLER_39_84 ();
 sg13g2_fill_2 FILLER_39_93 ();
 sg13g2_fill_1 FILLER_39_147 ();
 sg13g2_fill_2 FILLER_39_195 ();
 sg13g2_fill_2 FILLER_39_211 ();
 sg13g2_fill_1 FILLER_39_213 ();
 sg13g2_fill_2 FILLER_39_226 ();
 sg13g2_fill_1 FILLER_39_236 ();
 sg13g2_fill_2 FILLER_39_265 ();
 sg13g2_fill_1 FILLER_39_267 ();
 sg13g2_fill_2 FILLER_39_273 ();
 sg13g2_fill_1 FILLER_39_310 ();
 sg13g2_fill_1 FILLER_39_325 ();
 sg13g2_fill_2 FILLER_39_348 ();
 sg13g2_fill_2 FILLER_39_354 ();
 sg13g2_fill_2 FILLER_39_396 ();
 sg13g2_fill_2 FILLER_39_421 ();
 sg13g2_fill_1 FILLER_39_467 ();
 sg13g2_fill_2 FILLER_39_511 ();
 sg13g2_fill_1 FILLER_39_536 ();
 sg13g2_decap_4 FILLER_39_577 ();
 sg13g2_fill_1 FILLER_39_581 ();
 sg13g2_fill_1 FILLER_39_587 ();
 sg13g2_decap_4 FILLER_39_719 ();
 sg13g2_fill_2 FILLER_39_727 ();
 sg13g2_fill_1 FILLER_39_742 ();
 sg13g2_fill_1 FILLER_39_762 ();
 sg13g2_fill_1 FILLER_39_773 ();
 sg13g2_fill_2 FILLER_39_783 ();
 sg13g2_fill_1 FILLER_39_811 ();
 sg13g2_decap_4 FILLER_39_846 ();
 sg13g2_fill_1 FILLER_39_850 ();
 sg13g2_fill_1 FILLER_39_855 ();
 sg13g2_fill_1 FILLER_39_865 ();
 sg13g2_fill_2 FILLER_39_876 ();
 sg13g2_fill_2 FILLER_39_917 ();
 sg13g2_decap_8 FILLER_39_928 ();
 sg13g2_fill_2 FILLER_39_935 ();
 sg13g2_decap_8 FILLER_39_973 ();
 sg13g2_fill_2 FILLER_39_980 ();
 sg13g2_fill_1 FILLER_39_982 ();
 sg13g2_fill_1 FILLER_39_1019 ();
 sg13g2_decap_4 FILLER_39_1046 ();
 sg13g2_fill_2 FILLER_39_1081 ();
 sg13g2_fill_2 FILLER_39_1114 ();
 sg13g2_decap_8 FILLER_39_1128 ();
 sg13g2_decap_8 FILLER_39_1135 ();
 sg13g2_fill_2 FILLER_39_1142 ();
 sg13g2_fill_2 FILLER_39_1153 ();
 sg13g2_fill_1 FILLER_39_1155 ();
 sg13g2_fill_2 FILLER_39_1175 ();
 sg13g2_decap_8 FILLER_39_1224 ();
 sg13g2_decap_8 FILLER_39_1231 ();
 sg13g2_decap_8 FILLER_39_1238 ();
 sg13g2_decap_8 FILLER_39_1245 ();
 sg13g2_decap_8 FILLER_39_1252 ();
 sg13g2_decap_8 FILLER_39_1259 ();
 sg13g2_decap_8 FILLER_39_1266 ();
 sg13g2_decap_8 FILLER_39_1273 ();
 sg13g2_decap_8 FILLER_39_1280 ();
 sg13g2_decap_8 FILLER_39_1287 ();
 sg13g2_decap_8 FILLER_39_1294 ();
 sg13g2_decap_8 FILLER_39_1301 ();
 sg13g2_decap_8 FILLER_39_1308 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_4 FILLER_40_56 ();
 sg13g2_fill_1 FILLER_40_60 ();
 sg13g2_fill_2 FILLER_40_75 ();
 sg13g2_fill_1 FILLER_40_77 ();
 sg13g2_fill_1 FILLER_40_83 ();
 sg13g2_decap_8 FILLER_40_97 ();
 sg13g2_fill_2 FILLER_40_104 ();
 sg13g2_fill_2 FILLER_40_110 ();
 sg13g2_fill_2 FILLER_40_116 ();
 sg13g2_fill_2 FILLER_40_136 ();
 sg13g2_fill_1 FILLER_40_138 ();
 sg13g2_fill_1 FILLER_40_173 ();
 sg13g2_decap_4 FILLER_40_228 ();
 sg13g2_fill_1 FILLER_40_232 ();
 sg13g2_fill_2 FILLER_40_236 ();
 sg13g2_fill_2 FILLER_40_296 ();
 sg13g2_fill_2 FILLER_40_324 ();
 sg13g2_fill_1 FILLER_40_347 ();
 sg13g2_fill_2 FILLER_40_388 ();
 sg13g2_fill_2 FILLER_40_437 ();
 sg13g2_fill_1 FILLER_40_439 ();
 sg13g2_fill_2 FILLER_40_488 ();
 sg13g2_fill_1 FILLER_40_490 ();
 sg13g2_fill_1 FILLER_40_501 ();
 sg13g2_fill_2 FILLER_40_506 ();
 sg13g2_decap_8 FILLER_40_513 ();
 sg13g2_fill_1 FILLER_40_525 ();
 sg13g2_fill_2 FILLER_40_570 ();
 sg13g2_fill_1 FILLER_40_572 ();
 sg13g2_decap_8 FILLER_40_576 ();
 sg13g2_fill_2 FILLER_40_583 ();
 sg13g2_decap_8 FILLER_40_590 ();
 sg13g2_fill_1 FILLER_40_597 ();
 sg13g2_fill_2 FILLER_40_606 ();
 sg13g2_fill_1 FILLER_40_608 ();
 sg13g2_fill_1 FILLER_40_613 ();
 sg13g2_fill_1 FILLER_40_622 ();
 sg13g2_fill_1 FILLER_40_629 ();
 sg13g2_decap_8 FILLER_40_670 ();
 sg13g2_decap_8 FILLER_40_677 ();
 sg13g2_decap_4 FILLER_40_684 ();
 sg13g2_fill_1 FILLER_40_688 ();
 sg13g2_fill_2 FILLER_40_724 ();
 sg13g2_fill_1 FILLER_40_830 ();
 sg13g2_fill_2 FILLER_40_922 ();
 sg13g2_fill_1 FILLER_40_931 ();
 sg13g2_decap_8 FILLER_40_948 ();
 sg13g2_fill_1 FILLER_40_960 ();
 sg13g2_fill_1 FILLER_40_1020 ();
 sg13g2_fill_2 FILLER_40_1044 ();
 sg13g2_fill_2 FILLER_40_1093 ();
 sg13g2_fill_1 FILLER_40_1095 ();
 sg13g2_decap_8 FILLER_40_1122 ();
 sg13g2_decap_8 FILLER_40_1129 ();
 sg13g2_fill_2 FILLER_40_1136 ();
 sg13g2_decap_8 FILLER_40_1225 ();
 sg13g2_decap_8 FILLER_40_1232 ();
 sg13g2_decap_8 FILLER_40_1239 ();
 sg13g2_decap_8 FILLER_40_1246 ();
 sg13g2_decap_8 FILLER_40_1253 ();
 sg13g2_decap_8 FILLER_40_1260 ();
 sg13g2_decap_8 FILLER_40_1267 ();
 sg13g2_decap_8 FILLER_40_1274 ();
 sg13g2_decap_8 FILLER_40_1281 ();
 sg13g2_decap_8 FILLER_40_1288 ();
 sg13g2_decap_8 FILLER_40_1295 ();
 sg13g2_decap_8 FILLER_40_1302 ();
 sg13g2_decap_4 FILLER_40_1309 ();
 sg13g2_fill_2 FILLER_40_1313 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_fill_2 FILLER_41_56 ();
 sg13g2_fill_2 FILLER_41_67 ();
 sg13g2_fill_1 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_92 ();
 sg13g2_fill_2 FILLER_41_99 ();
 sg13g2_fill_2 FILLER_41_127 ();
 sg13g2_fill_1 FILLER_41_155 ();
 sg13g2_decap_4 FILLER_41_217 ();
 sg13g2_fill_1 FILLER_41_221 ();
 sg13g2_fill_2 FILLER_41_230 ();
 sg13g2_fill_1 FILLER_41_249 ();
 sg13g2_fill_2 FILLER_41_260 ();
 sg13g2_fill_1 FILLER_41_262 ();
 sg13g2_fill_2 FILLER_41_292 ();
 sg13g2_fill_2 FILLER_41_368 ();
 sg13g2_fill_1 FILLER_41_370 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_decap_8 FILLER_41_416 ();
 sg13g2_fill_2 FILLER_41_423 ();
 sg13g2_fill_1 FILLER_41_425 ();
 sg13g2_fill_2 FILLER_41_488 ();
 sg13g2_fill_1 FILLER_41_490 ();
 sg13g2_decap_4 FILLER_41_525 ();
 sg13g2_fill_2 FILLER_41_542 ();
 sg13g2_fill_1 FILLER_41_544 ();
 sg13g2_decap_4 FILLER_41_558 ();
 sg13g2_fill_1 FILLER_41_562 ();
 sg13g2_fill_1 FILLER_41_572 ();
 sg13g2_fill_1 FILLER_41_607 ();
 sg13g2_fill_2 FILLER_41_617 ();
 sg13g2_fill_1 FILLER_41_653 ();
 sg13g2_fill_1 FILLER_41_659 ();
 sg13g2_decap_4 FILLER_41_686 ();
 sg13g2_fill_2 FILLER_41_695 ();
 sg13g2_fill_1 FILLER_41_697 ();
 sg13g2_fill_1 FILLER_41_712 ();
 sg13g2_fill_1 FILLER_41_756 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_4 FILLER_41_777 ();
 sg13g2_fill_2 FILLER_41_781 ();
 sg13g2_decap_8 FILLER_41_792 ();
 sg13g2_decap_8 FILLER_41_799 ();
 sg13g2_fill_2 FILLER_41_811 ();
 sg13g2_fill_1 FILLER_41_817 ();
 sg13g2_fill_2 FILLER_41_832 ();
 sg13g2_fill_1 FILLER_41_834 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_41_847 ();
 sg13g2_decap_4 FILLER_41_854 ();
 sg13g2_fill_1 FILLER_41_858 ();
 sg13g2_decap_8 FILLER_41_868 ();
 sg13g2_fill_2 FILLER_41_875 ();
 sg13g2_fill_1 FILLER_41_877 ();
 sg13g2_decap_4 FILLER_41_945 ();
 sg13g2_fill_2 FILLER_41_959 ();
 sg13g2_fill_1 FILLER_41_961 ();
 sg13g2_fill_1 FILLER_41_979 ();
 sg13g2_fill_1 FILLER_41_997 ();
 sg13g2_fill_1 FILLER_41_1016 ();
 sg13g2_fill_1 FILLER_41_1052 ();
 sg13g2_fill_2 FILLER_41_1175 ();
 sg13g2_fill_2 FILLER_41_1182 ();
 sg13g2_fill_1 FILLER_41_1184 ();
 sg13g2_fill_2 FILLER_41_1208 ();
 sg13g2_decap_8 FILLER_41_1214 ();
 sg13g2_decap_8 FILLER_41_1221 ();
 sg13g2_decap_8 FILLER_41_1228 ();
 sg13g2_decap_8 FILLER_41_1235 ();
 sg13g2_decap_8 FILLER_41_1242 ();
 sg13g2_decap_8 FILLER_41_1249 ();
 sg13g2_decap_8 FILLER_41_1256 ();
 sg13g2_decap_8 FILLER_41_1263 ();
 sg13g2_decap_8 FILLER_41_1270 ();
 sg13g2_decap_8 FILLER_41_1277 ();
 sg13g2_decap_8 FILLER_41_1284 ();
 sg13g2_decap_8 FILLER_41_1291 ();
 sg13g2_decap_8 FILLER_41_1298 ();
 sg13g2_decap_8 FILLER_41_1305 ();
 sg13g2_fill_2 FILLER_41_1312 ();
 sg13g2_fill_1 FILLER_41_1314 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_4 FILLER_42_56 ();
 sg13g2_fill_1 FILLER_42_60 ();
 sg13g2_fill_2 FILLER_42_86 ();
 sg13g2_fill_1 FILLER_42_88 ();
 sg13g2_fill_1 FILLER_42_100 ();
 sg13g2_decap_8 FILLER_42_127 ();
 sg13g2_fill_2 FILLER_42_134 ();
 sg13g2_fill_2 FILLER_42_152 ();
 sg13g2_fill_1 FILLER_42_154 ();
 sg13g2_fill_1 FILLER_42_164 ();
 sg13g2_fill_1 FILLER_42_183 ();
 sg13g2_fill_2 FILLER_42_198 ();
 sg13g2_fill_1 FILLER_42_200 ();
 sg13g2_fill_2 FILLER_42_244 ();
 sg13g2_fill_1 FILLER_42_246 ();
 sg13g2_fill_2 FILLER_42_260 ();
 sg13g2_fill_1 FILLER_42_262 ();
 sg13g2_fill_2 FILLER_42_272 ();
 sg13g2_fill_2 FILLER_42_291 ();
 sg13g2_fill_2 FILLER_42_324 ();
 sg13g2_fill_1 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_358 ();
 sg13g2_decap_8 FILLER_42_365 ();
 sg13g2_decap_8 FILLER_42_372 ();
 sg13g2_fill_1 FILLER_42_382 ();
 sg13g2_fill_2 FILLER_42_416 ();
 sg13g2_fill_1 FILLER_42_486 ();
 sg13g2_fill_2 FILLER_42_492 ();
 sg13g2_decap_8 FILLER_42_499 ();
 sg13g2_fill_2 FILLER_42_506 ();
 sg13g2_fill_1 FILLER_42_508 ();
 sg13g2_fill_2 FILLER_42_532 ();
 sg13g2_decap_4 FILLER_42_560 ();
 sg13g2_fill_1 FILLER_42_583 ();
 sg13g2_decap_8 FILLER_42_633 ();
 sg13g2_fill_1 FILLER_42_640 ();
 sg13g2_decap_8 FILLER_42_663 ();
 sg13g2_fill_1 FILLER_42_670 ();
 sg13g2_decap_4 FILLER_42_675 ();
 sg13g2_fill_2 FILLER_42_679 ();
 sg13g2_fill_2 FILLER_42_698 ();
 sg13g2_fill_2 FILLER_42_726 ();
 sg13g2_fill_1 FILLER_42_728 ();
 sg13g2_fill_2 FILLER_42_742 ();
 sg13g2_fill_1 FILLER_42_744 ();
 sg13g2_decap_8 FILLER_42_761 ();
 sg13g2_decap_4 FILLER_42_768 ();
 sg13g2_fill_1 FILLER_42_772 ();
 sg13g2_fill_2 FILLER_42_799 ();
 sg13g2_decap_4 FILLER_42_809 ();
 sg13g2_fill_2 FILLER_42_836 ();
 sg13g2_fill_1 FILLER_42_891 ();
 sg13g2_fill_1 FILLER_42_931 ();
 sg13g2_fill_1 FILLER_42_981 ();
 sg13g2_decap_4 FILLER_42_1023 ();
 sg13g2_decap_8 FILLER_42_1031 ();
 sg13g2_decap_4 FILLER_42_1038 ();
 sg13g2_fill_1 FILLER_42_1042 ();
 sg13g2_fill_2 FILLER_42_1051 ();
 sg13g2_fill_1 FILLER_42_1063 ();
 sg13g2_decap_8 FILLER_42_1068 ();
 sg13g2_decap_8 FILLER_42_1075 ();
 sg13g2_fill_2 FILLER_42_1082 ();
 sg13g2_fill_1 FILLER_42_1093 ();
 sg13g2_decap_4 FILLER_42_1097 ();
 sg13g2_fill_2 FILLER_42_1101 ();
 sg13g2_decap_8 FILLER_42_1107 ();
 sg13g2_fill_2 FILLER_42_1119 ();
 sg13g2_fill_2 FILLER_42_1129 ();
 sg13g2_fill_1 FILLER_42_1167 ();
 sg13g2_decap_4 FILLER_42_1178 ();
 sg13g2_decap_8 FILLER_42_1208 ();
 sg13g2_decap_8 FILLER_42_1215 ();
 sg13g2_decap_8 FILLER_42_1222 ();
 sg13g2_decap_8 FILLER_42_1229 ();
 sg13g2_decap_8 FILLER_42_1236 ();
 sg13g2_decap_8 FILLER_42_1243 ();
 sg13g2_decap_8 FILLER_42_1250 ();
 sg13g2_decap_8 FILLER_42_1257 ();
 sg13g2_decap_8 FILLER_42_1264 ();
 sg13g2_decap_8 FILLER_42_1271 ();
 sg13g2_decap_8 FILLER_42_1278 ();
 sg13g2_decap_8 FILLER_42_1285 ();
 sg13g2_decap_8 FILLER_42_1292 ();
 sg13g2_decap_8 FILLER_42_1299 ();
 sg13g2_decap_8 FILLER_42_1306 ();
 sg13g2_fill_2 FILLER_42_1313 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_4 FILLER_43_21 ();
 sg13g2_fill_1 FILLER_43_25 ();
 sg13g2_fill_1 FILLER_43_52 ();
 sg13g2_fill_1 FILLER_43_57 ();
 sg13g2_fill_2 FILLER_43_74 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_fill_1 FILLER_43_105 ();
 sg13g2_fill_2 FILLER_43_181 ();
 sg13g2_fill_1 FILLER_43_183 ();
 sg13g2_fill_2 FILLER_43_210 ();
 sg13g2_fill_1 FILLER_43_212 ();
 sg13g2_fill_1 FILLER_43_232 ();
 sg13g2_decap_4 FILLER_43_305 ();
 sg13g2_decap_4 FILLER_43_313 ();
 sg13g2_fill_2 FILLER_43_317 ();
 sg13g2_fill_1 FILLER_43_335 ();
 sg13g2_fill_1 FILLER_43_388 ();
 sg13g2_fill_2 FILLER_43_437 ();
 sg13g2_fill_1 FILLER_43_474 ();
 sg13g2_fill_2 FILLER_43_510 ();
 sg13g2_fill_1 FILLER_43_512 ();
 sg13g2_fill_1 FILLER_43_531 ();
 sg13g2_fill_2 FILLER_43_562 ();
 sg13g2_decap_8 FILLER_43_585 ();
 sg13g2_decap_8 FILLER_43_592 ();
 sg13g2_decap_4 FILLER_43_599 ();
 sg13g2_fill_1 FILLER_43_603 ();
 sg13g2_decap_4 FILLER_43_608 ();
 sg13g2_fill_2 FILLER_43_612 ();
 sg13g2_decap_4 FILLER_43_678 ();
 sg13g2_fill_2 FILLER_43_682 ();
 sg13g2_fill_1 FILLER_43_697 ();
 sg13g2_fill_2 FILLER_43_703 ();
 sg13g2_fill_1 FILLER_43_709 ();
 sg13g2_fill_2 FILLER_43_719 ();
 sg13g2_fill_2 FILLER_43_738 ();
 sg13g2_fill_1 FILLER_43_740 ();
 sg13g2_fill_1 FILLER_43_821 ();
 sg13g2_fill_1 FILLER_43_833 ();
 sg13g2_decap_8 FILLER_43_860 ();
 sg13g2_fill_2 FILLER_43_871 ();
 sg13g2_fill_2 FILLER_43_916 ();
 sg13g2_fill_1 FILLER_43_931 ();
 sg13g2_fill_2 FILLER_43_940 ();
 sg13g2_fill_2 FILLER_43_968 ();
 sg13g2_fill_2 FILLER_43_1001 ();
 sg13g2_fill_1 FILLER_43_1003 ();
 sg13g2_fill_2 FILLER_43_1013 ();
 sg13g2_fill_1 FILLER_43_1046 ();
 sg13g2_decap_4 FILLER_43_1076 ();
 sg13g2_decap_4 FILLER_43_1173 ();
 sg13g2_fill_1 FILLER_43_1177 ();
 sg13g2_decap_8 FILLER_43_1183 ();
 sg13g2_fill_2 FILLER_43_1190 ();
 sg13g2_decap_8 FILLER_43_1201 ();
 sg13g2_decap_8 FILLER_43_1208 ();
 sg13g2_decap_8 FILLER_43_1215 ();
 sg13g2_decap_8 FILLER_43_1222 ();
 sg13g2_decap_8 FILLER_43_1229 ();
 sg13g2_decap_8 FILLER_43_1236 ();
 sg13g2_decap_8 FILLER_43_1243 ();
 sg13g2_decap_8 FILLER_43_1250 ();
 sg13g2_decap_8 FILLER_43_1257 ();
 sg13g2_decap_8 FILLER_43_1264 ();
 sg13g2_decap_8 FILLER_43_1271 ();
 sg13g2_decap_8 FILLER_43_1278 ();
 sg13g2_decap_8 FILLER_43_1285 ();
 sg13g2_decap_8 FILLER_43_1292 ();
 sg13g2_decap_8 FILLER_43_1299 ();
 sg13g2_decap_8 FILLER_43_1306 ();
 sg13g2_fill_2 FILLER_43_1313 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_fill_2 FILLER_44_35 ();
 sg13g2_fill_2 FILLER_44_41 ();
 sg13g2_fill_1 FILLER_44_48 ();
 sg13g2_fill_1 FILLER_44_80 ();
 sg13g2_fill_1 FILLER_44_91 ();
 sg13g2_fill_1 FILLER_44_127 ();
 sg13g2_fill_1 FILLER_44_142 ();
 sg13g2_fill_2 FILLER_44_210 ();
 sg13g2_fill_1 FILLER_44_220 ();
 sg13g2_decap_8 FILLER_44_226 ();
 sg13g2_decap_4 FILLER_44_233 ();
 sg13g2_fill_1 FILLER_44_247 ();
 sg13g2_decap_8 FILLER_44_252 ();
 sg13g2_fill_2 FILLER_44_259 ();
 sg13g2_decap_4 FILLER_44_310 ();
 sg13g2_fill_2 FILLER_44_314 ();
 sg13g2_fill_2 FILLER_44_341 ();
 sg13g2_fill_1 FILLER_44_343 ();
 sg13g2_fill_2 FILLER_44_397 ();
 sg13g2_fill_2 FILLER_44_412 ();
 sg13g2_fill_2 FILLER_44_423 ();
 sg13g2_fill_1 FILLER_44_425 ();
 sg13g2_decap_8 FILLER_44_478 ();
 sg13g2_decap_4 FILLER_44_485 ();
 sg13g2_fill_1 FILLER_44_498 ();
 sg13g2_fill_2 FILLER_44_545 ();
 sg13g2_fill_1 FILLER_44_572 ();
 sg13g2_fill_2 FILLER_44_580 ();
 sg13g2_fill_1 FILLER_44_582 ();
 sg13g2_fill_2 FILLER_44_614 ();
 sg13g2_fill_1 FILLER_44_616 ();
 sg13g2_fill_2 FILLER_44_652 ();
 sg13g2_fill_1 FILLER_44_659 ();
 sg13g2_fill_2 FILLER_44_669 ();
 sg13g2_fill_1 FILLER_44_671 ();
 sg13g2_decap_8 FILLER_44_677 ();
 sg13g2_decap_4 FILLER_44_684 ();
 sg13g2_fill_2 FILLER_44_688 ();
 sg13g2_fill_2 FILLER_44_694 ();
 sg13g2_fill_1 FILLER_44_696 ();
 sg13g2_decap_4 FILLER_44_723 ();
 sg13g2_fill_2 FILLER_44_727 ();
 sg13g2_fill_1 FILLER_44_769 ();
 sg13g2_fill_1 FILLER_44_790 ();
 sg13g2_fill_2 FILLER_44_795 ();
 sg13g2_fill_1 FILLER_44_814 ();
 sg13g2_fill_1 FILLER_44_820 ();
 sg13g2_decap_8 FILLER_44_829 ();
 sg13g2_decap_8 FILLER_44_836 ();
 sg13g2_fill_2 FILLER_44_843 ();
 sg13g2_decap_8 FILLER_44_849 ();
 sg13g2_fill_1 FILLER_44_856 ();
 sg13g2_decap_8 FILLER_44_862 ();
 sg13g2_decap_8 FILLER_44_869 ();
 sg13g2_fill_1 FILLER_44_876 ();
 sg13g2_fill_1 FILLER_44_886 ();
 sg13g2_fill_1 FILLER_44_892 ();
 sg13g2_fill_1 FILLER_44_911 ();
 sg13g2_fill_1 FILLER_44_927 ();
 sg13g2_fill_1 FILLER_44_936 ();
 sg13g2_fill_1 FILLER_44_945 ();
 sg13g2_decap_4 FILLER_44_977 ();
 sg13g2_fill_2 FILLER_44_999 ();
 sg13g2_fill_2 FILLER_44_1024 ();
 sg13g2_fill_1 FILLER_44_1038 ();
 sg13g2_decap_4 FILLER_44_1065 ();
 sg13g2_fill_2 FILLER_44_1104 ();
 sg13g2_fill_1 FILLER_44_1106 ();
 sg13g2_fill_1 FILLER_44_1138 ();
 sg13g2_fill_1 FILLER_44_1165 ();
 sg13g2_fill_1 FILLER_44_1192 ();
 sg13g2_decap_8 FILLER_44_1219 ();
 sg13g2_decap_8 FILLER_44_1226 ();
 sg13g2_decap_8 FILLER_44_1233 ();
 sg13g2_decap_8 FILLER_44_1240 ();
 sg13g2_decap_8 FILLER_44_1247 ();
 sg13g2_decap_8 FILLER_44_1254 ();
 sg13g2_decap_8 FILLER_44_1261 ();
 sg13g2_decap_8 FILLER_44_1268 ();
 sg13g2_decap_8 FILLER_44_1275 ();
 sg13g2_decap_8 FILLER_44_1282 ();
 sg13g2_decap_8 FILLER_44_1289 ();
 sg13g2_decap_8 FILLER_44_1296 ();
 sg13g2_decap_8 FILLER_44_1303 ();
 sg13g2_decap_4 FILLER_44_1310 ();
 sg13g2_fill_1 FILLER_44_1314 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_fill_1 FILLER_45_86 ();
 sg13g2_fill_2 FILLER_45_91 ();
 sg13g2_fill_1 FILLER_45_93 ();
 sg13g2_fill_2 FILLER_45_121 ();
 sg13g2_fill_2 FILLER_45_188 ();
 sg13g2_fill_1 FILLER_45_190 ();
 sg13g2_fill_2 FILLER_45_242 ();
 sg13g2_fill_1 FILLER_45_244 ();
 sg13g2_fill_2 FILLER_45_271 ();
 sg13g2_fill_2 FILLER_45_337 ();
 sg13g2_fill_2 FILLER_45_369 ();
 sg13g2_fill_1 FILLER_45_397 ();
 sg13g2_decap_4 FILLER_45_455 ();
 sg13g2_fill_2 FILLER_45_463 ();
 sg13g2_fill_1 FILLER_45_465 ();
 sg13g2_fill_1 FILLER_45_522 ();
 sg13g2_fill_1 FILLER_45_572 ();
 sg13g2_decap_4 FILLER_45_577 ();
 sg13g2_fill_2 FILLER_45_581 ();
 sg13g2_decap_8 FILLER_45_588 ();
 sg13g2_fill_1 FILLER_45_595 ();
 sg13g2_decap_4 FILLER_45_613 ();
 sg13g2_fill_1 FILLER_45_617 ();
 sg13g2_decap_4 FILLER_45_635 ();
 sg13g2_decap_4 FILLER_45_643 ();
 sg13g2_fill_2 FILLER_45_647 ();
 sg13g2_fill_2 FILLER_45_705 ();
 sg13g2_fill_2 FILLER_45_711 ();
 sg13g2_fill_1 FILLER_45_737 ();
 sg13g2_fill_2 FILLER_45_746 ();
 sg13g2_fill_1 FILLER_45_748 ();
 sg13g2_fill_1 FILLER_45_828 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_fill_1 FILLER_45_862 ();
 sg13g2_fill_2 FILLER_45_948 ();
 sg13g2_fill_1 FILLER_45_950 ();
 sg13g2_decap_8 FILLER_45_973 ();
 sg13g2_fill_1 FILLER_45_980 ();
 sg13g2_fill_1 FILLER_45_1064 ();
 sg13g2_fill_2 FILLER_45_1074 ();
 sg13g2_fill_1 FILLER_45_1094 ();
 sg13g2_fill_2 FILLER_45_1103 ();
 sg13g2_decap_8 FILLER_45_1139 ();
 sg13g2_decap_4 FILLER_45_1160 ();
 sg13g2_fill_2 FILLER_45_1187 ();
 sg13g2_decap_4 FILLER_45_1197 ();
 sg13g2_fill_1 FILLER_45_1201 ();
 sg13g2_decap_8 FILLER_45_1215 ();
 sg13g2_decap_8 FILLER_45_1222 ();
 sg13g2_decap_8 FILLER_45_1229 ();
 sg13g2_decap_8 FILLER_45_1236 ();
 sg13g2_decap_8 FILLER_45_1243 ();
 sg13g2_decap_8 FILLER_45_1250 ();
 sg13g2_decap_8 FILLER_45_1257 ();
 sg13g2_decap_8 FILLER_45_1264 ();
 sg13g2_decap_8 FILLER_45_1271 ();
 sg13g2_decap_8 FILLER_45_1278 ();
 sg13g2_decap_8 FILLER_45_1285 ();
 sg13g2_decap_8 FILLER_45_1292 ();
 sg13g2_decap_8 FILLER_45_1299 ();
 sg13g2_decap_8 FILLER_45_1306 ();
 sg13g2_fill_2 FILLER_45_1313 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_4 ();
 sg13g2_fill_1 FILLER_46_56 ();
 sg13g2_fill_2 FILLER_46_99 ();
 sg13g2_fill_1 FILLER_46_127 ();
 sg13g2_fill_2 FILLER_46_177 ();
 sg13g2_fill_1 FILLER_46_179 ();
 sg13g2_fill_1 FILLER_46_199 ();
 sg13g2_fill_2 FILLER_46_218 ();
 sg13g2_fill_1 FILLER_46_220 ();
 sg13g2_fill_1 FILLER_46_230 ();
 sg13g2_fill_1 FILLER_46_255 ();
 sg13g2_fill_2 FILLER_46_260 ();
 sg13g2_fill_1 FILLER_46_262 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_4 FILLER_46_308 ();
 sg13g2_fill_1 FILLER_46_312 ();
 sg13g2_fill_2 FILLER_46_317 ();
 sg13g2_fill_2 FILLER_46_324 ();
 sg13g2_fill_1 FILLER_46_326 ();
 sg13g2_fill_2 FILLER_46_337 ();
 sg13g2_fill_2 FILLER_46_352 ();
 sg13g2_fill_1 FILLER_46_380 ();
 sg13g2_fill_2 FILLER_46_395 ();
 sg13g2_fill_1 FILLER_46_397 ();
 sg13g2_fill_2 FILLER_46_449 ();
 sg13g2_fill_1 FILLER_46_461 ();
 sg13g2_decap_8 FILLER_46_466 ();
 sg13g2_decap_8 FILLER_46_473 ();
 sg13g2_decap_8 FILLER_46_511 ();
 sg13g2_fill_2 FILLER_46_527 ();
 sg13g2_fill_1 FILLER_46_569 ();
 sg13g2_fill_1 FILLER_46_589 ();
 sg13g2_fill_2 FILLER_46_616 ();
 sg13g2_fill_1 FILLER_46_631 ();
 sg13g2_decap_8 FILLER_46_645 ();
 sg13g2_fill_1 FILLER_46_652 ();
 sg13g2_fill_2 FILLER_46_658 ();
 sg13g2_fill_1 FILLER_46_660 ();
 sg13g2_fill_2 FILLER_46_664 ();
 sg13g2_fill_1 FILLER_46_666 ();
 sg13g2_fill_1 FILLER_46_689 ();
 sg13g2_fill_2 FILLER_46_707 ();
 sg13g2_fill_1 FILLER_46_709 ();
 sg13g2_fill_2 FILLER_46_728 ();
 sg13g2_fill_2 FILLER_46_756 ();
 sg13g2_fill_1 FILLER_46_758 ();
 sg13g2_fill_1 FILLER_46_768 ();
 sg13g2_fill_2 FILLER_46_783 ();
 sg13g2_fill_1 FILLER_46_785 ();
 sg13g2_fill_2 FILLER_46_795 ();
 sg13g2_fill_1 FILLER_46_802 ();
 sg13g2_fill_1 FILLER_46_834 ();
 sg13g2_decap_4 FILLER_46_839 ();
 sg13g2_fill_1 FILLER_46_843 ();
 sg13g2_fill_2 FILLER_46_852 ();
 sg13g2_fill_1 FILLER_46_859 ();
 sg13g2_fill_2 FILLER_46_873 ();
 sg13g2_fill_1 FILLER_46_881 ();
 sg13g2_decap_4 FILLER_46_981 ();
 sg13g2_fill_1 FILLER_46_985 ();
 sg13g2_fill_1 FILLER_46_1007 ();
 sg13g2_fill_2 FILLER_46_1031 ();
 sg13g2_decap_4 FILLER_46_1094 ();
 sg13g2_fill_2 FILLER_46_1124 ();
 sg13g2_fill_1 FILLER_46_1187 ();
 sg13g2_fill_1 FILLER_46_1193 ();
 sg13g2_decap_8 FILLER_46_1220 ();
 sg13g2_decap_8 FILLER_46_1227 ();
 sg13g2_decap_8 FILLER_46_1234 ();
 sg13g2_decap_8 FILLER_46_1241 ();
 sg13g2_decap_8 FILLER_46_1248 ();
 sg13g2_decap_8 FILLER_46_1255 ();
 sg13g2_decap_8 FILLER_46_1262 ();
 sg13g2_decap_8 FILLER_46_1269 ();
 sg13g2_decap_8 FILLER_46_1276 ();
 sg13g2_decap_8 FILLER_46_1283 ();
 sg13g2_decap_8 FILLER_46_1290 ();
 sg13g2_decap_8 FILLER_46_1297 ();
 sg13g2_decap_8 FILLER_46_1304 ();
 sg13g2_decap_4 FILLER_46_1311 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_7 ();
 sg13g2_fill_1 FILLER_47_40 ();
 sg13g2_fill_2 FILLER_47_48 ();
 sg13g2_fill_1 FILLER_47_77 ();
 sg13g2_fill_1 FILLER_47_111 ();
 sg13g2_fill_1 FILLER_47_121 ();
 sg13g2_fill_1 FILLER_47_152 ();
 sg13g2_fill_2 FILLER_47_171 ();
 sg13g2_fill_1 FILLER_47_173 ();
 sg13g2_fill_2 FILLER_47_223 ();
 sg13g2_fill_1 FILLER_47_250 ();
 sg13g2_fill_1 FILLER_47_308 ();
 sg13g2_fill_1 FILLER_47_333 ();
 sg13g2_fill_2 FILLER_47_403 ();
 sg13g2_fill_2 FILLER_47_423 ();
 sg13g2_fill_1 FILLER_47_425 ();
 sg13g2_fill_2 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_fill_1 FILLER_47_469 ();
 sg13g2_decap_4 FILLER_47_478 ();
 sg13g2_fill_1 FILLER_47_482 ();
 sg13g2_fill_1 FILLER_47_488 ();
 sg13g2_decap_4 FILLER_47_501 ();
 sg13g2_fill_2 FILLER_47_510 ();
 sg13g2_fill_1 FILLER_47_512 ();
 sg13g2_fill_2 FILLER_47_518 ();
 sg13g2_fill_1 FILLER_47_546 ();
 sg13g2_fill_2 FILLER_47_573 ();
 sg13g2_fill_1 FILLER_47_602 ();
 sg13g2_fill_2 FILLER_47_630 ();
 sg13g2_fill_1 FILLER_47_658 ();
 sg13g2_decap_8 FILLER_47_664 ();
 sg13g2_fill_2 FILLER_47_671 ();
 sg13g2_fill_1 FILLER_47_673 ();
 sg13g2_decap_8 FILLER_47_690 ();
 sg13g2_fill_2 FILLER_47_706 ();
 sg13g2_fill_1 FILLER_47_708 ();
 sg13g2_fill_1 FILLER_47_714 ();
 sg13g2_decap_8 FILLER_47_732 ();
 sg13g2_fill_1 FILLER_47_755 ();
 sg13g2_fill_2 FILLER_47_851 ();
 sg13g2_fill_1 FILLER_47_853 ();
 sg13g2_fill_2 FILLER_47_938 ();
 sg13g2_fill_1 FILLER_47_950 ();
 sg13g2_fill_1 FILLER_47_969 ();
 sg13g2_fill_2 FILLER_47_975 ();
 sg13g2_fill_1 FILLER_47_981 ();
 sg13g2_fill_1 FILLER_47_996 ();
 sg13g2_fill_2 FILLER_47_1001 ();
 sg13g2_fill_1 FILLER_47_1013 ();
 sg13g2_fill_2 FILLER_47_1022 ();
 sg13g2_fill_2 FILLER_47_1115 ();
 sg13g2_fill_2 FILLER_47_1122 ();
 sg13g2_decap_8 FILLER_47_1149 ();
 sg13g2_fill_1 FILLER_47_1156 ();
 sg13g2_fill_2 FILLER_47_1165 ();
 sg13g2_fill_1 FILLER_47_1167 ();
 sg13g2_fill_2 FILLER_47_1191 ();
 sg13g2_fill_2 FILLER_47_1198 ();
 sg13g2_decap_8 FILLER_47_1213 ();
 sg13g2_decap_8 FILLER_47_1220 ();
 sg13g2_decap_8 FILLER_47_1227 ();
 sg13g2_decap_8 FILLER_47_1234 ();
 sg13g2_decap_8 FILLER_47_1241 ();
 sg13g2_decap_8 FILLER_47_1248 ();
 sg13g2_decap_8 FILLER_47_1255 ();
 sg13g2_decap_8 FILLER_47_1262 ();
 sg13g2_decap_8 FILLER_47_1269 ();
 sg13g2_decap_8 FILLER_47_1276 ();
 sg13g2_decap_8 FILLER_47_1283 ();
 sg13g2_decap_8 FILLER_47_1290 ();
 sg13g2_decap_8 FILLER_47_1297 ();
 sg13g2_decap_8 FILLER_47_1304 ();
 sg13g2_decap_4 FILLER_47_1311 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_28 ();
 sg13g2_fill_1 FILLER_48_30 ();
 sg13g2_fill_2 FILLER_48_45 ();
 sg13g2_fill_2 FILLER_48_51 ();
 sg13g2_fill_2 FILLER_48_61 ();
 sg13g2_fill_1 FILLER_48_63 ();
 sg13g2_fill_2 FILLER_48_130 ();
 sg13g2_fill_2 FILLER_48_195 ();
 sg13g2_fill_2 FILLER_48_206 ();
 sg13g2_fill_1 FILLER_48_221 ();
 sg13g2_fill_1 FILLER_48_266 ();
 sg13g2_fill_2 FILLER_48_289 ();
 sg13g2_fill_1 FILLER_48_291 ();
 sg13g2_fill_2 FILLER_48_346 ();
 sg13g2_fill_1 FILLER_48_385 ();
 sg13g2_fill_1 FILLER_48_400 ();
 sg13g2_fill_1 FILLER_48_406 ();
 sg13g2_fill_2 FILLER_48_415 ();
 sg13g2_fill_1 FILLER_48_422 ();
 sg13g2_fill_2 FILLER_48_432 ();
 sg13g2_fill_2 FILLER_48_474 ();
 sg13g2_fill_2 FILLER_48_500 ();
 sg13g2_fill_1 FILLER_48_502 ();
 sg13g2_fill_2 FILLER_48_563 ();
 sg13g2_decap_4 FILLER_48_589 ();
 sg13g2_fill_2 FILLER_48_593 ();
 sg13g2_fill_2 FILLER_48_630 ();
 sg13g2_fill_2 FILLER_48_641 ();
 sg13g2_decap_4 FILLER_48_651 ();
 sg13g2_decap_4 FILLER_48_691 ();
 sg13g2_fill_1 FILLER_48_695 ();
 sg13g2_decap_4 FILLER_48_701 ();
 sg13g2_decap_8 FILLER_48_727 ();
 sg13g2_decap_8 FILLER_48_738 ();
 sg13g2_decap_4 FILLER_48_745 ();
 sg13g2_fill_2 FILLER_48_749 ();
 sg13g2_fill_2 FILLER_48_765 ();
 sg13g2_fill_1 FILLER_48_767 ();
 sg13g2_fill_2 FILLER_48_777 ();
 sg13g2_fill_1 FILLER_48_779 ();
 sg13g2_fill_2 FILLER_48_789 ();
 sg13g2_decap_4 FILLER_48_795 ();
 sg13g2_fill_1 FILLER_48_799 ();
 sg13g2_fill_1 FILLER_48_805 ();
 sg13g2_fill_2 FILLER_48_810 ();
 sg13g2_fill_1 FILLER_48_812 ();
 sg13g2_fill_2 FILLER_48_853 ();
 sg13g2_fill_1 FILLER_48_855 ();
 sg13g2_fill_2 FILLER_48_861 ();
 sg13g2_fill_1 FILLER_48_863 ();
 sg13g2_fill_1 FILLER_48_883 ();
 sg13g2_fill_2 FILLER_48_936 ();
 sg13g2_fill_1 FILLER_48_951 ();
 sg13g2_fill_2 FILLER_48_1047 ();
 sg13g2_fill_2 FILLER_48_1054 ();
 sg13g2_fill_1 FILLER_48_1079 ();
 sg13g2_fill_1 FILLER_48_1115 ();
 sg13g2_fill_1 FILLER_48_1125 ();
 sg13g2_fill_2 FILLER_48_1131 ();
 sg13g2_fill_2 FILLER_48_1181 ();
 sg13g2_decap_8 FILLER_48_1212 ();
 sg13g2_decap_8 FILLER_48_1219 ();
 sg13g2_decap_8 FILLER_48_1226 ();
 sg13g2_decap_8 FILLER_48_1233 ();
 sg13g2_decap_8 FILLER_48_1240 ();
 sg13g2_decap_8 FILLER_48_1247 ();
 sg13g2_decap_8 FILLER_48_1254 ();
 sg13g2_decap_8 FILLER_48_1261 ();
 sg13g2_decap_8 FILLER_48_1268 ();
 sg13g2_decap_8 FILLER_48_1275 ();
 sg13g2_decap_8 FILLER_48_1282 ();
 sg13g2_decap_8 FILLER_48_1289 ();
 sg13g2_decap_8 FILLER_48_1296 ();
 sg13g2_decap_8 FILLER_48_1303 ();
 sg13g2_decap_4 FILLER_48_1310 ();
 sg13g2_fill_1 FILLER_48_1314 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_4 FILLER_49_7 ();
 sg13g2_fill_2 FILLER_49_11 ();
 sg13g2_decap_8 FILLER_49_17 ();
 sg13g2_fill_2 FILLER_49_38 ();
 sg13g2_fill_2 FILLER_49_44 ();
 sg13g2_fill_1 FILLER_49_51 ();
 sg13g2_fill_2 FILLER_49_56 ();
 sg13g2_fill_1 FILLER_49_115 ();
 sg13g2_fill_2 FILLER_49_156 ();
 sg13g2_fill_1 FILLER_49_176 ();
 sg13g2_fill_2 FILLER_49_229 ();
 sg13g2_fill_2 FILLER_49_248 ();
 sg13g2_fill_1 FILLER_49_250 ();
 sg13g2_decap_4 FILLER_49_269 ();
 sg13g2_fill_1 FILLER_49_273 ();
 sg13g2_fill_1 FILLER_49_331 ();
 sg13g2_fill_1 FILLER_49_362 ();
 sg13g2_fill_2 FILLER_49_386 ();
 sg13g2_fill_1 FILLER_49_388 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_fill_2 FILLER_49_431 ();
 sg13g2_fill_1 FILLER_49_433 ();
 sg13g2_fill_1 FILLER_49_439 ();
 sg13g2_fill_2 FILLER_49_449 ();
 sg13g2_fill_1 FILLER_49_470 ();
 sg13g2_decap_4 FILLER_49_480 ();
 sg13g2_decap_4 FILLER_49_492 ();
 sg13g2_fill_2 FILLER_49_496 ();
 sg13g2_fill_2 FILLER_49_512 ();
 sg13g2_fill_2 FILLER_49_542 ();
 sg13g2_fill_1 FILLER_49_544 ();
 sg13g2_fill_2 FILLER_49_576 ();
 sg13g2_fill_2 FILLER_49_639 ();
 sg13g2_decap_8 FILLER_49_661 ();
 sg13g2_decap_8 FILLER_49_668 ();
 sg13g2_fill_1 FILLER_49_675 ();
 sg13g2_fill_2 FILLER_49_701 ();
 sg13g2_fill_1 FILLER_49_703 ();
 sg13g2_fill_1 FILLER_49_723 ();
 sg13g2_decap_8 FILLER_49_750 ();
 sg13g2_fill_2 FILLER_49_757 ();
 sg13g2_fill_1 FILLER_49_776 ();
 sg13g2_fill_2 FILLER_49_808 ();
 sg13g2_fill_1 FILLER_49_819 ();
 sg13g2_fill_2 FILLER_49_870 ();
 sg13g2_fill_2 FILLER_49_903 ();
 sg13g2_fill_1 FILLER_49_905 ();
 sg13g2_fill_2 FILLER_49_911 ();
 sg13g2_fill_2 FILLER_49_923 ();
 sg13g2_fill_1 FILLER_49_950 ();
 sg13g2_fill_1 FILLER_49_990 ();
 sg13g2_fill_1 FILLER_49_1045 ();
 sg13g2_fill_1 FILLER_49_1055 ();
 sg13g2_fill_1 FILLER_49_1143 ();
 sg13g2_fill_2 FILLER_49_1148 ();
 sg13g2_fill_1 FILLER_49_1150 ();
 sg13g2_decap_8 FILLER_49_1210 ();
 sg13g2_decap_8 FILLER_49_1217 ();
 sg13g2_decap_8 FILLER_49_1224 ();
 sg13g2_decap_8 FILLER_49_1231 ();
 sg13g2_decap_8 FILLER_49_1238 ();
 sg13g2_decap_8 FILLER_49_1245 ();
 sg13g2_decap_8 FILLER_49_1252 ();
 sg13g2_decap_8 FILLER_49_1259 ();
 sg13g2_decap_8 FILLER_49_1266 ();
 sg13g2_decap_8 FILLER_49_1273 ();
 sg13g2_decap_8 FILLER_49_1280 ();
 sg13g2_decap_8 FILLER_49_1287 ();
 sg13g2_decap_8 FILLER_49_1294 ();
 sg13g2_decap_8 FILLER_49_1301 ();
 sg13g2_decap_8 FILLER_49_1308 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_28 ();
 sg13g2_fill_1 FILLER_50_30 ();
 sg13g2_decap_4 FILLER_50_60 ();
 sg13g2_fill_1 FILLER_50_64 ();
 sg13g2_fill_1 FILLER_50_93 ();
 sg13g2_fill_1 FILLER_50_125 ();
 sg13g2_fill_2 FILLER_50_140 ();
 sg13g2_fill_2 FILLER_50_147 ();
 sg13g2_fill_1 FILLER_50_149 ();
 sg13g2_fill_2 FILLER_50_192 ();
 sg13g2_fill_1 FILLER_50_194 ();
 sg13g2_decap_8 FILLER_50_285 ();
 sg13g2_fill_2 FILLER_50_292 ();
 sg13g2_decap_8 FILLER_50_298 ();
 sg13g2_decap_8 FILLER_50_305 ();
 sg13g2_fill_2 FILLER_50_312 ();
 sg13g2_fill_1 FILLER_50_314 ();
 sg13g2_fill_2 FILLER_50_318 ();
 sg13g2_fill_2 FILLER_50_325 ();
 sg13g2_fill_1 FILLER_50_327 ();
 sg13g2_fill_2 FILLER_50_332 ();
 sg13g2_fill_1 FILLER_50_334 ();
 sg13g2_fill_1 FILLER_50_416 ();
 sg13g2_fill_1 FILLER_50_457 ();
 sg13g2_fill_2 FILLER_50_497 ();
 sg13g2_fill_1 FILLER_50_560 ();
 sg13g2_decap_8 FILLER_50_565 ();
 sg13g2_fill_2 FILLER_50_572 ();
 sg13g2_fill_1 FILLER_50_574 ();
 sg13g2_fill_1 FILLER_50_649 ();
 sg13g2_fill_2 FILLER_50_665 ();
 sg13g2_fill_1 FILLER_50_667 ();
 sg13g2_decap_4 FILLER_50_682 ();
 sg13g2_fill_2 FILLER_50_721 ();
 sg13g2_decap_4 FILLER_50_731 ();
 sg13g2_fill_2 FILLER_50_771 ();
 sg13g2_fill_1 FILLER_50_786 ();
 sg13g2_decap_8 FILLER_50_791 ();
 sg13g2_fill_2 FILLER_50_798 ();
 sg13g2_fill_1 FILLER_50_843 ();
 sg13g2_fill_2 FILLER_50_871 ();
 sg13g2_fill_1 FILLER_50_882 ();
 sg13g2_decap_8 FILLER_50_899 ();
 sg13g2_decap_8 FILLER_50_906 ();
 sg13g2_decap_4 FILLER_50_957 ();
 sg13g2_decap_4 FILLER_50_965 ();
 sg13g2_fill_2 FILLER_50_981 ();
 sg13g2_fill_2 FILLER_50_1070 ();
 sg13g2_fill_2 FILLER_50_1158 ();
 sg13g2_fill_1 FILLER_50_1165 ();
 sg13g2_decap_8 FILLER_50_1214 ();
 sg13g2_decap_8 FILLER_50_1221 ();
 sg13g2_decap_8 FILLER_50_1228 ();
 sg13g2_decap_8 FILLER_50_1235 ();
 sg13g2_decap_8 FILLER_50_1242 ();
 sg13g2_decap_8 FILLER_50_1249 ();
 sg13g2_decap_8 FILLER_50_1256 ();
 sg13g2_decap_8 FILLER_50_1263 ();
 sg13g2_decap_8 FILLER_50_1270 ();
 sg13g2_decap_8 FILLER_50_1277 ();
 sg13g2_decap_8 FILLER_50_1284 ();
 sg13g2_decap_8 FILLER_50_1291 ();
 sg13g2_decap_8 FILLER_50_1298 ();
 sg13g2_decap_8 FILLER_50_1305 ();
 sg13g2_fill_2 FILLER_50_1312 ();
 sg13g2_fill_1 FILLER_50_1314 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_7 ();
 sg13g2_fill_1 FILLER_51_11 ();
 sg13g2_decap_4 FILLER_51_25 ();
 sg13g2_fill_1 FILLER_51_42 ();
 sg13g2_fill_2 FILLER_51_73 ();
 sg13g2_fill_2 FILLER_51_80 ();
 sg13g2_fill_1 FILLER_51_82 ();
 sg13g2_fill_1 FILLER_51_105 ();
 sg13g2_fill_2 FILLER_51_155 ();
 sg13g2_fill_1 FILLER_51_191 ();
 sg13g2_fill_1 FILLER_51_218 ();
 sg13g2_fill_1 FILLER_51_231 ();
 sg13g2_decap_4 FILLER_51_244 ();
 sg13g2_fill_2 FILLER_51_248 ();
 sg13g2_decap_8 FILLER_51_254 ();
 sg13g2_fill_2 FILLER_51_261 ();
 sg13g2_fill_1 FILLER_51_312 ();
 sg13g2_decap_8 FILLER_51_337 ();
 sg13g2_fill_2 FILLER_51_344 ();
 sg13g2_fill_1 FILLER_51_377 ();
 sg13g2_fill_2 FILLER_51_381 ();
 sg13g2_fill_1 FILLER_51_387 ();
 sg13g2_fill_2 FILLER_51_411 ();
 sg13g2_fill_1 FILLER_51_413 ();
 sg13g2_decap_8 FILLER_51_423 ();
 sg13g2_fill_2 FILLER_51_496 ();
 sg13g2_fill_1 FILLER_51_498 ();
 sg13g2_fill_1 FILLER_51_534 ();
 sg13g2_fill_2 FILLER_51_558 ();
 sg13g2_fill_1 FILLER_51_560 ();
 sg13g2_decap_4 FILLER_51_566 ();
 sg13g2_fill_2 FILLER_51_577 ();
 sg13g2_fill_1 FILLER_51_579 ();
 sg13g2_fill_2 FILLER_51_584 ();
 sg13g2_fill_1 FILLER_51_586 ();
 sg13g2_fill_1 FILLER_51_594 ();
 sg13g2_fill_2 FILLER_51_626 ();
 sg13g2_fill_1 FILLER_51_628 ();
 sg13g2_decap_4 FILLER_51_642 ();
 sg13g2_fill_1 FILLER_51_646 ();
 sg13g2_fill_2 FILLER_51_665 ();
 sg13g2_fill_1 FILLER_51_719 ();
 sg13g2_fill_2 FILLER_51_728 ();
 sg13g2_fill_1 FILLER_51_730 ();
 sg13g2_fill_2 FILLER_51_762 ();
 sg13g2_fill_1 FILLER_51_764 ();
 sg13g2_decap_8 FILLER_51_791 ();
 sg13g2_decap_4 FILLER_51_798 ();
 sg13g2_fill_2 FILLER_51_807 ();
 sg13g2_fill_1 FILLER_51_809 ();
 sg13g2_fill_2 FILLER_51_814 ();
 sg13g2_fill_1 FILLER_51_821 ();
 sg13g2_fill_1 FILLER_51_834 ();
 sg13g2_fill_2 FILLER_51_879 ();
 sg13g2_fill_2 FILLER_51_999 ();
 sg13g2_fill_2 FILLER_51_1032 ();
 sg13g2_fill_1 FILLER_51_1054 ();
 sg13g2_fill_2 FILLER_51_1109 ();
 sg13g2_fill_1 FILLER_51_1151 ();
 sg13g2_fill_2 FILLER_51_1173 ();
 sg13g2_fill_1 FILLER_51_1175 ();
 sg13g2_decap_4 FILLER_51_1184 ();
 sg13g2_fill_2 FILLER_51_1188 ();
 sg13g2_decap_8 FILLER_51_1194 ();
 sg13g2_decap_8 FILLER_51_1201 ();
 sg13g2_decap_8 FILLER_51_1208 ();
 sg13g2_decap_8 FILLER_51_1215 ();
 sg13g2_decap_8 FILLER_51_1222 ();
 sg13g2_decap_8 FILLER_51_1229 ();
 sg13g2_decap_8 FILLER_51_1236 ();
 sg13g2_decap_8 FILLER_51_1243 ();
 sg13g2_decap_8 FILLER_51_1250 ();
 sg13g2_decap_8 FILLER_51_1257 ();
 sg13g2_decap_8 FILLER_51_1264 ();
 sg13g2_decap_8 FILLER_51_1271 ();
 sg13g2_decap_8 FILLER_51_1278 ();
 sg13g2_decap_8 FILLER_51_1285 ();
 sg13g2_decap_8 FILLER_51_1292 ();
 sg13g2_decap_8 FILLER_51_1299 ();
 sg13g2_decap_8 FILLER_51_1306 ();
 sg13g2_fill_2 FILLER_51_1313 ();
 sg13g2_fill_1 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_40 ();
 sg13g2_fill_2 FILLER_52_97 ();
 sg13g2_fill_1 FILLER_52_134 ();
 sg13g2_fill_2 FILLER_52_200 ();
 sg13g2_fill_1 FILLER_52_202 ();
 sg13g2_fill_1 FILLER_52_216 ();
 sg13g2_fill_2 FILLER_52_231 ();
 sg13g2_fill_1 FILLER_52_233 ();
 sg13g2_decap_8 FILLER_52_248 ();
 sg13g2_decap_4 FILLER_52_255 ();
 sg13g2_fill_2 FILLER_52_270 ();
 sg13g2_fill_1 FILLER_52_272 ();
 sg13g2_fill_2 FILLER_52_328 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_fill_1 FILLER_52_463 ();
 sg13g2_fill_2 FILLER_52_482 ();
 sg13g2_decap_4 FILLER_52_489 ();
 sg13g2_fill_1 FILLER_52_550 ();
 sg13g2_fill_2 FILLER_52_559 ();
 sg13g2_fill_1 FILLER_52_561 ();
 sg13g2_fill_1 FILLER_52_602 ();
 sg13g2_fill_2 FILLER_52_617 ();
 sg13g2_fill_2 FILLER_52_628 ();
 sg13g2_fill_2 FILLER_52_644 ();
 sg13g2_fill_1 FILLER_52_646 ();
 sg13g2_decap_4 FILLER_52_659 ();
 sg13g2_fill_1 FILLER_52_663 ();
 sg13g2_decap_4 FILLER_52_677 ();
 sg13g2_fill_2 FILLER_52_724 ();
 sg13g2_fill_1 FILLER_52_726 ();
 sg13g2_fill_1 FILLER_52_737 ();
 sg13g2_fill_2 FILLER_52_747 ();
 sg13g2_fill_1 FILLER_52_757 ();
 sg13g2_fill_1 FILLER_52_768 ();
 sg13g2_fill_1 FILLER_52_829 ();
 sg13g2_fill_2 FILLER_52_838 ();
 sg13g2_fill_1 FILLER_52_840 ();
 sg13g2_fill_2 FILLER_52_867 ();
 sg13g2_fill_2 FILLER_52_874 ();
 sg13g2_decap_4 FILLER_52_892 ();
 sg13g2_fill_1 FILLER_52_896 ();
 sg13g2_decap_8 FILLER_52_901 ();
 sg13g2_fill_1 FILLER_52_908 ();
 sg13g2_decap_8 FILLER_52_951 ();
 sg13g2_decap_8 FILLER_52_958 ();
 sg13g2_fill_1 FILLER_52_977 ();
 sg13g2_fill_2 FILLER_52_1001 ();
 sg13g2_fill_1 FILLER_52_1041 ();
 sg13g2_fill_2 FILLER_52_1051 ();
 sg13g2_fill_2 FILLER_52_1084 ();
 sg13g2_fill_1 FILLER_52_1121 ();
 sg13g2_fill_2 FILLER_52_1148 ();
 sg13g2_fill_1 FILLER_52_1150 ();
 sg13g2_fill_2 FILLER_52_1162 ();
 sg13g2_fill_1 FILLER_52_1164 ();
 sg13g2_decap_8 FILLER_52_1195 ();
 sg13g2_decap_8 FILLER_52_1202 ();
 sg13g2_decap_8 FILLER_52_1209 ();
 sg13g2_decap_8 FILLER_52_1216 ();
 sg13g2_decap_8 FILLER_52_1223 ();
 sg13g2_decap_8 FILLER_52_1230 ();
 sg13g2_decap_8 FILLER_52_1237 ();
 sg13g2_decap_8 FILLER_52_1244 ();
 sg13g2_decap_8 FILLER_52_1251 ();
 sg13g2_decap_8 FILLER_52_1258 ();
 sg13g2_decap_8 FILLER_52_1265 ();
 sg13g2_decap_8 FILLER_52_1272 ();
 sg13g2_decap_8 FILLER_52_1279 ();
 sg13g2_decap_8 FILLER_52_1286 ();
 sg13g2_decap_8 FILLER_52_1293 ();
 sg13g2_decap_8 FILLER_52_1300 ();
 sg13g2_decap_8 FILLER_52_1307 ();
 sg13g2_fill_1 FILLER_52_1314 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_9 ();
 sg13g2_fill_2 FILLER_53_23 ();
 sg13g2_fill_2 FILLER_53_45 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_fill_1 FILLER_53_63 ();
 sg13g2_fill_1 FILLER_53_74 ();
 sg13g2_fill_2 FILLER_53_80 ();
 sg13g2_fill_1 FILLER_53_82 ();
 sg13g2_decap_4 FILLER_53_100 ();
 sg13g2_fill_2 FILLER_53_104 ();
 sg13g2_fill_2 FILLER_53_114 ();
 sg13g2_fill_1 FILLER_53_116 ();
 sg13g2_fill_2 FILLER_53_147 ();
 sg13g2_fill_1 FILLER_53_180 ();
 sg13g2_fill_2 FILLER_53_298 ();
 sg13g2_fill_2 FILLER_53_316 ();
 sg13g2_fill_1 FILLER_53_318 ();
 sg13g2_fill_1 FILLER_53_331 ();
 sg13g2_fill_2 FILLER_53_336 ();
 sg13g2_fill_2 FILLER_53_346 ();
 sg13g2_fill_2 FILLER_53_367 ();
 sg13g2_fill_2 FILLER_53_404 ();
 sg13g2_decap_4 FILLER_53_419 ();
 sg13g2_fill_2 FILLER_53_423 ();
 sg13g2_decap_4 FILLER_53_429 ();
 sg13g2_fill_2 FILLER_53_433 ();
 sg13g2_fill_1 FILLER_53_448 ();
 sg13g2_fill_1 FILLER_53_478 ();
 sg13g2_fill_2 FILLER_53_494 ();
 sg13g2_fill_1 FILLER_53_496 ();
 sg13g2_fill_2 FILLER_53_511 ();
 sg13g2_fill_1 FILLER_53_559 ();
 sg13g2_fill_2 FILLER_53_584 ();
 sg13g2_fill_1 FILLER_53_683 ();
 sg13g2_fill_2 FILLER_53_716 ();
 sg13g2_fill_1 FILLER_53_718 ();
 sg13g2_fill_1 FILLER_53_736 ();
 sg13g2_fill_1 FILLER_53_768 ();
 sg13g2_decap_4 FILLER_53_796 ();
 sg13g2_fill_2 FILLER_53_800 ();
 sg13g2_decap_8 FILLER_53_806 ();
 sg13g2_fill_2 FILLER_53_813 ();
 sg13g2_fill_1 FILLER_53_839 ();
 sg13g2_fill_1 FILLER_53_895 ();
 sg13g2_fill_1 FILLER_53_922 ();
 sg13g2_fill_2 FILLER_53_974 ();
 sg13g2_fill_1 FILLER_53_994 ();
 sg13g2_fill_2 FILLER_53_1087 ();
 sg13g2_fill_1 FILLER_53_1089 ();
 sg13g2_fill_2 FILLER_53_1093 ();
 sg13g2_fill_1 FILLER_53_1095 ();
 sg13g2_fill_2 FILLER_53_1185 ();
 sg13g2_decap_8 FILLER_53_1200 ();
 sg13g2_decap_8 FILLER_53_1207 ();
 sg13g2_decap_8 FILLER_53_1214 ();
 sg13g2_decap_8 FILLER_53_1221 ();
 sg13g2_decap_8 FILLER_53_1228 ();
 sg13g2_decap_8 FILLER_53_1235 ();
 sg13g2_decap_8 FILLER_53_1242 ();
 sg13g2_decap_8 FILLER_53_1249 ();
 sg13g2_decap_8 FILLER_53_1256 ();
 sg13g2_decap_8 FILLER_53_1263 ();
 sg13g2_decap_8 FILLER_53_1270 ();
 sg13g2_decap_8 FILLER_53_1277 ();
 sg13g2_decap_8 FILLER_53_1284 ();
 sg13g2_decap_8 FILLER_53_1291 ();
 sg13g2_decap_8 FILLER_53_1298 ();
 sg13g2_decap_8 FILLER_53_1305 ();
 sg13g2_fill_2 FILLER_53_1312 ();
 sg13g2_fill_1 FILLER_53_1314 ();
 sg13g2_fill_2 FILLER_54_26 ();
 sg13g2_fill_2 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_69 ();
 sg13g2_fill_1 FILLER_54_76 ();
 sg13g2_fill_2 FILLER_54_125 ();
 sg13g2_fill_1 FILLER_54_127 ();
 sg13g2_fill_2 FILLER_54_221 ();
 sg13g2_fill_1 FILLER_54_223 ();
 sg13g2_decap_8 FILLER_54_242 ();
 sg13g2_decap_8 FILLER_54_249 ();
 sg13g2_fill_2 FILLER_54_256 ();
 sg13g2_fill_1 FILLER_54_258 ();
 sg13g2_fill_2 FILLER_54_265 ();
 sg13g2_fill_2 FILLER_54_279 ();
 sg13g2_fill_1 FILLER_54_281 ();
 sg13g2_fill_1 FILLER_54_308 ();
 sg13g2_fill_2 FILLER_54_375 ();
 sg13g2_fill_1 FILLER_54_377 ();
 sg13g2_fill_2 FILLER_54_383 ();
 sg13g2_fill_2 FILLER_54_394 ();
 sg13g2_fill_2 FILLER_54_401 ();
 sg13g2_fill_1 FILLER_54_422 ();
 sg13g2_fill_2 FILLER_54_448 ();
 sg13g2_fill_1 FILLER_54_454 ();
 sg13g2_fill_1 FILLER_54_467 ();
 sg13g2_fill_2 FILLER_54_472 ();
 sg13g2_fill_1 FILLER_54_474 ();
 sg13g2_fill_1 FILLER_54_489 ();
 sg13g2_fill_2 FILLER_54_595 ();
 sg13g2_decap_4 FILLER_54_602 ();
 sg13g2_fill_1 FILLER_54_606 ();
 sg13g2_fill_2 FILLER_54_615 ();
 sg13g2_decap_4 FILLER_54_622 ();
 sg13g2_fill_2 FILLER_54_626 ();
 sg13g2_fill_1 FILLER_54_642 ();
 sg13g2_decap_8 FILLER_54_665 ();
 sg13g2_fill_2 FILLER_54_672 ();
 sg13g2_fill_1 FILLER_54_674 ();
 sg13g2_fill_1 FILLER_54_706 ();
 sg13g2_fill_1 FILLER_54_726 ();
 sg13g2_fill_2 FILLER_54_740 ();
 sg13g2_fill_1 FILLER_54_742 ();
 sg13g2_fill_2 FILLER_54_757 ();
 sg13g2_fill_2 FILLER_54_849 ();
 sg13g2_fill_2 FILLER_54_855 ();
 sg13g2_fill_1 FILLER_54_865 ();
 sg13g2_decap_8 FILLER_54_888 ();
 sg13g2_fill_1 FILLER_54_895 ();
 sg13g2_fill_1 FILLER_54_918 ();
 sg13g2_fill_1 FILLER_54_945 ();
 sg13g2_decap_4 FILLER_54_951 ();
 sg13g2_fill_1 FILLER_54_955 ();
 sg13g2_fill_2 FILLER_54_1063 ();
 sg13g2_fill_2 FILLER_54_1170 ();
 sg13g2_fill_1 FILLER_54_1172 ();
 sg13g2_decap_8 FILLER_54_1199 ();
 sg13g2_decap_8 FILLER_54_1206 ();
 sg13g2_decap_8 FILLER_54_1213 ();
 sg13g2_decap_8 FILLER_54_1220 ();
 sg13g2_decap_8 FILLER_54_1227 ();
 sg13g2_decap_8 FILLER_54_1234 ();
 sg13g2_decap_8 FILLER_54_1241 ();
 sg13g2_decap_8 FILLER_54_1248 ();
 sg13g2_decap_8 FILLER_54_1255 ();
 sg13g2_decap_8 FILLER_54_1262 ();
 sg13g2_decap_8 FILLER_54_1269 ();
 sg13g2_decap_8 FILLER_54_1276 ();
 sg13g2_decap_8 FILLER_54_1283 ();
 sg13g2_decap_8 FILLER_54_1290 ();
 sg13g2_decap_8 FILLER_54_1297 ();
 sg13g2_decap_8 FILLER_54_1304 ();
 sg13g2_decap_4 FILLER_54_1311 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_28 ();
 sg13g2_fill_1 FILLER_55_33 ();
 sg13g2_fill_2 FILLER_55_80 ();
 sg13g2_fill_1 FILLER_55_108 ();
 sg13g2_fill_2 FILLER_55_149 ();
 sg13g2_fill_1 FILLER_55_151 ();
 sg13g2_fill_2 FILLER_55_182 ();
 sg13g2_fill_2 FILLER_55_235 ();
 sg13g2_fill_1 FILLER_55_263 ();
 sg13g2_decap_8 FILLER_55_285 ();
 sg13g2_decap_4 FILLER_55_296 ();
 sg13g2_fill_2 FILLER_55_418 ();
 sg13g2_fill_2 FILLER_55_428 ();
 sg13g2_decap_8 FILLER_55_482 ();
 sg13g2_decap_4 FILLER_55_489 ();
 sg13g2_fill_2 FILLER_55_503 ();
 sg13g2_fill_2 FILLER_55_513 ();
 sg13g2_fill_1 FILLER_55_530 ();
 sg13g2_decap_8 FILLER_55_548 ();
 sg13g2_fill_2 FILLER_55_559 ();
 sg13g2_fill_1 FILLER_55_561 ();
 sg13g2_fill_1 FILLER_55_580 ();
 sg13g2_decap_4 FILLER_55_607 ();
 sg13g2_fill_2 FILLER_55_645 ();
 sg13g2_fill_2 FILLER_55_673 ();
 sg13g2_decap_8 FILLER_55_680 ();
 sg13g2_fill_1 FILLER_55_687 ();
 sg13g2_fill_1 FILLER_55_701 ();
 sg13g2_fill_1 FILLER_55_715 ();
 sg13g2_fill_1 FILLER_55_733 ();
 sg13g2_fill_2 FILLER_55_739 ();
 sg13g2_fill_1 FILLER_55_741 ();
 sg13g2_fill_1 FILLER_55_796 ();
 sg13g2_fill_2 FILLER_55_806 ();
 sg13g2_fill_2 FILLER_55_835 ();
 sg13g2_fill_1 FILLER_55_837 ();
 sg13g2_fill_2 FILLER_55_851 ();
 sg13g2_decap_4 FILLER_55_858 ();
 sg13g2_fill_1 FILLER_55_862 ();
 sg13g2_fill_2 FILLER_55_867 ();
 sg13g2_fill_1 FILLER_55_869 ();
 sg13g2_fill_1 FILLER_55_922 ();
 sg13g2_fill_1 FILLER_55_951 ();
 sg13g2_fill_2 FILLER_55_959 ();
 sg13g2_fill_2 FILLER_55_978 ();
 sg13g2_fill_1 FILLER_55_980 ();
 sg13g2_fill_1 FILLER_55_990 ();
 sg13g2_fill_1 FILLER_55_1022 ();
 sg13g2_fill_1 FILLER_55_1070 ();
 sg13g2_fill_2 FILLER_55_1088 ();
 sg13g2_fill_1 FILLER_55_1090 ();
 sg13g2_fill_1 FILLER_55_1101 ();
 sg13g2_fill_1 FILLER_55_1128 ();
 sg13g2_fill_2 FILLER_55_1157 ();
 sg13g2_fill_1 FILLER_55_1159 ();
 sg13g2_fill_2 FILLER_55_1170 ();
 sg13g2_fill_2 FILLER_55_1185 ();
 sg13g2_decap_8 FILLER_55_1204 ();
 sg13g2_decap_8 FILLER_55_1211 ();
 sg13g2_decap_8 FILLER_55_1218 ();
 sg13g2_decap_8 FILLER_55_1225 ();
 sg13g2_decap_8 FILLER_55_1232 ();
 sg13g2_decap_8 FILLER_55_1239 ();
 sg13g2_decap_8 FILLER_55_1246 ();
 sg13g2_decap_8 FILLER_55_1253 ();
 sg13g2_decap_8 FILLER_55_1260 ();
 sg13g2_decap_8 FILLER_55_1267 ();
 sg13g2_decap_8 FILLER_55_1274 ();
 sg13g2_decap_8 FILLER_55_1281 ();
 sg13g2_decap_8 FILLER_55_1288 ();
 sg13g2_decap_8 FILLER_55_1295 ();
 sg13g2_decap_8 FILLER_55_1302 ();
 sg13g2_decap_4 FILLER_55_1309 ();
 sg13g2_fill_2 FILLER_55_1313 ();
 sg13g2_decap_8 FILLER_56_31 ();
 sg13g2_fill_1 FILLER_56_38 ();
 sg13g2_fill_1 FILLER_56_44 ();
 sg13g2_fill_1 FILLER_56_62 ();
 sg13g2_fill_1 FILLER_56_93 ();
 sg13g2_fill_2 FILLER_56_195 ();
 sg13g2_fill_1 FILLER_56_197 ();
 sg13g2_fill_1 FILLER_56_230 ();
 sg13g2_fill_2 FILLER_56_244 ();
 sg13g2_fill_1 FILLER_56_246 ();
 sg13g2_fill_1 FILLER_56_260 ();
 sg13g2_decap_4 FILLER_56_269 ();
 sg13g2_fill_1 FILLER_56_353 ();
 sg13g2_fill_2 FILLER_56_363 ();
 sg13g2_fill_1 FILLER_56_365 ();
 sg13g2_fill_1 FILLER_56_409 ();
 sg13g2_fill_2 FILLER_56_415 ();
 sg13g2_decap_8 FILLER_56_425 ();
 sg13g2_fill_2 FILLER_56_432 ();
 sg13g2_fill_1 FILLER_56_434 ();
 sg13g2_fill_2 FILLER_56_440 ();
 sg13g2_fill_1 FILLER_56_442 ();
 sg13g2_fill_2 FILLER_56_484 ();
 sg13g2_fill_2 FILLER_56_551 ();
 sg13g2_fill_1 FILLER_56_553 ();
 sg13g2_fill_2 FILLER_56_568 ();
 sg13g2_decap_4 FILLER_56_579 ();
 sg13g2_fill_1 FILLER_56_583 ();
 sg13g2_decap_4 FILLER_56_602 ();
 sg13g2_fill_2 FILLER_56_606 ();
 sg13g2_decap_8 FILLER_56_645 ();
 sg13g2_fill_1 FILLER_56_657 ();
 sg13g2_fill_1 FILLER_56_662 ();
 sg13g2_fill_2 FILLER_56_726 ();
 sg13g2_fill_2 FILLER_56_736 ();
 sg13g2_fill_1 FILLER_56_738 ();
 sg13g2_fill_1 FILLER_56_814 ();
 sg13g2_fill_2 FILLER_56_883 ();
 sg13g2_fill_2 FILLER_56_938 ();
 sg13g2_fill_1 FILLER_56_940 ();
 sg13g2_fill_1 FILLER_56_1087 ();
 sg13g2_fill_1 FILLER_56_1120 ();
 sg13g2_fill_1 FILLER_56_1135 ();
 sg13g2_decap_8 FILLER_56_1197 ();
 sg13g2_decap_8 FILLER_56_1204 ();
 sg13g2_decap_8 FILLER_56_1211 ();
 sg13g2_decap_8 FILLER_56_1218 ();
 sg13g2_decap_8 FILLER_56_1225 ();
 sg13g2_decap_8 FILLER_56_1232 ();
 sg13g2_decap_8 FILLER_56_1239 ();
 sg13g2_decap_8 FILLER_56_1246 ();
 sg13g2_decap_8 FILLER_56_1253 ();
 sg13g2_decap_8 FILLER_56_1260 ();
 sg13g2_decap_8 FILLER_56_1267 ();
 sg13g2_decap_8 FILLER_56_1274 ();
 sg13g2_decap_8 FILLER_56_1281 ();
 sg13g2_decap_8 FILLER_56_1288 ();
 sg13g2_decap_8 FILLER_56_1295 ();
 sg13g2_decap_8 FILLER_56_1302 ();
 sg13g2_decap_4 FILLER_56_1309 ();
 sg13g2_fill_2 FILLER_56_1313 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_7 ();
 sg13g2_fill_2 FILLER_57_22 ();
 sg13g2_fill_1 FILLER_57_24 ();
 sg13g2_fill_2 FILLER_57_102 ();
 sg13g2_fill_1 FILLER_57_170 ();
 sg13g2_fill_1 FILLER_57_201 ();
 sg13g2_fill_2 FILLER_57_232 ();
 sg13g2_fill_1 FILLER_57_234 ();
 sg13g2_fill_1 FILLER_57_247 ();
 sg13g2_fill_2 FILLER_57_261 ();
 sg13g2_fill_1 FILLER_57_292 ();
 sg13g2_fill_1 FILLER_57_326 ();
 sg13g2_fill_2 FILLER_57_337 ();
 sg13g2_fill_1 FILLER_57_339 ();
 sg13g2_fill_1 FILLER_57_413 ();
 sg13g2_fill_2 FILLER_57_428 ();
 sg13g2_fill_1 FILLER_57_430 ();
 sg13g2_fill_2 FILLER_57_441 ();
 sg13g2_fill_1 FILLER_57_471 ();
 sg13g2_fill_2 FILLER_57_480 ();
 sg13g2_fill_2 FILLER_57_497 ();
 sg13g2_fill_1 FILLER_57_503 ();
 sg13g2_fill_2 FILLER_57_544 ();
 sg13g2_fill_1 FILLER_57_585 ();
 sg13g2_decap_4 FILLER_57_607 ();
 sg13g2_fill_1 FILLER_57_611 ();
 sg13g2_decap_8 FILLER_57_616 ();
 sg13g2_fill_1 FILLER_57_641 ();
 sg13g2_fill_2 FILLER_57_667 ();
 sg13g2_fill_1 FILLER_57_669 ();
 sg13g2_decap_8 FILLER_57_701 ();
 sg13g2_decap_4 FILLER_57_708 ();
 sg13g2_fill_2 FILLER_57_728 ();
 sg13g2_fill_1 FILLER_57_730 ();
 sg13g2_fill_1 FILLER_57_778 ();
 sg13g2_fill_2 FILLER_57_788 ();
 sg13g2_fill_1 FILLER_57_808 ();
 sg13g2_decap_4 FILLER_57_860 ();
 sg13g2_fill_2 FILLER_57_864 ();
 sg13g2_fill_2 FILLER_57_1047 ();
 sg13g2_decap_4 FILLER_57_1070 ();
 sg13g2_fill_1 FILLER_57_1074 ();
 sg13g2_fill_2 FILLER_57_1107 ();
 sg13g2_fill_1 FILLER_57_1189 ();
 sg13g2_decap_8 FILLER_57_1203 ();
 sg13g2_decap_8 FILLER_57_1210 ();
 sg13g2_decap_8 FILLER_57_1217 ();
 sg13g2_decap_8 FILLER_57_1224 ();
 sg13g2_decap_8 FILLER_57_1231 ();
 sg13g2_decap_8 FILLER_57_1238 ();
 sg13g2_decap_8 FILLER_57_1245 ();
 sg13g2_decap_8 FILLER_57_1252 ();
 sg13g2_decap_8 FILLER_57_1259 ();
 sg13g2_decap_8 FILLER_57_1266 ();
 sg13g2_decap_8 FILLER_57_1273 ();
 sg13g2_decap_8 FILLER_57_1280 ();
 sg13g2_decap_8 FILLER_57_1287 ();
 sg13g2_decap_8 FILLER_57_1294 ();
 sg13g2_decap_8 FILLER_57_1301 ();
 sg13g2_decap_8 FILLER_57_1308 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_fill_2 FILLER_58_14 ();
 sg13g2_fill_1 FILLER_58_16 ();
 sg13g2_fill_1 FILLER_58_44 ();
 sg13g2_fill_1 FILLER_58_63 ();
 sg13g2_fill_2 FILLER_58_107 ();
 sg13g2_fill_1 FILLER_58_137 ();
 sg13g2_fill_2 FILLER_58_164 ();
 sg13g2_fill_1 FILLER_58_209 ();
 sg13g2_fill_1 FILLER_58_228 ();
 sg13g2_fill_2 FILLER_58_237 ();
 sg13g2_fill_1 FILLER_58_239 ();
 sg13g2_fill_2 FILLER_58_271 ();
 sg13g2_fill_1 FILLER_58_273 ();
 sg13g2_fill_1 FILLER_58_317 ();
 sg13g2_fill_2 FILLER_58_353 ();
 sg13g2_fill_2 FILLER_58_412 ();
 sg13g2_fill_2 FILLER_58_480 ();
 sg13g2_fill_1 FILLER_58_524 ();
 sg13g2_fill_1 FILLER_58_534 ();
 sg13g2_fill_1 FILLER_58_540 ();
 sg13g2_fill_1 FILLER_58_551 ();
 sg13g2_fill_1 FILLER_58_557 ();
 sg13g2_fill_1 FILLER_58_566 ();
 sg13g2_fill_2 FILLER_58_627 ();
 sg13g2_fill_1 FILLER_58_629 ();
 sg13g2_fill_2 FILLER_58_639 ();
 sg13g2_fill_1 FILLER_58_646 ();
 sg13g2_fill_1 FILLER_58_662 ();
 sg13g2_decap_8 FILLER_58_667 ();
 sg13g2_decap_4 FILLER_58_674 ();
 sg13g2_fill_2 FILLER_58_678 ();
 sg13g2_fill_1 FILLER_58_685 ();
 sg13g2_decap_8 FILLER_58_690 ();
 sg13g2_fill_2 FILLER_58_697 ();
 sg13g2_fill_1 FILLER_58_699 ();
 sg13g2_fill_2 FILLER_58_722 ();
 sg13g2_fill_1 FILLER_58_750 ();
 sg13g2_fill_2 FILLER_58_777 ();
 sg13g2_decap_8 FILLER_58_827 ();
 sg13g2_fill_2 FILLER_58_834 ();
 sg13g2_fill_1 FILLER_58_836 ();
 sg13g2_fill_1 FILLER_58_850 ();
 sg13g2_fill_1 FILLER_58_877 ();
 sg13g2_fill_2 FILLER_58_929 ();
 sg13g2_fill_2 FILLER_58_1049 ();
 sg13g2_fill_1 FILLER_58_1103 ();
 sg13g2_decap_8 FILLER_58_1201 ();
 sg13g2_decap_8 FILLER_58_1208 ();
 sg13g2_decap_8 FILLER_58_1215 ();
 sg13g2_decap_8 FILLER_58_1222 ();
 sg13g2_decap_8 FILLER_58_1229 ();
 sg13g2_decap_8 FILLER_58_1236 ();
 sg13g2_decap_8 FILLER_58_1243 ();
 sg13g2_decap_8 FILLER_58_1250 ();
 sg13g2_decap_8 FILLER_58_1257 ();
 sg13g2_decap_8 FILLER_58_1264 ();
 sg13g2_decap_8 FILLER_58_1271 ();
 sg13g2_decap_8 FILLER_58_1278 ();
 sg13g2_decap_8 FILLER_58_1285 ();
 sg13g2_decap_8 FILLER_58_1292 ();
 sg13g2_decap_8 FILLER_58_1299 ();
 sg13g2_decap_8 FILLER_58_1306 ();
 sg13g2_fill_2 FILLER_58_1313 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_4 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_45 ();
 sg13g2_fill_1 FILLER_59_55 ();
 sg13g2_fill_2 FILLER_59_107 ();
 sg13g2_fill_2 FILLER_59_113 ();
 sg13g2_fill_1 FILLER_59_141 ();
 sg13g2_fill_1 FILLER_59_185 ();
 sg13g2_fill_1 FILLER_59_244 ();
 sg13g2_decap_8 FILLER_59_258 ();
 sg13g2_decap_4 FILLER_59_265 ();
 sg13g2_fill_2 FILLER_59_269 ();
 sg13g2_fill_2 FILLER_59_288 ();
 sg13g2_fill_1 FILLER_59_290 ();
 sg13g2_fill_1 FILLER_59_335 ();
 sg13g2_fill_1 FILLER_59_381 ();
 sg13g2_fill_1 FILLER_59_400 ();
 sg13g2_fill_1 FILLER_59_475 ();
 sg13g2_fill_2 FILLER_59_572 ();
 sg13g2_fill_2 FILLER_59_593 ();
 sg13g2_fill_1 FILLER_59_595 ();
 sg13g2_decap_8 FILLER_59_600 ();
 sg13g2_fill_2 FILLER_59_607 ();
 sg13g2_fill_2 FILLER_59_625 ();
 sg13g2_fill_2 FILLER_59_635 ();
 sg13g2_fill_1 FILLER_59_647 ();
 sg13g2_fill_1 FILLER_59_684 ();
 sg13g2_fill_2 FILLER_59_689 ();
 sg13g2_fill_1 FILLER_59_691 ();
 sg13g2_decap_8 FILLER_59_728 ();
 sg13g2_fill_2 FILLER_59_739 ();
 sg13g2_fill_1 FILLER_59_741 ();
 sg13g2_fill_2 FILLER_59_747 ();
 sg13g2_fill_1 FILLER_59_771 ();
 sg13g2_fill_1 FILLER_59_810 ();
 sg13g2_decap_8 FILLER_59_848 ();
 sg13g2_fill_1 FILLER_59_855 ();
 sg13g2_fill_2 FILLER_59_860 ();
 sg13g2_fill_1 FILLER_59_866 ();
 sg13g2_decap_4 FILLER_59_906 ();
 sg13g2_fill_1 FILLER_59_936 ();
 sg13g2_fill_2 FILLER_59_942 ();
 sg13g2_decap_4 FILLER_59_957 ();
 sg13g2_fill_2 FILLER_59_1046 ();
 sg13g2_fill_1 FILLER_59_1073 ();
 sg13g2_fill_2 FILLER_59_1088 ();
 sg13g2_fill_2 FILLER_59_1104 ();
 sg13g2_fill_1 FILLER_59_1106 ();
 sg13g2_fill_2 FILLER_59_1123 ();
 sg13g2_fill_1 FILLER_59_1125 ();
 sg13g2_decap_8 FILLER_59_1203 ();
 sg13g2_decap_8 FILLER_59_1210 ();
 sg13g2_decap_8 FILLER_59_1217 ();
 sg13g2_decap_8 FILLER_59_1224 ();
 sg13g2_decap_8 FILLER_59_1231 ();
 sg13g2_decap_8 FILLER_59_1238 ();
 sg13g2_decap_8 FILLER_59_1245 ();
 sg13g2_decap_8 FILLER_59_1252 ();
 sg13g2_decap_8 FILLER_59_1259 ();
 sg13g2_decap_8 FILLER_59_1266 ();
 sg13g2_decap_8 FILLER_59_1273 ();
 sg13g2_decap_8 FILLER_59_1280 ();
 sg13g2_decap_8 FILLER_59_1287 ();
 sg13g2_decap_8 FILLER_59_1294 ();
 sg13g2_decap_8 FILLER_59_1301 ();
 sg13g2_decap_8 FILLER_59_1308 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_39 ();
 sg13g2_fill_2 FILLER_60_70 ();
 sg13g2_fill_2 FILLER_60_107 ();
 sg13g2_fill_1 FILLER_60_109 ();
 sg13g2_fill_2 FILLER_60_128 ();
 sg13g2_fill_1 FILLER_60_130 ();
 sg13g2_fill_2 FILLER_60_135 ();
 sg13g2_decap_4 FILLER_60_156 ();
 sg13g2_fill_1 FILLER_60_216 ();
 sg13g2_fill_2 FILLER_60_226 ();
 sg13g2_fill_1 FILLER_60_276 ();
 sg13g2_fill_2 FILLER_60_291 ();
 sg13g2_fill_1 FILLER_60_319 ();
 sg13g2_fill_2 FILLER_60_329 ();
 sg13g2_fill_1 FILLER_60_407 ();
 sg13g2_fill_2 FILLER_60_421 ();
 sg13g2_decap_8 FILLER_60_497 ();
 sg13g2_fill_2 FILLER_60_504 ();
 sg13g2_fill_1 FILLER_60_506 ();
 sg13g2_decap_4 FILLER_60_512 ();
 sg13g2_fill_1 FILLER_60_516 ();
 sg13g2_fill_2 FILLER_60_530 ();
 sg13g2_fill_1 FILLER_60_570 ();
 sg13g2_fill_1 FILLER_60_577 ();
 sg13g2_fill_2 FILLER_60_583 ();
 sg13g2_fill_1 FILLER_60_664 ();
 sg13g2_fill_1 FILLER_60_700 ();
 sg13g2_fill_2 FILLER_60_733 ();
 sg13g2_fill_1 FILLER_60_806 ();
 sg13g2_fill_2 FILLER_60_820 ();
 sg13g2_fill_2 FILLER_60_827 ();
 sg13g2_fill_1 FILLER_60_829 ();
 sg13g2_fill_1 FILLER_60_834 ();
 sg13g2_fill_1 FILLER_60_844 ();
 sg13g2_decap_4 FILLER_60_850 ();
 sg13g2_fill_1 FILLER_60_854 ();
 sg13g2_fill_1 FILLER_60_864 ();
 sg13g2_decap_8 FILLER_60_902 ();
 sg13g2_decap_8 FILLER_60_909 ();
 sg13g2_fill_1 FILLER_60_920 ();
 sg13g2_fill_1 FILLER_60_930 ();
 sg13g2_fill_2 FILLER_60_934 ();
 sg13g2_fill_1 FILLER_60_1007 ();
 sg13g2_fill_1 FILLER_60_1034 ();
 sg13g2_decap_8 FILLER_60_1064 ();
 sg13g2_decap_8 FILLER_60_1071 ();
 sg13g2_decap_8 FILLER_60_1193 ();
 sg13g2_decap_8 FILLER_60_1200 ();
 sg13g2_decap_8 FILLER_60_1207 ();
 sg13g2_decap_8 FILLER_60_1214 ();
 sg13g2_decap_8 FILLER_60_1221 ();
 sg13g2_decap_8 FILLER_60_1228 ();
 sg13g2_decap_8 FILLER_60_1235 ();
 sg13g2_decap_8 FILLER_60_1242 ();
 sg13g2_decap_8 FILLER_60_1249 ();
 sg13g2_decap_8 FILLER_60_1256 ();
 sg13g2_decap_8 FILLER_60_1263 ();
 sg13g2_decap_8 FILLER_60_1270 ();
 sg13g2_decap_8 FILLER_60_1277 ();
 sg13g2_decap_8 FILLER_60_1284 ();
 sg13g2_decap_8 FILLER_60_1291 ();
 sg13g2_decap_8 FILLER_60_1298 ();
 sg13g2_decap_8 FILLER_60_1305 ();
 sg13g2_fill_2 FILLER_60_1312 ();
 sg13g2_fill_1 FILLER_60_1314 ();
 sg13g2_fill_1 FILLER_61_26 ();
 sg13g2_fill_1 FILLER_61_35 ();
 sg13g2_fill_2 FILLER_61_121 ();
 sg13g2_fill_1 FILLER_61_123 ();
 sg13g2_fill_2 FILLER_61_133 ();
 sg13g2_decap_8 FILLER_61_156 ();
 sg13g2_fill_2 FILLER_61_163 ();
 sg13g2_fill_1 FILLER_61_165 ();
 sg13g2_fill_2 FILLER_61_175 ();
 sg13g2_fill_1 FILLER_61_177 ();
 sg13g2_fill_1 FILLER_61_203 ();
 sg13g2_decap_4 FILLER_61_248 ();
 sg13g2_fill_2 FILLER_61_265 ();
 sg13g2_fill_1 FILLER_61_267 ();
 sg13g2_fill_1 FILLER_61_286 ();
 sg13g2_fill_2 FILLER_61_301 ();
 sg13g2_fill_2 FILLER_61_338 ();
 sg13g2_fill_1 FILLER_61_340 ();
 sg13g2_fill_2 FILLER_61_350 ();
 sg13g2_decap_4 FILLER_61_373 ();
 sg13g2_fill_2 FILLER_61_396 ();
 sg13g2_fill_1 FILLER_61_409 ();
 sg13g2_fill_1 FILLER_61_418 ();
 sg13g2_fill_2 FILLER_61_434 ();
 sg13g2_fill_1 FILLER_61_436 ();
 sg13g2_decap_4 FILLER_61_445 ();
 sg13g2_fill_1 FILLER_61_449 ();
 sg13g2_fill_1 FILLER_61_459 ();
 sg13g2_fill_2 FILLER_61_474 ();
 sg13g2_decap_4 FILLER_61_484 ();
 sg13g2_fill_1 FILLER_61_488 ();
 sg13g2_fill_2 FILLER_61_497 ();
 sg13g2_fill_1 FILLER_61_499 ();
 sg13g2_fill_2 FILLER_61_531 ();
 sg13g2_fill_1 FILLER_61_565 ();
 sg13g2_fill_1 FILLER_61_585 ();
 sg13g2_fill_1 FILLER_61_621 ();
 sg13g2_decap_4 FILLER_61_685 ();
 sg13g2_fill_2 FILLER_61_758 ();
 sg13g2_fill_2 FILLER_61_765 ();
 sg13g2_fill_2 FILLER_61_772 ();
 sg13g2_fill_1 FILLER_61_866 ();
 sg13g2_decap_4 FILLER_61_901 ();
 sg13g2_fill_2 FILLER_61_965 ();
 sg13g2_fill_1 FILLER_61_975 ();
 sg13g2_fill_1 FILLER_61_989 ();
 sg13g2_fill_1 FILLER_61_1020 ();
 sg13g2_fill_2 FILLER_61_1028 ();
 sg13g2_decap_8 FILLER_61_1072 ();
 sg13g2_fill_2 FILLER_61_1079 ();
 sg13g2_fill_1 FILLER_61_1081 ();
 sg13g2_fill_1 FILLER_61_1087 ();
 sg13g2_fill_2 FILLER_61_1119 ();
 sg13g2_decap_8 FILLER_61_1201 ();
 sg13g2_decap_8 FILLER_61_1208 ();
 sg13g2_decap_8 FILLER_61_1215 ();
 sg13g2_decap_8 FILLER_61_1222 ();
 sg13g2_decap_8 FILLER_61_1229 ();
 sg13g2_decap_8 FILLER_61_1236 ();
 sg13g2_decap_8 FILLER_61_1243 ();
 sg13g2_decap_8 FILLER_61_1250 ();
 sg13g2_decap_8 FILLER_61_1257 ();
 sg13g2_decap_8 FILLER_61_1264 ();
 sg13g2_decap_8 FILLER_61_1271 ();
 sg13g2_decap_8 FILLER_61_1278 ();
 sg13g2_decap_8 FILLER_61_1285 ();
 sg13g2_decap_8 FILLER_61_1292 ();
 sg13g2_decap_8 FILLER_61_1299 ();
 sg13g2_decap_8 FILLER_61_1306 ();
 sg13g2_fill_2 FILLER_61_1313 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_43 ();
 sg13g2_fill_2 FILLER_62_50 ();
 sg13g2_fill_1 FILLER_62_67 ();
 sg13g2_fill_2 FILLER_62_75 ();
 sg13g2_decap_4 FILLER_62_82 ();
 sg13g2_fill_2 FILLER_62_86 ();
 sg13g2_fill_1 FILLER_62_96 ();
 sg13g2_fill_2 FILLER_62_127 ();
 sg13g2_fill_2 FILLER_62_181 ();
 sg13g2_fill_1 FILLER_62_183 ();
 sg13g2_fill_2 FILLER_62_188 ();
 sg13g2_fill_2 FILLER_62_229 ();
 sg13g2_fill_1 FILLER_62_231 ();
 sg13g2_fill_2 FILLER_62_251 ();
 sg13g2_fill_1 FILLER_62_253 ();
 sg13g2_fill_1 FILLER_62_280 ();
 sg13g2_fill_2 FILLER_62_330 ();
 sg13g2_fill_1 FILLER_62_332 ();
 sg13g2_fill_1 FILLER_62_337 ();
 sg13g2_fill_1 FILLER_62_346 ();
 sg13g2_fill_2 FILLER_62_351 ();
 sg13g2_fill_1 FILLER_62_419 ();
 sg13g2_decap_4 FILLER_62_446 ();
 sg13g2_fill_1 FILLER_62_450 ();
 sg13g2_fill_1 FILLER_62_460 ();
 sg13g2_fill_1 FILLER_62_503 ();
 sg13g2_decap_4 FILLER_62_509 ();
 sg13g2_fill_2 FILLER_62_526 ();
 sg13g2_decap_4 FILLER_62_538 ();
 sg13g2_fill_2 FILLER_62_542 ();
 sg13g2_decap_8 FILLER_62_548 ();
 sg13g2_decap_4 FILLER_62_555 ();
 sg13g2_fill_2 FILLER_62_559 ();
 sg13g2_fill_2 FILLER_62_566 ();
 sg13g2_fill_1 FILLER_62_568 ();
 sg13g2_fill_2 FILLER_62_575 ();
 sg13g2_fill_1 FILLER_62_596 ();
 sg13g2_fill_1 FILLER_62_634 ();
 sg13g2_decap_8 FILLER_62_665 ();
 sg13g2_fill_1 FILLER_62_672 ();
 sg13g2_fill_2 FILLER_62_699 ();
 sg13g2_fill_1 FILLER_62_715 ();
 sg13g2_fill_1 FILLER_62_729 ();
 sg13g2_fill_1 FILLER_62_740 ();
 sg13g2_decap_4 FILLER_62_752 ();
 sg13g2_fill_1 FILLER_62_756 ();
 sg13g2_fill_2 FILLER_62_761 ();
 sg13g2_fill_1 FILLER_62_821 ();
 sg13g2_fill_2 FILLER_62_845 ();
 sg13g2_fill_2 FILLER_62_883 ();
 sg13g2_fill_1 FILLER_62_928 ();
 sg13g2_fill_1 FILLER_62_1087 ();
 sg13g2_fill_1 FILLER_62_1108 ();
 sg13g2_fill_2 FILLER_62_1127 ();
 sg13g2_fill_1 FILLER_62_1147 ();
 sg13g2_decap_8 FILLER_62_1196 ();
 sg13g2_decap_8 FILLER_62_1203 ();
 sg13g2_decap_8 FILLER_62_1210 ();
 sg13g2_decap_8 FILLER_62_1217 ();
 sg13g2_decap_8 FILLER_62_1224 ();
 sg13g2_decap_8 FILLER_62_1231 ();
 sg13g2_decap_8 FILLER_62_1238 ();
 sg13g2_decap_8 FILLER_62_1245 ();
 sg13g2_decap_8 FILLER_62_1252 ();
 sg13g2_decap_8 FILLER_62_1259 ();
 sg13g2_decap_8 FILLER_62_1266 ();
 sg13g2_decap_8 FILLER_62_1273 ();
 sg13g2_decap_8 FILLER_62_1280 ();
 sg13g2_decap_8 FILLER_62_1287 ();
 sg13g2_decap_8 FILLER_62_1294 ();
 sg13g2_decap_8 FILLER_62_1301 ();
 sg13g2_decap_8 FILLER_62_1308 ();
 sg13g2_decap_4 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_25 ();
 sg13g2_fill_1 FILLER_63_51 ();
 sg13g2_fill_1 FILLER_63_71 ();
 sg13g2_fill_1 FILLER_63_103 ();
 sg13g2_fill_2 FILLER_63_137 ();
 sg13g2_fill_1 FILLER_63_139 ();
 sg13g2_fill_2 FILLER_63_145 ();
 sg13g2_fill_1 FILLER_63_151 ();
 sg13g2_fill_2 FILLER_63_156 ();
 sg13g2_fill_2 FILLER_63_171 ();
 sg13g2_fill_2 FILLER_63_213 ();
 sg13g2_fill_1 FILLER_63_220 ();
 sg13g2_fill_2 FILLER_63_226 ();
 sg13g2_fill_1 FILLER_63_228 ();
 sg13g2_fill_2 FILLER_63_234 ();
 sg13g2_decap_4 FILLER_63_240 ();
 sg13g2_fill_1 FILLER_63_244 ();
 sg13g2_fill_2 FILLER_63_258 ();
 sg13g2_fill_2 FILLER_63_273 ();
 sg13g2_fill_2 FILLER_63_292 ();
 sg13g2_fill_2 FILLER_63_308 ();
 sg13g2_fill_1 FILLER_63_335 ();
 sg13g2_fill_2 FILLER_63_380 ();
 sg13g2_fill_1 FILLER_63_407 ();
 sg13g2_fill_2 FILLER_63_428 ();
 sg13g2_fill_1 FILLER_63_430 ();
 sg13g2_decap_4 FILLER_63_435 ();
 sg13g2_fill_2 FILLER_63_444 ();
 sg13g2_fill_2 FILLER_63_485 ();
 sg13g2_fill_1 FILLER_63_534 ();
 sg13g2_fill_1 FILLER_63_570 ();
 sg13g2_fill_2 FILLER_63_646 ();
 sg13g2_fill_2 FILLER_63_662 ();
 sg13g2_fill_2 FILLER_63_673 ();
 sg13g2_fill_1 FILLER_63_688 ();
 sg13g2_fill_1 FILLER_63_716 ();
 sg13g2_fill_2 FILLER_63_735 ();
 sg13g2_fill_1 FILLER_63_745 ();
 sg13g2_fill_1 FILLER_63_888 ();
 sg13g2_fill_2 FILLER_63_919 ();
 sg13g2_fill_2 FILLER_63_1019 ();
 sg13g2_fill_2 FILLER_63_1029 ();
 sg13g2_decap_8 FILLER_63_1101 ();
 sg13g2_fill_1 FILLER_63_1108 ();
 sg13g2_fill_1 FILLER_63_1114 ();
 sg13g2_decap_8 FILLER_63_1118 ();
 sg13g2_fill_1 FILLER_63_1125 ();
 sg13g2_fill_2 FILLER_63_1153 ();
 sg13g2_fill_1 FILLER_63_1155 ();
 sg13g2_fill_1 FILLER_63_1164 ();
 sg13g2_fill_2 FILLER_63_1179 ();
 sg13g2_decap_8 FILLER_63_1194 ();
 sg13g2_decap_8 FILLER_63_1201 ();
 sg13g2_decap_8 FILLER_63_1208 ();
 sg13g2_decap_8 FILLER_63_1215 ();
 sg13g2_decap_8 FILLER_63_1222 ();
 sg13g2_decap_8 FILLER_63_1229 ();
 sg13g2_decap_8 FILLER_63_1236 ();
 sg13g2_decap_8 FILLER_63_1243 ();
 sg13g2_decap_8 FILLER_63_1250 ();
 sg13g2_decap_8 FILLER_63_1257 ();
 sg13g2_decap_8 FILLER_63_1264 ();
 sg13g2_decap_8 FILLER_63_1271 ();
 sg13g2_decap_8 FILLER_63_1278 ();
 sg13g2_decap_8 FILLER_63_1285 ();
 sg13g2_decap_8 FILLER_63_1292 ();
 sg13g2_decap_8 FILLER_63_1299 ();
 sg13g2_decap_8 FILLER_63_1306 ();
 sg13g2_fill_2 FILLER_63_1313 ();
 sg13g2_fill_2 FILLER_64_44 ();
 sg13g2_fill_1 FILLER_64_46 ();
 sg13g2_fill_2 FILLER_64_82 ();
 sg13g2_fill_1 FILLER_64_98 ();
 sg13g2_fill_1 FILLER_64_125 ();
 sg13g2_fill_2 FILLER_64_172 ();
 sg13g2_fill_1 FILLER_64_174 ();
 sg13g2_fill_2 FILLER_64_179 ();
 sg13g2_decap_4 FILLER_64_195 ();
 sg13g2_decap_8 FILLER_64_225 ();
 sg13g2_fill_2 FILLER_64_232 ();
 sg13g2_fill_1 FILLER_64_249 ();
 sg13g2_fill_2 FILLER_64_268 ();
 sg13g2_fill_1 FILLER_64_270 ();
 sg13g2_fill_1 FILLER_64_296 ();
 sg13g2_fill_2 FILLER_64_355 ();
 sg13g2_fill_1 FILLER_64_357 ();
 sg13g2_fill_1 FILLER_64_411 ();
 sg13g2_fill_1 FILLER_64_419 ();
 sg13g2_fill_2 FILLER_64_438 ();
 sg13g2_fill_1 FILLER_64_440 ();
 sg13g2_decap_8 FILLER_64_451 ();
 sg13g2_fill_2 FILLER_64_458 ();
 sg13g2_fill_2 FILLER_64_465 ();
 sg13g2_fill_1 FILLER_64_485 ();
 sg13g2_fill_1 FILLER_64_499 ();
 sg13g2_decap_4 FILLER_64_518 ();
 sg13g2_fill_1 FILLER_64_522 ();
 sg13g2_fill_2 FILLER_64_611 ();
 sg13g2_fill_1 FILLER_64_613 ();
 sg13g2_fill_2 FILLER_64_626 ();
 sg13g2_fill_1 FILLER_64_628 ();
 sg13g2_fill_2 FILLER_64_634 ();
 sg13g2_fill_2 FILLER_64_640 ();
 sg13g2_fill_1 FILLER_64_642 ();
 sg13g2_fill_1 FILLER_64_739 ();
 sg13g2_fill_2 FILLER_64_769 ();
 sg13g2_fill_2 FILLER_64_781 ();
 sg13g2_fill_1 FILLER_64_863 ();
 sg13g2_fill_2 FILLER_64_874 ();
 sg13g2_fill_1 FILLER_64_876 ();
 sg13g2_fill_1 FILLER_64_936 ();
 sg13g2_fill_2 FILLER_64_948 ();
 sg13g2_fill_1 FILLER_64_1049 ();
 sg13g2_decap_4 FILLER_64_1074 ();
 sg13g2_fill_1 FILLER_64_1083 ();
 sg13g2_fill_2 FILLER_64_1116 ();
 sg13g2_fill_1 FILLER_64_1118 ();
 sg13g2_fill_2 FILLER_64_1149 ();
 sg13g2_fill_2 FILLER_64_1169 ();
 sg13g2_fill_1 FILLER_64_1171 ();
 sg13g2_decap_8 FILLER_64_1189 ();
 sg13g2_decap_8 FILLER_64_1196 ();
 sg13g2_decap_8 FILLER_64_1203 ();
 sg13g2_decap_8 FILLER_64_1210 ();
 sg13g2_decap_8 FILLER_64_1217 ();
 sg13g2_decap_8 FILLER_64_1224 ();
 sg13g2_decap_8 FILLER_64_1231 ();
 sg13g2_decap_8 FILLER_64_1238 ();
 sg13g2_decap_8 FILLER_64_1245 ();
 sg13g2_decap_8 FILLER_64_1252 ();
 sg13g2_decap_8 FILLER_64_1259 ();
 sg13g2_decap_8 FILLER_64_1266 ();
 sg13g2_decap_8 FILLER_64_1273 ();
 sg13g2_decap_8 FILLER_64_1280 ();
 sg13g2_decap_8 FILLER_64_1287 ();
 sg13g2_decap_8 FILLER_64_1294 ();
 sg13g2_decap_8 FILLER_64_1301 ();
 sg13g2_decap_8 FILLER_64_1308 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_14 ();
 sg13g2_fill_1 FILLER_65_46 ();
 sg13g2_decap_8 FILLER_65_101 ();
 sg13g2_decap_4 FILLER_65_108 ();
 sg13g2_fill_2 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_118 ();
 sg13g2_decap_4 FILLER_65_135 ();
 sg13g2_fill_2 FILLER_65_139 ();
 sg13g2_fill_2 FILLER_65_151 ();
 sg13g2_fill_2 FILLER_65_162 ();
 sg13g2_fill_1 FILLER_65_190 ();
 sg13g2_decap_8 FILLER_65_217 ();
 sg13g2_fill_1 FILLER_65_256 ();
 sg13g2_fill_2 FILLER_65_306 ();
 sg13g2_fill_2 FILLER_65_312 ();
 sg13g2_fill_2 FILLER_65_375 ();
 sg13g2_decap_4 FILLER_65_445 ();
 sg13g2_fill_1 FILLER_65_475 ();
 sg13g2_decap_4 FILLER_65_513 ();
 sg13g2_fill_1 FILLER_65_517 ();
 sg13g2_fill_2 FILLER_65_523 ();
 sg13g2_fill_1 FILLER_65_611 ();
 sg13g2_decap_4 FILLER_65_616 ();
 sg13g2_fill_1 FILLER_65_620 ();
 sg13g2_fill_2 FILLER_65_656 ();
 sg13g2_fill_2 FILLER_65_663 ();
 sg13g2_decap_8 FILLER_65_693 ();
 sg13g2_fill_2 FILLER_65_700 ();
 sg13g2_fill_2 FILLER_65_709 ();
 sg13g2_fill_1 FILLER_65_711 ();
 sg13g2_fill_2 FILLER_65_743 ();
 sg13g2_fill_2 FILLER_65_816 ();
 sg13g2_fill_1 FILLER_65_818 ();
 sg13g2_fill_1 FILLER_65_849 ();
 sg13g2_decap_8 FILLER_65_881 ();
 sg13g2_fill_1 FILLER_65_900 ();
 sg13g2_fill_1 FILLER_65_995 ();
 sg13g2_fill_2 FILLER_65_1041 ();
 sg13g2_fill_2 FILLER_65_1046 ();
 sg13g2_fill_1 FILLER_65_1056 ();
 sg13g2_fill_1 FILLER_65_1071 ();
 sg13g2_fill_2 FILLER_65_1077 ();
 sg13g2_fill_2 FILLER_65_1118 ();
 sg13g2_fill_1 FILLER_65_1133 ();
 sg13g2_fill_2 FILLER_65_1148 ();
 sg13g2_decap_8 FILLER_65_1185 ();
 sg13g2_decap_8 FILLER_65_1192 ();
 sg13g2_decap_8 FILLER_65_1199 ();
 sg13g2_decap_8 FILLER_65_1206 ();
 sg13g2_decap_8 FILLER_65_1213 ();
 sg13g2_decap_8 FILLER_65_1220 ();
 sg13g2_decap_8 FILLER_65_1227 ();
 sg13g2_decap_8 FILLER_65_1234 ();
 sg13g2_decap_8 FILLER_65_1241 ();
 sg13g2_decap_8 FILLER_65_1248 ();
 sg13g2_decap_8 FILLER_65_1255 ();
 sg13g2_decap_8 FILLER_65_1262 ();
 sg13g2_decap_8 FILLER_65_1269 ();
 sg13g2_decap_8 FILLER_65_1276 ();
 sg13g2_decap_8 FILLER_65_1283 ();
 sg13g2_decap_8 FILLER_65_1290 ();
 sg13g2_decap_8 FILLER_65_1297 ();
 sg13g2_decap_8 FILLER_65_1304 ();
 sg13g2_decap_4 FILLER_65_1311 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_7 ();
 sg13g2_fill_2 FILLER_66_51 ();
 sg13g2_fill_2 FILLER_66_79 ();
 sg13g2_fill_1 FILLER_66_81 ();
 sg13g2_fill_2 FILLER_66_121 ();
 sg13g2_fill_1 FILLER_66_123 ();
 sg13g2_fill_2 FILLER_66_134 ();
 sg13g2_fill_1 FILLER_66_136 ();
 sg13g2_fill_2 FILLER_66_176 ();
 sg13g2_fill_1 FILLER_66_178 ();
 sg13g2_fill_2 FILLER_66_188 ();
 sg13g2_fill_1 FILLER_66_190 ();
 sg13g2_decap_4 FILLER_66_217 ();
 sg13g2_fill_2 FILLER_66_243 ();
 sg13g2_fill_1 FILLER_66_245 ();
 sg13g2_fill_2 FILLER_66_263 ();
 sg13g2_fill_1 FILLER_66_265 ();
 sg13g2_fill_1 FILLER_66_280 ();
 sg13g2_fill_1 FILLER_66_324 ();
 sg13g2_fill_1 FILLER_66_339 ();
 sg13g2_fill_1 FILLER_66_349 ();
 sg13g2_fill_2 FILLER_66_358 ();
 sg13g2_fill_1 FILLER_66_360 ();
 sg13g2_fill_1 FILLER_66_384 ();
 sg13g2_fill_2 FILLER_66_398 ();
 sg13g2_fill_2 FILLER_66_405 ();
 sg13g2_fill_1 FILLER_66_415 ();
 sg13g2_fill_2 FILLER_66_444 ();
 sg13g2_fill_1 FILLER_66_446 ();
 sg13g2_decap_8 FILLER_66_452 ();
 sg13g2_fill_1 FILLER_66_459 ();
 sg13g2_decap_4 FILLER_66_468 ();
 sg13g2_fill_2 FILLER_66_495 ();
 sg13g2_fill_1 FILLER_66_497 ();
 sg13g2_decap_4 FILLER_66_507 ();
 sg13g2_fill_1 FILLER_66_523 ();
 sg13g2_fill_1 FILLER_66_528 ();
 sg13g2_fill_1 FILLER_66_538 ();
 sg13g2_fill_2 FILLER_66_552 ();
 sg13g2_fill_2 FILLER_66_572 ();
 sg13g2_fill_1 FILLER_66_587 ();
 sg13g2_fill_2 FILLER_66_627 ();
 sg13g2_fill_2 FILLER_66_646 ();
 sg13g2_fill_2 FILLER_66_667 ();
 sg13g2_fill_1 FILLER_66_669 ();
 sg13g2_decap_4 FILLER_66_703 ();
 sg13g2_decap_4 FILLER_66_712 ();
 sg13g2_fill_2 FILLER_66_723 ();
 sg13g2_fill_1 FILLER_66_725 ();
 sg13g2_fill_2 FILLER_66_794 ();
 sg13g2_decap_4 FILLER_66_823 ();
 sg13g2_fill_1 FILLER_66_834 ();
 sg13g2_fill_1 FILLER_66_855 ();
 sg13g2_fill_1 FILLER_66_910 ();
 sg13g2_fill_1 FILLER_66_957 ();
 sg13g2_fill_2 FILLER_66_989 ();
 sg13g2_fill_1 FILLER_66_1052 ();
 sg13g2_fill_1 FILLER_66_1077 ();
 sg13g2_decap_4 FILLER_66_1085 ();
 sg13g2_fill_2 FILLER_66_1089 ();
 sg13g2_fill_1 FILLER_66_1095 ();
 sg13g2_decap_8 FILLER_66_1162 ();
 sg13g2_fill_1 FILLER_66_1169 ();
 sg13g2_decap_8 FILLER_66_1174 ();
 sg13g2_decap_8 FILLER_66_1181 ();
 sg13g2_decap_8 FILLER_66_1188 ();
 sg13g2_decap_8 FILLER_66_1195 ();
 sg13g2_decap_8 FILLER_66_1202 ();
 sg13g2_decap_8 FILLER_66_1209 ();
 sg13g2_decap_8 FILLER_66_1216 ();
 sg13g2_decap_8 FILLER_66_1223 ();
 sg13g2_decap_8 FILLER_66_1230 ();
 sg13g2_decap_8 FILLER_66_1237 ();
 sg13g2_decap_8 FILLER_66_1244 ();
 sg13g2_decap_8 FILLER_66_1251 ();
 sg13g2_decap_8 FILLER_66_1258 ();
 sg13g2_decap_8 FILLER_66_1265 ();
 sg13g2_decap_8 FILLER_66_1272 ();
 sg13g2_decap_8 FILLER_66_1279 ();
 sg13g2_decap_8 FILLER_66_1286 ();
 sg13g2_decap_8 FILLER_66_1293 ();
 sg13g2_decap_8 FILLER_66_1300 ();
 sg13g2_decap_8 FILLER_66_1307 ();
 sg13g2_fill_1 FILLER_66_1314 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_4 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_15 ();
 sg13g2_decap_8 FILLER_67_22 ();
 sg13g2_fill_2 FILLER_67_29 ();
 sg13g2_fill_1 FILLER_67_31 ();
 sg13g2_fill_2 FILLER_67_55 ();
 sg13g2_fill_1 FILLER_67_57 ();
 sg13g2_fill_2 FILLER_67_62 ();
 sg13g2_fill_2 FILLER_67_72 ();
 sg13g2_fill_1 FILLER_67_74 ();
 sg13g2_decap_4 FILLER_67_83 ();
 sg13g2_decap_4 FILLER_67_113 ();
 sg13g2_fill_2 FILLER_67_117 ();
 sg13g2_fill_1 FILLER_67_128 ();
 sg13g2_fill_2 FILLER_67_134 ();
 sg13g2_fill_2 FILLER_67_180 ();
 sg13g2_fill_1 FILLER_67_191 ();
 sg13g2_decap_8 FILLER_67_218 ();
 sg13g2_fill_1 FILLER_67_225 ();
 sg13g2_fill_2 FILLER_67_260 ();
 sg13g2_decap_4 FILLER_67_313 ();
 sg13g2_fill_2 FILLER_67_317 ();
 sg13g2_fill_2 FILLER_67_334 ();
 sg13g2_fill_2 FILLER_67_396 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_fill_2 FILLER_67_425 ();
 sg13g2_fill_2 FILLER_67_435 ();
 sg13g2_fill_1 FILLER_67_504 ();
 sg13g2_decap_8 FILLER_67_518 ();
 sg13g2_fill_2 FILLER_67_525 ();
 sg13g2_fill_1 FILLER_67_527 ();
 sg13g2_fill_2 FILLER_67_569 ();
 sg13g2_fill_1 FILLER_67_587 ();
 sg13g2_decap_8 FILLER_67_614 ();
 sg13g2_fill_1 FILLER_67_621 ();
 sg13g2_decap_4 FILLER_67_626 ();
 sg13g2_fill_2 FILLER_67_677 ();
 sg13g2_fill_1 FILLER_67_679 ();
 sg13g2_fill_2 FILLER_67_693 ();
 sg13g2_fill_1 FILLER_67_764 ();
 sg13g2_fill_2 FILLER_67_770 ();
 sg13g2_fill_2 FILLER_67_876 ();
 sg13g2_fill_2 FILLER_67_925 ();
 sg13g2_fill_1 FILLER_67_982 ();
 sg13g2_fill_2 FILLER_67_1002 ();
 sg13g2_fill_2 FILLER_67_1018 ();
 sg13g2_fill_1 FILLER_67_1020 ();
 sg13g2_decap_4 FILLER_67_1067 ();
 sg13g2_fill_2 FILLER_67_1107 ();
 sg13g2_fill_2 FILLER_67_1117 ();
 sg13g2_fill_2 FILLER_67_1123 ();
 sg13g2_fill_1 FILLER_67_1125 ();
 sg13g2_fill_1 FILLER_67_1135 ();
 sg13g2_fill_1 FILLER_67_1144 ();
 sg13g2_decap_8 FILLER_67_1162 ();
 sg13g2_decap_8 FILLER_67_1169 ();
 sg13g2_decap_8 FILLER_67_1176 ();
 sg13g2_decap_8 FILLER_67_1183 ();
 sg13g2_decap_8 FILLER_67_1190 ();
 sg13g2_decap_8 FILLER_67_1197 ();
 sg13g2_decap_8 FILLER_67_1204 ();
 sg13g2_decap_8 FILLER_67_1211 ();
 sg13g2_decap_8 FILLER_67_1218 ();
 sg13g2_decap_8 FILLER_67_1225 ();
 sg13g2_decap_8 FILLER_67_1232 ();
 sg13g2_decap_8 FILLER_67_1239 ();
 sg13g2_decap_8 FILLER_67_1246 ();
 sg13g2_decap_8 FILLER_67_1253 ();
 sg13g2_decap_8 FILLER_67_1260 ();
 sg13g2_decap_8 FILLER_67_1267 ();
 sg13g2_decap_8 FILLER_67_1274 ();
 sg13g2_decap_8 FILLER_67_1281 ();
 sg13g2_decap_8 FILLER_67_1288 ();
 sg13g2_decap_8 FILLER_67_1295 ();
 sg13g2_decap_8 FILLER_67_1302 ();
 sg13g2_decap_4 FILLER_67_1309 ();
 sg13g2_fill_2 FILLER_67_1313 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_27 ();
 sg13g2_fill_2 FILLER_68_50 ();
 sg13g2_fill_2 FILLER_68_66 ();
 sg13g2_fill_1 FILLER_68_99 ();
 sg13g2_fill_1 FILLER_68_126 ();
 sg13g2_fill_2 FILLER_68_147 ();
 sg13g2_fill_2 FILLER_68_201 ();
 sg13g2_fill_1 FILLER_68_278 ();
 sg13g2_fill_1 FILLER_68_340 ();
 sg13g2_fill_2 FILLER_68_384 ();
 sg13g2_fill_2 FILLER_68_497 ();
 sg13g2_fill_1 FILLER_68_504 ();
 sg13g2_decap_8 FILLER_68_535 ();
 sg13g2_fill_1 FILLER_68_552 ();
 sg13g2_fill_1 FILLER_68_566 ();
 sg13g2_fill_2 FILLER_68_596 ();
 sg13g2_fill_2 FILLER_68_645 ();
 sg13g2_fill_1 FILLER_68_647 ();
 sg13g2_fill_2 FILLER_68_657 ();
 sg13g2_fill_2 FILLER_68_682 ();
 sg13g2_fill_1 FILLER_68_699 ();
 sg13g2_fill_1 FILLER_68_769 ();
 sg13g2_fill_1 FILLER_68_783 ();
 sg13g2_decap_8 FILLER_68_813 ();
 sg13g2_decap_4 FILLER_68_820 ();
 sg13g2_fill_1 FILLER_68_954 ();
 sg13g2_fill_1 FILLER_68_1004 ();
 sg13g2_fill_2 FILLER_68_1038 ();
 sg13g2_decap_8 FILLER_68_1084 ();
 sg13g2_fill_2 FILLER_68_1091 ();
 sg13g2_decap_4 FILLER_68_1102 ();
 sg13g2_fill_1 FILLER_68_1106 ();
 sg13g2_decap_4 FILLER_68_1111 ();
 sg13g2_fill_2 FILLER_68_1115 ();
 sg13g2_decap_8 FILLER_68_1125 ();
 sg13g2_fill_1 FILLER_68_1158 ();
 sg13g2_decap_8 FILLER_68_1171 ();
 sg13g2_decap_8 FILLER_68_1178 ();
 sg13g2_decap_8 FILLER_68_1185 ();
 sg13g2_decap_8 FILLER_68_1192 ();
 sg13g2_decap_8 FILLER_68_1199 ();
 sg13g2_decap_8 FILLER_68_1206 ();
 sg13g2_decap_8 FILLER_68_1213 ();
 sg13g2_decap_8 FILLER_68_1220 ();
 sg13g2_decap_8 FILLER_68_1227 ();
 sg13g2_decap_8 FILLER_68_1234 ();
 sg13g2_decap_8 FILLER_68_1241 ();
 sg13g2_decap_8 FILLER_68_1248 ();
 sg13g2_decap_8 FILLER_68_1255 ();
 sg13g2_decap_8 FILLER_68_1262 ();
 sg13g2_decap_8 FILLER_68_1269 ();
 sg13g2_decap_8 FILLER_68_1276 ();
 sg13g2_decap_8 FILLER_68_1283 ();
 sg13g2_decap_8 FILLER_68_1290 ();
 sg13g2_decap_8 FILLER_68_1297 ();
 sg13g2_decap_8 FILLER_68_1304 ();
 sg13g2_decap_4 FILLER_68_1311 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_7 ();
 sg13g2_fill_2 FILLER_69_38 ();
 sg13g2_fill_2 FILLER_69_43 ();
 sg13g2_fill_2 FILLER_69_50 ();
 sg13g2_fill_2 FILLER_69_57 ();
 sg13g2_fill_1 FILLER_69_82 ();
 sg13g2_fill_1 FILLER_69_87 ();
 sg13g2_decap_4 FILLER_69_105 ();
 sg13g2_fill_2 FILLER_69_109 ();
 sg13g2_decap_4 FILLER_69_115 ();
 sg13g2_fill_2 FILLER_69_119 ();
 sg13g2_fill_2 FILLER_69_135 ();
 sg13g2_fill_1 FILLER_69_175 ();
 sg13g2_fill_1 FILLER_69_180 ();
 sg13g2_fill_2 FILLER_69_185 ();
 sg13g2_fill_1 FILLER_69_187 ();
 sg13g2_fill_1 FILLER_69_233 ();
 sg13g2_fill_2 FILLER_69_249 ();
 sg13g2_fill_1 FILLER_69_251 ();
 sg13g2_fill_2 FILLER_69_257 ();
 sg13g2_fill_2 FILLER_69_264 ();
 sg13g2_decap_8 FILLER_69_316 ();
 sg13g2_fill_2 FILLER_69_333 ();
 sg13g2_fill_1 FILLER_69_361 ();
 sg13g2_fill_1 FILLER_69_393 ();
 sg13g2_fill_2 FILLER_69_420 ();
 sg13g2_fill_2 FILLER_69_430 ();
 sg13g2_fill_2 FILLER_69_441 ();
 sg13g2_fill_1 FILLER_69_452 ();
 sg13g2_fill_1 FILLER_69_505 ();
 sg13g2_fill_2 FILLER_69_516 ();
 sg13g2_fill_2 FILLER_69_522 ();
 sg13g2_fill_1 FILLER_69_524 ();
 sg13g2_fill_2 FILLER_69_530 ();
 sg13g2_decap_8 FILLER_69_536 ();
 sg13g2_fill_1 FILLER_69_572 ();
 sg13g2_fill_2 FILLER_69_579 ();
 sg13g2_fill_1 FILLER_69_589 ();
 sg13g2_decap_8 FILLER_69_616 ();
 sg13g2_decap_4 FILLER_69_623 ();
 sg13g2_fill_2 FILLER_69_627 ();
 sg13g2_fill_1 FILLER_69_664 ();
 sg13g2_fill_2 FILLER_69_708 ();
 sg13g2_fill_1 FILLER_69_736 ();
 sg13g2_fill_1 FILLER_69_745 ();
 sg13g2_decap_4 FILLER_69_772 ();
 sg13g2_fill_1 FILLER_69_776 ();
 sg13g2_fill_2 FILLER_69_786 ();
 sg13g2_fill_2 FILLER_69_801 ();
 sg13g2_fill_1 FILLER_69_803 ();
 sg13g2_fill_1 FILLER_69_886 ();
 sg13g2_decap_4 FILLER_69_903 ();
 sg13g2_fill_2 FILLER_69_907 ();
 sg13g2_fill_2 FILLER_69_944 ();
 sg13g2_fill_1 FILLER_69_983 ();
 sg13g2_fill_2 FILLER_69_989 ();
 sg13g2_fill_1 FILLER_69_991 ();
 sg13g2_fill_2 FILLER_69_1001 ();
 sg13g2_fill_2 FILLER_69_1035 ();
 sg13g2_fill_1 FILLER_69_1037 ();
 sg13g2_fill_2 FILLER_69_1065 ();
 sg13g2_fill_1 FILLER_69_1067 ();
 sg13g2_fill_2 FILLER_69_1072 ();
 sg13g2_fill_1 FILLER_69_1074 ();
 sg13g2_fill_2 FILLER_69_1150 ();
 sg13g2_decap_8 FILLER_69_1178 ();
 sg13g2_decap_8 FILLER_69_1185 ();
 sg13g2_decap_8 FILLER_69_1192 ();
 sg13g2_decap_8 FILLER_69_1199 ();
 sg13g2_decap_8 FILLER_69_1206 ();
 sg13g2_decap_8 FILLER_69_1213 ();
 sg13g2_decap_8 FILLER_69_1220 ();
 sg13g2_decap_8 FILLER_69_1227 ();
 sg13g2_decap_8 FILLER_69_1234 ();
 sg13g2_decap_8 FILLER_69_1241 ();
 sg13g2_decap_8 FILLER_69_1248 ();
 sg13g2_decap_8 FILLER_69_1255 ();
 sg13g2_decap_8 FILLER_69_1262 ();
 sg13g2_decap_8 FILLER_69_1269 ();
 sg13g2_decap_8 FILLER_69_1276 ();
 sg13g2_decap_8 FILLER_69_1283 ();
 sg13g2_decap_8 FILLER_69_1290 ();
 sg13g2_decap_8 FILLER_69_1297 ();
 sg13g2_decap_8 FILLER_69_1304 ();
 sg13g2_decap_4 FILLER_69_1311 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_4 FILLER_70_14 ();
 sg13g2_fill_2 FILLER_70_18 ();
 sg13g2_fill_2 FILLER_70_59 ();
 sg13g2_fill_1 FILLER_70_61 ();
 sg13g2_fill_2 FILLER_70_71 ();
 sg13g2_fill_1 FILLER_70_87 ();
 sg13g2_fill_2 FILLER_70_97 ();
 sg13g2_fill_1 FILLER_70_99 ();
 sg13g2_fill_2 FILLER_70_104 ();
 sg13g2_fill_2 FILLER_70_170 ();
 sg13g2_fill_1 FILLER_70_172 ();
 sg13g2_fill_2 FILLER_70_178 ();
 sg13g2_fill_1 FILLER_70_180 ();
 sg13g2_fill_2 FILLER_70_212 ();
 sg13g2_fill_1 FILLER_70_214 ();
 sg13g2_fill_1 FILLER_70_223 ();
 sg13g2_fill_2 FILLER_70_258 ();
 sg13g2_fill_1 FILLER_70_260 ();
 sg13g2_fill_1 FILLER_70_325 ();
 sg13g2_fill_1 FILLER_70_421 ();
 sg13g2_fill_1 FILLER_70_458 ();
 sg13g2_fill_1 FILLER_70_468 ();
 sg13g2_decap_4 FILLER_70_473 ();
 sg13g2_fill_1 FILLER_70_505 ();
 sg13g2_fill_2 FILLER_70_514 ();
 sg13g2_fill_2 FILLER_70_609 ();
 sg13g2_fill_1 FILLER_70_611 ();
 sg13g2_fill_1 FILLER_70_701 ();
 sg13g2_fill_2 FILLER_70_711 ();
 sg13g2_fill_2 FILLER_70_745 ();
 sg13g2_fill_1 FILLER_70_747 ();
 sg13g2_fill_1 FILLER_70_757 ();
 sg13g2_fill_1 FILLER_70_793 ();
 sg13g2_decap_8 FILLER_70_797 ();
 sg13g2_fill_1 FILLER_70_804 ();
 sg13g2_fill_2 FILLER_70_865 ();
 sg13g2_fill_2 FILLER_70_893 ();
 sg13g2_fill_1 FILLER_70_895 ();
 sg13g2_fill_2 FILLER_70_1061 ();
 sg13g2_fill_1 FILLER_70_1063 ();
 sg13g2_fill_2 FILLER_70_1087 ();
 sg13g2_fill_1 FILLER_70_1089 ();
 sg13g2_fill_2 FILLER_70_1111 ();
 sg13g2_fill_1 FILLER_70_1113 ();
 sg13g2_fill_1 FILLER_70_1119 ();
 sg13g2_fill_1 FILLER_70_1129 ();
 sg13g2_fill_1 FILLER_70_1144 ();
 sg13g2_fill_2 FILLER_70_1158 ();
 sg13g2_decap_8 FILLER_70_1178 ();
 sg13g2_decap_8 FILLER_70_1185 ();
 sg13g2_decap_8 FILLER_70_1192 ();
 sg13g2_decap_8 FILLER_70_1199 ();
 sg13g2_decap_8 FILLER_70_1206 ();
 sg13g2_decap_8 FILLER_70_1213 ();
 sg13g2_decap_8 FILLER_70_1220 ();
 sg13g2_decap_8 FILLER_70_1227 ();
 sg13g2_decap_8 FILLER_70_1234 ();
 sg13g2_decap_8 FILLER_70_1241 ();
 sg13g2_decap_8 FILLER_70_1248 ();
 sg13g2_decap_8 FILLER_70_1255 ();
 sg13g2_decap_8 FILLER_70_1262 ();
 sg13g2_decap_8 FILLER_70_1269 ();
 sg13g2_decap_8 FILLER_70_1276 ();
 sg13g2_decap_8 FILLER_70_1283 ();
 sg13g2_decap_8 FILLER_70_1290 ();
 sg13g2_decap_8 FILLER_70_1297 ();
 sg13g2_decap_8 FILLER_70_1304 ();
 sg13g2_decap_4 FILLER_70_1311 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_4 FILLER_71_7 ();
 sg13g2_fill_1 FILLER_71_11 ();
 sg13g2_fill_1 FILLER_71_38 ();
 sg13g2_fill_1 FILLER_71_57 ();
 sg13g2_fill_1 FILLER_71_123 ();
 sg13g2_fill_2 FILLER_71_168 ();
 sg13g2_fill_1 FILLER_71_170 ();
 sg13g2_fill_1 FILLER_71_176 ();
 sg13g2_fill_1 FILLER_71_185 ();
 sg13g2_decap_8 FILLER_71_217 ();
 sg13g2_decap_8 FILLER_71_233 ();
 sg13g2_decap_8 FILLER_71_240 ();
 sg13g2_fill_2 FILLER_71_247 ();
 sg13g2_fill_1 FILLER_71_249 ();
 sg13g2_fill_1 FILLER_71_304 ();
 sg13g2_fill_1 FILLER_71_319 ();
 sg13g2_fill_2 FILLER_71_330 ();
 sg13g2_fill_1 FILLER_71_332 ();
 sg13g2_fill_2 FILLER_71_359 ();
 sg13g2_fill_2 FILLER_71_375 ();
 sg13g2_fill_2 FILLER_71_434 ();
 sg13g2_fill_1 FILLER_71_453 ();
 sg13g2_fill_2 FILLER_71_512 ();
 sg13g2_fill_2 FILLER_71_530 ();
 sg13g2_fill_1 FILLER_71_532 ();
 sg13g2_fill_2 FILLER_71_585 ();
 sg13g2_decap_4 FILLER_71_613 ();
 sg13g2_fill_1 FILLER_71_648 ();
 sg13g2_decap_8 FILLER_71_659 ();
 sg13g2_fill_1 FILLER_71_666 ();
 sg13g2_fill_1 FILLER_71_672 ();
 sg13g2_fill_2 FILLER_71_687 ();
 sg13g2_fill_1 FILLER_71_709 ();
 sg13g2_fill_1 FILLER_71_736 ();
 sg13g2_fill_2 FILLER_71_774 ();
 sg13g2_fill_2 FILLER_71_821 ();
 sg13g2_fill_1 FILLER_71_823 ();
 sg13g2_fill_2 FILLER_71_836 ();
 sg13g2_fill_1 FILLER_71_838 ();
 sg13g2_fill_1 FILLER_71_852 ();
 sg13g2_fill_2 FILLER_71_912 ();
 sg13g2_fill_1 FILLER_71_918 ();
 sg13g2_fill_1 FILLER_71_942 ();
 sg13g2_fill_2 FILLER_71_960 ();
 sg13g2_fill_2 FILLER_71_967 ();
 sg13g2_fill_1 FILLER_71_969 ();
 sg13g2_fill_1 FILLER_71_978 ();
 sg13g2_fill_1 FILLER_71_988 ();
 sg13g2_fill_1 FILLER_71_1014 ();
 sg13g2_fill_1 FILLER_71_1054 ();
 sg13g2_fill_2 FILLER_71_1084 ();
 sg13g2_fill_1 FILLER_71_1086 ();
 sg13g2_fill_1 FILLER_71_1126 ();
 sg13g2_fill_2 FILLER_71_1137 ();
 sg13g2_fill_1 FILLER_71_1139 ();
 sg13g2_decap_8 FILLER_71_1179 ();
 sg13g2_decap_8 FILLER_71_1186 ();
 sg13g2_decap_8 FILLER_71_1193 ();
 sg13g2_decap_8 FILLER_71_1200 ();
 sg13g2_decap_8 FILLER_71_1207 ();
 sg13g2_decap_8 FILLER_71_1214 ();
 sg13g2_decap_8 FILLER_71_1221 ();
 sg13g2_decap_8 FILLER_71_1228 ();
 sg13g2_decap_8 FILLER_71_1235 ();
 sg13g2_decap_8 FILLER_71_1242 ();
 sg13g2_decap_8 FILLER_71_1249 ();
 sg13g2_decap_8 FILLER_71_1256 ();
 sg13g2_decap_8 FILLER_71_1263 ();
 sg13g2_decap_8 FILLER_71_1270 ();
 sg13g2_decap_8 FILLER_71_1277 ();
 sg13g2_decap_8 FILLER_71_1284 ();
 sg13g2_decap_8 FILLER_71_1291 ();
 sg13g2_decap_8 FILLER_71_1298 ();
 sg13g2_decap_8 FILLER_71_1305 ();
 sg13g2_fill_2 FILLER_71_1312 ();
 sg13g2_fill_1 FILLER_71_1314 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_fill_1 FILLER_72_21 ();
 sg13g2_fill_2 FILLER_72_35 ();
 sg13g2_fill_1 FILLER_72_45 ();
 sg13g2_fill_2 FILLER_72_67 ();
 sg13g2_decap_4 FILLER_72_88 ();
 sg13g2_fill_2 FILLER_72_92 ();
 sg13g2_fill_2 FILLER_72_126 ();
 sg13g2_fill_1 FILLER_72_128 ();
 sg13g2_fill_2 FILLER_72_138 ();
 sg13g2_fill_1 FILLER_72_180 ();
 sg13g2_fill_1 FILLER_72_238 ();
 sg13g2_fill_1 FILLER_72_247 ();
 sg13g2_fill_1 FILLER_72_278 ();
 sg13g2_decap_4 FILLER_72_283 ();
 sg13g2_fill_2 FILLER_72_287 ();
 sg13g2_fill_1 FILLER_72_294 ();
 sg13g2_fill_2 FILLER_72_322 ();
 sg13g2_fill_1 FILLER_72_324 ();
 sg13g2_fill_2 FILLER_72_404 ();
 sg13g2_fill_1 FILLER_72_415 ();
 sg13g2_decap_4 FILLER_72_438 ();
 sg13g2_fill_2 FILLER_72_442 ();
 sg13g2_fill_1 FILLER_72_493 ();
 sg13g2_decap_4 FILLER_72_499 ();
 sg13g2_decap_4 FILLER_72_510 ();
 sg13g2_fill_2 FILLER_72_522 ();
 sg13g2_fill_2 FILLER_72_533 ();
 sg13g2_fill_1 FILLER_72_557 ();
 sg13g2_fill_1 FILLER_72_567 ();
 sg13g2_fill_2 FILLER_72_573 ();
 sg13g2_fill_1 FILLER_72_586 ();
 sg13g2_fill_1 FILLER_72_655 ();
 sg13g2_fill_1 FILLER_72_662 ();
 sg13g2_decap_4 FILLER_72_668 ();
 sg13g2_fill_1 FILLER_72_688 ();
 sg13g2_decap_8 FILLER_72_705 ();
 sg13g2_fill_1 FILLER_72_712 ();
 sg13g2_fill_2 FILLER_72_718 ();
 sg13g2_fill_1 FILLER_72_720 ();
 sg13g2_decap_8 FILLER_72_728 ();
 sg13g2_fill_1 FILLER_72_738 ();
 sg13g2_fill_1 FILLER_72_749 ();
 sg13g2_fill_1 FILLER_72_791 ();
 sg13g2_fill_1 FILLER_72_797 ();
 sg13g2_decap_4 FILLER_72_802 ();
 sg13g2_fill_2 FILLER_72_819 ();
 sg13g2_fill_2 FILLER_72_831 ();
 sg13g2_decap_8 FILLER_72_896 ();
 sg13g2_fill_2 FILLER_72_903 ();
 sg13g2_fill_1 FILLER_72_905 ();
 sg13g2_fill_2 FILLER_72_910 ();
 sg13g2_fill_2 FILLER_72_917 ();
 sg13g2_decap_4 FILLER_72_958 ();
 sg13g2_fill_2 FILLER_72_1011 ();
 sg13g2_fill_2 FILLER_72_1048 ();
 sg13g2_fill_1 FILLER_72_1059 ();
 sg13g2_fill_2 FILLER_72_1072 ();
 sg13g2_decap_8 FILLER_72_1098 ();
 sg13g2_fill_2 FILLER_72_1105 ();
 sg13g2_fill_1 FILLER_72_1107 ();
 sg13g2_fill_1 FILLER_72_1120 ();
 sg13g2_decap_4 FILLER_72_1126 ();
 sg13g2_fill_2 FILLER_72_1130 ();
 sg13g2_fill_2 FILLER_72_1155 ();
 sg13g2_decap_8 FILLER_72_1174 ();
 sg13g2_decap_8 FILLER_72_1181 ();
 sg13g2_decap_8 FILLER_72_1188 ();
 sg13g2_decap_8 FILLER_72_1195 ();
 sg13g2_decap_8 FILLER_72_1202 ();
 sg13g2_decap_8 FILLER_72_1209 ();
 sg13g2_decap_8 FILLER_72_1216 ();
 sg13g2_decap_8 FILLER_72_1223 ();
 sg13g2_decap_8 FILLER_72_1230 ();
 sg13g2_decap_8 FILLER_72_1237 ();
 sg13g2_decap_8 FILLER_72_1244 ();
 sg13g2_decap_8 FILLER_72_1251 ();
 sg13g2_decap_8 FILLER_72_1258 ();
 sg13g2_decap_8 FILLER_72_1265 ();
 sg13g2_decap_8 FILLER_72_1272 ();
 sg13g2_decap_8 FILLER_72_1279 ();
 sg13g2_decap_8 FILLER_72_1286 ();
 sg13g2_decap_8 FILLER_72_1293 ();
 sg13g2_decap_8 FILLER_72_1300 ();
 sg13g2_decap_8 FILLER_72_1307 ();
 sg13g2_fill_1 FILLER_72_1314 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_fill_2 FILLER_73_160 ();
 sg13g2_fill_1 FILLER_73_162 ();
 sg13g2_fill_1 FILLER_73_172 ();
 sg13g2_decap_4 FILLER_73_223 ();
 sg13g2_fill_1 FILLER_73_244 ();
 sg13g2_fill_1 FILLER_73_258 ();
 sg13g2_fill_1 FILLER_73_263 ();
 sg13g2_decap_4 FILLER_73_277 ();
 sg13g2_fill_1 FILLER_73_281 ();
 sg13g2_decap_4 FILLER_73_286 ();
 sg13g2_fill_2 FILLER_73_290 ();
 sg13g2_fill_2 FILLER_73_310 ();
 sg13g2_fill_1 FILLER_73_338 ();
 sg13g2_fill_1 FILLER_73_343 ();
 sg13g2_fill_1 FILLER_73_436 ();
 sg13g2_fill_1 FILLER_73_453 ();
 sg13g2_decap_8 FILLER_73_464 ();
 sg13g2_decap_4 FILLER_73_471 ();
 sg13g2_decap_8 FILLER_73_681 ();
 sg13g2_fill_1 FILLER_73_688 ();
 sg13g2_fill_1 FILLER_73_692 ();
 sg13g2_fill_2 FILLER_73_701 ();
 sg13g2_fill_1 FILLER_73_738 ();
 sg13g2_fill_2 FILLER_73_768 ();
 sg13g2_fill_1 FILLER_73_809 ();
 sg13g2_decap_4 FILLER_73_826 ();
 sg13g2_fill_2 FILLER_73_830 ();
 sg13g2_fill_1 FILLER_73_836 ();
 sg13g2_fill_2 FILLER_73_882 ();
 sg13g2_decap_4 FILLER_73_888 ();
 sg13g2_fill_2 FILLER_73_892 ();
 sg13g2_fill_2 FILLER_73_944 ();
 sg13g2_fill_2 FILLER_73_972 ();
 sg13g2_fill_1 FILLER_73_998 ();
 sg13g2_fill_2 FILLER_73_1025 ();
 sg13g2_fill_2 FILLER_73_1109 ();
 sg13g2_fill_1 FILLER_73_1111 ();
 sg13g2_decap_8 FILLER_73_1181 ();
 sg13g2_decap_8 FILLER_73_1188 ();
 sg13g2_decap_8 FILLER_73_1195 ();
 sg13g2_decap_8 FILLER_73_1202 ();
 sg13g2_decap_8 FILLER_73_1209 ();
 sg13g2_decap_8 FILLER_73_1216 ();
 sg13g2_decap_8 FILLER_73_1223 ();
 sg13g2_decap_8 FILLER_73_1230 ();
 sg13g2_decap_8 FILLER_73_1237 ();
 sg13g2_decap_8 FILLER_73_1244 ();
 sg13g2_decap_8 FILLER_73_1251 ();
 sg13g2_decap_8 FILLER_73_1258 ();
 sg13g2_decap_8 FILLER_73_1265 ();
 sg13g2_decap_8 FILLER_73_1272 ();
 sg13g2_decap_8 FILLER_73_1279 ();
 sg13g2_decap_8 FILLER_73_1286 ();
 sg13g2_decap_8 FILLER_73_1293 ();
 sg13g2_decap_8 FILLER_73_1300 ();
 sg13g2_decap_8 FILLER_73_1307 ();
 sg13g2_fill_1 FILLER_73_1314 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_4 FILLER_74_35 ();
 sg13g2_fill_2 FILLER_74_39 ();
 sg13g2_fill_1 FILLER_74_54 ();
 sg13g2_fill_1 FILLER_74_84 ();
 sg13g2_fill_2 FILLER_74_146 ();
 sg13g2_fill_1 FILLER_74_210 ();
 sg13g2_fill_1 FILLER_74_330 ();
 sg13g2_fill_2 FILLER_74_388 ();
 sg13g2_fill_2 FILLER_74_421 ();
 sg13g2_fill_2 FILLER_74_469 ();
 sg13g2_fill_2 FILLER_74_520 ();
 sg13g2_fill_2 FILLER_74_551 ();
 sg13g2_fill_1 FILLER_74_569 ();
 sg13g2_fill_2 FILLER_74_594 ();
 sg13g2_fill_1 FILLER_74_596 ();
 sg13g2_fill_2 FILLER_74_612 ();
 sg13g2_fill_2 FILLER_74_656 ();
 sg13g2_fill_1 FILLER_74_663 ();
 sg13g2_fill_1 FILLER_74_670 ();
 sg13g2_decap_8 FILLER_74_675 ();
 sg13g2_fill_1 FILLER_74_682 ();
 sg13g2_decap_4 FILLER_74_708 ();
 sg13g2_fill_1 FILLER_74_712 ();
 sg13g2_decap_8 FILLER_74_721 ();
 sg13g2_fill_2 FILLER_74_728 ();
 sg13g2_fill_2 FILLER_74_756 ();
 sg13g2_decap_4 FILLER_74_795 ();
 sg13g2_fill_2 FILLER_74_799 ();
 sg13g2_fill_2 FILLER_74_806 ();
 sg13g2_fill_1 FILLER_74_816 ();
 sg13g2_fill_1 FILLER_74_849 ();
 sg13g2_fill_2 FILLER_74_864 ();
 sg13g2_fill_1 FILLER_74_892 ();
 sg13g2_fill_2 FILLER_74_898 ();
 sg13g2_fill_1 FILLER_74_915 ();
 sg13g2_fill_2 FILLER_74_921 ();
 sg13g2_fill_1 FILLER_74_923 ();
 sg13g2_fill_2 FILLER_74_945 ();
 sg13g2_decap_4 FILLER_74_961 ();
 sg13g2_fill_2 FILLER_74_1000 ();
 sg13g2_fill_2 FILLER_74_1043 ();
 sg13g2_fill_1 FILLER_74_1074 ();
 sg13g2_decap_4 FILLER_74_1089 ();
 sg13g2_fill_1 FILLER_74_1093 ();
 sg13g2_decap_8 FILLER_74_1098 ();
 sg13g2_decap_8 FILLER_74_1105 ();
 sg13g2_fill_1 FILLER_74_1112 ();
 sg13g2_fill_1 FILLER_74_1118 ();
 sg13g2_decap_8 FILLER_74_1181 ();
 sg13g2_decap_8 FILLER_74_1188 ();
 sg13g2_decap_8 FILLER_74_1195 ();
 sg13g2_decap_8 FILLER_74_1202 ();
 sg13g2_decap_8 FILLER_74_1209 ();
 sg13g2_decap_8 FILLER_74_1216 ();
 sg13g2_decap_8 FILLER_74_1223 ();
 sg13g2_decap_8 FILLER_74_1230 ();
 sg13g2_decap_8 FILLER_74_1237 ();
 sg13g2_decap_8 FILLER_74_1244 ();
 sg13g2_decap_8 FILLER_74_1251 ();
 sg13g2_decap_8 FILLER_74_1258 ();
 sg13g2_decap_8 FILLER_74_1265 ();
 sg13g2_decap_8 FILLER_74_1272 ();
 sg13g2_decap_8 FILLER_74_1279 ();
 sg13g2_decap_8 FILLER_74_1286 ();
 sg13g2_decap_8 FILLER_74_1293 ();
 sg13g2_decap_8 FILLER_74_1300 ();
 sg13g2_decap_8 FILLER_74_1307 ();
 sg13g2_fill_1 FILLER_74_1314 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_fill_2 FILLER_75_42 ();
 sg13g2_fill_1 FILLER_75_44 ();
 sg13g2_decap_8 FILLER_75_75 ();
 sg13g2_decap_8 FILLER_75_82 ();
 sg13g2_decap_8 FILLER_75_89 ();
 sg13g2_decap_4 FILLER_75_96 ();
 sg13g2_fill_1 FILLER_75_126 ();
 sg13g2_fill_2 FILLER_75_145 ();
 sg13g2_fill_1 FILLER_75_165 ();
 sg13g2_fill_2 FILLER_75_171 ();
 sg13g2_fill_1 FILLER_75_185 ();
 sg13g2_fill_1 FILLER_75_190 ();
 sg13g2_decap_4 FILLER_75_203 ();
 sg13g2_fill_1 FILLER_75_207 ();
 sg13g2_fill_2 FILLER_75_243 ();
 sg13g2_fill_2 FILLER_75_254 ();
 sg13g2_fill_2 FILLER_75_297 ();
 sg13g2_fill_1 FILLER_75_299 ();
 sg13g2_decap_4 FILLER_75_318 ();
 sg13g2_fill_2 FILLER_75_322 ();
 sg13g2_fill_1 FILLER_75_350 ();
 sg13g2_fill_2 FILLER_75_401 ();
 sg13g2_fill_2 FILLER_75_443 ();
 sg13g2_fill_1 FILLER_75_458 ();
 sg13g2_fill_2 FILLER_75_577 ();
 sg13g2_fill_1 FILLER_75_605 ();
 sg13g2_fill_2 FILLER_75_615 ();
 sg13g2_decap_4 FILLER_75_685 ();
 sg13g2_decap_8 FILLER_75_694 ();
 sg13g2_fill_2 FILLER_75_736 ();
 sg13g2_fill_2 FILLER_75_748 ();
 sg13g2_fill_1 FILLER_75_754 ();
 sg13g2_fill_2 FILLER_75_802 ();
 sg13g2_fill_1 FILLER_75_804 ();
 sg13g2_fill_1 FILLER_75_826 ();
 sg13g2_fill_2 FILLER_75_844 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_fill_1 FILLER_75_882 ();
 sg13g2_fill_2 FILLER_75_910 ();
 sg13g2_fill_1 FILLER_75_912 ();
 sg13g2_fill_2 FILLER_75_972 ();
 sg13g2_fill_1 FILLER_75_974 ();
 sg13g2_fill_2 FILLER_75_980 ();
 sg13g2_fill_1 FILLER_75_1016 ();
 sg13g2_fill_1 FILLER_75_1043 ();
 sg13g2_fill_2 FILLER_75_1052 ();
 sg13g2_fill_1 FILLER_75_1054 ();
 sg13g2_fill_2 FILLER_75_1114 ();
 sg13g2_fill_1 FILLER_75_1116 ();
 sg13g2_fill_1 FILLER_75_1129 ();
 sg13g2_decap_8 FILLER_75_1177 ();
 sg13g2_decap_8 FILLER_75_1184 ();
 sg13g2_decap_8 FILLER_75_1191 ();
 sg13g2_decap_8 FILLER_75_1198 ();
 sg13g2_decap_8 FILLER_75_1205 ();
 sg13g2_decap_8 FILLER_75_1212 ();
 sg13g2_decap_8 FILLER_75_1219 ();
 sg13g2_decap_8 FILLER_75_1226 ();
 sg13g2_decap_8 FILLER_75_1233 ();
 sg13g2_decap_8 FILLER_75_1240 ();
 sg13g2_decap_8 FILLER_75_1247 ();
 sg13g2_decap_8 FILLER_75_1254 ();
 sg13g2_decap_8 FILLER_75_1261 ();
 sg13g2_decap_8 FILLER_75_1268 ();
 sg13g2_decap_8 FILLER_75_1275 ();
 sg13g2_decap_8 FILLER_75_1282 ();
 sg13g2_decap_8 FILLER_75_1289 ();
 sg13g2_decap_8 FILLER_75_1296 ();
 sg13g2_decap_8 FILLER_75_1303 ();
 sg13g2_decap_4 FILLER_75_1310 ();
 sg13g2_fill_1 FILLER_75_1314 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_4 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_64 ();
 sg13g2_decap_8 FILLER_76_71 ();
 sg13g2_decap_8 FILLER_76_78 ();
 sg13g2_decap_8 FILLER_76_85 ();
 sg13g2_decap_8 FILLER_76_92 ();
 sg13g2_decap_8 FILLER_76_99 ();
 sg13g2_fill_2 FILLER_76_132 ();
 sg13g2_fill_1 FILLER_76_134 ();
 sg13g2_fill_2 FILLER_76_210 ();
 sg13g2_fill_1 FILLER_76_212 ();
 sg13g2_fill_1 FILLER_76_218 ();
 sg13g2_fill_1 FILLER_76_402 ();
 sg13g2_fill_2 FILLER_76_452 ();
 sg13g2_fill_2 FILLER_76_467 ();
 sg13g2_fill_1 FILLER_76_469 ();
 sg13g2_fill_1 FILLER_76_474 ();
 sg13g2_fill_1 FILLER_76_484 ();
 sg13g2_fill_1 FILLER_76_508 ();
 sg13g2_fill_1 FILLER_76_514 ();
 sg13g2_fill_2 FILLER_76_551 ();
 sg13g2_fill_2 FILLER_76_580 ();
 sg13g2_fill_2 FILLER_76_596 ();
 sg13g2_fill_1 FILLER_76_665 ();
 sg13g2_decap_4 FILLER_76_697 ();
 sg13g2_fill_2 FILLER_76_701 ();
 sg13g2_decap_4 FILLER_76_706 ();
 sg13g2_fill_1 FILLER_76_710 ();
 sg13g2_fill_2 FILLER_76_719 ();
 sg13g2_fill_1 FILLER_76_783 ();
 sg13g2_fill_2 FILLER_76_802 ();
 sg13g2_fill_1 FILLER_76_816 ();
 sg13g2_decap_8 FILLER_76_877 ();
 sg13g2_decap_4 FILLER_76_896 ();
 sg13g2_fill_2 FILLER_76_939 ();
 sg13g2_fill_1 FILLER_76_941 ();
 sg13g2_fill_2 FILLER_76_1035 ();
 sg13g2_fill_2 FILLER_76_1066 ();
 sg13g2_fill_2 FILLER_76_1075 ();
 sg13g2_fill_2 FILLER_76_1101 ();
 sg13g2_fill_1 FILLER_76_1103 ();
 sg13g2_fill_1 FILLER_76_1130 ();
 sg13g2_fill_2 FILLER_76_1150 ();
 sg13g2_fill_1 FILLER_76_1152 ();
 sg13g2_decap_8 FILLER_76_1169 ();
 sg13g2_decap_8 FILLER_76_1176 ();
 sg13g2_decap_8 FILLER_76_1183 ();
 sg13g2_decap_8 FILLER_76_1190 ();
 sg13g2_decap_8 FILLER_76_1197 ();
 sg13g2_decap_8 FILLER_76_1204 ();
 sg13g2_decap_8 FILLER_76_1211 ();
 sg13g2_decap_8 FILLER_76_1218 ();
 sg13g2_decap_8 FILLER_76_1225 ();
 sg13g2_decap_8 FILLER_76_1232 ();
 sg13g2_decap_8 FILLER_76_1239 ();
 sg13g2_decap_8 FILLER_76_1246 ();
 sg13g2_decap_8 FILLER_76_1253 ();
 sg13g2_decap_8 FILLER_76_1260 ();
 sg13g2_decap_8 FILLER_76_1267 ();
 sg13g2_decap_8 FILLER_76_1274 ();
 sg13g2_decap_8 FILLER_76_1281 ();
 sg13g2_decap_8 FILLER_76_1288 ();
 sg13g2_decap_8 FILLER_76_1295 ();
 sg13g2_decap_8 FILLER_76_1302 ();
 sg13g2_decap_4 FILLER_76_1309 ();
 sg13g2_fill_2 FILLER_76_1313 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_4 FILLER_77_105 ();
 sg13g2_fill_2 FILLER_77_109 ();
 sg13g2_fill_2 FILLER_77_115 ();
 sg13g2_decap_8 FILLER_77_121 ();
 sg13g2_fill_2 FILLER_77_128 ();
 sg13g2_fill_1 FILLER_77_130 ();
 sg13g2_fill_1 FILLER_77_208 ();
 sg13g2_fill_2 FILLER_77_227 ();
 sg13g2_fill_1 FILLER_77_229 ();
 sg13g2_fill_2 FILLER_77_238 ();
 sg13g2_fill_2 FILLER_77_259 ();
 sg13g2_fill_1 FILLER_77_265 ();
 sg13g2_fill_2 FILLER_77_291 ();
 sg13g2_fill_1 FILLER_77_293 ();
 sg13g2_decap_4 FILLER_77_308 ();
 sg13g2_fill_1 FILLER_77_312 ();
 sg13g2_decap_8 FILLER_77_317 ();
 sg13g2_fill_1 FILLER_77_343 ();
 sg13g2_fill_2 FILLER_77_414 ();
 sg13g2_fill_2 FILLER_77_460 ();
 sg13g2_fill_1 FILLER_77_488 ();
 sg13g2_fill_2 FILLER_77_512 ();
 sg13g2_fill_1 FILLER_77_534 ();
 sg13g2_fill_1 FILLER_77_624 ();
 sg13g2_fill_1 FILLER_77_640 ();
 sg13g2_fill_2 FILLER_77_671 ();
 sg13g2_decap_4 FILLER_77_694 ();
 sg13g2_fill_2 FILLER_77_698 ();
 sg13g2_fill_1 FILLER_77_740 ();
 sg13g2_decap_8 FILLER_77_745 ();
 sg13g2_fill_1 FILLER_77_752 ();
 sg13g2_fill_1 FILLER_77_785 ();
 sg13g2_fill_2 FILLER_77_804 ();
 sg13g2_fill_2 FILLER_77_818 ();
 sg13g2_fill_2 FILLER_77_829 ();
 sg13g2_fill_1 FILLER_77_834 ();
 sg13g2_fill_2 FILLER_77_847 ();
 sg13g2_decap_4 FILLER_77_859 ();
 sg13g2_fill_2 FILLER_77_863 ();
 sg13g2_decap_8 FILLER_77_875 ();
 sg13g2_fill_2 FILLER_77_909 ();
 sg13g2_fill_2 FILLER_77_915 ();
 sg13g2_fill_2 FILLER_77_925 ();
 sg13g2_fill_1 FILLER_77_927 ();
 sg13g2_fill_2 FILLER_77_934 ();
 sg13g2_fill_1 FILLER_77_979 ();
 sg13g2_fill_1 FILLER_77_994 ();
 sg13g2_fill_2 FILLER_77_1074 ();
 sg13g2_fill_1 FILLER_77_1076 ();
 sg13g2_fill_2 FILLER_77_1108 ();
 sg13g2_fill_2 FILLER_77_1113 ();
 sg13g2_fill_1 FILLER_77_1119 ();
 sg13g2_decap_8 FILLER_77_1170 ();
 sg13g2_decap_8 FILLER_77_1177 ();
 sg13g2_decap_8 FILLER_77_1184 ();
 sg13g2_decap_8 FILLER_77_1191 ();
 sg13g2_decap_8 FILLER_77_1198 ();
 sg13g2_decap_8 FILLER_77_1205 ();
 sg13g2_decap_8 FILLER_77_1212 ();
 sg13g2_decap_8 FILLER_77_1219 ();
 sg13g2_decap_8 FILLER_77_1226 ();
 sg13g2_decap_8 FILLER_77_1233 ();
 sg13g2_decap_8 FILLER_77_1240 ();
 sg13g2_decap_8 FILLER_77_1247 ();
 sg13g2_decap_8 FILLER_77_1254 ();
 sg13g2_decap_8 FILLER_77_1261 ();
 sg13g2_decap_8 FILLER_77_1268 ();
 sg13g2_decap_8 FILLER_77_1275 ();
 sg13g2_decap_8 FILLER_77_1282 ();
 sg13g2_decap_8 FILLER_77_1289 ();
 sg13g2_decap_8 FILLER_77_1296 ();
 sg13g2_decap_8 FILLER_77_1303 ();
 sg13g2_decap_4 FILLER_77_1310 ();
 sg13g2_fill_1 FILLER_77_1314 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_fill_1 FILLER_78_142 ();
 sg13g2_fill_2 FILLER_78_148 ();
 sg13g2_fill_1 FILLER_78_155 ();
 sg13g2_fill_2 FILLER_78_179 ();
 sg13g2_fill_1 FILLER_78_181 ();
 sg13g2_fill_1 FILLER_78_199 ();
 sg13g2_fill_2 FILLER_78_232 ();
 sg13g2_fill_1 FILLER_78_234 ();
 sg13g2_fill_2 FILLER_78_251 ();
 sg13g2_fill_1 FILLER_78_274 ();
 sg13g2_fill_2 FILLER_78_302 ();
 sg13g2_fill_1 FILLER_78_304 ();
 sg13g2_fill_2 FILLER_78_434 ();
 sg13g2_fill_1 FILLER_78_436 ();
 sg13g2_decap_4 FILLER_78_479 ();
 sg13g2_fill_2 FILLER_78_526 ();
 sg13g2_fill_1 FILLER_78_581 ();
 sg13g2_fill_2 FILLER_78_616 ();
 sg13g2_fill_2 FILLER_78_632 ();
 sg13g2_fill_1 FILLER_78_674 ();
 sg13g2_decap_8 FILLER_78_706 ();
 sg13g2_decap_8 FILLER_78_713 ();
 sg13g2_decap_8 FILLER_78_720 ();
 sg13g2_fill_2 FILLER_78_727 ();
 sg13g2_fill_1 FILLER_78_729 ();
 sg13g2_fill_2 FILLER_78_774 ();
 sg13g2_fill_1 FILLER_78_798 ();
 sg13g2_fill_2 FILLER_78_822 ();
 sg13g2_fill_1 FILLER_78_824 ();
 sg13g2_fill_2 FILLER_78_843 ();
 sg13g2_decap_8 FILLER_78_955 ();
 sg13g2_decap_8 FILLER_78_962 ();
 sg13g2_fill_2 FILLER_78_978 ();
 sg13g2_fill_1 FILLER_78_999 ();
 sg13g2_fill_1 FILLER_78_1039 ();
 sg13g2_fill_1 FILLER_78_1047 ();
 sg13g2_fill_1 FILLER_78_1064 ();
 sg13g2_fill_2 FILLER_78_1089 ();
 sg13g2_fill_1 FILLER_78_1112 ();
 sg13g2_fill_1 FILLER_78_1139 ();
 sg13g2_decap_8 FILLER_78_1170 ();
 sg13g2_decap_8 FILLER_78_1177 ();
 sg13g2_decap_8 FILLER_78_1184 ();
 sg13g2_decap_8 FILLER_78_1191 ();
 sg13g2_decap_8 FILLER_78_1198 ();
 sg13g2_decap_8 FILLER_78_1205 ();
 sg13g2_decap_8 FILLER_78_1212 ();
 sg13g2_decap_8 FILLER_78_1219 ();
 sg13g2_decap_8 FILLER_78_1226 ();
 sg13g2_decap_8 FILLER_78_1233 ();
 sg13g2_decap_8 FILLER_78_1240 ();
 sg13g2_decap_8 FILLER_78_1247 ();
 sg13g2_decap_8 FILLER_78_1254 ();
 sg13g2_decap_8 FILLER_78_1261 ();
 sg13g2_decap_8 FILLER_78_1268 ();
 sg13g2_decap_8 FILLER_78_1275 ();
 sg13g2_decap_8 FILLER_78_1282 ();
 sg13g2_decap_8 FILLER_78_1289 ();
 sg13g2_decap_8 FILLER_78_1296 ();
 sg13g2_decap_8 FILLER_78_1303 ();
 sg13g2_decap_4 FILLER_78_1310 ();
 sg13g2_fill_1 FILLER_78_1314 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_fill_1 FILLER_79_171 ();
 sg13g2_fill_1 FILLER_79_231 ();
 sg13g2_fill_2 FILLER_79_236 ();
 sg13g2_fill_1 FILLER_79_280 ();
 sg13g2_decap_4 FILLER_79_307 ();
 sg13g2_fill_1 FILLER_79_311 ();
 sg13g2_fill_2 FILLER_79_316 ();
 sg13g2_fill_1 FILLER_79_318 ();
 sg13g2_decap_4 FILLER_79_427 ();
 sg13g2_fill_2 FILLER_79_431 ();
 sg13g2_fill_2 FILLER_79_459 ();
 sg13g2_fill_1 FILLER_79_526 ();
 sg13g2_fill_2 FILLER_79_682 ();
 sg13g2_fill_1 FILLER_79_684 ();
 sg13g2_decap_8 FILLER_79_703 ();
 sg13g2_decap_8 FILLER_79_710 ();
 sg13g2_decap_8 FILLER_79_717 ();
 sg13g2_decap_8 FILLER_79_724 ();
 sg13g2_decap_8 FILLER_79_731 ();
 sg13g2_decap_8 FILLER_79_738 ();
 sg13g2_decap_8 FILLER_79_745 ();
 sg13g2_fill_1 FILLER_79_752 ();
 sg13g2_decap_8 FILLER_79_894 ();
 sg13g2_decap_8 FILLER_79_901 ();
 sg13g2_decap_8 FILLER_79_920 ();
 sg13g2_decap_8 FILLER_79_943 ();
 sg13g2_decap_4 FILLER_79_950 ();
 sg13g2_fill_1 FILLER_79_954 ();
 sg13g2_decap_8 FILLER_79_959 ();
 sg13g2_decap_8 FILLER_79_966 ();
 sg13g2_fill_2 FILLER_79_1060 ();
 sg13g2_fill_1 FILLER_79_1062 ();
 sg13g2_fill_2 FILLER_79_1090 ();
 sg13g2_fill_1 FILLER_79_1092 ();
 sg13g2_fill_2 FILLER_79_1097 ();
 sg13g2_fill_2 FILLER_79_1107 ();
 sg13g2_fill_1 FILLER_79_1135 ();
 sg13g2_decap_8 FILLER_79_1162 ();
 sg13g2_decap_8 FILLER_79_1169 ();
 sg13g2_decap_8 FILLER_79_1176 ();
 sg13g2_decap_8 FILLER_79_1183 ();
 sg13g2_decap_8 FILLER_79_1190 ();
 sg13g2_decap_8 FILLER_79_1197 ();
 sg13g2_decap_8 FILLER_79_1204 ();
 sg13g2_decap_8 FILLER_79_1211 ();
 sg13g2_decap_8 FILLER_79_1218 ();
 sg13g2_decap_8 FILLER_79_1225 ();
 sg13g2_decap_8 FILLER_79_1232 ();
 sg13g2_decap_8 FILLER_79_1239 ();
 sg13g2_decap_8 FILLER_79_1246 ();
 sg13g2_decap_8 FILLER_79_1253 ();
 sg13g2_decap_8 FILLER_79_1260 ();
 sg13g2_decap_8 FILLER_79_1267 ();
 sg13g2_decap_8 FILLER_79_1274 ();
 sg13g2_decap_8 FILLER_79_1281 ();
 sg13g2_decap_8 FILLER_79_1288 ();
 sg13g2_decap_8 FILLER_79_1295 ();
 sg13g2_decap_8 FILLER_79_1302 ();
 sg13g2_decap_4 FILLER_79_1309 ();
 sg13g2_fill_2 FILLER_79_1313 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_fill_1 FILLER_80_116 ();
 sg13g2_fill_1 FILLER_80_203 ();
 sg13g2_fill_1 FILLER_80_212 ();
 sg13g2_fill_1 FILLER_80_247 ();
 sg13g2_fill_2 FILLER_80_257 ();
 sg13g2_fill_2 FILLER_80_294 ();
 sg13g2_decap_4 FILLER_80_327 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_decap_4 FILLER_80_406 ();
 sg13g2_decap_8 FILLER_80_414 ();
 sg13g2_decap_8 FILLER_80_421 ();
 sg13g2_decap_8 FILLER_80_428 ();
 sg13g2_decap_4 FILLER_80_435 ();
 sg13g2_fill_2 FILLER_80_439 ();
 sg13g2_decap_4 FILLER_80_476 ();
 sg13g2_fill_2 FILLER_80_484 ();
 sg13g2_fill_2 FILLER_80_539 ();
 sg13g2_fill_1 FILLER_80_577 ();
 sg13g2_fill_1 FILLER_80_629 ();
 sg13g2_fill_2 FILLER_80_666 ();
 sg13g2_fill_1 FILLER_80_668 ();
 sg13g2_decap_8 FILLER_80_699 ();
 sg13g2_decap_8 FILLER_80_706 ();
 sg13g2_decap_8 FILLER_80_713 ();
 sg13g2_decap_8 FILLER_80_720 ();
 sg13g2_decap_8 FILLER_80_727 ();
 sg13g2_decap_8 FILLER_80_734 ();
 sg13g2_decap_8 FILLER_80_741 ();
 sg13g2_decap_8 FILLER_80_748 ();
 sg13g2_decap_8 FILLER_80_755 ();
 sg13g2_decap_8 FILLER_80_762 ();
 sg13g2_fill_1 FILLER_80_769 ();
 sg13g2_decap_8 FILLER_80_778 ();
 sg13g2_decap_4 FILLER_80_785 ();
 sg13g2_decap_8 FILLER_80_793 ();
 sg13g2_fill_2 FILLER_80_830 ();
 sg13g2_decap_8 FILLER_80_880 ();
 sg13g2_decap_8 FILLER_80_887 ();
 sg13g2_decap_8 FILLER_80_894 ();
 sg13g2_decap_8 FILLER_80_901 ();
 sg13g2_decap_8 FILLER_80_908 ();
 sg13g2_decap_8 FILLER_80_915 ();
 sg13g2_decap_8 FILLER_80_922 ();
 sg13g2_decap_8 FILLER_80_929 ();
 sg13g2_decap_8 FILLER_80_936 ();
 sg13g2_decap_8 FILLER_80_943 ();
 sg13g2_decap_8 FILLER_80_950 ();
 sg13g2_decap_8 FILLER_80_957 ();
 sg13g2_fill_2 FILLER_80_964 ();
 sg13g2_fill_2 FILLER_80_1001 ();
 sg13g2_decap_8 FILLER_80_1029 ();
 sg13g2_decap_4 FILLER_80_1036 ();
 sg13g2_decap_8 FILLER_80_1066 ();
 sg13g2_fill_2 FILLER_80_1073 ();
 sg13g2_decap_4 FILLER_80_1114 ();
 sg13g2_fill_2 FILLER_80_1118 ();
 sg13g2_fill_2 FILLER_80_1127 ();
 sg13g2_fill_1 FILLER_80_1129 ();
 sg13g2_fill_1 FILLER_80_1134 ();
 sg13g2_decap_8 FILLER_80_1157 ();
 sg13g2_decap_8 FILLER_80_1164 ();
 sg13g2_decap_8 FILLER_80_1171 ();
 sg13g2_decap_8 FILLER_80_1178 ();
 sg13g2_decap_8 FILLER_80_1185 ();
 sg13g2_decap_8 FILLER_80_1192 ();
 sg13g2_decap_8 FILLER_80_1199 ();
 sg13g2_decap_8 FILLER_80_1206 ();
 sg13g2_decap_8 FILLER_80_1213 ();
 sg13g2_decap_8 FILLER_80_1220 ();
 sg13g2_decap_8 FILLER_80_1227 ();
 sg13g2_decap_8 FILLER_80_1234 ();
 sg13g2_decap_8 FILLER_80_1241 ();
 sg13g2_decap_8 FILLER_80_1248 ();
 sg13g2_decap_8 FILLER_80_1255 ();
 sg13g2_decap_8 FILLER_80_1262 ();
 sg13g2_decap_8 FILLER_80_1269 ();
 sg13g2_decap_8 FILLER_80_1276 ();
 sg13g2_decap_8 FILLER_80_1283 ();
 sg13g2_decap_8 FILLER_80_1290 ();
 sg13g2_decap_8 FILLER_80_1297 ();
 sg13g2_decap_8 FILLER_80_1304 ();
 sg13g2_decap_4 FILLER_80_1311 ();
 assign uio_oe[0] = net5;
 assign uio_oe[1] = net6;
 assign uio_oe[2] = net7;
 assign uio_oe[3] = net8;
 assign uio_oe[4] = net9;
 assign uio_oe[5] = net10;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[0] = net13;
 assign uio_out[1] = net14;
 assign uio_out[2] = net15;
 assign uio_out[3] = net16;
 assign uio_out[4] = net17;
 assign uio_out[5] = net18;
 assign uio_out[6] = net19;
 assign uio_out[7] = net20;
 assign uo_out[2] = net21;
 assign uo_out[3] = net22;
 assign uo_out[4] = net23;
 assign uo_out[5] = net24;
 assign uo_out[6] = net25;
 assign uo_out[7] = net26;
endmodule

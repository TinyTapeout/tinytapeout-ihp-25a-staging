module tt_um_db_MAC (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire \a1.fa[0].fa0.A ;
 wire \a1.fa[0].fa0.S ;
 wire \a1.fa[0].fa1.A ;
 wire \a1.fa[0].fa1.S ;
 wire \a1.fa[0].fa2.A ;
 wire \a1.fa[0].fa2.S ;
 wire \a1.fa[0].fa3.A ;
 wire \a1.fa[0].fa3.S ;
 wire \a1.fa[1].fa0.A ;
 wire \a1.fa[1].fa0.S ;
 wire \a1.fa[1].fa1.A ;
 wire \a1.fa[1].fa1.S ;
 wire \a1.fa[1].fa2.A ;
 wire \a1.fa[1].fa2.S ;
 wire \a1.fa[1].fa3.A ;
 wire \a1.fa[1].fa3.S ;
 wire \a1.fa[2].fa0.A ;
 wire \a1.fa[2].fa0.S ;
 wire \a1.fa[2].fa1.A ;
 wire \a1.fa[2].fa1.S ;
 wire \a1.fa[2].fa2.A ;
 wire \a1.fa[2].fa2.S ;
 wire \a1.fa[2].fa3.A ;
 wire \a1.fa[2].fa3.S ;
 wire \a1.fa[3].fa0.A ;
 wire \a1.fa[3].fa0.S ;
 wire \a1.fa[3].fa1.A ;
 wire \a1.fa[3].fa1.S ;
 wire \a1.fa[3].fa2.A ;
 wire \a1.fa[3].fa2.S ;
 wire \a1.fa[3].fa3.A ;
 wire \a1.fa[3].fa3.S ;
 wire \m1.U0.U0.b1.A ;
 wire \m1.U0.U0.b1.B ;
 wire \m1.U0.U0.b1.D ;
 wire \m1.U0.U0.p1.A ;
 wire \m1.U0.U1.b1.B ;
 wire \m1.U0.U1.b1.D ;
 wire \m1.U0.U2.b1.A ;
 wire \m1.U0.U2.p1.A ;
 wire \m1.U1.U0.b1.B ;
 wire \m1.U1.U0.b1.D ;
 wire \m1.U1.U1.b1.B ;
 wire \m1.U1.U1.b1.D ;
 wire \m1.U2.U0.b1.A ;
 wire \m1.U2.U0.p1.A ;
 wire \m1.U2.U2.b1.A ;
 wire \m1.U2.U2.p1.A ;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;

 sg13g2_inv_1 _409_ (.Y(_344_),
    .A(net52));
 sg13g2_inv_1 _410_ (.Y(_345_),
    .A(net51));
 sg13g2_inv_1 _787__2 (.Y(net18),
    .A(clk));
 sg13g2_nand2_1 _412_ (.Y(_346_),
    .A(net96),
    .B(net86));
 sg13g2_nand4_1 _413_ (.B(net86),
    .C(net84),
    .A(net96),
    .Y(_347_),
    .D(net95));
 sg13g2_inv_1 _414_ (.Y(_348_),
    .A(_347_));
 sg13g2_a22oi_1 _415_ (.Y(_349_),
    .B1(net95),
    .B2(net86),
    .A2(net84),
    .A1(net96));
 sg13g2_nor2_1 _416_ (.A(_348_),
    .B(_349_),
    .Y(_350_));
 sg13g2_nand2_1 _417_ (.Y(_351_),
    .A(net87),
    .B(net102));
 sg13g2_nand4_1 _418_ (.B(net100),
    .C(net102),
    .A(net87),
    .Y(_352_),
    .D(net85));
 sg13g2_inv_1 _419_ (.Y(_353_),
    .A(_352_));
 sg13g2_nand2_1 _420_ (.Y(_354_),
    .A(\m1.U2.U2.b1.A ),
    .B(net102));
 sg13g2_and4_2 _421_ (.A(\m1.U2.U2.b1.A ),
    .B(\m1.U2.U2.p1.A ),
    .C(net100),
    .D(net102),
    .X(_355_));
 sg13g2_a22oi_1 _422_ (.Y(_356_),
    .B1(net102),
    .B2(\m1.U2.U2.p1.A ),
    .A2(net100),
    .A1(net83));
 sg13g2_nor3_1 _423_ (.A(_352_),
    .B(_355_),
    .C(_356_),
    .Y(_357_));
 sg13g2_nand2_1 _424_ (.Y(_358_),
    .A(net87),
    .B(net99));
 sg13g2_and4_1 _425_ (.A(net87),
    .B(net99),
    .C(net98),
    .D(net85),
    .X(_359_));
 sg13g2_a22oi_1 _426_ (.Y(_360_),
    .B1(net85),
    .B2(net99),
    .A2(\m1.U0.U1.b1.D ),
    .A1(net86));
 sg13g2_nor2_1 _427_ (.A(_359_),
    .B(_360_),
    .Y(_361_));
 sg13g2_o21ai_1 _428_ (.B1(_352_),
    .Y(_362_),
    .A1(_355_),
    .A2(_356_));
 sg13g2_nor2b_1 _429_ (.A(_357_),
    .B_N(_362_),
    .Y(_363_));
 sg13g2_a21oi_2 _430_ (.B1(_357_),
    .Y(_364_),
    .A2(_362_),
    .A1(_361_));
 sg13g2_nand3_1 _431_ (.B(net85),
    .C(_358_),
    .A(net98),
    .Y(_365_));
 sg13g2_nand2_2 _432_ (.Y(_366_),
    .A(net83),
    .B(net99));
 sg13g2_and3_1 _433_ (.X(_367_),
    .A(net82),
    .B(net100),
    .C(_354_));
 sg13g2_nand2b_1 _434_ (.Y(_368_),
    .B(_367_),
    .A_N(_366_));
 sg13g2_xnor2_1 _435_ (.Y(_369_),
    .A(_366_),
    .B(_367_));
 sg13g2_nand2b_1 _436_ (.Y(_370_),
    .B(_369_),
    .A_N(_365_));
 sg13g2_xor2_1 _437_ (.B(_369_),
    .A(_365_),
    .X(_371_));
 sg13g2_nor2_1 _438_ (.A(_364_),
    .B(_371_),
    .Y(_372_));
 sg13g2_xnor2_1 _439_ (.Y(_373_),
    .A(_361_),
    .B(_363_));
 sg13g2_nand3_1 _440_ (.B(net84),
    .C(_351_),
    .A(net100),
    .Y(_374_));
 sg13g2_or2_1 _441_ (.X(_375_),
    .B(_374_),
    .A(_354_));
 sg13g2_xor2_1 _442_ (.B(_374_),
    .A(_354_),
    .X(_376_));
 sg13g2_nand2b_1 _443_ (.Y(_016_),
    .B(_376_),
    .A_N(_358_));
 sg13g2_a21oi_2 _444_ (.B1(_373_),
    .Y(_017_),
    .A2(_016_),
    .A1(_375_));
 sg13g2_xor2_1 _445_ (.B(_371_),
    .A(_364_),
    .X(_018_));
 sg13g2_a21oi_1 _446_ (.A1(_017_),
    .A2(_018_),
    .Y(_019_),
    .B1(_372_));
 sg13g2_and2_1 _447_ (.A(_368_),
    .B(_370_),
    .X(_020_));
 sg13g2_nand2_1 _448_ (.Y(_021_),
    .A(net82),
    .B(net98));
 sg13g2_nor2_1 _449_ (.A(_366_),
    .B(_021_),
    .Y(_022_));
 sg13g2_a22oi_1 _450_ (.Y(_023_),
    .B1(net98),
    .B2(net83),
    .A2(net99),
    .A1(net82));
 sg13g2_nor2_1 _451_ (.A(_022_),
    .B(_023_),
    .Y(_024_));
 sg13g2_and2_1 _452_ (.A(_355_),
    .B(_024_),
    .X(_025_));
 sg13g2_xor2_1 _453_ (.B(_024_),
    .A(_355_),
    .X(_026_));
 sg13g2_xor2_1 _454_ (.B(_026_),
    .A(_359_),
    .X(_027_));
 sg13g2_nand2b_1 _455_ (.Y(_028_),
    .B(_027_),
    .A_N(_020_));
 sg13g2_xnor2_1 _456_ (.Y(_029_),
    .A(_020_),
    .B(_027_));
 sg13g2_nand2b_1 _457_ (.Y(_030_),
    .B(_029_),
    .A_N(_019_));
 sg13g2_xnor2_1 _458_ (.Y(_031_),
    .A(_019_),
    .B(_029_));
 sg13g2_xnor2_1 _459_ (.Y(_032_),
    .A(_350_),
    .B(_031_));
 sg13g2_and2_1 _460_ (.A(net97),
    .B(net92),
    .X(_033_));
 sg13g2_nand2_1 _461_ (.Y(_034_),
    .A(net97),
    .B(net92));
 sg13g2_nand2_1 _462_ (.Y(_035_),
    .A(net95),
    .B(net91));
 sg13g2_nor2_2 _463_ (.A(_034_),
    .B(_035_),
    .Y(_036_));
 sg13g2_nand2_1 _464_ (.Y(_037_),
    .A(net97),
    .B(net89));
 sg13g2_and4_1 _465_ (.A(net96),
    .B(net89),
    .C(\m1.U1.U0.b1.D ),
    .D(net88),
    .X(_038_));
 sg13g2_a22oi_1 _466_ (.Y(_039_),
    .B1(net88),
    .B2(net96),
    .A2(\m1.U1.U0.b1.D ),
    .A1(net89));
 sg13g2_nor2_1 _467_ (.A(_038_),
    .B(_039_),
    .Y(_040_));
 sg13g2_and2_1 _468_ (.A(\m1.U1.U1.b1.B ),
    .B(net92),
    .X(_041_));
 sg13g2_and3_1 _469_ (.X(_042_),
    .A(\m1.U1.U1.b1.D ),
    .B(net91),
    .C(_041_));
 sg13g2_a22oi_1 _470_ (.Y(_043_),
    .B1(net91),
    .B2(net94),
    .A2(net92),
    .A1(\m1.U1.U1.b1.D ));
 sg13g2_nor2_1 _471_ (.A(_042_),
    .B(_043_),
    .Y(_044_));
 sg13g2_xor2_1 _472_ (.B(_040_),
    .A(_036_),
    .X(_045_));
 sg13g2_and2_1 _473_ (.A(_044_),
    .B(_045_),
    .X(_046_));
 sg13g2_a21oi_1 _474_ (.A1(_036_),
    .A2(_040_),
    .Y(_047_),
    .B1(_046_));
 sg13g2_nand3b_1 _475_ (.B(net91),
    .C(net93),
    .Y(_048_),
    .A_N(_041_));
 sg13g2_nand2_2 _476_ (.Y(_049_),
    .A(net94),
    .B(net89));
 sg13g2_and3_1 _477_ (.X(_050_),
    .A(\m1.U1.U0.b1.D ),
    .B(net88),
    .C(_037_));
 sg13g2_nand2b_1 _478_ (.Y(_051_),
    .B(_050_),
    .A_N(_049_));
 sg13g2_xnor2_1 _479_ (.Y(_052_),
    .A(_049_),
    .B(_050_));
 sg13g2_nand2b_1 _480_ (.Y(_053_),
    .B(_052_),
    .A_N(_048_));
 sg13g2_xor2_1 _481_ (.B(_052_),
    .A(_048_),
    .X(_054_));
 sg13g2_nor2_1 _482_ (.A(_047_),
    .B(_054_),
    .Y(_055_));
 sg13g2_xnor2_1 _483_ (.Y(_056_),
    .A(_044_),
    .B(_045_));
 sg13g2_nor3_1 _484_ (.A(_033_),
    .B(_035_),
    .C(_037_),
    .Y(_057_));
 sg13g2_o21ai_1 _485_ (.B1(_037_),
    .Y(_058_),
    .A1(_033_),
    .A2(_035_));
 sg13g2_nor2b_1 _486_ (.A(_057_),
    .B_N(_058_),
    .Y(_059_));
 sg13g2_a21oi_1 _487_ (.A1(_041_),
    .A2(_058_),
    .Y(_060_),
    .B1(_057_));
 sg13g2_nor2_1 _488_ (.A(_056_),
    .B(_060_),
    .Y(_061_));
 sg13g2_xor2_1 _489_ (.B(_054_),
    .A(_047_),
    .X(_062_));
 sg13g2_a21oi_1 _490_ (.A1(_061_),
    .A2(_062_),
    .Y(_063_),
    .B1(_055_));
 sg13g2_and2_1 _491_ (.A(_051_),
    .B(_053_),
    .X(_064_));
 sg13g2_nand2_1 _492_ (.Y(_065_),
    .A(net93),
    .B(net88));
 sg13g2_nor2_1 _493_ (.A(_049_),
    .B(_065_),
    .Y(_066_));
 sg13g2_a22oi_1 _494_ (.Y(_067_),
    .B1(net88),
    .B2(net94),
    .A2(net89),
    .A1(net93));
 sg13g2_nor2_1 _495_ (.A(_066_),
    .B(_067_),
    .Y(_068_));
 sg13g2_and2_1 _496_ (.A(_038_),
    .B(_068_),
    .X(_069_));
 sg13g2_xor2_1 _497_ (.B(_068_),
    .A(_038_),
    .X(_070_));
 sg13g2_xor2_1 _498_ (.B(_070_),
    .A(_042_),
    .X(_071_));
 sg13g2_inv_1 _499_ (.Y(_072_),
    .A(_071_));
 sg13g2_xnor2_1 _500_ (.Y(_073_),
    .A(_064_),
    .B(_071_));
 sg13g2_nand2b_1 _501_ (.Y(_074_),
    .B(_073_),
    .A_N(_063_));
 sg13g2_xnor2_1 _502_ (.Y(_075_),
    .A(_063_),
    .B(_073_));
 sg13g2_nor2b_1 _503_ (.A(_032_),
    .B_N(_075_),
    .Y(_076_));
 sg13g2_xnor2_1 _504_ (.Y(_077_),
    .A(_032_),
    .B(_075_));
 sg13g2_xnor2_1 _505_ (.Y(_078_),
    .A(_017_),
    .B(_018_));
 sg13g2_nor2_1 _506_ (.A(_346_),
    .B(_078_),
    .Y(_079_));
 sg13g2_xor2_1 _507_ (.B(_078_),
    .A(_346_),
    .X(_080_));
 sg13g2_xor2_1 _508_ (.B(_062_),
    .A(_061_),
    .X(_081_));
 sg13g2_a21oi_1 _509_ (.A1(_080_),
    .A2(_081_),
    .Y(_082_),
    .B1(_079_));
 sg13g2_nor2b_1 _510_ (.A(_082_),
    .B_N(_077_),
    .Y(_083_));
 sg13g2_a21o_1 _511_ (.A2(_031_),
    .A1(_350_),
    .B1(_076_),
    .X(_084_));
 sg13g2_nor2b_1 _512_ (.A(_065_),
    .B_N(_049_),
    .Y(_085_));
 sg13g2_a21oi_1 _513_ (.A1(_042_),
    .A2(_070_),
    .Y(_086_),
    .B1(_069_));
 sg13g2_xnor2_1 _514_ (.Y(_087_),
    .A(_085_),
    .B(_086_));
 sg13g2_o21ai_1 _515_ (.B1(_074_),
    .Y(_088_),
    .A1(_064_),
    .A2(_072_));
 sg13g2_xor2_1 _516_ (.B(_088_),
    .A(_087_),
    .X(_089_));
 sg13g2_inv_1 _517_ (.Y(_090_),
    .A(_089_));
 sg13g2_nand2_1 _518_ (.Y(_091_),
    .A(net94),
    .B(net86));
 sg13g2_nand2_1 _519_ (.Y(_092_),
    .A(net83),
    .B(net96));
 sg13g2_nand3_1 _520_ (.B(net95),
    .C(_346_),
    .A(net84),
    .Y(_093_));
 sg13g2_or2_1 _521_ (.X(_094_),
    .B(_093_),
    .A(_092_));
 sg13g2_xor2_1 _522_ (.B(_093_),
    .A(_092_),
    .X(_095_));
 sg13g2_nand2b_1 _523_ (.Y(_096_),
    .B(_095_),
    .A_N(_091_));
 sg13g2_xnor2_1 _524_ (.Y(_097_),
    .A(_091_),
    .B(_095_));
 sg13g2_nor2b_1 _525_ (.A(_021_),
    .B_N(_366_),
    .Y(_098_));
 sg13g2_a21oi_1 _526_ (.A1(_359_),
    .A2(_026_),
    .Y(_099_),
    .B1(_025_));
 sg13g2_xnor2_1 _527_ (.Y(_100_),
    .A(_098_),
    .B(_099_));
 sg13g2_nand2_1 _528_ (.Y(_101_),
    .A(_028_),
    .B(_030_));
 sg13g2_xor2_1 _529_ (.B(_101_),
    .A(_100_),
    .X(_102_));
 sg13g2_xnor2_1 _530_ (.Y(_103_),
    .A(_097_),
    .B(_102_));
 sg13g2_nor2_1 _531_ (.A(_090_),
    .B(_103_),
    .Y(_104_));
 sg13g2_xor2_1 _532_ (.B(_103_),
    .A(_089_),
    .X(_105_));
 sg13g2_nor2b_1 _533_ (.A(_105_),
    .B_N(_084_),
    .Y(_106_));
 sg13g2_xor2_1 _534_ (.B(_105_),
    .A(_084_),
    .X(_107_));
 sg13g2_inv_1 _535_ (.Y(_108_),
    .A(_107_));
 sg13g2_xnor2_1 _536_ (.Y(_109_),
    .A(_083_),
    .B(_107_));
 sg13g2_xnor2_1 _537_ (.Y(_110_),
    .A(_080_),
    .B(_081_));
 sg13g2_nand3_1 _538_ (.B(_375_),
    .C(_016_),
    .A(_373_),
    .Y(_111_));
 sg13g2_nand2b_1 _539_ (.Y(_112_),
    .B(_111_),
    .A_N(_017_));
 sg13g2_nand2_2 _540_ (.Y(_113_),
    .A(net99),
    .B(net90));
 sg13g2_nand2_1 _541_ (.Y(_114_),
    .A(net98),
    .B(\m1.U0.U2.p1.A ));
 sg13g2_nand2b_1 _542_ (.Y(_115_),
    .B(_113_),
    .A_N(_114_));
 sg13g2_nand2_2 _543_ (.Y(_116_),
    .A(net103),
    .B(net90));
 sg13g2_and2_1 _544_ (.A(net101),
    .B(\m1.U0.U2.p1.A ),
    .X(_117_));
 sg13g2_and4_2 _545_ (.A(net100),
    .B(net102),
    .C(net90),
    .D(net88),
    .X(_118_));
 sg13g2_nand2_1 _546_ (.Y(_119_),
    .A(\m1.U0.U1.b1.D ),
    .B(net90));
 sg13g2_nand2_1 _547_ (.Y(_120_),
    .A(net99),
    .B(net88));
 sg13g2_xor2_1 _548_ (.B(_120_),
    .A(_119_),
    .X(_121_));
 sg13g2_and2_2 _549_ (.A(\m1.U0.U1.b1.B ),
    .B(\m1.U0.U0.b1.A ),
    .X(_122_));
 sg13g2_and2_1 _550_ (.A(net98),
    .B(\m1.U0.U0.p1.A ),
    .X(_123_));
 sg13g2_nand2_1 _551_ (.Y(_124_),
    .A(net98),
    .B(\m1.U0.U0.p1.A ));
 sg13g2_nand2_1 _552_ (.Y(_125_),
    .A(_122_),
    .B(_123_));
 sg13g2_xor2_1 _553_ (.B(_121_),
    .A(_118_),
    .X(_126_));
 sg13g2_nor2b_1 _554_ (.A(_125_),
    .B_N(_126_),
    .Y(_127_));
 sg13g2_a21oi_1 _555_ (.A1(_118_),
    .A2(_121_),
    .Y(_128_),
    .B1(_127_));
 sg13g2_xor2_1 _556_ (.B(_128_),
    .A(_115_),
    .X(_129_));
 sg13g2_and4_1 _557_ (.A(\m1.U0.U1.b1.B ),
    .B(net89),
    .C(_116_),
    .D(_117_),
    .X(_130_));
 sg13g2_nor2_1 _558_ (.A(_122_),
    .B(_124_),
    .Y(_131_));
 sg13g2_a22oi_1 _559_ (.Y(_132_),
    .B1(_116_),
    .B2(_117_),
    .A2(net89),
    .A1(\m1.U0.U1.b1.B ));
 sg13g2_a21oi_1 _560_ (.A1(_116_),
    .A2(_117_),
    .Y(_133_),
    .B1(_113_));
 sg13g2_and3_1 _561_ (.X(_134_),
    .A(_113_),
    .B(_116_),
    .C(_117_));
 sg13g2_nor4_2 _562_ (.A(_122_),
    .B(_124_),
    .C(_130_),
    .Y(_135_),
    .D(_132_));
 sg13g2_nor2_1 _563_ (.A(_130_),
    .B(_135_),
    .Y(_136_));
 sg13g2_xnor2_1 _564_ (.Y(_137_),
    .A(_125_),
    .B(_126_));
 sg13g2_nand2b_1 _565_ (.Y(_138_),
    .B(_137_),
    .A_N(_136_));
 sg13g2_and2_1 _566_ (.A(net103),
    .B(net92),
    .X(_139_));
 sg13g2_nand2_1 _567_ (.Y(_140_),
    .A(net101),
    .B(\m1.U0.U0.p1.A ));
 sg13g2_nand4_1 _568_ (.B(net103),
    .C(\m1.U0.U0.b1.A ),
    .A(net101),
    .Y(_141_),
    .D(net91));
 sg13g2_inv_1 _569_ (.Y(_142_),
    .A(_141_));
 sg13g2_a22oi_1 _570_ (.Y(_143_),
    .B1(net88),
    .B2(net103),
    .A2(net89),
    .A1(net101));
 sg13g2_nor3_1 _571_ (.A(_118_),
    .B(_141_),
    .C(_143_),
    .Y(_144_));
 sg13g2_or3_1 _572_ (.A(_118_),
    .B(_141_),
    .C(_143_),
    .X(_145_));
 sg13g2_a22oi_1 _573_ (.Y(_146_),
    .B1(net91),
    .B2(net99),
    .A2(net92),
    .A1(net98));
 sg13g2_a21oi_1 _574_ (.A1(_122_),
    .A2(_123_),
    .Y(_147_),
    .B1(_146_));
 sg13g2_o21ai_1 _575_ (.B1(_141_),
    .Y(_148_),
    .A1(_118_),
    .A2(_143_));
 sg13g2_and3_1 _576_ (.X(_149_),
    .A(_145_),
    .B(_147_),
    .C(_148_));
 sg13g2_a21oi_1 _577_ (.A1(_147_),
    .A2(_148_),
    .Y(_150_),
    .B1(_144_));
 sg13g2_nor3_1 _578_ (.A(_131_),
    .B(_133_),
    .C(_134_),
    .Y(_151_));
 sg13g2_nor3_1 _579_ (.A(_135_),
    .B(_150_),
    .C(_151_),
    .Y(_152_));
 sg13g2_a21oi_1 _580_ (.A1(_145_),
    .A2(_148_),
    .Y(_153_),
    .B1(_147_));
 sg13g2_nor3_1 _581_ (.A(_116_),
    .B(_139_),
    .C(_140_),
    .Y(_154_));
 sg13g2_o21ai_1 _582_ (.B1(_116_),
    .Y(_155_),
    .A1(_139_),
    .A2(_140_));
 sg13g2_nor2b_1 _583_ (.A(_154_),
    .B_N(_155_),
    .Y(_156_));
 sg13g2_a21oi_1 _584_ (.A1(_122_),
    .A2(_155_),
    .Y(_157_),
    .B1(_154_));
 sg13g2_nor3_2 _585_ (.A(_149_),
    .B(_153_),
    .C(_157_),
    .Y(_158_));
 sg13g2_o21ai_1 _586_ (.B1(_150_),
    .Y(_159_),
    .A1(_135_),
    .A2(_151_));
 sg13g2_nor2b_1 _587_ (.A(_152_),
    .B_N(_159_),
    .Y(_160_));
 sg13g2_a21oi_2 _588_ (.B1(_152_),
    .Y(_161_),
    .A2(_159_),
    .A1(_158_));
 sg13g2_nor2b_1 _589_ (.A(_137_),
    .B_N(_136_),
    .Y(_162_));
 sg13g2_xnor2_1 _590_ (.Y(_163_),
    .A(_136_),
    .B(_137_));
 sg13g2_o21ai_1 _591_ (.B1(_138_),
    .Y(_164_),
    .A1(_161_),
    .A2(_162_));
 sg13g2_a21oi_1 _592_ (.A1(_113_),
    .A2(_128_),
    .Y(_165_),
    .B1(_114_));
 sg13g2_a21oi_2 _593_ (.B1(_165_),
    .Y(_166_),
    .A2(_164_),
    .A1(_129_));
 sg13g2_nor2_1 _594_ (.A(_112_),
    .B(_166_),
    .Y(_167_));
 sg13g2_xnor2_1 _595_ (.Y(_168_),
    .A(_056_),
    .B(_060_));
 sg13g2_inv_1 _596_ (.Y(_169_),
    .A(_168_));
 sg13g2_xor2_1 _597_ (.B(_166_),
    .A(_112_),
    .X(_170_));
 sg13g2_a21oi_2 _598_ (.B1(_167_),
    .Y(_171_),
    .A2(_170_),
    .A1(_169_));
 sg13g2_nor2_1 _599_ (.A(_110_),
    .B(_171_),
    .Y(_172_));
 sg13g2_xnor2_1 _600_ (.Y(_173_),
    .A(_077_),
    .B(_082_));
 sg13g2_and2_1 _601_ (.A(_172_),
    .B(_173_),
    .X(_174_));
 sg13g2_xnor2_1 _602_ (.Y(_175_),
    .A(_168_),
    .B(_170_));
 sg13g2_xnor2_1 _603_ (.Y(_176_),
    .A(_358_),
    .B(_376_));
 sg13g2_xor2_1 _604_ (.B(_164_),
    .A(_129_),
    .X(_177_));
 sg13g2_nand2_1 _605_ (.Y(_178_),
    .A(_176_),
    .B(_177_));
 sg13g2_xnor2_1 _606_ (.Y(_179_),
    .A(_041_),
    .B(_059_));
 sg13g2_xnor2_1 _607_ (.Y(_180_),
    .A(_176_),
    .B(_177_));
 sg13g2_o21ai_1 _608_ (.B1(_178_),
    .Y(_181_),
    .A1(_179_),
    .A2(_180_));
 sg13g2_nand2_1 _609_ (.Y(_182_),
    .A(_175_),
    .B(_181_));
 sg13g2_xnor2_1 _610_ (.Y(_183_),
    .A(_110_),
    .B(_171_));
 sg13g2_or2_1 _611_ (.X(_184_),
    .B(_183_),
    .A(_182_));
 sg13g2_xnor2_1 _612_ (.Y(_185_),
    .A(_179_),
    .B(_180_));
 sg13g2_a22oi_1 _613_ (.Y(_186_),
    .B1(net102),
    .B2(net84),
    .A2(net100),
    .A1(net86));
 sg13g2_nor2_1 _614_ (.A(_353_),
    .B(_186_),
    .Y(_187_));
 sg13g2_xnor2_1 _615_ (.Y(_188_),
    .A(_161_),
    .B(_163_));
 sg13g2_a22oi_1 _616_ (.Y(_189_),
    .B1(net91),
    .B2(net97),
    .A2(net92),
    .A1(net95));
 sg13g2_nor2_1 _617_ (.A(_036_),
    .B(_189_),
    .Y(_190_));
 sg13g2_xnor2_1 _618_ (.Y(_191_),
    .A(_187_),
    .B(_188_));
 sg13g2_nor3_1 _619_ (.A(_036_),
    .B(_189_),
    .C(_191_),
    .Y(_192_));
 sg13g2_a21o_1 _620_ (.A2(_188_),
    .A1(_187_),
    .B1(_192_),
    .X(_193_));
 sg13g2_nand2b_1 _621_ (.Y(_194_),
    .B(_193_),
    .A_N(_185_));
 sg13g2_xnor2_1 _622_ (.Y(_195_),
    .A(_175_),
    .B(_181_));
 sg13g2_nor2_1 _623_ (.A(_194_),
    .B(_195_),
    .Y(_196_));
 sg13g2_xor2_1 _624_ (.B(_193_),
    .A(_185_),
    .X(_197_));
 sg13g2_xnor2_1 _625_ (.Y(_198_),
    .A(_158_),
    .B(_160_));
 sg13g2_nor2_1 _626_ (.A(_351_),
    .B(_198_),
    .Y(_199_));
 sg13g2_xor2_1 _627_ (.B(_198_),
    .A(_351_),
    .X(_200_));
 sg13g2_a21oi_1 _628_ (.A1(_033_),
    .A2(_200_),
    .Y(_201_),
    .B1(_199_));
 sg13g2_xor2_1 _629_ (.B(_191_),
    .A(_190_),
    .X(_202_));
 sg13g2_nor2_1 _630_ (.A(_201_),
    .B(_202_),
    .Y(_203_));
 sg13g2_inv_1 _631_ (.Y(_204_),
    .A(_203_));
 sg13g2_nor3_1 _632_ (.A(_195_),
    .B(_197_),
    .C(_204_),
    .Y(_205_));
 sg13g2_xor2_1 _633_ (.B(_183_),
    .A(_182_),
    .X(_206_));
 sg13g2_o21ai_1 _634_ (.B1(_206_),
    .Y(_207_),
    .A1(_196_),
    .A2(_205_));
 sg13g2_xnor2_1 _635_ (.Y(_208_),
    .A(_172_),
    .B(_173_));
 sg13g2_a21oi_1 _636_ (.A1(_184_),
    .A2(_207_),
    .Y(_209_),
    .B1(_208_));
 sg13g2_nor2_1 _637_ (.A(_174_),
    .B(_209_),
    .Y(_210_));
 sg13g2_o21ai_1 _638_ (.B1(_109_),
    .Y(_211_),
    .A1(_174_),
    .A2(_209_));
 sg13g2_a21oi_1 _639_ (.A1(_083_),
    .A2(_108_),
    .Y(_212_),
    .B1(_106_));
 sg13g2_a21oi_1 _640_ (.A1(_097_),
    .A2(_102_),
    .Y(_213_),
    .B1(_104_));
 sg13g2_a21oi_1 _641_ (.A1(_049_),
    .A2(_086_),
    .Y(_214_),
    .B1(_065_));
 sg13g2_a21oi_2 _642_ (.B1(_214_),
    .Y(_215_),
    .A2(_088_),
    .A1(_087_));
 sg13g2_a22oi_1 _643_ (.Y(_216_),
    .B1(net84),
    .B2(net94),
    .A2(net86),
    .A1(net93));
 sg13g2_nand4_1 _644_ (.B(net94),
    .C(net86),
    .A(net93),
    .Y(_217_),
    .D(net84));
 sg13g2_nor2b_1 _645_ (.A(_216_),
    .B_N(_217_),
    .Y(_218_));
 sg13g2_a22oi_1 _646_ (.Y(_219_),
    .B1(net95),
    .B2(net83),
    .A2(net96),
    .A1(net82));
 sg13g2_nand4_1 _647_ (.B(net82),
    .C(net96),
    .A(net83),
    .Y(_220_),
    .D(net95));
 sg13g2_nor2b_1 _648_ (.A(_219_),
    .B_N(_220_),
    .Y(_221_));
 sg13g2_xnor2_1 _649_ (.Y(_222_),
    .A(_347_),
    .B(_221_));
 sg13g2_and2_1 _650_ (.A(_218_),
    .B(_222_),
    .X(_223_));
 sg13g2_xnor2_1 _651_ (.Y(_224_),
    .A(_218_),
    .B(_222_));
 sg13g2_a21oi_2 _652_ (.B1(_224_),
    .Y(_225_),
    .A2(_096_),
    .A1(_094_));
 sg13g2_nand3_1 _653_ (.B(_096_),
    .C(_224_),
    .A(_094_),
    .Y(_226_));
 sg13g2_nand2b_1 _654_ (.Y(_227_),
    .B(_226_),
    .A_N(_225_));
 sg13g2_a21oi_1 _655_ (.A1(_366_),
    .A2(_099_),
    .Y(_228_),
    .B1(_021_));
 sg13g2_a21oi_2 _656_ (.B1(_228_),
    .Y(_229_),
    .A2(_101_),
    .A1(_100_));
 sg13g2_or2_1 _657_ (.X(_230_),
    .B(_229_),
    .A(_227_));
 sg13g2_xnor2_1 _658_ (.Y(_231_),
    .A(_227_),
    .B(_229_));
 sg13g2_xnor2_1 _659_ (.Y(_232_),
    .A(_215_),
    .B(_231_));
 sg13g2_nor2_1 _660_ (.A(_213_),
    .B(_232_),
    .Y(_233_));
 sg13g2_xnor2_1 _661_ (.Y(_234_),
    .A(_213_),
    .B(_232_));
 sg13g2_a21oi_1 _662_ (.A1(_211_),
    .A2(_212_),
    .Y(_235_),
    .B1(_234_));
 sg13g2_nand3_1 _663_ (.B(_212_),
    .C(_234_),
    .A(_211_),
    .Y(_236_));
 sg13g2_nand2b_1 _664_ (.Y(_237_),
    .B(_236_),
    .A_N(_235_));
 sg13g2_or2_1 _665_ (.X(_238_),
    .B(_237_),
    .A(_344_));
 sg13g2_xor2_1 _666_ (.B(_210_),
    .A(_109_),
    .X(_239_));
 sg13g2_nor2_1 _667_ (.A(_345_),
    .B(_239_),
    .Y(_240_));
 sg13g2_nand3_1 _668_ (.B(_207_),
    .C(_208_),
    .A(_184_),
    .Y(_241_));
 sg13g2_nor2b_1 _669_ (.A(_209_),
    .B_N(_241_),
    .Y(_242_));
 sg13g2_nand2_1 _670_ (.Y(_243_),
    .A(net43),
    .B(_242_));
 sg13g2_or3_1 _671_ (.A(_196_),
    .B(_205_),
    .C(_206_),
    .X(_244_));
 sg13g2_and2_1 _672_ (.A(_207_),
    .B(_244_),
    .X(_245_));
 sg13g2_and2_1 _673_ (.A(\a1.fa[2].fa0.A ),
    .B(_245_),
    .X(_246_));
 sg13g2_o21ai_1 _674_ (.B1(_194_),
    .Y(_247_),
    .A1(_197_),
    .A2(_204_));
 sg13g2_xnor2_1 _675_ (.Y(_248_),
    .A(_195_),
    .B(_247_));
 sg13g2_and2_1 _676_ (.A(net49),
    .B(_248_),
    .X(_249_));
 sg13g2_xnor2_1 _677_ (.Y(_250_),
    .A(_197_),
    .B(_203_));
 sg13g2_and2_1 _678_ (.A(net46),
    .B(_250_),
    .X(_251_));
 sg13g2_xor2_1 _679_ (.B(_202_),
    .A(_201_),
    .X(_252_));
 sg13g2_xnor2_1 _680_ (.Y(_253_),
    .A(_034_),
    .B(_200_));
 sg13g2_nand2_1 _681_ (.Y(_254_),
    .A(\a1.fa[1].fa0.A ),
    .B(_253_));
 sg13g2_o21ai_1 _682_ (.B1(_157_),
    .Y(_255_),
    .A1(_149_),
    .A2(_153_));
 sg13g2_nor2b_1 _683_ (.A(_158_),
    .B_N(_255_),
    .Y(_256_));
 sg13g2_xor2_1 _684_ (.B(_156_),
    .A(_122_),
    .X(_257_));
 sg13g2_nand2_1 _685_ (.Y(_258_),
    .A(\a1.fa[0].fa2.A ),
    .B(_257_));
 sg13g2_a22oi_1 _686_ (.Y(_259_),
    .B1(net91),
    .B2(net102),
    .A2(net92),
    .A1(net100));
 sg13g2_nor2_1 _687_ (.A(_142_),
    .B(_259_),
    .Y(_260_));
 sg13g2_nand2_1 _688_ (.Y(_261_),
    .A(net33),
    .B(_139_));
 sg13g2_xnor2_1 _689_ (.Y(_262_),
    .A(net34),
    .B(_260_));
 sg13g2_nor2_1 _690_ (.A(_261_),
    .B(_262_),
    .Y(_263_));
 sg13g2_a21oi_1 _691_ (.A1(net34),
    .A2(_260_),
    .Y(_264_),
    .B1(_263_));
 sg13g2_xnor2_1 _692_ (.Y(_265_),
    .A(net42),
    .B(_257_));
 sg13g2_o21ai_1 _693_ (.B1(_258_),
    .Y(_266_),
    .A1(_264_),
    .A2(_265_));
 sg13g2_xnor2_1 _694_ (.Y(_267_),
    .A(net39),
    .B(_256_));
 sg13g2_nor2b_1 _695_ (.A(_267_),
    .B_N(_266_),
    .Y(_268_));
 sg13g2_a21oi_1 _696_ (.A1(net39),
    .A2(_256_),
    .Y(_269_),
    .B1(_268_));
 sg13g2_xnor2_1 _697_ (.Y(_270_),
    .A(net41),
    .B(_253_));
 sg13g2_o21ai_1 _698_ (.B1(_254_),
    .Y(_271_),
    .A1(_269_),
    .A2(_270_));
 sg13g2_xnor2_1 _699_ (.Y(_272_),
    .A(net35),
    .B(_252_));
 sg13g2_nor2b_1 _700_ (.A(_272_),
    .B_N(_271_),
    .Y(_273_));
 sg13g2_a21o_1 _701_ (.A2(_252_),
    .A1(net35),
    .B1(_273_),
    .X(_274_));
 sg13g2_xor2_1 _702_ (.B(_250_),
    .A(net46),
    .X(_275_));
 sg13g2_a21o_1 _703_ (.A2(_275_),
    .A1(_274_),
    .B1(_251_),
    .X(_276_));
 sg13g2_xor2_1 _704_ (.B(_248_),
    .A(net49),
    .X(_277_));
 sg13g2_a21o_1 _705_ (.A2(_277_),
    .A1(_276_),
    .B1(_249_),
    .X(_278_));
 sg13g2_xor2_1 _706_ (.B(_245_),
    .A(net50),
    .X(_279_));
 sg13g2_a21oi_1 _707_ (.A1(_278_),
    .A2(_279_),
    .Y(_280_),
    .B1(_246_));
 sg13g2_xnor2_1 _708_ (.Y(_281_),
    .A(net43),
    .B(_242_));
 sg13g2_o21ai_1 _709_ (.B1(_243_),
    .Y(_282_),
    .A1(_280_),
    .A2(_281_));
 sg13g2_nand2_1 _710_ (.Y(_283_),
    .A(_345_),
    .B(_239_));
 sg13g2_nand2b_1 _711_ (.Y(_284_),
    .B(_283_),
    .A_N(_240_));
 sg13g2_a21oi_1 _712_ (.A1(_282_),
    .A2(_283_),
    .Y(_285_),
    .B1(_240_));
 sg13g2_xnor2_1 _713_ (.Y(_286_),
    .A(_344_),
    .B(_237_));
 sg13g2_o21ai_1 _714_ (.B1(_238_),
    .Y(_287_),
    .A1(_285_),
    .A2(_286_));
 sg13g2_a21oi_2 _715_ (.B1(_223_),
    .Y(_288_),
    .A2(_221_),
    .A1(_348_));
 sg13g2_nand3_1 _716_ (.B(net84),
    .C(_091_),
    .A(net93),
    .Y(_289_));
 sg13g2_nand2_2 _717_ (.Y(_290_),
    .A(net83),
    .B(net94));
 sg13g2_and3_1 _718_ (.X(_291_),
    .A(net82),
    .B(net95),
    .C(_092_));
 sg13g2_nand2b_1 _719_ (.Y(_292_),
    .B(_291_),
    .A_N(_290_));
 sg13g2_xnor2_1 _720_ (.Y(_293_),
    .A(_290_),
    .B(_291_));
 sg13g2_nand2b_1 _721_ (.Y(_294_),
    .B(_293_),
    .A_N(_289_));
 sg13g2_xor2_1 _722_ (.B(_293_),
    .A(_289_),
    .X(_295_));
 sg13g2_nor2_1 _723_ (.A(_288_),
    .B(_295_),
    .Y(_296_));
 sg13g2_xor2_1 _724_ (.B(_295_),
    .A(_288_),
    .X(_297_));
 sg13g2_xnor2_1 _725_ (.Y(_298_),
    .A(_225_),
    .B(_297_));
 sg13g2_o21ai_1 _726_ (.B1(_230_),
    .Y(_299_),
    .A1(_215_),
    .A2(_231_));
 sg13g2_nand2b_1 _727_ (.Y(_300_),
    .B(_299_),
    .A_N(_298_));
 sg13g2_xnor2_1 _728_ (.Y(_301_),
    .A(_298_),
    .B(_299_));
 sg13g2_o21ai_1 _729_ (.B1(_301_),
    .Y(_302_),
    .A1(_233_),
    .A2(_235_));
 sg13g2_or3_1 _730_ (.A(_233_),
    .B(_235_),
    .C(_301_),
    .X(_303_));
 sg13g2_and2_1 _731_ (.A(_302_),
    .B(_303_),
    .X(_304_));
 sg13g2_and2_1 _732_ (.A(\a1.fa[3].fa0.A ),
    .B(_304_),
    .X(_305_));
 sg13g2_xor2_1 _733_ (.B(_304_),
    .A(net45),
    .X(_306_));
 sg13g2_xor2_1 _734_ (.B(_306_),
    .A(_287_),
    .X(\a1.fa[3].fa0.S ));
 sg13g2_a21oi_1 _735_ (.A1(_287_),
    .A2(_306_),
    .Y(_307_),
    .B1(_305_));
 sg13g2_a21oi_1 _736_ (.A1(_225_),
    .A2(_297_),
    .Y(_308_),
    .B1(_296_));
 sg13g2_and2_1 _737_ (.A(_292_),
    .B(_294_),
    .X(_309_));
 sg13g2_nand2_1 _738_ (.Y(_310_),
    .A(net93),
    .B(net82));
 sg13g2_nor2_1 _739_ (.A(_290_),
    .B(_310_),
    .Y(_311_));
 sg13g2_a22oi_1 _740_ (.Y(_312_),
    .B1(net82),
    .B2(net94),
    .A2(net83),
    .A1(net93));
 sg13g2_nor3_1 _741_ (.A(_220_),
    .B(_311_),
    .C(_312_),
    .Y(_313_));
 sg13g2_o21ai_1 _742_ (.B1(_220_),
    .Y(_314_),
    .A1(_311_),
    .A2(_312_));
 sg13g2_nor2b_1 _743_ (.A(_313_),
    .B_N(_314_),
    .Y(_315_));
 sg13g2_nor2b_1 _744_ (.A(_217_),
    .B_N(_315_),
    .Y(_316_));
 sg13g2_xnor2_1 _745_ (.Y(_317_),
    .A(_217_),
    .B(_315_));
 sg13g2_inv_1 _746_ (.Y(_318_),
    .A(_317_));
 sg13g2_xnor2_1 _747_ (.Y(_319_),
    .A(_309_),
    .B(_317_));
 sg13g2_nand2b_1 _748_ (.Y(_320_),
    .B(_319_),
    .A_N(_308_));
 sg13g2_xnor2_1 _749_ (.Y(_321_),
    .A(_308_),
    .B(_319_));
 sg13g2_nand2_2 _750_ (.Y(_322_),
    .A(_300_),
    .B(_302_));
 sg13g2_xor2_1 _751_ (.B(_322_),
    .A(_321_),
    .X(_323_));
 sg13g2_nand2_1 _752_ (.Y(_324_),
    .A(net37),
    .B(_323_));
 sg13g2_nor2_1 _753_ (.A(net53),
    .B(_323_),
    .Y(_325_));
 sg13g2_xor2_1 _754_ (.B(_323_),
    .A(net37),
    .X(_326_));
 sg13g2_xnor2_1 _755_ (.Y(\a1.fa[3].fa1.S ),
    .A(_307_),
    .B(_326_));
 sg13g2_o21ai_1 _756_ (.B1(_324_),
    .Y(_327_),
    .A1(_307_),
    .A2(_325_));
 sg13g2_o21ai_1 _757_ (.B1(_320_),
    .Y(_328_),
    .A1(_309_),
    .A2(_318_));
 sg13g2_nor2b_1 _758_ (.A(_310_),
    .B_N(_290_),
    .Y(_329_));
 sg13g2_nor2_1 _759_ (.A(_313_),
    .B(_316_),
    .Y(_330_));
 sg13g2_xnor2_1 _760_ (.Y(_331_),
    .A(_329_),
    .B(_330_));
 sg13g2_xor2_1 _761_ (.B(_331_),
    .A(_328_),
    .X(_332_));
 sg13g2_nand2_1 _762_ (.Y(_333_),
    .A(_321_),
    .B(_322_));
 sg13g2_nand3_1 _763_ (.B(_322_),
    .C(_332_),
    .A(_321_),
    .Y(_334_));
 sg13g2_xnor2_1 _764_ (.Y(_335_),
    .A(_332_),
    .B(_333_));
 sg13g2_and2_1 _765_ (.A(net47),
    .B(_335_),
    .X(_336_));
 sg13g2_or2_1 _766_ (.X(_337_),
    .B(_335_),
    .A(net47));
 sg13g2_nand2b_1 _767_ (.Y(_338_),
    .B(_337_),
    .A_N(_336_));
 sg13g2_xnor2_1 _768_ (.Y(\a1.fa[3].fa2.S ),
    .A(_327_),
    .B(_338_));
 sg13g2_a21oi_1 _769_ (.A1(_327_),
    .A2(_337_),
    .Y(_339_),
    .B1(_336_));
 sg13g2_a21oi_1 _770_ (.A1(_290_),
    .A2(_330_),
    .Y(_340_),
    .B1(_310_));
 sg13g2_a21oi_1 _771_ (.A1(_328_),
    .A2(_331_),
    .Y(_341_),
    .B1(_340_));
 sg13g2_xnor2_1 _772_ (.Y(_342_),
    .A(\a1.fa[3].fa3.A ),
    .B(_341_));
 sg13g2_xnor2_1 _773_ (.Y(_343_),
    .A(_334_),
    .B(_342_));
 sg13g2_xnor2_1 _774_ (.Y(\a1.fa[3].fa3.S ),
    .A(_339_),
    .B(_343_));
 sg13g2_xor2_1 _775_ (.B(_139_),
    .A(net33),
    .X(\a1.fa[0].fa0.S ));
 sg13g2_xor2_1 _776_ (.B(_279_),
    .A(_278_),
    .X(\a1.fa[2].fa0.S ));
 sg13g2_xor2_1 _777_ (.B(_281_),
    .A(_280_),
    .X(\a1.fa[2].fa1.S ));
 sg13g2_xnor2_1 _778_ (.Y(\a1.fa[2].fa2.S ),
    .A(_282_),
    .B(_284_));
 sg13g2_xor2_1 _779_ (.B(_286_),
    .A(_285_),
    .X(\a1.fa[2].fa3.S ));
 sg13g2_xor2_1 _780_ (.B(_270_),
    .A(_269_),
    .X(\a1.fa[1].fa0.S ));
 sg13g2_xnor2_1 _781_ (.Y(\a1.fa[1].fa1.S ),
    .A(_271_),
    .B(_272_));
 sg13g2_xor2_1 _782_ (.B(_275_),
    .A(_274_),
    .X(\a1.fa[1].fa2.S ));
 sg13g2_xor2_1 _783_ (.B(_277_),
    .A(_276_),
    .X(\a1.fa[1].fa3.S ));
 sg13g2_xor2_1 _784_ (.B(_262_),
    .A(_261_),
    .X(\a1.fa[0].fa1.S ));
 sg13g2_xor2_1 _785_ (.B(_265_),
    .A(_264_),
    .X(\a1.fa[0].fa2.S ));
 sg13g2_xnor2_1 _786_ (.Y(\a1.fa[0].fa3.S ),
    .A(_266_),
    .B(_267_));
 sg13g2_inv_1 _788__3 (.Y(net19),
    .A(clk));
 sg13g2_inv_1 _789__4 (.Y(net20),
    .A(clk));
 sg13g2_inv_1 _790__5 (.Y(net21),
    .A(clk));
 sg13g2_inv_1 _791__6 (.Y(net22),
    .A(clk));
 sg13g2_inv_1 _792__7 (.Y(net23),
    .A(clk));
 sg13g2_inv_1 _793__8 (.Y(net24),
    .A(clk));
 sg13g2_inv_1 _794__9 (.Y(net25),
    .A(clk));
 sg13g2_inv_1 _795__10 (.Y(net26),
    .A(clk));
 sg13g2_inv_1 _796__11 (.Y(net27),
    .A(clk));
 sg13g2_inv_1 _797__12 (.Y(net28),
    .A(clk));
 sg13g2_inv_1 _798__13 (.Y(net29),
    .A(clk));
 sg13g2_inv_1 _799__14 (.Y(net30),
    .A(clk));
 sg13g2_inv_1 _800__15 (.Y(net31),
    .A(clk));
 sg13g2_inv_1 _801__16 (.Y(net32),
    .A(clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\a1.fa[0].fa0.A ),
    .X(net33));
 sg13g2_dfrbp_1 _802_ (.CLK(clk),
    .RESET_B(net106),
    .D(net9),
    .Q_N(_394_),
    .Q(\m1.U0.U0.b1.B ));
 sg13g2_dfrbp_1 _803_ (.CLK(clk),
    .RESET_B(net106),
    .D(net10),
    .Q_N(_395_),
    .Q(\m1.U0.U0.b1.D ));
 sg13g2_dfrbp_1 _804_ (.CLK(clk),
    .RESET_B(net106),
    .D(net11),
    .Q_N(_396_),
    .Q(\m1.U0.U1.b1.B ));
 sg13g2_dfrbp_1 _805_ (.CLK(clk),
    .RESET_B(net107),
    .D(net12),
    .Q_N(_397_),
    .Q(\m1.U0.U1.b1.D ));
 sg13g2_dfrbp_1 _806_ (.CLK(clk),
    .RESET_B(net107),
    .D(net13),
    .Q_N(_398_),
    .Q(\m1.U1.U0.b1.B ));
 sg13g2_dfrbp_1 _807_ (.CLK(clk),
    .RESET_B(net107),
    .D(net14),
    .Q_N(_399_),
    .Q(\m1.U1.U0.b1.D ));
 sg13g2_dfrbp_1 _808_ (.CLK(clk),
    .RESET_B(net107),
    .D(net15),
    .Q_N(_400_),
    .Q(\m1.U1.U1.b1.B ));
 sg13g2_dfrbp_1 _809_ (.CLK(clk),
    .RESET_B(net107),
    .D(net16),
    .Q_N(_393_),
    .Q(\m1.U1.U1.b1.D ));
 sg13g2_dfrbp_1 _810_ (.CLK(net17),
    .RESET_B(net107),
    .D(\a1.fa[0].fa0.S ),
    .Q_N(_392_),
    .Q(\a1.fa[0].fa0.A ));
 sg13g2_dfrbp_1 _811_ (.CLK(net18),
    .RESET_B(net107),
    .D(\a1.fa[0].fa1.S ),
    .Q_N(_391_),
    .Q(\a1.fa[0].fa1.A ));
 sg13g2_dfrbp_1 _812_ (.CLK(net19),
    .RESET_B(net107),
    .D(\a1.fa[0].fa2.S ),
    .Q_N(_390_),
    .Q(\a1.fa[0].fa2.A ));
 sg13g2_dfrbp_1 _813_ (.CLK(net20),
    .RESET_B(net105),
    .D(net40),
    .Q_N(_389_),
    .Q(\a1.fa[0].fa3.A ));
 sg13g2_dfrbp_1 _814_ (.CLK(net21),
    .RESET_B(net105),
    .D(\a1.fa[1].fa0.S ),
    .Q_N(_388_),
    .Q(\a1.fa[1].fa0.A ));
 sg13g2_dfrbp_1 _815_ (.CLK(net22),
    .RESET_B(net105),
    .D(net36),
    .Q_N(_387_),
    .Q(\a1.fa[1].fa1.A ));
 sg13g2_dfrbp_1 _816_ (.CLK(net23),
    .RESET_B(net105),
    .D(\a1.fa[1].fa2.S ),
    .Q_N(_386_),
    .Q(\a1.fa[1].fa2.A ));
 sg13g2_dfrbp_1 _817_ (.CLK(net24),
    .RESET_B(net105),
    .D(\a1.fa[1].fa3.S ),
    .Q_N(_385_),
    .Q(\a1.fa[1].fa3.A ));
 sg13g2_dfrbp_1 _818_ (.CLK(net25),
    .RESET_B(net104),
    .D(\a1.fa[2].fa0.S ),
    .Q_N(_384_),
    .Q(\a1.fa[2].fa0.A ));
 sg13g2_dfrbp_1 _819_ (.CLK(net26),
    .RESET_B(net104),
    .D(net44),
    .Q_N(_383_),
    .Q(\a1.fa[2].fa1.A ));
 sg13g2_dfrbp_1 _820_ (.CLK(net27),
    .RESET_B(net104),
    .D(\a1.fa[2].fa2.S ),
    .Q_N(_382_),
    .Q(\a1.fa[2].fa2.A ));
 sg13g2_dfrbp_1 _821_ (.CLK(net28),
    .RESET_B(net104),
    .D(\a1.fa[2].fa3.S ),
    .Q_N(_381_),
    .Q(\a1.fa[2].fa3.A ));
 sg13g2_dfrbp_1 _822_ (.CLK(net29),
    .RESET_B(net104),
    .D(\a1.fa[3].fa0.S ),
    .Q_N(_380_),
    .Q(\a1.fa[3].fa0.A ));
 sg13g2_dfrbp_1 _823_ (.CLK(net30),
    .RESET_B(net104),
    .D(net38),
    .Q_N(_379_),
    .Q(\a1.fa[3].fa1.A ));
 sg13g2_dfrbp_1 _824_ (.CLK(net31),
    .RESET_B(net104),
    .D(\a1.fa[3].fa2.S ),
    .Q_N(_378_),
    .Q(\a1.fa[3].fa2.A ));
 sg13g2_dfrbp_1 _825_ (.CLK(net32),
    .RESET_B(net104),
    .D(net48),
    .Q_N(_401_),
    .Q(\a1.fa[3].fa3.A ));
 sg13g2_dfrbp_1 _826_ (.CLK(clk),
    .RESET_B(net108),
    .D(net1),
    .Q_N(_402_),
    .Q(\m1.U0.U0.b1.A ));
 sg13g2_dfrbp_1 _827_ (.CLK(clk),
    .RESET_B(net108),
    .D(net2),
    .Q_N(_403_),
    .Q(\m1.U0.U0.p1.A ));
 sg13g2_dfrbp_1 _828_ (.CLK(clk),
    .RESET_B(net106),
    .D(net3),
    .Q_N(_404_),
    .Q(\m1.U0.U2.b1.A ));
 sg13g2_dfrbp_1 _829_ (.CLK(clk),
    .RESET_B(net106),
    .D(net4),
    .Q_N(_405_),
    .Q(\m1.U0.U2.p1.A ));
 sg13g2_dfrbp_1 _830_ (.CLK(clk),
    .RESET_B(net106),
    .D(net5),
    .Q_N(_406_),
    .Q(\m1.U2.U0.b1.A ));
 sg13g2_dfrbp_1 _831_ (.CLK(clk),
    .RESET_B(net108),
    .D(net6),
    .Q_N(_407_),
    .Q(\m1.U2.U0.p1.A ));
 sg13g2_dfrbp_1 _832_ (.CLK(clk),
    .RESET_B(net106),
    .D(net7),
    .Q_N(_408_),
    .Q(\m1.U2.U2.b1.A ));
 sg13g2_dfrbp_1 _833_ (.CLK(clk),
    .RESET_B(net106),
    .D(net8),
    .Q_N(_377_),
    .Q(\m1.U2.U2.p1.A ));
 sg13g2_buf_1 _834_ (.A(clk),
    .X(uio_oe[0]));
 sg13g2_buf_1 _835_ (.A(clk),
    .X(uio_oe[1]));
 sg13g2_buf_1 _836_ (.A(clk),
    .X(uio_oe[2]));
 sg13g2_buf_1 _837_ (.A(clk),
    .X(uio_oe[3]));
 sg13g2_buf_1 _838_ (.A(clk),
    .X(uio_oe[4]));
 sg13g2_buf_1 _839_ (.A(clk),
    .X(uio_oe[5]));
 sg13g2_buf_1 _840_ (.A(clk),
    .X(uio_oe[6]));
 sg13g2_buf_1 _841_ (.A(clk),
    .X(uio_oe[7]));
 sg13g2_buf_1 _842_ (.A(\a1.fa[2].fa0.A ),
    .X(uio_out[0]));
 sg13g2_buf_1 _843_ (.A(\a1.fa[2].fa1.A ),
    .X(uio_out[1]));
 sg13g2_buf_1 _844_ (.A(\a1.fa[2].fa2.A ),
    .X(uio_out[2]));
 sg13g2_buf_1 _845_ (.A(\a1.fa[2].fa3.A ),
    .X(uio_out[3]));
 sg13g2_buf_1 _846_ (.A(\a1.fa[3].fa0.A ),
    .X(uio_out[4]));
 sg13g2_buf_1 _847_ (.A(\a1.fa[3].fa1.A ),
    .X(uio_out[5]));
 sg13g2_buf_1 _848_ (.A(\a1.fa[3].fa2.A ),
    .X(uio_out[6]));
 sg13g2_buf_1 _849_ (.A(\a1.fa[3].fa3.A ),
    .X(uio_out[7]));
 sg13g2_buf_1 _850_ (.A(\a1.fa[0].fa0.A ),
    .X(uo_out[0]));
 sg13g2_buf_1 _851_ (.A(\a1.fa[0].fa1.A ),
    .X(uo_out[1]));
 sg13g2_buf_1 _852_ (.A(\a1.fa[0].fa2.A ),
    .X(uo_out[2]));
 sg13g2_buf_1 _853_ (.A(\a1.fa[0].fa3.A ),
    .X(uo_out[3]));
 sg13g2_buf_1 _854_ (.A(\a1.fa[1].fa0.A ),
    .X(uo_out[4]));
 sg13g2_buf_1 _855_ (.A(\a1.fa[1].fa1.A ),
    .X(uo_out[5]));
 sg13g2_buf_1 _856_ (.A(\a1.fa[1].fa2.A ),
    .X(uo_out[6]));
 sg13g2_buf_1 _857_ (.A(\a1.fa[1].fa3.A ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout82 (.A(\m1.U2.U2.p1.A ),
    .X(net82));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(\m1.U2.U2.b1.A ));
 sg13g2_buf_2 fanout84 (.A(\m1.U2.U0.p1.A ),
    .X(net84));
 sg13g2_buf_1 fanout85 (.A(\m1.U2.U0.p1.A ),
    .X(net85));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(\m1.U2.U0.b1.A ));
 sg13g2_buf_1 fanout87 (.A(\m1.U2.U0.b1.A ),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(\m1.U0.U2.p1.A ),
    .X(net88));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(\m1.U0.U2.b1.A ));
 sg13g2_buf_2 fanout90 (.A(\m1.U0.U2.b1.A ),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(\m1.U0.U0.p1.A ),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(\m1.U0.U0.b1.A ),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(\m1.U1.U1.b1.D ),
    .X(net93));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(\m1.U1.U1.b1.B ));
 sg13g2_buf_2 fanout95 (.A(\m1.U1.U0.b1.D ),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(\m1.U1.U0.b1.B ),
    .X(net96));
 sg13g2_buf_1 fanout97 (.A(\m1.U1.U0.b1.B ),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(\m1.U0.U1.b1.D ),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(\m1.U0.U1.b1.B ),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(\m1.U0.U0.b1.D ),
    .X(net100));
 sg13g2_buf_1 fanout101 (.A(\m1.U0.U0.b1.D ),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(\m1.U0.U0.b1.B ),
    .X(net102));
 sg13g2_buf_1 fanout103 (.A(\m1.U0.U0.b1.B ),
    .X(net103));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(net109));
 sg13g2_buf_2 fanout105 (.A(net109),
    .X(net105));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(net108));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(net109));
 sg13g2_buf_2 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(rst_n),
    .X(net109));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_inv_1 _411__1 (.Y(net17),
    .A(clk));
 sg13g2_dlygate4sd3_1 hold2 (.A(\a1.fa[0].fa1.A ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold3 (.A(\a1.fa[1].fa1.A ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold4 (.A(\a1.fa[1].fa1.S ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold5 (.A(\a1.fa[3].fa1.A ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold6 (.A(\a1.fa[3].fa1.S ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold7 (.A(\a1.fa[0].fa3.A ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold8 (.A(\a1.fa[0].fa3.S ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold9 (.A(\a1.fa[1].fa0.A ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold10 (.A(\a1.fa[0].fa2.A ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold11 (.A(\a1.fa[2].fa1.A ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold12 (.A(\a1.fa[2].fa1.S ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold13 (.A(\a1.fa[3].fa0.A ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold14 (.A(\a1.fa[1].fa2.A ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold15 (.A(\a1.fa[3].fa2.A ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold16 (.A(\a1.fa[3].fa3.S ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold17 (.A(\a1.fa[1].fa3.A ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold18 (.A(\a1.fa[2].fa0.A ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold19 (.A(\a1.fa[2].fa2.A ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold20 (.A(\a1.fa[2].fa3.A ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold21 (.A(\a1.fa[3].fa1.A ),
    .X(net53));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_fill_2 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_157 ();
 sg13g2_decap_4 FILLER_22_164 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_decap_4 FILLER_22_180 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_decap_4 FILLER_22_194 ();
 sg13g2_fill_2 FILLER_22_198 ();
 sg13g2_decap_8 FILLER_22_205 ();
 sg13g2_decap_8 FILLER_22_212 ();
 sg13g2_fill_1 FILLER_22_219 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_235 ();
 sg13g2_fill_2 FILLER_22_242 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_fill_1 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_279 ();
 sg13g2_decap_8 FILLER_22_286 ();
 sg13g2_decap_8 FILLER_22_293 ();
 sg13g2_decap_8 FILLER_22_300 ();
 sg13g2_decap_8 FILLER_22_307 ();
 sg13g2_decap_8 FILLER_22_314 ();
 sg13g2_decap_8 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_fill_1 FILLER_23_134 ();
 sg13g2_fill_1 FILLER_23_148 ();
 sg13g2_fill_2 FILLER_23_157 ();
 sg13g2_fill_1 FILLER_23_159 ();
 sg13g2_fill_2 FILLER_23_204 ();
 sg13g2_fill_1 FILLER_23_206 ();
 sg13g2_fill_2 FILLER_23_215 ();
 sg13g2_decap_8 FILLER_23_233 ();
 sg13g2_fill_2 FILLER_23_256 ();
 sg13g2_decap_4 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_297 ();
 sg13g2_decap_8 FILLER_23_304 ();
 sg13g2_decap_8 FILLER_23_311 ();
 sg13g2_decap_8 FILLER_23_318 ();
 sg13g2_decap_8 FILLER_23_325 ();
 sg13g2_decap_8 FILLER_23_332 ();
 sg13g2_decap_8 FILLER_23_339 ();
 sg13g2_decap_8 FILLER_23_346 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_8 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_88 ();
 sg13g2_fill_1 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_104 ();
 sg13g2_decap_4 FILLER_24_111 ();
 sg13g2_fill_2 FILLER_24_115 ();
 sg13g2_decap_8 FILLER_24_129 ();
 sg13g2_decap_4 FILLER_24_136 ();
 sg13g2_fill_2 FILLER_24_140 ();
 sg13g2_fill_2 FILLER_24_146 ();
 sg13g2_decap_4 FILLER_24_164 ();
 sg13g2_fill_1 FILLER_24_173 ();
 sg13g2_decap_8 FILLER_24_179 ();
 sg13g2_decap_4 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_fill_1 FILLER_24_196 ();
 sg13g2_decap_4 FILLER_24_210 ();
 sg13g2_fill_1 FILLER_24_214 ();
 sg13g2_fill_1 FILLER_24_220 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_254 ();
 sg13g2_fill_2 FILLER_24_261 ();
 sg13g2_fill_1 FILLER_24_263 ();
 sg13g2_decap_8 FILLER_24_274 ();
 sg13g2_fill_2 FILLER_24_285 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_52 ();
 sg13g2_decap_8 FILLER_25_59 ();
 sg13g2_decap_4 FILLER_25_66 ();
 sg13g2_fill_2 FILLER_25_70 ();
 sg13g2_fill_2 FILLER_25_85 ();
 sg13g2_decap_4 FILLER_25_110 ();
 sg13g2_decap_4 FILLER_25_160 ();
 sg13g2_decap_8 FILLER_25_188 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_fill_2 FILLER_25_210 ();
 sg13g2_fill_1 FILLER_25_212 ();
 sg13g2_decap_8 FILLER_25_229 ();
 sg13g2_fill_1 FILLER_25_236 ();
 sg13g2_decap_4 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_fill_1 FILLER_25_284 ();
 sg13g2_decap_8 FILLER_25_299 ();
 sg13g2_decap_8 FILLER_25_306 ();
 sg13g2_decap_8 FILLER_25_313 ();
 sg13g2_decap_8 FILLER_25_320 ();
 sg13g2_decap_8 FILLER_25_327 ();
 sg13g2_decap_8 FILLER_25_334 ();
 sg13g2_decap_8 FILLER_25_341 ();
 sg13g2_decap_8 FILLER_25_348 ();
 sg13g2_decap_8 FILLER_25_355 ();
 sg13g2_decap_8 FILLER_25_362 ();
 sg13g2_decap_8 FILLER_25_369 ();
 sg13g2_decap_8 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_fill_2 FILLER_26_42 ();
 sg13g2_fill_1 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_88 ();
 sg13g2_decap_4 FILLER_26_108 ();
 sg13g2_fill_1 FILLER_26_112 ();
 sg13g2_fill_2 FILLER_26_118 ();
 sg13g2_fill_1 FILLER_26_120 ();
 sg13g2_decap_4 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_138 ();
 sg13g2_fill_2 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_decap_8 FILLER_26_156 ();
 sg13g2_decap_4 FILLER_26_163 ();
 sg13g2_fill_2 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_fill_2 FILLER_26_189 ();
 sg13g2_fill_1 FILLER_26_191 ();
 sg13g2_fill_1 FILLER_26_221 ();
 sg13g2_decap_4 FILLER_26_238 ();
 sg13g2_fill_2 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_fill_1 FILLER_26_256 ();
 sg13g2_fill_2 FILLER_26_262 ();
 sg13g2_fill_1 FILLER_26_264 ();
 sg13g2_decap_4 FILLER_26_270 ();
 sg13g2_fill_2 FILLER_26_274 ();
 sg13g2_fill_2 FILLER_26_340 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_26_348 ();
 sg13g2_decap_8 FILLER_26_355 ();
 sg13g2_decap_8 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_46 ();
 sg13g2_decap_8 FILLER_27_53 ();
 sg13g2_decap_4 FILLER_27_86 ();
 sg13g2_fill_1 FILLER_27_90 ();
 sg13g2_fill_2 FILLER_27_108 ();
 sg13g2_fill_2 FILLER_27_126 ();
 sg13g2_decap_4 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_140 ();
 sg13g2_decap_4 FILLER_27_154 ();
 sg13g2_fill_1 FILLER_27_168 ();
 sg13g2_fill_1 FILLER_27_209 ();
 sg13g2_fill_2 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_229 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_decap_4 FILLER_27_240 ();
 sg13g2_fill_2 FILLER_27_249 ();
 sg13g2_fill_1 FILLER_27_264 ();
 sg13g2_fill_2 FILLER_27_281 ();
 sg13g2_fill_1 FILLER_27_283 ();
 sg13g2_fill_1 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_307 ();
 sg13g2_decap_4 FILLER_27_314 ();
 sg13g2_fill_1 FILLER_27_318 ();
 sg13g2_decap_4 FILLER_27_355 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_37 ();
 sg13g2_fill_2 FILLER_28_64 ();
 sg13g2_fill_1 FILLER_28_75 ();
 sg13g2_fill_1 FILLER_28_81 ();
 sg13g2_decap_4 FILLER_28_111 ();
 sg13g2_fill_2 FILLER_28_125 ();
 sg13g2_fill_1 FILLER_28_127 ();
 sg13g2_decap_8 FILLER_28_163 ();
 sg13g2_decap_8 FILLER_28_170 ();
 sg13g2_decap_8 FILLER_28_177 ();
 sg13g2_decap_8 FILLER_28_184 ();
 sg13g2_fill_1 FILLER_28_191 ();
 sg13g2_fill_2 FILLER_28_207 ();
 sg13g2_fill_1 FILLER_28_209 ();
 sg13g2_fill_1 FILLER_28_239 ();
 sg13g2_fill_2 FILLER_28_252 ();
 sg13g2_fill_1 FILLER_28_254 ();
 sg13g2_fill_1 FILLER_28_271 ();
 sg13g2_decap_8 FILLER_28_276 ();
 sg13g2_fill_1 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_304 ();
 sg13g2_fill_1 FILLER_28_311 ();
 sg13g2_fill_2 FILLER_28_333 ();
 sg13g2_fill_1 FILLER_28_335 ();
 sg13g2_decap_4 FILLER_28_341 ();
 sg13g2_decap_8 FILLER_28_351 ();
 sg13g2_fill_1 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_372 ();
 sg13g2_decap_8 FILLER_28_379 ();
 sg13g2_decap_8 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_4 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_49 ();
 sg13g2_decap_4 FILLER_29_85 ();
 sg13g2_fill_1 FILLER_29_89 ();
 sg13g2_fill_2 FILLER_29_99 ();
 sg13g2_fill_1 FILLER_29_101 ();
 sg13g2_decap_4 FILLER_29_110 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_134 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_142 ();
 sg13g2_fill_1 FILLER_29_149 ();
 sg13g2_decap_8 FILLER_29_155 ();
 sg13g2_decap_4 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_166 ();
 sg13g2_decap_8 FILLER_29_212 ();
 sg13g2_decap_4 FILLER_29_228 ();
 sg13g2_fill_2 FILLER_29_232 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_fill_2 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_297 ();
 sg13g2_decap_8 FILLER_29_306 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_decap_4 FILLER_29_329 ();
 sg13g2_fill_2 FILLER_29_339 ();
 sg13g2_fill_2 FILLER_29_346 ();
 sg13g2_decap_4 FILLER_29_357 ();
 sg13g2_fill_2 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_4 FILLER_30_35 ();
 sg13g2_fill_2 FILLER_30_39 ();
 sg13g2_fill_1 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_93 ();
 sg13g2_fill_1 FILLER_30_95 ();
 sg13g2_fill_2 FILLER_30_109 ();
 sg13g2_fill_1 FILLER_30_124 ();
 sg13g2_fill_1 FILLER_30_152 ();
 sg13g2_decap_4 FILLER_30_165 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_4 FILLER_30_189 ();
 sg13g2_fill_1 FILLER_30_193 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_214 ();
 sg13g2_decap_4 FILLER_30_233 ();
 sg13g2_fill_2 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_fill_2 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_314 ();
 sg13g2_fill_1 FILLER_30_339 ();
 sg13g2_decap_4 FILLER_30_349 ();
 sg13g2_fill_2 FILLER_30_353 ();
 sg13g2_decap_4 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_fill_2 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_109 ();
 sg13g2_decap_8 FILLER_31_113 ();
 sg13g2_decap_4 FILLER_31_137 ();
 sg13g2_fill_2 FILLER_31_141 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_fill_2 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_169 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_fill_1 FILLER_31_198 ();
 sg13g2_decap_4 FILLER_31_204 ();
 sg13g2_fill_1 FILLER_31_208 ();
 sg13g2_decap_4 FILLER_31_228 ();
 sg13g2_decap_4 FILLER_31_236 ();
 sg13g2_fill_1 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_4 FILLER_31_280 ();
 sg13g2_fill_2 FILLER_31_284 ();
 sg13g2_decap_8 FILLER_31_312 ();
 sg13g2_decap_4 FILLER_31_319 ();
 sg13g2_fill_2 FILLER_31_329 ();
 sg13g2_fill_2 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_345 ();
 sg13g2_decap_4 FILLER_31_352 ();
 sg13g2_fill_2 FILLER_31_356 ();
 sg13g2_decap_4 FILLER_31_379 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_63 ();
 sg13g2_fill_2 FILLER_32_102 ();
 sg13g2_fill_1 FILLER_32_104 ();
 sg13g2_fill_1 FILLER_32_152 ();
 sg13g2_fill_2 FILLER_32_170 ();
 sg13g2_fill_1 FILLER_32_172 ();
 sg13g2_fill_2 FILLER_32_204 ();
 sg13g2_fill_1 FILLER_32_206 ();
 sg13g2_fill_2 FILLER_32_211 ();
 sg13g2_fill_1 FILLER_32_213 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_239 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_327 ();
 sg13g2_fill_2 FILLER_32_354 ();
 sg13g2_fill_1 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_32_396 ();
 sg13g2_decap_4 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_fill_2 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_116 ();
 sg13g2_fill_1 FILLER_33_140 ();
 sg13g2_fill_2 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_160 ();
 sg13g2_decap_8 FILLER_33_184 ();
 sg13g2_decap_4 FILLER_33_191 ();
 sg13g2_decap_8 FILLER_33_212 ();
 sg13g2_fill_2 FILLER_33_219 ();
 sg13g2_fill_2 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_253 ();
 sg13g2_fill_1 FILLER_33_260 ();
 sg13g2_decap_8 FILLER_33_274 ();
 sg13g2_decap_8 FILLER_33_281 ();
 sg13g2_decap_8 FILLER_33_288 ();
 sg13g2_decap_8 FILLER_33_295 ();
 sg13g2_decap_8 FILLER_33_302 ();
 sg13g2_fill_2 FILLER_33_309 ();
 sg13g2_fill_1 FILLER_33_311 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_fill_2 FILLER_33_332 ();
 sg13g2_fill_1 FILLER_33_334 ();
 sg13g2_fill_2 FILLER_33_364 ();
 sg13g2_fill_1 FILLER_33_366 ();
 sg13g2_decap_4 FILLER_33_373 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_4 FILLER_34_102 ();
 sg13g2_fill_2 FILLER_34_106 ();
 sg13g2_fill_1 FILLER_34_134 ();
 sg13g2_fill_1 FILLER_34_153 ();
 sg13g2_decap_8 FILLER_34_166 ();
 sg13g2_decap_8 FILLER_34_173 ();
 sg13g2_decap_8 FILLER_34_180 ();
 sg13g2_decap_8 FILLER_34_187 ();
 sg13g2_fill_1 FILLER_34_194 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_4 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_228 ();
 sg13g2_fill_2 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_247 ();
 sg13g2_decap_4 FILLER_34_266 ();
 sg13g2_fill_1 FILLER_34_270 ();
 sg13g2_decap_4 FILLER_34_326 ();
 sg13g2_fill_1 FILLER_34_330 ();
 sg13g2_decap_4 FILLER_34_334 ();
 sg13g2_fill_1 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_344 ();
 sg13g2_fill_2 FILLER_34_360 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_decap_8 FILLER_34_375 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_4 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_57 ();
 sg13g2_decap_8 FILLER_35_64 ();
 sg13g2_decap_8 FILLER_35_71 ();
 sg13g2_decap_8 FILLER_35_78 ();
 sg13g2_decap_8 FILLER_35_85 ();
 sg13g2_decap_8 FILLER_35_92 ();
 sg13g2_decap_8 FILLER_35_99 ();
 sg13g2_decap_8 FILLER_35_106 ();
 sg13g2_decap_8 FILLER_35_113 ();
 sg13g2_decap_8 FILLER_35_120 ();
 sg13g2_fill_2 FILLER_35_165 ();
 sg13g2_fill_1 FILLER_35_193 ();
 sg13g2_fill_2 FILLER_35_253 ();
 sg13g2_decap_8 FILLER_35_281 ();
 sg13g2_decap_8 FILLER_35_288 ();
 sg13g2_decap_4 FILLER_35_295 ();
 sg13g2_fill_1 FILLER_35_299 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_fill_2 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_122 ();
 sg13g2_decap_8 FILLER_36_129 ();
 sg13g2_fill_2 FILLER_36_136 ();
 sg13g2_decap_8 FILLER_36_144 ();
 sg13g2_fill_2 FILLER_36_151 ();
 sg13g2_fill_1 FILLER_36_171 ();
 sg13g2_decap_4 FILLER_36_175 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_decap_4 FILLER_36_207 ();
 sg13g2_decap_8 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_269 ();
 sg13g2_fill_2 FILLER_36_276 ();
 sg13g2_decap_8 FILLER_36_285 ();
 sg13g2_decap_4 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_343 ();
 sg13g2_fill_1 FILLER_36_349 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_fill_2 FILLER_37_42 ();
 sg13g2_fill_2 FILLER_37_48 ();
 sg13g2_decap_8 FILLER_37_54 ();
 sg13g2_decap_8 FILLER_37_61 ();
 sg13g2_decap_8 FILLER_37_68 ();
 sg13g2_decap_8 FILLER_37_75 ();
 sg13g2_decap_8 FILLER_37_82 ();
 sg13g2_decap_8 FILLER_37_89 ();
 sg13g2_decap_8 FILLER_37_96 ();
 sg13g2_decap_8 FILLER_37_103 ();
 sg13g2_decap_8 FILLER_37_110 ();
 sg13g2_decap_8 FILLER_37_117 ();
 sg13g2_decap_8 FILLER_37_124 ();
 sg13g2_decap_8 FILLER_37_131 ();
 sg13g2_decap_8 FILLER_37_138 ();
 sg13g2_decap_8 FILLER_37_145 ();
 sg13g2_fill_2 FILLER_37_152 ();
 sg13g2_decap_8 FILLER_37_158 ();
 sg13g2_decap_8 FILLER_37_165 ();
 sg13g2_decap_8 FILLER_37_172 ();
 sg13g2_decap_8 FILLER_37_179 ();
 sg13g2_fill_1 FILLER_37_186 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_4 FILLER_37_203 ();
 sg13g2_fill_1 FILLER_37_207 ();
 sg13g2_fill_1 FILLER_37_234 ();
 sg13g2_fill_1 FILLER_37_251 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_fill_2 FILLER_38_210 ();
 sg13g2_fill_1 FILLER_38_212 ();
 sg13g2_decap_8 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_223 ();
 sg13g2_fill_2 FILLER_38_252 ();
 sg13g2_fill_2 FILLER_38_297 ();
 sg13g2_fill_2 FILLER_38_331 ();
 sg13g2_fill_1 FILLER_38_333 ();
 sg13g2_fill_1 FILLER_38_365 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
endmodule

module tt_um_simon_cipher (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire clknet_leaf_0_clk;
 wire \bitserial_cipher.bit_counter[0] ;
 wire \bitserial_cipher.bit_counter[1] ;
 wire \bitserial_cipher.bit_counter[2] ;
 wire \bitserial_cipher.bit_counter[3] ;
 wire \bitserial_cipher.bit_counter[4] ;
 wire \bitserial_cipher.bit_counter[5] ;
 wire \bitserial_cipher.cipher_data ;
 wire \bitserial_cipher.datapath.fifo_ff56 ;
 wire \bitserial_cipher.datapath.fifo_ff57 ;
 wire \bitserial_cipher.datapath.fifo_ff58 ;
 wire \bitserial_cipher.datapath.fifo_ff59 ;
 wire \bitserial_cipher.datapath.fifo_ff60 ;
 wire \bitserial_cipher.datapath.fifo_ff61 ;
 wire \bitserial_cipher.datapath.fifo_ff62 ;
 wire \bitserial_cipher.datapath.fifo_ff63 ;
 wire \bitserial_cipher.datapath.key_in ;
 wire \bitserial_cipher.datapath.lut_ff56 ;
 wire \bitserial_cipher.datapath.lut_ff57 ;
 wire \bitserial_cipher.datapath.lut_ff58 ;
 wire \bitserial_cipher.datapath.lut_ff59 ;
 wire \bitserial_cipher.datapath.lut_ff60 ;
 wire \bitserial_cipher.datapath.lut_ff61 ;
 wire \bitserial_cipher.datapath.lut_ff62 ;
 wire \bitserial_cipher.datapath.lut_ff63 ;
 wire \bitserial_cipher.datapath.round_counter[0] ;
 wire \bitserial_cipher.datapath.round_counter[1] ;
 wire \bitserial_cipher.datapath.round_counter[2] ;
 wire \bitserial_cipher.datapath.round_counter[3] ;
 wire \bitserial_cipher.datapath.round_counter[4] ;
 wire \bitserial_cipher.datapath.round_counter[5] ;
 wire \bitserial_cipher.datapath.round_counter[6] ;
 wire \bitserial_cipher.datapath.shift_in2 ;
 wire \bitserial_cipher.datapath.shifter1[10] ;
 wire \bitserial_cipher.datapath.shifter1[11] ;
 wire \bitserial_cipher.datapath.shifter1[12] ;
 wire \bitserial_cipher.datapath.shifter1[13] ;
 wire \bitserial_cipher.datapath.shifter1[14] ;
 wire \bitserial_cipher.datapath.shifter1[15] ;
 wire \bitserial_cipher.datapath.shifter1[16] ;
 wire \bitserial_cipher.datapath.shifter1[17] ;
 wire \bitserial_cipher.datapath.shifter1[18] ;
 wire \bitserial_cipher.datapath.shifter1[19] ;
 wire \bitserial_cipher.datapath.shifter1[1] ;
 wire \bitserial_cipher.datapath.shifter1[20] ;
 wire \bitserial_cipher.datapath.shifter1[21] ;
 wire \bitserial_cipher.datapath.shifter1[22] ;
 wire \bitserial_cipher.datapath.shifter1[23] ;
 wire \bitserial_cipher.datapath.shifter1[24] ;
 wire \bitserial_cipher.datapath.shifter1[25] ;
 wire \bitserial_cipher.datapath.shifter1[26] ;
 wire \bitserial_cipher.datapath.shifter1[27] ;
 wire \bitserial_cipher.datapath.shifter1[28] ;
 wire \bitserial_cipher.datapath.shifter1[29] ;
 wire \bitserial_cipher.datapath.shifter1[2] ;
 wire \bitserial_cipher.datapath.shifter1[30] ;
 wire \bitserial_cipher.datapath.shifter1[31] ;
 wire \bitserial_cipher.datapath.shifter1[32] ;
 wire \bitserial_cipher.datapath.shifter1[33] ;
 wire \bitserial_cipher.datapath.shifter1[34] ;
 wire \bitserial_cipher.datapath.shifter1[35] ;
 wire \bitserial_cipher.datapath.shifter1[36] ;
 wire \bitserial_cipher.datapath.shifter1[37] ;
 wire \bitserial_cipher.datapath.shifter1[38] ;
 wire \bitserial_cipher.datapath.shifter1[39] ;
 wire \bitserial_cipher.datapath.shifter1[3] ;
 wire \bitserial_cipher.datapath.shifter1[40] ;
 wire \bitserial_cipher.datapath.shifter1[41] ;
 wire \bitserial_cipher.datapath.shifter1[42] ;
 wire \bitserial_cipher.datapath.shifter1[43] ;
 wire \bitserial_cipher.datapath.shifter1[44] ;
 wire \bitserial_cipher.datapath.shifter1[45] ;
 wire \bitserial_cipher.datapath.shifter1[46] ;
 wire \bitserial_cipher.datapath.shifter1[47] ;
 wire \bitserial_cipher.datapath.shifter1[48] ;
 wire \bitserial_cipher.datapath.shifter1[49] ;
 wire \bitserial_cipher.datapath.shifter1[4] ;
 wire \bitserial_cipher.datapath.shifter1[50] ;
 wire \bitserial_cipher.datapath.shifter1[51] ;
 wire \bitserial_cipher.datapath.shifter1[52] ;
 wire \bitserial_cipher.datapath.shifter1[53] ;
 wire \bitserial_cipher.datapath.shifter1[54] ;
 wire \bitserial_cipher.datapath.shifter1[55] ;
 wire \bitserial_cipher.datapath.shifter1[5] ;
 wire \bitserial_cipher.datapath.shifter1[6] ;
 wire \bitserial_cipher.datapath.shifter1[7] ;
 wire \bitserial_cipher.datapath.shifter1[8] ;
 wire \bitserial_cipher.datapath.shifter1[9] ;
 wire \bitserial_cipher.datapath.shifter2[10] ;
 wire \bitserial_cipher.datapath.shifter2[11] ;
 wire \bitserial_cipher.datapath.shifter2[12] ;
 wire \bitserial_cipher.datapath.shifter2[13] ;
 wire \bitserial_cipher.datapath.shifter2[14] ;
 wire \bitserial_cipher.datapath.shifter2[15] ;
 wire \bitserial_cipher.datapath.shifter2[16] ;
 wire \bitserial_cipher.datapath.shifter2[17] ;
 wire \bitserial_cipher.datapath.shifter2[18] ;
 wire \bitserial_cipher.datapath.shifter2[19] ;
 wire \bitserial_cipher.datapath.shifter2[1] ;
 wire \bitserial_cipher.datapath.shifter2[20] ;
 wire \bitserial_cipher.datapath.shifter2[21] ;
 wire \bitserial_cipher.datapath.shifter2[22] ;
 wire \bitserial_cipher.datapath.shifter2[23] ;
 wire \bitserial_cipher.datapath.shifter2[24] ;
 wire \bitserial_cipher.datapath.shifter2[25] ;
 wire \bitserial_cipher.datapath.shifter2[26] ;
 wire \bitserial_cipher.datapath.shifter2[27] ;
 wire \bitserial_cipher.datapath.shifter2[28] ;
 wire \bitserial_cipher.datapath.shifter2[29] ;
 wire \bitserial_cipher.datapath.shifter2[2] ;
 wire \bitserial_cipher.datapath.shifter2[30] ;
 wire \bitserial_cipher.datapath.shifter2[31] ;
 wire \bitserial_cipher.datapath.shifter2[32] ;
 wire \bitserial_cipher.datapath.shifter2[33] ;
 wire \bitserial_cipher.datapath.shifter2[34] ;
 wire \bitserial_cipher.datapath.shifter2[35] ;
 wire \bitserial_cipher.datapath.shifter2[36] ;
 wire \bitserial_cipher.datapath.shifter2[37] ;
 wire \bitserial_cipher.datapath.shifter2[38] ;
 wire \bitserial_cipher.datapath.shifter2[39] ;
 wire \bitserial_cipher.datapath.shifter2[3] ;
 wire \bitserial_cipher.datapath.shifter2[40] ;
 wire \bitserial_cipher.datapath.shifter2[41] ;
 wire \bitserial_cipher.datapath.shifter2[42] ;
 wire \bitserial_cipher.datapath.shifter2[43] ;
 wire \bitserial_cipher.datapath.shifter2[44] ;
 wire \bitserial_cipher.datapath.shifter2[45] ;
 wire \bitserial_cipher.datapath.shifter2[46] ;
 wire \bitserial_cipher.datapath.shifter2[47] ;
 wire \bitserial_cipher.datapath.shifter2[48] ;
 wire \bitserial_cipher.datapath.shifter2[49] ;
 wire \bitserial_cipher.datapath.shifter2[4] ;
 wire \bitserial_cipher.datapath.shifter2[50] ;
 wire \bitserial_cipher.datapath.shifter2[51] ;
 wire \bitserial_cipher.datapath.shifter2[52] ;
 wire \bitserial_cipher.datapath.shifter2[53] ;
 wire \bitserial_cipher.datapath.shifter2[54] ;
 wire \bitserial_cipher.datapath.shifter2[55] ;
 wire \bitserial_cipher.datapath.shifter2[56] ;
 wire \bitserial_cipher.datapath.shifter2[57] ;
 wire \bitserial_cipher.datapath.shifter2[58] ;
 wire \bitserial_cipher.datapath.shifter2[59] ;
 wire \bitserial_cipher.datapath.shifter2[5] ;
 wire \bitserial_cipher.datapath.shifter2[60] ;
 wire \bitserial_cipher.datapath.shifter2[61] ;
 wire \bitserial_cipher.datapath.shifter2[62] ;
 wire \bitserial_cipher.datapath.shifter2[63] ;
 wire \bitserial_cipher.datapath.shifter2[6] ;
 wire \bitserial_cipher.datapath.shifter2[7] ;
 wire \bitserial_cipher.datapath.shifter2[8] ;
 wire \bitserial_cipher.datapath.shifter2[9] ;
 wire \bitserial_cipher.datapath.valid ;
 wire \bitserial_cipher.key_exp.fifo_ff0 ;
 wire \bitserial_cipher.key_exp.fifo_ff1 ;
 wire \bitserial_cipher.key_exp.fifo_ff2 ;
 wire \bitserial_cipher.key_exp.fifo_ff3 ;
 wire \bitserial_cipher.key_exp.lut_ff0 ;
 wire \bitserial_cipher.key_exp.lut_ff1 ;
 wire \bitserial_cipher.key_exp.lut_ff2 ;
 wire \bitserial_cipher.key_exp.lut_ff3 ;
 wire \bitserial_cipher.key_exp.shift_out1 ;
 wire \bitserial_cipher.key_exp.shifter1[10] ;
 wire \bitserial_cipher.key_exp.shifter1[11] ;
 wire \bitserial_cipher.key_exp.shifter1[12] ;
 wire \bitserial_cipher.key_exp.shifter1[13] ;
 wire \bitserial_cipher.key_exp.shifter1[14] ;
 wire \bitserial_cipher.key_exp.shifter1[15] ;
 wire \bitserial_cipher.key_exp.shifter1[16] ;
 wire \bitserial_cipher.key_exp.shifter1[17] ;
 wire \bitserial_cipher.key_exp.shifter1[18] ;
 wire \bitserial_cipher.key_exp.shifter1[19] ;
 wire \bitserial_cipher.key_exp.shifter1[1] ;
 wire \bitserial_cipher.key_exp.shifter1[20] ;
 wire \bitserial_cipher.key_exp.shifter1[21] ;
 wire \bitserial_cipher.key_exp.shifter1[22] ;
 wire \bitserial_cipher.key_exp.shifter1[23] ;
 wire \bitserial_cipher.key_exp.shifter1[24] ;
 wire \bitserial_cipher.key_exp.shifter1[25] ;
 wire \bitserial_cipher.key_exp.shifter1[26] ;
 wire \bitserial_cipher.key_exp.shifter1[27] ;
 wire \bitserial_cipher.key_exp.shifter1[28] ;
 wire \bitserial_cipher.key_exp.shifter1[29] ;
 wire \bitserial_cipher.key_exp.shifter1[2] ;
 wire \bitserial_cipher.key_exp.shifter1[30] ;
 wire \bitserial_cipher.key_exp.shifter1[31] ;
 wire \bitserial_cipher.key_exp.shifter1[32] ;
 wire \bitserial_cipher.key_exp.shifter1[33] ;
 wire \bitserial_cipher.key_exp.shifter1[34] ;
 wire \bitserial_cipher.key_exp.shifter1[35] ;
 wire \bitserial_cipher.key_exp.shifter1[36] ;
 wire \bitserial_cipher.key_exp.shifter1[37] ;
 wire \bitserial_cipher.key_exp.shifter1[38] ;
 wire \bitserial_cipher.key_exp.shifter1[39] ;
 wire \bitserial_cipher.key_exp.shifter1[3] ;
 wire \bitserial_cipher.key_exp.shifter1[40] ;
 wire \bitserial_cipher.key_exp.shifter1[41] ;
 wire \bitserial_cipher.key_exp.shifter1[42] ;
 wire \bitserial_cipher.key_exp.shifter1[43] ;
 wire \bitserial_cipher.key_exp.shifter1[44] ;
 wire \bitserial_cipher.key_exp.shifter1[45] ;
 wire \bitserial_cipher.key_exp.shifter1[46] ;
 wire \bitserial_cipher.key_exp.shifter1[47] ;
 wire \bitserial_cipher.key_exp.shifter1[48] ;
 wire \bitserial_cipher.key_exp.shifter1[49] ;
 wire \bitserial_cipher.key_exp.shifter1[4] ;
 wire \bitserial_cipher.key_exp.shifter1[50] ;
 wire \bitserial_cipher.key_exp.shifter1[51] ;
 wire \bitserial_cipher.key_exp.shifter1[52] ;
 wire \bitserial_cipher.key_exp.shifter1[53] ;
 wire \bitserial_cipher.key_exp.shifter1[54] ;
 wire \bitserial_cipher.key_exp.shifter1[55] ;
 wire \bitserial_cipher.key_exp.shifter1[56] ;
 wire \bitserial_cipher.key_exp.shifter1[57] ;
 wire \bitserial_cipher.key_exp.shifter1[58] ;
 wire \bitserial_cipher.key_exp.shifter1[59] ;
 wire \bitserial_cipher.key_exp.shifter1[5] ;
 wire \bitserial_cipher.key_exp.shifter1[6] ;
 wire \bitserial_cipher.key_exp.shifter1[7] ;
 wire \bitserial_cipher.key_exp.shifter1[8] ;
 wire \bitserial_cipher.key_exp.shifter1[9] ;
 wire \bitserial_cipher.key_exp.shifter2[10] ;
 wire \bitserial_cipher.key_exp.shifter2[11] ;
 wire \bitserial_cipher.key_exp.shifter2[12] ;
 wire \bitserial_cipher.key_exp.shifter2[13] ;
 wire \bitserial_cipher.key_exp.shifter2[14] ;
 wire \bitserial_cipher.key_exp.shifter2[15] ;
 wire \bitserial_cipher.key_exp.shifter2[16] ;
 wire \bitserial_cipher.key_exp.shifter2[17] ;
 wire \bitserial_cipher.key_exp.shifter2[18] ;
 wire \bitserial_cipher.key_exp.shifter2[19] ;
 wire \bitserial_cipher.key_exp.shifter2[1] ;
 wire \bitserial_cipher.key_exp.shifter2[20] ;
 wire \bitserial_cipher.key_exp.shifter2[21] ;
 wire \bitserial_cipher.key_exp.shifter2[22] ;
 wire \bitserial_cipher.key_exp.shifter2[23] ;
 wire \bitserial_cipher.key_exp.shifter2[24] ;
 wire \bitserial_cipher.key_exp.shifter2[25] ;
 wire \bitserial_cipher.key_exp.shifter2[26] ;
 wire \bitserial_cipher.key_exp.shifter2[27] ;
 wire \bitserial_cipher.key_exp.shifter2[28] ;
 wire \bitserial_cipher.key_exp.shifter2[29] ;
 wire \bitserial_cipher.key_exp.shifter2[2] ;
 wire \bitserial_cipher.key_exp.shifter2[30] ;
 wire \bitserial_cipher.key_exp.shifter2[31] ;
 wire \bitserial_cipher.key_exp.shifter2[32] ;
 wire \bitserial_cipher.key_exp.shifter2[33] ;
 wire \bitserial_cipher.key_exp.shifter2[34] ;
 wire \bitserial_cipher.key_exp.shifter2[35] ;
 wire \bitserial_cipher.key_exp.shifter2[36] ;
 wire \bitserial_cipher.key_exp.shifter2[37] ;
 wire \bitserial_cipher.key_exp.shifter2[38] ;
 wire \bitserial_cipher.key_exp.shifter2[39] ;
 wire \bitserial_cipher.key_exp.shifter2[3] ;
 wire \bitserial_cipher.key_exp.shifter2[40] ;
 wire \bitserial_cipher.key_exp.shifter2[41] ;
 wire \bitserial_cipher.key_exp.shifter2[42] ;
 wire \bitserial_cipher.key_exp.shifter2[43] ;
 wire \bitserial_cipher.key_exp.shifter2[44] ;
 wire \bitserial_cipher.key_exp.shifter2[45] ;
 wire \bitserial_cipher.key_exp.shifter2[46] ;
 wire \bitserial_cipher.key_exp.shifter2[47] ;
 wire \bitserial_cipher.key_exp.shifter2[48] ;
 wire \bitserial_cipher.key_exp.shifter2[49] ;
 wire \bitserial_cipher.key_exp.shifter2[4] ;
 wire \bitserial_cipher.key_exp.shifter2[50] ;
 wire \bitserial_cipher.key_exp.shifter2[51] ;
 wire \bitserial_cipher.key_exp.shifter2[52] ;
 wire \bitserial_cipher.key_exp.shifter2[53] ;
 wire \bitserial_cipher.key_exp.shifter2[54] ;
 wire \bitserial_cipher.key_exp.shifter2[55] ;
 wire \bitserial_cipher.key_exp.shifter2[56] ;
 wire \bitserial_cipher.key_exp.shifter2[57] ;
 wire \bitserial_cipher.key_exp.shifter2[58] ;
 wire \bitserial_cipher.key_exp.shifter2[59] ;
 wire \bitserial_cipher.key_exp.shifter2[5] ;
 wire \bitserial_cipher.key_exp.shifter2[60] ;
 wire \bitserial_cipher.key_exp.shifter2[61] ;
 wire \bitserial_cipher.key_exp.shifter2[62] ;
 wire \bitserial_cipher.key_exp.shifter2[63] ;
 wire \bitserial_cipher.key_exp.shifter2[6] ;
 wire \bitserial_cipher.key_exp.shifter2[7] ;
 wire \bitserial_cipher.key_exp.shifter2[8] ;
 wire \bitserial_cipher.key_exp.shifter2[9] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net1;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;

 sg13g2_inv_1 _1481_ (.Y(_0576_),
    .A(net434));
 sg13g2_inv_1 _1482_ (.Y(_0577_),
    .A(net808));
 sg13g2_inv_1 _1483_ (.Y(_0578_),
    .A(net625));
 sg13g2_inv_1 _1484_ (.Y(_0579_),
    .A(net608));
 sg13g2_inv_1 _1485_ (.Y(_0580_),
    .A(net368));
 sg13g2_inv_1 _1486_ (.Y(_0581_),
    .A(net689));
 sg13g2_inv_1 _1487_ (.Y(_0582_),
    .A(net378));
 sg13g2_inv_1 _1488_ (.Y(_0583_),
    .A(net766));
 sg13g2_inv_1 _1489_ (.Y(_0584_),
    .A(net727));
 sg13g2_inv_1 _1490_ (.Y(_0585_),
    .A(net782));
 sg13g2_inv_1 _1491_ (.Y(_0586_),
    .A(net333));
 sg13g2_inv_1 _1492_ (.Y(_0587_),
    .A(net692));
 sg13g2_inv_1 _1493_ (.Y(_0588_),
    .A(net587));
 sg13g2_inv_1 _1494_ (.Y(_0589_),
    .A(net620));
 sg13g2_inv_1 _1495_ (.Y(_0590_),
    .A(net602));
 sg13g2_inv_1 _1496_ (.Y(_0591_),
    .A(net684));
 sg13g2_inv_1 _1497_ (.Y(_0592_),
    .A(net714));
 sg13g2_inv_1 _1498_ (.Y(_0593_),
    .A(net674));
 sg13g2_inv_1 _1499_ (.Y(_0594_),
    .A(net805));
 sg13g2_inv_1 _1500_ (.Y(_0595_),
    .A(net663));
 sg13g2_inv_1 _1501_ (.Y(_0596_),
    .A(net813));
 sg13g2_inv_1 _1502_ (.Y(_0597_),
    .A(net314));
 sg13g2_inv_1 _1503_ (.Y(_0598_),
    .A(net773));
 sg13g2_inv_1 _1504_ (.Y(_0599_),
    .A(net654));
 sg13g2_inv_1 _1505_ (.Y(_0600_),
    .A(net720));
 sg13g2_inv_1 _1506_ (.Y(_0601_),
    .A(net844));
 sg13g2_inv_1 _1507_ (.Y(_0602_),
    .A(net310));
 sg13g2_inv_1 _1508_ (.Y(_0603_),
    .A(net833));
 sg13g2_inv_1 _1509_ (.Y(_0604_),
    .A(net704));
 sg13g2_inv_1 _1510_ (.Y(_0605_),
    .A(net600));
 sg13g2_inv_1 _1511_ (.Y(_0606_),
    .A(net832));
 sg13g2_inv_1 _1512_ (.Y(_0607_),
    .A(net768));
 sg13g2_inv_1 _1513_ (.Y(_0608_),
    .A(net763));
 sg13g2_inv_1 _1514_ (.Y(_0609_),
    .A(net671));
 sg13g2_inv_1 _1515_ (.Y(_0610_),
    .A(net627));
 sg13g2_inv_1 _1516_ (.Y(_0611_),
    .A(net711));
 sg13g2_inv_1 _1517_ (.Y(_0612_),
    .A(net436));
 sg13g2_inv_1 _1518_ (.Y(_0613_),
    .A(net794));
 sg13g2_inv_1 _1519_ (.Y(_0614_),
    .A(net841));
 sg13g2_inv_1 _1520_ (.Y(_0615_),
    .A(net636));
 sg13g2_inv_1 _1521_ (.Y(_0616_),
    .A(net335));
 sg13g2_inv_1 _1522_ (.Y(_0617_),
    .A(net746));
 sg13g2_inv_1 _1523_ (.Y(_0618_),
    .A(net756));
 sg13g2_inv_1 _1524_ (.Y(_0619_),
    .A(net786));
 sg13g2_inv_1 _1525_ (.Y(_0620_),
    .A(net838));
 sg13g2_inv_1 _1526_ (.Y(_0621_),
    .A(net440));
 sg13g2_inv_1 _1527_ (.Y(_0622_),
    .A(net611));
 sg13g2_inv_1 _1528_ (.Y(_0623_),
    .A(net834));
 sg13g2_inv_1 _1529_ (.Y(_0624_),
    .A(net823));
 sg13g2_inv_1 _1530_ (.Y(_0625_),
    .A(net646));
 sg13g2_inv_1 _1531_ (.Y(_0626_),
    .A(net355));
 sg13g2_inv_1 _1532_ (.Y(_0627_),
    .A(net845));
 sg13g2_inv_1 _1533_ (.Y(_0628_),
    .A(net416));
 sg13g2_inv_1 _1534_ (.Y(_0629_),
    .A(net761));
 sg13g2_inv_1 _1535_ (.Y(_0630_),
    .A(net793));
 sg13g2_inv_1 _1536_ (.Y(_0631_),
    .A(net347));
 sg13g2_inv_1 _1537_ (.Y(_0632_),
    .A(net680));
 sg13g2_inv_1 _1538_ (.Y(_0633_),
    .A(net785));
 sg13g2_inv_1 _1539_ (.Y(_0634_),
    .A(net394));
 sg13g2_inv_1 _1540_ (.Y(_0635_),
    .A(net801));
 sg13g2_inv_1 _1541_ (.Y(_0636_),
    .A(net609));
 sg13g2_inv_1 _1542_ (.Y(_0637_),
    .A(net329));
 sg13g2_inv_1 _1543_ (.Y(_0638_),
    .A(net583));
 sg13g2_inv_1 _1544_ (.Y(_0639_),
    .A(net764));
 sg13g2_inv_1 _1545_ (.Y(_0640_),
    .A(net826));
 sg13g2_inv_1 _1546_ (.Y(_0641_),
    .A(net807));
 sg13g2_inv_1 _1547_ (.Y(_0642_),
    .A(net312));
 sg13g2_inv_1 _1548_ (.Y(_0643_),
    .A(net776));
 sg13g2_inv_1 _1549_ (.Y(_0644_),
    .A(net837));
 sg13g2_inv_1 _1550_ (.Y(_0645_),
    .A(net737));
 sg13g2_inv_1 _1551_ (.Y(_0646_),
    .A(net345));
 sg13g2_inv_1 _1552_ (.Y(_0647_),
    .A(net732));
 sg13g2_inv_1 _1553_ (.Y(_0648_),
    .A(net339));
 sg13g2_inv_1 _1554_ (.Y(_0649_),
    .A(net406));
 sg13g2_inv_1 _1555_ (.Y(_0650_),
    .A(net769));
 sg13g2_inv_1 _1556_ (.Y(_0651_),
    .A(net729));
 sg13g2_inv_1 _1557_ (.Y(_0652_),
    .A(net814));
 sg13g2_inv_1 _1558_ (.Y(_0653_),
    .A(net715));
 sg13g2_inv_1 _1559_ (.Y(_0654_),
    .A(net725));
 sg13g2_inv_1 _1560_ (.Y(_0655_),
    .A(net640));
 sg13g2_inv_1 _1561_ (.Y(_0656_),
    .A(net364));
 sg13g2_inv_1 _1562_ (.Y(_0657_),
    .A(net425));
 sg13g2_inv_1 _1563_ (.Y(_0658_),
    .A(net733));
 sg13g2_inv_1 _1564_ (.Y(_0659_),
    .A(net656));
 sg13g2_inv_1 _1565_ (.Y(_0660_),
    .A(net806));
 sg13g2_inv_1 _1566_ (.Y(_0661_),
    .A(net755));
 sg13g2_inv_1 _1567_ (.Y(_0662_),
    .A(net414));
 sg13g2_inv_1 _1568_ (.Y(_0663_),
    .A(net771));
 sg13g2_inv_1 _1569_ (.Y(_0664_),
    .A(net612));
 sg13g2_inv_1 _1570_ (.Y(_0665_),
    .A(net392));
 sg13g2_inv_1 _1571_ (.Y(_0666_),
    .A(net706));
 sg13g2_inv_1 _1572_ (.Y(_0667_),
    .A(net710));
 sg13g2_inv_1 _1573_ (.Y(_0668_),
    .A(net380));
 sg13g2_inv_1 _1574_ (.Y(_0669_),
    .A(net408));
 sg13g2_inv_1 _1575_ (.Y(_0670_),
    .A(net731));
 sg13g2_inv_1 _1576_ (.Y(_0671_),
    .A(net623));
 sg13g2_inv_1 _1577_ (.Y(_0672_),
    .A(net633));
 sg13g2_inv_1 _1578_ (.Y(_0673_),
    .A(net351));
 sg13g2_inv_1 _1579_ (.Y(_0674_),
    .A(net666));
 sg13g2_inv_1 _1580_ (.Y(_0675_),
    .A(net422));
 sg13g2_inv_1 _1581_ (.Y(_0676_),
    .A(net758));
 sg13g2_inv_1 _1582_ (.Y(_0677_),
    .A(net676));
 sg13g2_inv_1 _1583_ (.Y(_0678_),
    .A(net712));
 sg13g2_inv_1 _1584_ (.Y(_0679_),
    .A(net384));
 sg13g2_inv_1 _1585_ (.Y(_0680_),
    .A(net695));
 sg13g2_inv_1 _1586_ (.Y(_0681_),
    .A(net741));
 sg13g2_inv_1 _1587_ (.Y(_0682_),
    .A(net661));
 sg13g2_inv_1 _1588_ (.Y(_0683_),
    .A(net386));
 sg13g2_inv_1 _1589_ (.Y(_0684_),
    .A(net366));
 sg13g2_inv_1 _1590_ (.Y(_0685_),
    .A(net400));
 sg13g2_inv_1 _1591_ (.Y(_0686_),
    .A(net701));
 sg13g2_inv_1 _1592_ (.Y(_0687_),
    .A(net420));
 sg13g2_inv_1 _1593_ (.Y(_0688_),
    .A(net752));
 sg13g2_inv_1 _1594_ (.Y(_0689_),
    .A(net579));
 sg13g2_inv_1 _1595_ (.Y(_0690_),
    .A(net708));
 sg13g2_inv_1 _1596_ (.Y(_0691_),
    .A(net323));
 sg13g2_inv_1 _1597_ (.Y(_0692_),
    .A(net815));
 sg13g2_inv_1 _1598_ (.Y(_0693_),
    .A(net374));
 sg13g2_inv_1 _1599_ (.Y(_0694_),
    .A(net396));
 sg13g2_inv_1 _1600_ (.Y(_0695_),
    .A(net618));
 sg13g2_inv_1 _1601_ (.Y(_0696_),
    .A(net693));
 sg13g2_inv_1 _1602_ (.Y(_0697_),
    .A(net734));
 sg13g2_inv_1 _1603_ (.Y(_0698_),
    .A(net790));
 sg13g2_inv_1 _1604_ (.Y(_0699_),
    .A(net798));
 sg13g2_inv_1 _1605_ (.Y(_0700_),
    .A(net717));
 sg13g2_inv_1 _1606_ (.Y(_0701_),
    .A(net349));
 sg13g2_inv_1 _1607_ (.Y(_0702_),
    .A(net722));
 sg13g2_inv_1 _1608_ (.Y(_0703_),
    .A(net639));
 sg13g2_inv_1 _1609_ (.Y(_0704_),
    .A(net325));
 sg13g2_inv_1 _1610_ (.Y(_0705_),
    .A(net418));
 sg13g2_inv_1 _1611_ (.Y(_0706_),
    .A(net780));
 sg13g2_inv_1 _1612_ (.Y(_0707_),
    .A(net795));
 sg13g2_inv_1 _1613_ (.Y(_0708_),
    .A(net822));
 sg13g2_inv_1 _1614_ (.Y(_0709_),
    .A(net800));
 sg13g2_inv_1 _1615_ (.Y(_0710_),
    .A(net626));
 sg13g2_inv_1 _1616_ (.Y(_0711_),
    .A(net591));
 sg13g2_inv_1 _1617_ (.Y(_0712_),
    .A(net772));
 sg13g2_inv_1 _1618_ (.Y(_0713_),
    .A(net760));
 sg13g2_inv_1 _1619_ (.Y(_0714_),
    .A(net745));
 sg13g2_inv_1 _1620_ (.Y(_0715_),
    .A(net353));
 sg13g2_inv_1 _1621_ (.Y(_0716_),
    .A(net775));
 sg13g2_inv_1 _1622_ (.Y(_0717_),
    .A(net432));
 sg13g2_inv_1 _1623_ (.Y(_0718_),
    .A(net698));
 sg13g2_inv_1 _1624_ (.Y(_0719_),
    .A(net783));
 sg13g2_inv_1 _1625_ (.Y(_0720_),
    .A(net341));
 sg13g2_inv_1 _1626_ (.Y(_0721_),
    .A(net840));
 sg13g2_inv_1 _1627_ (.Y(_0722_),
    .A(net682));
 sg13g2_inv_1 _1628_ (.Y(_0723_),
    .A(net779));
 sg13g2_inv_1 _1629_ (.Y(_0724_),
    .A(net412));
 sg13g2_inv_1 _1630_ (.Y(_0725_),
    .A(net660));
 sg13g2_inv_1 _1631_ (.Y(_0726_),
    .A(net316));
 sg13g2_inv_1 _1632_ (.Y(_0727_),
    .A(net753));
 sg13g2_inv_1 _1633_ (.Y(_0728_),
    .A(net658));
 sg13g2_inv_1 _1634_ (.Y(_0729_),
    .A(net724));
 sg13g2_inv_1 _1635_ (.Y(_0730_),
    .A(net629));
 sg13g2_inv_1 _1636_ (.Y(_0731_),
    .A(net604));
 sg13g2_inv_1 _1637_ (.Y(_0732_),
    .A(net630));
 sg13g2_inv_1 _1638_ (.Y(_0733_),
    .A(net665));
 sg13g2_inv_1 _1639_ (.Y(_0734_),
    .A(net645));
 sg13g2_inv_1 _1640_ (.Y(_0735_),
    .A(net362));
 sg13g2_inv_1 _1641_ (.Y(_0736_),
    .A(net754));
 sg13g2_inv_1 _1642_ (.Y(_0737_),
    .A(net376));
 sg13g2_inv_1 _1643_ (.Y(_0738_),
    .A(net606));
 sg13g2_inv_1 _1644_ (.Y(_0739_),
    .A(net718));
 sg13g2_inv_1 _1645_ (.Y(_0740_),
    .A(net810));
 sg13g2_inv_1 _1646_ (.Y(_0741_),
    .A(net825));
 sg13g2_inv_1 _1647_ (.Y(_0742_),
    .A(net778));
 sg13g2_inv_1 _1648_ (.Y(_0743_),
    .A(net669));
 sg13g2_inv_1 _1649_ (.Y(_0744_),
    .A(net337));
 sg13g2_inv_1 _1650_ (.Y(_0745_),
    .A(net388));
 sg13g2_inv_1 _1651_ (.Y(_0746_),
    .A(net641));
 sg13g2_inv_1 _1652_ (.Y(_0747_),
    .A(net821));
 sg13g2_inv_1 _1653_ (.Y(_0748_),
    .A(net424));
 sg13g2_inv_1 _1654_ (.Y(_0749_),
    .A(net357));
 sg13g2_inv_1 _1655_ (.Y(_0750_),
    .A(net662));
 sg13g2_inv_1 _1656_ (.Y(_0751_),
    .A(net430));
 sg13g2_inv_1 _1657_ (.Y(_0752_),
    .A(net829));
 sg13g2_inv_1 _1658_ (.Y(_0753_),
    .A(net598));
 sg13g2_inv_1 _1659_ (.Y(_0754_),
    .A(net713));
 sg13g2_inv_1 _1660_ (.Y(_0755_),
    .A(net703));
 sg13g2_inv_1 _1661_ (.Y(_0756_),
    .A(net382));
 sg13g2_inv_1 _1662_ (.Y(_0757_),
    .A(net427));
 sg13g2_inv_1 _1663_ (.Y(_0758_),
    .A(net743));
 sg13g2_inv_1 _1664_ (.Y(_0759_),
    .A(net700));
 sg13g2_inv_1 _1665_ (.Y(_0760_),
    .A(net589));
 sg13g2_inv_1 _1666_ (.Y(_0761_),
    .A(net697));
 sg13g2_inv_1 _1667_ (.Y(_0762_),
    .A(net402));
 sg13g2_inv_1 _1668_ (.Y(_0763_),
    .A(net812));
 sg13g2_inv_1 _1669_ (.Y(_0764_),
    .A(net690));
 sg13g2_inv_1 _1670_ (.Y(_0765_),
    .A(net370));
 sg13g2_inv_1 _1671_ (.Y(_0766_),
    .A(net830));
 sg13g2_inv_1 _1672_ (.Y(_0767_),
    .A(net751));
 sg13g2_inv_1 _1673_ (.Y(_0768_),
    .A(net691));
 sg13g2_inv_1 _1674_ (.Y(_0769_),
    .A(net321));
 sg13g2_inv_1 _1675_ (.Y(_0770_),
    .A(net804));
 sg13g2_inv_1 _1676_ (.Y(_0771_),
    .A(net726));
 sg13g2_inv_1 _1677_ (.Y(_0772_),
    .A(net360));
 sg13g2_inv_1 _1678_ (.Y(_0773_),
    .A(net831));
 sg13g2_inv_1 _1679_ (.Y(_0774_),
    .A(net803));
 sg13g2_inv_1 _1680_ (.Y(_0775_),
    .A(net688));
 sg13g2_inv_1 _1681_ (.Y(_0776_),
    .A(net686));
 sg13g2_inv_1 _1682_ (.Y(_0777_),
    .A(net702));
 sg13g2_inv_1 _1683_ (.Y(_0778_),
    .A(net632));
 sg13g2_inv_1 _1684_ (.Y(_0779_),
    .A(net318));
 sg13g2_inv_1 _1685_ (.Y(_0780_),
    .A(net797));
 sg13g2_inv_1 _1686_ (.Y(_0781_),
    .A(net610));
 sg13g2_inv_1 _1687_ (.Y(_0782_),
    .A(net593));
 sg13g2_inv_1 _1688_ (.Y(_0783_),
    .A(net809));
 sg13g2_inv_1 _1689_ (.Y(_0784_),
    .A(net759));
 sg13g2_inv_1 _1690_ (.Y(_0785_),
    .A(net740));
 sg13g2_inv_1 _1691_ (.Y(_0786_),
    .A(net387));
 sg13g2_inv_1 _1692_ (.Y(_0787_),
    .A(net331));
 sg13g2_inv_1 _1693_ (.Y(_0788_),
    .A(net595));
 sg13g2_inv_1 _1694_ (.Y(_0789_),
    .A(net637));
 sg13g2_inv_1 _1695_ (.Y(_0790_),
    .A(net742));
 sg13g2_inv_1 _1696_ (.Y(_0791_),
    .A(net327));
 sg13g2_inv_1 _1697_ (.Y(_0792_),
    .A(net738));
 sg13g2_inv_1 _1698_ (.Y(_0793_),
    .A(net390));
 sg13g2_inv_1 _1699_ (.Y(_0794_),
    .A(net770));
 sg13g2_inv_1 _1700_ (.Y(_0795_),
    .A(net615));
 sg13g2_inv_1 _1701_ (.Y(_0796_),
    .A(net650));
 sg13g2_inv_1 _1702_ (.Y(_0797_),
    .A(net767));
 sg13g2_inv_1 _1703_ (.Y(_0798_),
    .A(net621));
 sg13g2_inv_1 _1704_ (.Y(_0799_),
    .A(net643));
 sg13g2_inv_1 _1705_ (.Y(_0800_),
    .A(net784));
 sg13g2_inv_1 _1706_ (.Y(_0801_),
    .A(net748));
 sg13g2_inv_1 _1707_ (.Y(_0802_),
    .A(net819));
 sg13g2_inv_1 _1708_ (.Y(_0803_),
    .A(net723));
 sg13g2_inv_1 _1709_ (.Y(_0804_),
    .A(net343));
 sg13g2_inv_1 _1710_ (.Y(_0805_),
    .A(net672));
 sg13g2_inv_1 _1711_ (.Y(_0806_),
    .A(net372));
 sg13g2_inv_1 _1712_ (.Y(_0807_),
    .A(net799));
 sg13g2_inv_1 _1713_ (.Y(_0808_),
    .A(net617));
 sg13g2_inv_1 _1714_ (.Y(_0809_),
    .A(net410));
 sg13g2_inv_1 _1715_ (.Y(_0810_),
    .A(net613));
 sg13g2_inv_1 _1716_ (.Y(_0811_),
    .A(net827));
 sg13g2_inv_1 _1717_ (.Y(_0812_),
    .A(net750));
 sg13g2_inv_1 _1718_ (.Y(_0813_),
    .A(net581));
 sg13g2_inv_1 _1719_ (.Y(_0814_),
    .A(net828));
 sg13g2_inv_1 _1720_ (.Y(_0815_),
    .A(net705));
 sg13g2_inv_1 _1721_ (.Y(_0816_),
    .A(net585));
 sg13g2_inv_1 _1722_ (.Y(_0817_),
    .A(net802));
 sg13g2_inv_1 _1723_ (.Y(_0818_),
    .A(net667));
 sg13g2_inv_1 _1724_ (.Y(_0819_),
    .A(net736));
 sg13g2_inv_1 _1725_ (.Y(_0820_),
    .A(net398));
 sg13g2_inv_1 _1726_ (.Y(_0821_),
    .A(net652));
 sg13g2_inv_1 _1727_ (.Y(_0822_),
    .A(net774));
 sg13g2_inv_1 _1728_ (.Y(_0823_),
    .A(net739));
 sg13g2_inv_1 _1729_ (.Y(_0824_),
    .A(net648));
 sg13g2_inv_1 _1730_ (.Y(_0825_),
    .A(net744));
 sg13g2_inv_1 _1731_ (.Y(_0826_),
    .A(net597));
 sg13g2_inv_1 _1732_ (.Y(_0827_),
    .A(net429));
 sg13g2_inv_1 _1733_ (.Y(_0828_),
    .A(net404));
 sg13g2_inv_1 _1734_ (.Y(_0829_),
    .A(net634));
 sg13g2_inv_1 _1735_ (.Y(_0830_),
    .A(net792));
 sg13g2_inv_1 _1736_ (.Y(_0831_),
    .A(net678));
 sg13g2_inv_1 _1737_ (.Y(_0832_),
    .A(net528));
 sg13g2_inv_2 _1738_ (.Y(_0833_),
    .A(net487));
 sg13g2_inv_1 _1739_ (.Y(_0834_),
    .A(net574));
 sg13g2_inv_1 _1740_ (.Y(_0835_),
    .A(\bitserial_cipher.datapath.lut_ff56 ));
 sg13g2_inv_1 _1741_ (.Y(_0836_),
    .A(_0003_));
 sg13g2_nand2_1 _1742_ (.Y(_0837_),
    .A(\bitserial_cipher.datapath.round_counter[6] ),
    .B(net439));
 sg13g2_nor4_1 _1743_ (.A(\bitserial_cipher.datapath.round_counter[5] ),
    .B(\bitserial_cipher.datapath.round_counter[4] ),
    .C(\bitserial_cipher.datapath.round_counter[3] ),
    .D(\bitserial_cipher.datapath.round_counter[1] ),
    .Y(_0838_));
 sg13g2_nor2b_1 _1744_ (.A(_0837_),
    .B_N(_0838_),
    .Y(\bitserial_cipher.datapath.valid ));
 sg13g2_o21ai_1 _1745_ (.B1(net540),
    .Y(_0839_),
    .A1(\bitserial_cipher.key_exp.shifter2[37] ),
    .A2(net462));
 sg13g2_a21oi_1 _1746_ (.A1(_0831_),
    .A2(net462),
    .Y(_0006_),
    .B1(_0839_));
 sg13g2_o21ai_1 _1747_ (.B1(net540),
    .Y(_0840_),
    .A1(net678),
    .A2(net458));
 sg13g2_a21oi_1 _1748_ (.A1(_0830_),
    .A2(net457),
    .Y(_0007_),
    .B1(_0840_));
 sg13g2_o21ai_1 _1749_ (.B1(net539),
    .Y(_0841_),
    .A1(\bitserial_cipher.key_exp.shifter2[39] ),
    .A2(net457));
 sg13g2_a21oi_1 _1750_ (.A1(_0829_),
    .A2(net457),
    .Y(_0008_),
    .B1(_0841_));
 sg13g2_o21ai_1 _1751_ (.B1(net539),
    .Y(_0842_),
    .A1(\bitserial_cipher.key_exp.shifter2[40] ),
    .A2(net457));
 sg13g2_a21oi_1 _1752_ (.A1(_0828_),
    .A2(net451),
    .Y(_0009_),
    .B1(_0842_));
 sg13g2_o21ai_1 _1753_ (.B1(net535),
    .Y(_0843_),
    .A1(net404),
    .A2(net452));
 sg13g2_a21oi_1 _1754_ (.A1(_0827_),
    .A2(net451),
    .Y(_0010_),
    .B1(_0843_));
 sg13g2_o21ai_1 _1755_ (.B1(net535),
    .Y(_0844_),
    .A1(net429),
    .A2(net451));
 sg13g2_a21oi_1 _1756_ (.A1(_0826_),
    .A2(net451),
    .Y(_0011_),
    .B1(_0844_));
 sg13g2_o21ai_1 _1757_ (.B1(net535),
    .Y(_0845_),
    .A1(net597),
    .A2(net447));
 sg13g2_a21oi_1 _1758_ (.A1(_0825_),
    .A2(net447),
    .Y(_0012_),
    .B1(_0845_));
 sg13g2_o21ai_1 _1759_ (.B1(net535),
    .Y(_0846_),
    .A1(\bitserial_cipher.key_exp.shifter2[44] ),
    .A2(net450));
 sg13g2_a21oi_1 _1760_ (.A1(_0824_),
    .A2(net447),
    .Y(_0013_),
    .B1(_0846_));
 sg13g2_o21ai_1 _1761_ (.B1(net534),
    .Y(_0847_),
    .A1(net648),
    .A2(net446));
 sg13g2_a21oi_1 _1762_ (.A1(_0823_),
    .A2(net448),
    .Y(_0014_),
    .B1(_0847_));
 sg13g2_o21ai_1 _1763_ (.B1(net536),
    .Y(_0848_),
    .A1(net739),
    .A2(net448));
 sg13g2_a21oi_1 _1764_ (.A1(_0822_),
    .A2(net448),
    .Y(_0015_),
    .B1(_0848_));
 sg13g2_o21ai_1 _1765_ (.B1(net536),
    .Y(_0849_),
    .A1(\bitserial_cipher.key_exp.shifter2[47] ),
    .A2(net448));
 sg13g2_a21oi_1 _1766_ (.A1(_0821_),
    .A2(net448),
    .Y(_0016_),
    .B1(_0849_));
 sg13g2_o21ai_1 _1767_ (.B1(net534),
    .Y(_0850_),
    .A1(\bitserial_cipher.key_exp.shifter2[48] ),
    .A2(net448));
 sg13g2_a21oi_1 _1768_ (.A1(_0820_),
    .A2(net448),
    .Y(_0017_),
    .B1(_0850_));
 sg13g2_o21ai_1 _1769_ (.B1(net537),
    .Y(_0851_),
    .A1(net398),
    .A2(net449));
 sg13g2_a21oi_1 _1770_ (.A1(_0819_),
    .A2(net448),
    .Y(_0018_),
    .B1(_0851_));
 sg13g2_o21ai_1 _1771_ (.B1(net538),
    .Y(_0852_),
    .A1(\bitserial_cipher.key_exp.shifter2[50] ),
    .A2(net449));
 sg13g2_a21oi_1 _1772_ (.A1(_0818_),
    .A2(net449),
    .Y(_0019_),
    .B1(_0852_));
 sg13g2_o21ai_1 _1773_ (.B1(net538),
    .Y(_0853_),
    .A1(net667),
    .A2(net453));
 sg13g2_a21oi_1 _1774_ (.A1(_0817_),
    .A2(net453),
    .Y(_0020_),
    .B1(_0853_));
 sg13g2_o21ai_1 _1775_ (.B1(net543),
    .Y(_0854_),
    .A1(\bitserial_cipher.key_exp.shifter2[52] ),
    .A2(net455));
 sg13g2_a21oi_1 _1776_ (.A1(_0816_),
    .A2(net455),
    .Y(_0021_),
    .B1(_0854_));
 sg13g2_o21ai_1 _1777_ (.B1(net543),
    .Y(_0855_),
    .A1(net585),
    .A2(net466));
 sg13g2_a21oi_1 _1778_ (.A1(_0815_),
    .A2(net466),
    .Y(_0022_),
    .B1(_0855_));
 sg13g2_o21ai_1 _1779_ (.B1(net543),
    .Y(_0856_),
    .A1(net705),
    .A2(net466));
 sg13g2_a21oi_1 _1780_ (.A1(_0814_),
    .A2(net467),
    .Y(_0023_),
    .B1(_0856_));
 sg13g2_o21ai_1 _1781_ (.B1(net543),
    .Y(_0857_),
    .A1(\bitserial_cipher.key_exp.shifter2[55] ),
    .A2(net467));
 sg13g2_a21oi_1 _1782_ (.A1(_0813_),
    .A2(net467),
    .Y(_0024_),
    .B1(_0857_));
 sg13g2_o21ai_1 _1783_ (.B1(net544),
    .Y(_0858_),
    .A1(net581),
    .A2(net468));
 sg13g2_a21oi_1 _1784_ (.A1(_0812_),
    .A2(net468),
    .Y(_0025_),
    .B1(_0858_));
 sg13g2_o21ai_1 _1785_ (.B1(net542),
    .Y(_0859_),
    .A1(net750),
    .A2(net468));
 sg13g2_a21oi_1 _1786_ (.A1(_0811_),
    .A2(net469),
    .Y(_0026_),
    .B1(_0859_));
 sg13g2_o21ai_1 _1787_ (.B1(net562),
    .Y(_0860_),
    .A1(\bitserial_cipher.key_exp.shifter2[58] ),
    .A2(net475));
 sg13g2_a21oi_1 _1788_ (.A1(_0810_),
    .A2(net475),
    .Y(_0027_),
    .B1(_0860_));
 sg13g2_o21ai_1 _1789_ (.B1(net569),
    .Y(_0861_),
    .A1(\bitserial_cipher.key_exp.shifter2[59] ),
    .A2(net475));
 sg13g2_a21oi_1 _1790_ (.A1(_0809_),
    .A2(net475),
    .Y(_0028_),
    .B1(_0861_));
 sg13g2_o21ai_1 _1791_ (.B1(net562),
    .Y(_0862_),
    .A1(net410),
    .A2(net475));
 sg13g2_a21oi_1 _1792_ (.A1(_0808_),
    .A2(net471),
    .Y(_0029_),
    .B1(_0862_));
 sg13g2_o21ai_1 _1793_ (.B1(net562),
    .Y(_0863_),
    .A1(net617),
    .A2(net476));
 sg13g2_a21oi_1 _1794_ (.A1(_0807_),
    .A2(net476),
    .Y(_0030_),
    .B1(_0863_));
 sg13g2_o21ai_1 _1795_ (.B1(net562),
    .Y(_0864_),
    .A1(\bitserial_cipher.key_exp.shifter2[62] ),
    .A2(net475));
 sg13g2_a21oi_1 _1796_ (.A1(_0806_),
    .A2(net476),
    .Y(_0031_),
    .B1(_0864_));
 sg13g2_nor3_2 _1797_ (.A(\bitserial_cipher.bit_counter[5] ),
    .B(\bitserial_cipher.bit_counter[4] ),
    .C(\bitserial_cipher.bit_counter[3] ),
    .Y(_0865_));
 sg13g2_nor2b_2 _1798_ (.A(net820),
    .B_N(_0865_),
    .Y(_0866_));
 sg13g2_nor2_2 _1799_ (.A(\bitserial_cipher.datapath.round_counter[3] ),
    .B(\bitserial_cipher.datapath.round_counter[2] ),
    .Y(_0867_));
 sg13g2_or4_2 _1800_ (.A(\bitserial_cipher.datapath.round_counter[5] ),
    .B(\bitserial_cipher.datapath.round_counter[4] ),
    .C(\bitserial_cipher.datapath.round_counter[3] ),
    .D(net439),
    .X(_0868_));
 sg13g2_or2_1 _1801_ (.X(_0869_),
    .B(net441),
    .A(net440));
 sg13g2_or3_1 _1802_ (.A(\bitserial_cipher.datapath.round_counter[6] ),
    .B(_0868_),
    .C(_0869_),
    .X(_0870_));
 sg13g2_nand2_1 _1803_ (.Y(_0871_),
    .A(_0866_),
    .B(_0870_));
 sg13g2_a21oi_1 _1804_ (.A1(net444),
    .A2(net487),
    .Y(_0872_),
    .B1(_0871_));
 sg13g2_o21ai_1 _1805_ (.B1(net486),
    .Y(_0873_),
    .A1(\bitserial_cipher.key_exp.fifo_ff0 ),
    .A2(_0872_));
 sg13g2_a21oi_1 _1806_ (.A1(_0620_),
    .A2(_0872_),
    .Y(_0874_),
    .B1(_0873_));
 sg13g2_a21oi_1 _1807_ (.A1(net372),
    .A2(_0833_),
    .Y(_0875_),
    .B1(net839));
 sg13g2_nor2_1 _1808_ (.A(net443),
    .B(_0875_),
    .Y(_0032_));
 sg13g2_o21ai_1 _1809_ (.B1(net568),
    .Y(_0876_),
    .A1(\bitserial_cipher.key_exp.shift_out1 ),
    .A2(net488));
 sg13g2_a21oi_1 _1810_ (.A1(_0805_),
    .A2(net488),
    .Y(_0033_),
    .B1(_0876_));
 sg13g2_o21ai_1 _1811_ (.B1(net568),
    .Y(_0877_),
    .A1(\bitserial_cipher.key_exp.shifter1[1] ),
    .A2(net483));
 sg13g2_a21oi_1 _1812_ (.A1(_0804_),
    .A2(net484),
    .Y(_0034_),
    .B1(_0877_));
 sg13g2_o21ai_1 _1813_ (.B1(net568),
    .Y(_0878_),
    .A1(net343),
    .A2(net483));
 sg13g2_a21oi_1 _1814_ (.A1(_0803_),
    .A2(net483),
    .Y(_0035_),
    .B1(_0878_));
 sg13g2_o21ai_1 _1815_ (.B1(net565),
    .Y(_0879_),
    .A1(net723),
    .A2(net484));
 sg13g2_a21oi_1 _1816_ (.A1(_0802_),
    .A2(net484),
    .Y(_0036_),
    .B1(_0879_));
 sg13g2_o21ai_1 _1817_ (.B1(net565),
    .Y(_0880_),
    .A1(\bitserial_cipher.key_exp.shifter1[4] ),
    .A2(net484));
 sg13g2_a21oi_1 _1818_ (.A1(_0801_),
    .A2(net484),
    .Y(_0037_),
    .B1(_0880_));
 sg13g2_o21ai_1 _1819_ (.B1(net566),
    .Y(_0881_),
    .A1(net748),
    .A2(net479));
 sg13g2_a21oi_1 _1820_ (.A1(_0800_),
    .A2(net479),
    .Y(_0038_),
    .B1(_0881_));
 sg13g2_o21ai_1 _1821_ (.B1(net566),
    .Y(_0882_),
    .A1(\bitserial_cipher.key_exp.shifter1[6] ),
    .A2(net479));
 sg13g2_a21oi_1 _1822_ (.A1(_0799_),
    .A2(net479),
    .Y(_0039_),
    .B1(_0882_));
 sg13g2_o21ai_1 _1823_ (.B1(net563),
    .Y(_0883_),
    .A1(\bitserial_cipher.key_exp.shifter1[7] ),
    .A2(net479));
 sg13g2_a21oi_1 _1824_ (.A1(_0798_),
    .A2(net479),
    .Y(_0040_),
    .B1(_0883_));
 sg13g2_o21ai_1 _1825_ (.B1(net561),
    .Y(_0884_),
    .A1(net621),
    .A2(net473));
 sg13g2_a21oi_1 _1826_ (.A1(_0797_),
    .A2(net473),
    .Y(_0041_),
    .B1(_0884_));
 sg13g2_o21ai_1 _1827_ (.B1(net561),
    .Y(_0885_),
    .A1(\bitserial_cipher.key_exp.shifter1[9] ),
    .A2(net473));
 sg13g2_a21oi_1 _1828_ (.A1(_0796_),
    .A2(net473),
    .Y(_0042_),
    .B1(_0885_));
 sg13g2_o21ai_1 _1829_ (.B1(net561),
    .Y(_0886_),
    .A1(\bitserial_cipher.key_exp.shifter1[10] ),
    .A2(net473));
 sg13g2_a21oi_1 _1830_ (.A1(_0795_),
    .A2(net473),
    .Y(_0043_),
    .B1(_0886_));
 sg13g2_o21ai_1 _1831_ (.B1(net560),
    .Y(_0887_),
    .A1(net615),
    .A2(net471));
 sg13g2_a21oi_1 _1832_ (.A1(_0794_),
    .A2(net471),
    .Y(_0044_),
    .B1(_0887_));
 sg13g2_o21ai_1 _1833_ (.B1(net560),
    .Y(_0888_),
    .A1(\bitserial_cipher.key_exp.shifter1[12] ),
    .A2(net471));
 sg13g2_a21oi_1 _1834_ (.A1(_0793_),
    .A2(net471),
    .Y(_0045_),
    .B1(_0888_));
 sg13g2_o21ai_1 _1835_ (.B1(net561),
    .Y(_0889_),
    .A1(net390),
    .A2(net471));
 sg13g2_a21oi_1 _1836_ (.A1(_0792_),
    .A2(net471),
    .Y(_0046_),
    .B1(_0889_));
 sg13g2_o21ai_1 _1837_ (.B1(net569),
    .Y(_0890_),
    .A1(\bitserial_cipher.key_exp.shifter1[14] ),
    .A2(net463));
 sg13g2_a21oi_1 _1838_ (.A1(_0791_),
    .A2(net464),
    .Y(_0047_),
    .B1(_0890_));
 sg13g2_o21ai_1 _1839_ (.B1(net542),
    .Y(_0891_),
    .A1(net327),
    .A2(net464));
 sg13g2_a21oi_1 _1840_ (.A1(_0790_),
    .A2(net464),
    .Y(_0048_),
    .B1(_0891_));
 sg13g2_o21ai_1 _1841_ (.B1(net542),
    .Y(_0892_),
    .A1(\bitserial_cipher.key_exp.shifter1[16] ),
    .A2(net463));
 sg13g2_a21oi_1 _1842_ (.A1(_0789_),
    .A2(net463),
    .Y(_0049_),
    .B1(_0892_));
 sg13g2_o21ai_1 _1843_ (.B1(net542),
    .Y(_0893_),
    .A1(\bitserial_cipher.key_exp.shifter1[17] ),
    .A2(net459));
 sg13g2_a21oi_1 _1844_ (.A1(_0788_),
    .A2(net459),
    .Y(_0050_),
    .B1(_0893_));
 sg13g2_o21ai_1 _1845_ (.B1(net542),
    .Y(_0894_),
    .A1(\bitserial_cipher.key_exp.shifter1[18] ),
    .A2(net459));
 sg13g2_a21oi_1 _1846_ (.A1(_0787_),
    .A2(net459),
    .Y(_0051_),
    .B1(_0894_));
 sg13g2_o21ai_1 _1847_ (.B1(net539),
    .Y(_0895_),
    .A1(net331),
    .A2(net459));
 sg13g2_a21oi_1 _1848_ (.A1(_0786_),
    .A2(net459),
    .Y(_0052_),
    .B1(_0895_));
 sg13g2_o21ai_1 _1849_ (.B1(net541),
    .Y(_0896_),
    .A1(net387),
    .A2(net459));
 sg13g2_a21oi_1 _1850_ (.A1(_0785_),
    .A2(net463),
    .Y(_0053_),
    .B1(_0896_));
 sg13g2_o21ai_1 _1851_ (.B1(net541),
    .Y(_0897_),
    .A1(net740),
    .A2(net463));
 sg13g2_a21oi_1 _1852_ (.A1(_0784_),
    .A2(net463),
    .Y(_0054_),
    .B1(_0897_));
 sg13g2_o21ai_1 _1853_ (.B1(net560),
    .Y(_0898_),
    .A1(net759),
    .A2(net464));
 sg13g2_a21oi_1 _1854_ (.A1(_0783_),
    .A2(net464),
    .Y(_0055_),
    .B1(_0898_));
 sg13g2_o21ai_1 _1855_ (.B1(net560),
    .Y(_0899_),
    .A1(\bitserial_cipher.key_exp.shifter1[23] ),
    .A2(net470));
 sg13g2_a21oi_1 _1856_ (.A1(_0782_),
    .A2(net470),
    .Y(_0056_),
    .B1(_0899_));
 sg13g2_o21ai_1 _1857_ (.B1(net562),
    .Y(_0900_),
    .A1(net593),
    .A2(net470));
 sg13g2_a21oi_1 _1858_ (.A1(_0781_),
    .A2(net472),
    .Y(_0057_),
    .B1(_0900_));
 sg13g2_o21ai_1 _1859_ (.B1(net562),
    .Y(_0901_),
    .A1(net610),
    .A2(net472));
 sg13g2_a21oi_1 _1860_ (.A1(_0780_),
    .A2(net472),
    .Y(_0058_),
    .B1(_0901_));
 sg13g2_o21ai_1 _1861_ (.B1(net563),
    .Y(_0902_),
    .A1(\bitserial_cipher.key_exp.shifter1[26] ),
    .A2(net477));
 sg13g2_a21oi_1 _1862_ (.A1(_0779_),
    .A2(net477),
    .Y(_0059_),
    .B1(_0902_));
 sg13g2_o21ai_1 _1863_ (.B1(net563),
    .Y(_0903_),
    .A1(net318),
    .A2(net478));
 sg13g2_a21oi_1 _1864_ (.A1(_0778_),
    .A2(net478),
    .Y(_0060_),
    .B1(_0903_));
 sg13g2_o21ai_1 _1865_ (.B1(net564),
    .Y(_0904_),
    .A1(net632),
    .A2(net482));
 sg13g2_a21oi_1 _1866_ (.A1(_0777_),
    .A2(net482),
    .Y(_0061_),
    .B1(_0904_));
 sg13g2_o21ai_1 _1867_ (.B1(net564),
    .Y(_0905_),
    .A1(\bitserial_cipher.key_exp.shifter1[29] ),
    .A2(net480));
 sg13g2_a21oi_1 _1868_ (.A1(_0776_),
    .A2(net480),
    .Y(_0062_),
    .B1(_0905_));
 sg13g2_o21ai_1 _1869_ (.B1(net564),
    .Y(_0906_),
    .A1(net686),
    .A2(net480));
 sg13g2_a21oi_1 _1870_ (.A1(_0775_),
    .A2(net480),
    .Y(_0063_),
    .B1(_0906_));
 sg13g2_o21ai_1 _1871_ (.B1(net564),
    .Y(_0907_),
    .A1(net688),
    .A2(net482));
 sg13g2_a21oi_1 _1872_ (.A1(_0774_),
    .A2(net482),
    .Y(_0064_),
    .B1(_0907_));
 sg13g2_o21ai_1 _1873_ (.B1(net563),
    .Y(_0908_),
    .A1(net803),
    .A2(net477));
 sg13g2_a21oi_1 _1874_ (.A1(_0773_),
    .A2(net477),
    .Y(_0065_),
    .B1(_0908_));
 sg13g2_o21ai_1 _1875_ (.B1(net563),
    .Y(_0909_),
    .A1(\bitserial_cipher.key_exp.shifter1[33] ),
    .A2(net477));
 sg13g2_a21oi_1 _1876_ (.A1(_0772_),
    .A2(net477),
    .Y(_0066_),
    .B1(_0909_));
 sg13g2_o21ai_1 _1877_ (.B1(net561),
    .Y(_0910_),
    .A1(net360),
    .A2(net472));
 sg13g2_a21oi_1 _1878_ (.A1(_0771_),
    .A2(net472),
    .Y(_0067_),
    .B1(_0910_));
 sg13g2_o21ai_1 _1879_ (.B1(net561),
    .Y(_0911_),
    .A1(net726),
    .A2(net472));
 sg13g2_a21oi_1 _1880_ (.A1(_0770_),
    .A2(net470),
    .Y(_0068_),
    .B1(_0911_));
 sg13g2_o21ai_1 _1881_ (.B1(net560),
    .Y(_0912_),
    .A1(\bitserial_cipher.key_exp.shifter1[36] ),
    .A2(net470));
 sg13g2_a21oi_1 _1882_ (.A1(_0769_),
    .A2(net470),
    .Y(_0069_),
    .B1(_0912_));
 sg13g2_o21ai_1 _1883_ (.B1(net560),
    .Y(_0913_),
    .A1(net321),
    .A2(net465));
 sg13g2_a21oi_1 _1884_ (.A1(_0768_),
    .A2(net465),
    .Y(_0070_),
    .B1(_0913_));
 sg13g2_o21ai_1 _1885_ (.B1(net541),
    .Y(_0914_),
    .A1(net691),
    .A2(net463));
 sg13g2_a21oi_1 _1886_ (.A1(_0767_),
    .A2(net463),
    .Y(_0071_),
    .B1(_0914_));
 sg13g2_o21ai_1 _1887_ (.B1(net541),
    .Y(_0915_),
    .A1(net751),
    .A2(net460));
 sg13g2_a21oi_1 _1888_ (.A1(_0766_),
    .A2(net459),
    .Y(_0072_),
    .B1(_0915_));
 sg13g2_o21ai_1 _1889_ (.B1(net539),
    .Y(_0916_),
    .A1(\bitserial_cipher.key_exp.shifter1[40] ),
    .A2(net453));
 sg13g2_a21oi_1 _1890_ (.A1(_0765_),
    .A2(net453),
    .Y(_0073_),
    .B1(_0916_));
 sg13g2_o21ai_1 _1891_ (.B1(net536),
    .Y(_0917_),
    .A1(net370),
    .A2(net453));
 sg13g2_a21oi_1 _1892_ (.A1(_0764_),
    .A2(net453),
    .Y(_0074_),
    .B1(_0917_));
 sg13g2_o21ai_1 _1893_ (.B1(net538),
    .Y(_0918_),
    .A1(net690),
    .A2(net449));
 sg13g2_a21oi_1 _1894_ (.A1(_0763_),
    .A2(net449),
    .Y(_0075_),
    .B1(_0918_));
 sg13g2_o21ai_1 _1895_ (.B1(net537),
    .Y(_0919_),
    .A1(\bitserial_cipher.key_exp.shifter1[43] ),
    .A2(net449));
 sg13g2_a21oi_1 _1896_ (.A1(_0762_),
    .A2(net449),
    .Y(_0076_),
    .B1(_0919_));
 sg13g2_o21ai_1 _1897_ (.B1(net537),
    .Y(_0920_),
    .A1(net402),
    .A2(net454));
 sg13g2_a21oi_1 _1898_ (.A1(_0761_),
    .A2(net454),
    .Y(_0077_),
    .B1(_0920_));
 sg13g2_o21ai_1 _1899_ (.B1(net537),
    .Y(_0921_),
    .A1(\bitserial_cipher.key_exp.shifter1[45] ),
    .A2(net454));
 sg13g2_a21oi_1 _1900_ (.A1(_0760_),
    .A2(net454),
    .Y(_0078_),
    .B1(_0921_));
 sg13g2_o21ai_1 _1901_ (.B1(net537),
    .Y(_0922_),
    .A1(net589),
    .A2(net454));
 sg13g2_a21oi_1 _1902_ (.A1(_0759_),
    .A2(net454),
    .Y(_0079_),
    .B1(_0922_));
 sg13g2_o21ai_1 _1903_ (.B1(net537),
    .Y(_0923_),
    .A1(net700),
    .A2(net454));
 sg13g2_a21oi_1 _1904_ (.A1(_0758_),
    .A2(net454),
    .Y(_0080_),
    .B1(_0923_));
 sg13g2_o21ai_1 _1905_ (.B1(net537),
    .Y(_0924_),
    .A1(\bitserial_cipher.key_exp.shifter1[48] ),
    .A2(net455));
 sg13g2_a21oi_1 _1906_ (.A1(_0757_),
    .A2(net455),
    .Y(_0081_),
    .B1(_0924_));
 sg13g2_o21ai_1 _1907_ (.B1(net538),
    .Y(_0287_),
    .A1(\bitserial_cipher.key_exp.shifter1[49] ),
    .A2(net456));
 sg13g2_a21oi_1 _1908_ (.A1(_0756_),
    .A2(net455),
    .Y(_0082_),
    .B1(_0287_));
 sg13g2_o21ai_1 _1909_ (.B1(net537),
    .Y(_0288_),
    .A1(net382),
    .A2(net456));
 sg13g2_a21oi_1 _1910_ (.A1(_0755_),
    .A2(net456),
    .Y(_0083_),
    .B1(_0288_));
 sg13g2_o21ai_1 _1911_ (.B1(net543),
    .Y(_0289_),
    .A1(net703),
    .A2(net455));
 sg13g2_a21oi_1 _1912_ (.A1(_0754_),
    .A2(net455),
    .Y(_0084_),
    .B1(_0289_));
 sg13g2_o21ai_1 _1913_ (.B1(net543),
    .Y(_0290_),
    .A1(\bitserial_cipher.key_exp.shifter1[52] ),
    .A2(net466));
 sg13g2_a21oi_1 _1914_ (.A1(_0753_),
    .A2(net466),
    .Y(_0085_),
    .B1(_0290_));
 sg13g2_o21ai_1 _1915_ (.B1(net543),
    .Y(_0291_),
    .A1(net598),
    .A2(net466));
 sg13g2_a21oi_1 _1916_ (.A1(_0752_),
    .A2(net466),
    .Y(_0086_),
    .B1(_0291_));
 sg13g2_o21ai_1 _1917_ (.B1(net542),
    .Y(_0292_),
    .A1(\bitserial_cipher.key_exp.shifter1[54] ),
    .A2(net466));
 sg13g2_a21oi_1 _1918_ (.A1(_0751_),
    .A2(net468),
    .Y(_0087_),
    .B1(_0292_));
 sg13g2_o21ai_1 _1919_ (.B1(net542),
    .Y(_0293_),
    .A1(net430),
    .A2(net468));
 sg13g2_a21oi_1 _1920_ (.A1(_0750_),
    .A2(net468),
    .Y(_0088_),
    .B1(_0293_));
 sg13g2_o21ai_1 _1921_ (.B1(net542),
    .Y(_0294_),
    .A1(\bitserial_cipher.key_exp.shifter1[56] ),
    .A2(net468));
 sg13g2_a21oi_1 _1922_ (.A1(_0749_),
    .A2(net468),
    .Y(_0089_),
    .B1(_0294_));
 sg13g2_o21ai_1 _1923_ (.B1(net562),
    .Y(_0295_),
    .A1(net357),
    .A2(net475));
 sg13g2_a21oi_1 _1924_ (.A1(_0748_),
    .A2(net475),
    .Y(_0090_),
    .B1(_0295_));
 sg13g2_o21ai_1 _1925_ (.B1(net573),
    .Y(_0296_),
    .A1(net424),
    .A2(net476));
 sg13g2_a21oi_1 _1926_ (.A1(_0747_),
    .A2(net476),
    .Y(_0091_),
    .B1(_0296_));
 sg13g2_nor2_2 _1927_ (.A(net444),
    .B(_0833_),
    .Y(_0297_));
 sg13g2_and2_2 _1928_ (.A(_0866_),
    .B(_0297_),
    .X(_0298_));
 sg13g2_nand2_1 _1929_ (.Y(_0299_),
    .A(_0866_),
    .B(_0297_));
 sg13g2_nor3_1 _1930_ (.A(_0836_),
    .B(_0868_),
    .C(_0869_),
    .Y(_0300_));
 sg13g2_nor2_1 _1931_ (.A(_0299_),
    .B(_0300_),
    .Y(_0301_));
 sg13g2_nor2b_1 _1932_ (.A(\bitserial_cipher.bit_counter[1] ),
    .B_N(_0866_),
    .Y(_0302_));
 sg13g2_xnor2_1 _1933_ (.Y(_0303_),
    .A(_0836_),
    .B(_0868_));
 sg13g2_nand2_1 _1934_ (.Y(_0304_),
    .A(\bitserial_cipher.datapath.round_counter[6] ),
    .B(_0868_));
 sg13g2_a21oi_1 _1935_ (.A1(\bitserial_cipher.datapath.round_counter[6] ),
    .A2(_0868_),
    .Y(_0305_),
    .B1(_0000_));
 sg13g2_nor2_1 _1936_ (.A(\bitserial_cipher.datapath.round_counter[1] ),
    .B(_0305_),
    .Y(_0306_));
 sg13g2_a21oi_1 _1937_ (.A1(\bitserial_cipher.datapath.round_counter[6] ),
    .A2(_0868_),
    .Y(_0307_),
    .B1(net441));
 sg13g2_o21ai_1 _1938_ (.B1(net439),
    .Y(_0308_),
    .A1(_0621_),
    .A2(_0307_));
 sg13g2_nand2_1 _1939_ (.Y(_0309_),
    .A(\bitserial_cipher.datapath.round_counter[3] ),
    .B(net439));
 sg13g2_nor2b_1 _1940_ (.A(_0867_),
    .B_N(_0309_),
    .Y(_0310_));
 sg13g2_nand2b_1 _1941_ (.Y(_0311_),
    .B(_0309_),
    .A_N(_0867_));
 sg13g2_or2_1 _1942_ (.X(_0312_),
    .B(net440),
    .A(net439));
 sg13g2_a21oi_1 _1943_ (.A1(\bitserial_cipher.datapath.round_counter[6] ),
    .A2(_0868_),
    .Y(_0313_),
    .B1(_0312_));
 sg13g2_nor2_1 _1944_ (.A(_0311_),
    .B(_0313_),
    .Y(_0314_));
 sg13g2_o21ai_1 _1945_ (.B1(_0314_),
    .Y(_0315_),
    .A1(_0306_),
    .A2(_0308_));
 sg13g2_nand2_1 _1946_ (.Y(_0316_),
    .A(_0002_),
    .B(_0867_));
 sg13g2_xor2_1 _1947_ (.B(_0867_),
    .A(_0002_),
    .X(_0317_));
 sg13g2_xnor2_1 _1948_ (.Y(_0318_),
    .A(_0002_),
    .B(_0867_));
 sg13g2_nor2_1 _1949_ (.A(_0307_),
    .B(_0310_),
    .Y(_0319_));
 sg13g2_nand2_1 _1950_ (.Y(_0320_),
    .A(net439),
    .B(net440));
 sg13g2_nand3_1 _1951_ (.B(_0312_),
    .C(_0320_),
    .A(_0304_),
    .Y(_0321_));
 sg13g2_a21oi_1 _1952_ (.A1(_0319_),
    .A2(_0321_),
    .Y(_0322_),
    .B1(_0317_));
 sg13g2_o21ai_1 _1953_ (.B1(_0869_),
    .Y(_0323_),
    .A1(_0621_),
    .A2(_0000_));
 sg13g2_a21oi_1 _1954_ (.A1(_0304_),
    .A2(_0323_),
    .Y(_0324_),
    .B1(net439));
 sg13g2_nand2_1 _1955_ (.Y(_0325_),
    .A(_0837_),
    .B(_0311_));
 sg13g2_nand3b_1 _1956_ (.B(_0305_),
    .C(_0310_),
    .Y(_0326_),
    .A_N(_0004_));
 sg13g2_o21ai_1 _1957_ (.B1(_0326_),
    .Y(_0327_),
    .A1(_0324_),
    .A2(_0325_));
 sg13g2_xor2_1 _1958_ (.B(_0316_),
    .A(\bitserial_cipher.datapath.round_counter[5] ),
    .X(_0328_));
 sg13g2_inv_1 _1959_ (.Y(_0329_),
    .A(_0328_));
 sg13g2_a221oi_1 _1960_ (.B2(_0317_),
    .C1(_0328_),
    .B1(_0327_),
    .A1(_0315_),
    .Y(_0330_),
    .A2(_0322_));
 sg13g2_nor2_1 _1961_ (.A(\bitserial_cipher.datapath.round_counter[3] ),
    .B(_0305_),
    .Y(_0331_));
 sg13g2_o21ai_1 _1962_ (.B1(_0310_),
    .Y(_0332_),
    .A1(_0324_),
    .A2(_0331_));
 sg13g2_nor2b_1 _1963_ (.A(_0319_),
    .B_N(_0320_),
    .Y(_0333_));
 sg13g2_nand3_1 _1964_ (.B(_0332_),
    .C(_0333_),
    .A(_0318_),
    .Y(_0334_));
 sg13g2_o21ai_1 _1965_ (.B1(_0311_),
    .Y(_0335_),
    .A1(_0002_),
    .A2(_0004_));
 sg13g2_o21ai_1 _1966_ (.B1(_0304_),
    .Y(_0336_),
    .A1(_0002_),
    .A2(_0867_));
 sg13g2_a21oi_1 _1967_ (.A1(\bitserial_cipher.datapath.round_counter[3] ),
    .A2(_0306_),
    .Y(_0337_),
    .B1(_0336_));
 sg13g2_a21oi_1 _1968_ (.A1(_0335_),
    .A2(_0337_),
    .Y(_0338_),
    .B1(_0329_));
 sg13g2_a21oi_1 _1969_ (.A1(_0334_),
    .A2(_0338_),
    .Y(_0339_),
    .B1(_0330_));
 sg13g2_nor2b_1 _1970_ (.A(\bitserial_cipher.bit_counter[0] ),
    .B_N(_0302_),
    .Y(_0340_));
 sg13g2_nand4_1 _1971_ (.B(_0307_),
    .C(_0311_),
    .A(_0001_),
    .Y(_0341_),
    .D(_0318_));
 sg13g2_o21ai_1 _1972_ (.B1(_0303_),
    .Y(_0342_),
    .A1(_0328_),
    .A2(_0341_));
 sg13g2_and2_1 _1973_ (.A(_0340_),
    .B(_0342_),
    .X(_0343_));
 sg13g2_o21ai_1 _1974_ (.B1(_0343_),
    .Y(_0344_),
    .A1(_0303_),
    .A2(_0339_));
 sg13g2_nand2_1 _1975_ (.Y(_0345_),
    .A(_0870_),
    .B(_0340_));
 sg13g2_mux2_1 _1976_ (.A0(\bitserial_cipher.key_exp.lut_ff3 ),
    .A1(\bitserial_cipher.key_exp.fifo_ff3 ),
    .S(_0345_),
    .X(_0346_));
 sg13g2_xnor2_1 _1977_ (.Y(_0347_),
    .A(\bitserial_cipher.datapath.key_in ),
    .B(\bitserial_cipher.key_exp.shift_out1 ));
 sg13g2_xnor2_1 _1978_ (.Y(_0348_),
    .A(_0346_),
    .B(_0347_));
 sg13g2_xnor2_1 _1979_ (.Y(_0349_),
    .A(_0344_),
    .B(_0348_));
 sg13g2_xnor2_1 _1980_ (.Y(_0350_),
    .A(_0302_),
    .B(_0349_));
 sg13g2_nor2_1 _1981_ (.A(_0870_),
    .B(_0299_),
    .Y(_0351_));
 sg13g2_a221oi_1 _1982_ (.B2(_0620_),
    .C1(_0351_),
    .B1(_0301_),
    .A1(net444),
    .Y(_0352_),
    .A2(net487));
 sg13g2_o21ai_1 _1983_ (.B1(_0352_),
    .Y(_0353_),
    .A1(_0301_),
    .A2(_0350_));
 sg13g2_a21oi_1 _1984_ (.A1(net853),
    .A2(_0351_),
    .Y(_0354_),
    .B1(_0833_));
 sg13g2_a221oi_1 _1985_ (.B2(_0354_),
    .C1(net443),
    .B1(_0353_),
    .A1(_0747_),
    .Y(_0092_),
    .A2(_0833_));
 sg13g2_o21ai_1 _1986_ (.B1(net575),
    .Y(_0355_),
    .A1(\bitserial_cipher.datapath.fifo_ff57 ),
    .A2(net529));
 sg13g2_a21oi_1 _1987_ (.A1(_0746_),
    .A2(net529),
    .Y(_0093_),
    .B1(_0355_));
 sg13g2_o21ai_1 _1988_ (.B1(net576),
    .Y(_0356_),
    .A1(\bitserial_cipher.datapath.fifo_ff58 ),
    .A2(net531));
 sg13g2_a21oi_1 _1989_ (.A1(_0745_),
    .A2(net531),
    .Y(_0094_),
    .B1(_0356_));
 sg13g2_o21ai_1 _1990_ (.B1(net576),
    .Y(_0357_),
    .A1(\bitserial_cipher.datapath.fifo_ff59 ),
    .A2(net531));
 sg13g2_a21oi_1 _1991_ (.A1(_0744_),
    .A2(net529),
    .Y(_0095_),
    .B1(_0357_));
 sg13g2_o21ai_1 _1992_ (.B1(net575),
    .Y(_0358_),
    .A1(net337),
    .A2(net529));
 sg13g2_a21oi_1 _1993_ (.A1(_0622_),
    .A2(net529),
    .Y(_0096_),
    .B1(_0358_));
 sg13g2_o21ai_1 _1994_ (.B1(net576),
    .Y(_0359_),
    .A1(\bitserial_cipher.datapath.shift_in2 ),
    .A2(net530));
 sg13g2_a21oi_1 _1995_ (.A1(_0743_),
    .A2(net530),
    .Y(_0097_),
    .B1(_0359_));
 sg13g2_o21ai_1 _1996_ (.B1(net576),
    .Y(_0360_),
    .A1(net669),
    .A2(net530));
 sg13g2_a21oi_1 _1997_ (.A1(_0742_),
    .A2(net530),
    .Y(_0098_),
    .B1(_0360_));
 sg13g2_o21ai_1 _1998_ (.B1(net576),
    .Y(_0361_),
    .A1(net778),
    .A2(net530));
 sg13g2_a21oi_1 _1999_ (.A1(_0741_),
    .A2(net530),
    .Y(_0099_),
    .B1(_0361_));
 sg13g2_o21ai_1 _2000_ (.B1(net576),
    .Y(_0362_),
    .A1(\bitserial_cipher.datapath.shifter1[3] ),
    .A2(net530));
 sg13g2_a21oi_1 _2001_ (.A1(_0740_),
    .A2(net530),
    .Y(_0100_),
    .B1(_0362_));
 sg13g2_o21ai_1 _2002_ (.B1(net571),
    .Y(_0363_),
    .A1(\bitserial_cipher.datapath.shifter1[4] ),
    .A2(net525));
 sg13g2_a21oi_1 _2003_ (.A1(_0739_),
    .A2(net526),
    .Y(_0101_),
    .B1(_0363_));
 sg13g2_o21ai_1 _2004_ (.B1(net573),
    .Y(_0364_),
    .A1(\bitserial_cipher.datapath.shifter1[5] ),
    .A2(net525));
 sg13g2_a21oi_1 _2005_ (.A1(_0738_),
    .A2(net525),
    .Y(_0102_),
    .B1(_0364_));
 sg13g2_o21ai_1 _2006_ (.B1(net572),
    .Y(_0365_),
    .A1(\bitserial_cipher.datapath.shifter1[6] ),
    .A2(net527));
 sg13g2_a21oi_1 _2007_ (.A1(_0737_),
    .A2(net522),
    .Y(_0103_),
    .B1(_0365_));
 sg13g2_o21ai_1 _2008_ (.B1(net572),
    .Y(_0366_),
    .A1(net376),
    .A2(net522));
 sg13g2_a21oi_1 _2009_ (.A1(_0736_),
    .A2(net522),
    .Y(_0104_),
    .B1(_0366_));
 sg13g2_o21ai_1 _2010_ (.B1(net556),
    .Y(_0367_),
    .A1(\bitserial_cipher.datapath.shifter1[8] ),
    .A2(net516));
 sg13g2_a21oi_1 _2011_ (.A1(_0735_),
    .A2(net516),
    .Y(_0105_),
    .B1(_0367_));
 sg13g2_o21ai_1 _2012_ (.B1(net557),
    .Y(_0368_),
    .A1(net362),
    .A2(net515));
 sg13g2_a21oi_1 _2013_ (.A1(_0734_),
    .A2(net515),
    .Y(_0106_),
    .B1(_0368_));
 sg13g2_o21ai_1 _2014_ (.B1(net555),
    .Y(_0369_),
    .A1(net645),
    .A2(net512));
 sg13g2_a21oi_1 _2015_ (.A1(_0733_),
    .A2(net512),
    .Y(_0107_),
    .B1(_0369_));
 sg13g2_o21ai_1 _2016_ (.B1(net555),
    .Y(_0370_),
    .A1(\bitserial_cipher.datapath.shifter1[11] ),
    .A2(net511));
 sg13g2_a21oi_1 _2017_ (.A1(_0732_),
    .A2(net511),
    .Y(_0108_),
    .B1(_0370_));
 sg13g2_o21ai_1 _2018_ (.B1(net558),
    .Y(_0371_),
    .A1(\bitserial_cipher.datapath.shifter1[12] ),
    .A2(net511));
 sg13g2_a21oi_1 _2019_ (.A1(_0731_),
    .A2(net505),
    .Y(_0109_),
    .B1(_0371_));
 sg13g2_o21ai_1 _2020_ (.B1(net552),
    .Y(_0372_),
    .A1(net604),
    .A2(net504));
 sg13g2_a21oi_1 _2021_ (.A1(_0730_),
    .A2(net504),
    .Y(_0110_),
    .B1(_0372_));
 sg13g2_o21ai_1 _2022_ (.B1(net552),
    .Y(_0373_),
    .A1(net629),
    .A2(net504));
 sg13g2_a21oi_1 _2023_ (.A1(_0729_),
    .A2(net504),
    .Y(_0111_),
    .B1(_0373_));
 sg13g2_o21ai_1 _2024_ (.B1(net550),
    .Y(_0374_),
    .A1(\bitserial_cipher.datapath.shifter1[15] ),
    .A2(net502));
 sg13g2_a21oi_1 _2025_ (.A1(_0728_),
    .A2(net502),
    .Y(_0112_),
    .B1(_0374_));
 sg13g2_o21ai_1 _2026_ (.B1(net551),
    .Y(_0375_),
    .A1(net658),
    .A2(net503));
 sg13g2_a21oi_1 _2027_ (.A1(_0727_),
    .A2(net502),
    .Y(_0113_),
    .B1(_0375_));
 sg13g2_o21ai_1 _2028_ (.B1(net550),
    .Y(_0376_),
    .A1(\bitserial_cipher.datapath.shifter1[17] ),
    .A2(net502));
 sg13g2_a21oi_1 _2029_ (.A1(_0726_),
    .A2(net502),
    .Y(_0114_),
    .B1(_0376_));
 sg13g2_o21ai_1 _2030_ (.B1(net549),
    .Y(_0377_),
    .A1(net316),
    .A2(net500));
 sg13g2_a21oi_1 _2031_ (.A1(_0725_),
    .A2(net500),
    .Y(_0115_),
    .B1(_0377_));
 sg13g2_o21ai_1 _2032_ (.B1(net549),
    .Y(_0378_),
    .A1(\bitserial_cipher.datapath.shifter1[19] ),
    .A2(net500));
 sg13g2_a21oi_1 _2033_ (.A1(_0724_),
    .A2(net500),
    .Y(_0116_),
    .B1(_0378_));
 sg13g2_o21ai_1 _2034_ (.B1(net547),
    .Y(_0379_),
    .A1(net412),
    .A2(net496));
 sg13g2_a21oi_1 _2035_ (.A1(_0723_),
    .A2(net496),
    .Y(_0117_),
    .B1(_0379_));
 sg13g2_o21ai_1 _2036_ (.B1(net547),
    .Y(_0380_),
    .A1(\bitserial_cipher.datapath.shifter1[21] ),
    .A2(net496));
 sg13g2_a21oi_1 _2037_ (.A1(_0722_),
    .A2(net496),
    .Y(_0118_),
    .B1(_0380_));
 sg13g2_o21ai_1 _2038_ (.B1(net547),
    .Y(_0381_),
    .A1(net682),
    .A2(net497));
 sg13g2_a21oi_1 _2039_ (.A1(_0721_),
    .A2(net497),
    .Y(_0119_),
    .B1(_0381_));
 sg13g2_o21ai_1 _2040_ (.B1(net553),
    .Y(_0382_),
    .A1(\bitserial_cipher.datapath.shifter1[23] ),
    .A2(net508));
 sg13g2_a21oi_1 _2041_ (.A1(_0720_),
    .A2(net508),
    .Y(_0120_),
    .B1(_0382_));
 sg13g2_o21ai_1 _2042_ (.B1(net553),
    .Y(_0383_),
    .A1(net341),
    .A2(net508));
 sg13g2_a21oi_1 _2043_ (.A1(_0719_),
    .A2(net508),
    .Y(_0121_),
    .B1(_0383_));
 sg13g2_o21ai_1 _2044_ (.B1(net553),
    .Y(_0384_),
    .A1(\bitserial_cipher.datapath.shifter1[25] ),
    .A2(net510));
 sg13g2_a21oi_1 _2045_ (.A1(_0718_),
    .A2(net510),
    .Y(_0122_),
    .B1(_0384_));
 sg13g2_o21ai_1 _2046_ (.B1(net553),
    .Y(_0385_),
    .A1(\bitserial_cipher.datapath.shifter1[26] ),
    .A2(net508));
 sg13g2_a21oi_1 _2047_ (.A1(_0717_),
    .A2(net508),
    .Y(_0123_),
    .B1(_0385_));
 sg13g2_o21ai_1 _2048_ (.B1(net554),
    .Y(_0386_),
    .A1(net432),
    .A2(net518));
 sg13g2_a21oi_1 _2049_ (.A1(_0716_),
    .A2(net518),
    .Y(_0124_),
    .B1(_0386_));
 sg13g2_o21ai_1 _2050_ (.B1(net553),
    .Y(_0387_),
    .A1(\bitserial_cipher.datapath.shifter1[28] ),
    .A2(net508));
 sg13g2_a21oi_1 _2051_ (.A1(_0715_),
    .A2(net508),
    .Y(_0125_),
    .B1(_0387_));
 sg13g2_o21ai_1 _2052_ (.B1(net553),
    .Y(_0388_),
    .A1(net353),
    .A2(net510));
 sg13g2_a21oi_1 _2053_ (.A1(_0714_),
    .A2(net510),
    .Y(_0126_),
    .B1(_0388_));
 sg13g2_o21ai_1 _2054_ (.B1(net553),
    .Y(_0389_),
    .A1(net745),
    .A2(net509));
 sg13g2_a21oi_1 _2055_ (.A1(_0713_),
    .A2(net509),
    .Y(_0127_),
    .B1(_0389_));
 sg13g2_o21ai_1 _2056_ (.B1(net553),
    .Y(_0390_),
    .A1(net760),
    .A2(net509));
 sg13g2_a21oi_1 _2057_ (.A1(_0712_),
    .A2(net509),
    .Y(_0128_),
    .B1(_0390_));
 sg13g2_o21ai_1 _2058_ (.B1(net547),
    .Y(_0391_),
    .A1(\bitserial_cipher.datapath.shifter1[32] ),
    .A2(net496));
 sg13g2_a21oi_1 _2059_ (.A1(_0711_),
    .A2(net506),
    .Y(_0129_),
    .B1(_0391_));
 sg13g2_o21ai_1 _2060_ (.B1(net552),
    .Y(_0392_),
    .A1(net591),
    .A2(net506));
 sg13g2_a21oi_1 _2061_ (.A1(_0710_),
    .A2(net506),
    .Y(_0130_),
    .B1(_0392_));
 sg13g2_o21ai_1 _2062_ (.B1(net552),
    .Y(_0393_),
    .A1(net626),
    .A2(net506));
 sg13g2_a21oi_1 _2063_ (.A1(_0709_),
    .A2(net500),
    .Y(_0131_),
    .B1(_0393_));
 sg13g2_o21ai_1 _2064_ (.B1(net550),
    .Y(_0394_),
    .A1(net800),
    .A2(net502));
 sg13g2_a21oi_1 _2065_ (.A1(_0708_),
    .A2(net502),
    .Y(_0132_),
    .B1(_0394_));
 sg13g2_o21ai_1 _2066_ (.B1(net550),
    .Y(_0395_),
    .A1(\bitserial_cipher.datapath.shifter1[36] ),
    .A2(net501));
 sg13g2_a21oi_1 _2067_ (.A1(_0707_),
    .A2(net501),
    .Y(_0133_),
    .B1(_0395_));
 sg13g2_o21ai_1 _2068_ (.B1(net550),
    .Y(_0396_),
    .A1(\bitserial_cipher.datapath.shifter1[37] ),
    .A2(net501));
 sg13g2_a21oi_1 _2069_ (.A1(_0706_),
    .A2(net501),
    .Y(_0134_),
    .B1(_0396_));
 sg13g2_o21ai_1 _2070_ (.B1(net550),
    .Y(_0397_),
    .A1(\bitserial_cipher.datapath.shifter1[38] ),
    .A2(net501));
 sg13g2_a21oi_1 _2071_ (.A1(_0705_),
    .A2(net501),
    .Y(_0135_),
    .B1(_0397_));
 sg13g2_o21ai_1 _2072_ (.B1(net550),
    .Y(_0398_),
    .A1(\bitserial_cipher.datapath.shifter1[39] ),
    .A2(net501));
 sg13g2_a21oi_1 _2073_ (.A1(_0704_),
    .A2(net501),
    .Y(_0136_),
    .B1(_0398_));
 sg13g2_o21ai_1 _2074_ (.B1(net550),
    .Y(_0399_),
    .A1(net325),
    .A2(net503));
 sg13g2_a21oi_1 _2075_ (.A1(_0703_),
    .A2(net503),
    .Y(_0137_),
    .B1(_0399_));
 sg13g2_o21ai_1 _2076_ (.B1(net551),
    .Y(_0400_),
    .A1(net639),
    .A2(net503));
 sg13g2_a21oi_1 _2077_ (.A1(_0702_),
    .A2(net503),
    .Y(_0138_),
    .B1(_0400_));
 sg13g2_o21ai_1 _2078_ (.B1(net552),
    .Y(_0401_),
    .A1(\bitserial_cipher.datapath.shifter1[42] ),
    .A2(net504));
 sg13g2_a21oi_1 _2079_ (.A1(_0701_),
    .A2(net504),
    .Y(_0139_),
    .B1(_0401_));
 sg13g2_o21ai_1 _2080_ (.B1(net559),
    .Y(_0402_),
    .A1(net349),
    .A2(net505));
 sg13g2_a21oi_1 _2081_ (.A1(_0700_),
    .A2(net511),
    .Y(_0140_),
    .B1(_0402_));
 sg13g2_o21ai_1 _2082_ (.B1(net555),
    .Y(_0403_),
    .A1(net717),
    .A2(net512));
 sg13g2_a21oi_1 _2083_ (.A1(_0699_),
    .A2(net512),
    .Y(_0141_),
    .B1(_0403_));
 sg13g2_o21ai_1 _2084_ (.B1(net557),
    .Y(_0404_),
    .A1(\bitserial_cipher.datapath.shifter1[45] ),
    .A2(net515));
 sg13g2_a21oi_1 _2085_ (.A1(_0698_),
    .A2(net515),
    .Y(_0142_),
    .B1(_0404_));
 sg13g2_o21ai_1 _2086_ (.B1(net557),
    .Y(_0405_),
    .A1(\bitserial_cipher.datapath.shifter1[46] ),
    .A2(net516));
 sg13g2_a21oi_1 _2087_ (.A1(_0697_),
    .A2(net516),
    .Y(_0143_),
    .B1(_0405_));
 sg13g2_o21ai_1 _2088_ (.B1(net572),
    .Y(_0406_),
    .A1(\bitserial_cipher.datapath.shifter1[47] ),
    .A2(net522));
 sg13g2_a21oi_1 _2089_ (.A1(_0696_),
    .A2(net522),
    .Y(_0144_),
    .B1(_0406_));
 sg13g2_o21ai_1 _2090_ (.B1(net572),
    .Y(_0407_),
    .A1(\bitserial_cipher.datapath.shifter1[48] ),
    .A2(net522));
 sg13g2_a21oi_1 _2091_ (.A1(_0695_),
    .A2(net522),
    .Y(_0145_),
    .B1(_0407_));
 sg13g2_o21ai_1 _2092_ (.B1(net573),
    .Y(_0408_),
    .A1(\bitserial_cipher.datapath.shifter1[49] ),
    .A2(net525));
 sg13g2_a21oi_1 _2093_ (.A1(_0694_),
    .A2(net525),
    .Y(_0146_),
    .B1(_0408_));
 sg13g2_o21ai_1 _2094_ (.B1(net571),
    .Y(_0409_),
    .A1(\bitserial_cipher.datapath.shifter1[50] ),
    .A2(net525));
 sg13g2_a21oi_1 _2095_ (.A1(_0693_),
    .A2(net525),
    .Y(_0147_),
    .B1(_0409_));
 sg13g2_o21ai_1 _2096_ (.B1(net571),
    .Y(_0410_),
    .A1(net374),
    .A2(net525));
 sg13g2_a21oi_1 _2097_ (.A1(_0692_),
    .A2(net526),
    .Y(_0148_),
    .B1(_0410_));
 sg13g2_o21ai_1 _2098_ (.B1(net571),
    .Y(_0411_),
    .A1(\bitserial_cipher.datapath.shifter1[52] ),
    .A2(net524));
 sg13g2_a21oi_1 _2099_ (.A1(_0691_),
    .A2(net524),
    .Y(_0149_),
    .B1(_0411_));
 sg13g2_o21ai_1 _2100_ (.B1(net571),
    .Y(_0412_),
    .A1(net323),
    .A2(net524));
 sg13g2_a21oi_1 _2101_ (.A1(_0690_),
    .A2(net528),
    .Y(_0150_),
    .B1(_0412_));
 sg13g2_o21ai_1 _2102_ (.B1(net574),
    .Y(_0413_),
    .A1(\bitserial_cipher.datapath.shifter1[55] ),
    .A2(net444));
 sg13g2_a21oi_1 _2103_ (.A1(_0690_),
    .A2(net444),
    .Y(_0151_),
    .B1(_0413_));
 sg13g2_nor2_1 _2104_ (.A(_0832_),
    .B(net486),
    .Y(_0414_));
 sg13g2_xor2_1 _2105_ (.B(_0865_),
    .A(net441),
    .X(_0415_));
 sg13g2_nor2_1 _2106_ (.A(_0414_),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_o21ai_1 _2107_ (.B1(net528),
    .Y(_0417_),
    .A1(\bitserial_cipher.datapath.fifo_ff56 ),
    .A2(_0416_));
 sg13g2_a21oi_1 _2108_ (.A1(_0835_),
    .A2(_0416_),
    .Y(_0418_),
    .B1(_0417_));
 sg13g2_a21oi_1 _2109_ (.A1(net788),
    .A2(_0832_),
    .Y(_0419_),
    .B1(_0418_));
 sg13g2_nor2_1 _2110_ (.A(_0834_),
    .B(net789),
    .Y(_0152_));
 sg13g2_o21ai_1 _2111_ (.B1(net577),
    .Y(_0420_),
    .A1(\bitserial_cipher.cipher_data ),
    .A2(net532));
 sg13g2_a21oi_1 _2112_ (.A1(_0689_),
    .A2(net532),
    .Y(_0153_),
    .B1(_0420_));
 sg13g2_o21ai_1 _2113_ (.B1(net573),
    .Y(_0421_),
    .A1(net579),
    .A2(net521));
 sg13g2_a21oi_1 _2114_ (.A1(_0688_),
    .A2(net521),
    .Y(_0154_),
    .B1(_0421_));
 sg13g2_o21ai_1 _2115_ (.B1(net573),
    .Y(_0422_),
    .A1(\bitserial_cipher.datapath.shifter2[2] ),
    .A2(net521));
 sg13g2_a21oi_1 _2116_ (.A1(_0687_),
    .A2(net521),
    .Y(_0155_),
    .B1(_0422_));
 sg13g2_o21ai_1 _2117_ (.B1(net570),
    .Y(_0423_),
    .A1(net420),
    .A2(net519));
 sg13g2_a21oi_1 _2118_ (.A1(_0686_),
    .A2(net519),
    .Y(_0156_),
    .B1(_0423_));
 sg13g2_o21ai_1 _2119_ (.B1(net570),
    .Y(_0424_),
    .A1(\bitserial_cipher.datapath.shifter2[4] ),
    .A2(net519));
 sg13g2_a21oi_1 _2120_ (.A1(_0685_),
    .A2(net519),
    .Y(_0157_),
    .B1(_0424_));
 sg13g2_o21ai_1 _2121_ (.B1(net570),
    .Y(_0425_),
    .A1(\bitserial_cipher.datapath.shifter2[5] ),
    .A2(net519));
 sg13g2_a21oi_1 _2122_ (.A1(_0684_),
    .A2(net519),
    .Y(_0158_),
    .B1(_0425_));
 sg13g2_o21ai_1 _2123_ (.B1(net570),
    .Y(_0426_),
    .A1(net366),
    .A2(net519));
 sg13g2_a21oi_1 _2124_ (.A1(_0683_),
    .A2(net519),
    .Y(_0159_),
    .B1(_0426_));
 sg13g2_o21ai_1 _2125_ (.B1(net570),
    .Y(_0427_),
    .A1(net386),
    .A2(net520));
 sg13g2_a21oi_1 _2126_ (.A1(_0682_),
    .A2(net520),
    .Y(_0160_),
    .B1(_0427_));
 sg13g2_o21ai_1 _2127_ (.B1(net570),
    .Y(_0428_),
    .A1(net661),
    .A2(net520));
 sg13g2_a21oi_1 _2128_ (.A1(_0681_),
    .A2(net520),
    .Y(_0161_),
    .B1(_0428_));
 sg13g2_o21ai_1 _2129_ (.B1(net570),
    .Y(_0429_),
    .A1(\bitserial_cipher.datapath.shifter2[9] ),
    .A2(net520));
 sg13g2_a21oi_1 _2130_ (.A1(_0680_),
    .A2(net520),
    .Y(_0162_),
    .B1(_0429_));
 sg13g2_o21ai_1 _2131_ (.B1(net570),
    .Y(_0430_),
    .A1(\bitserial_cipher.datapath.shifter2[10] ),
    .A2(net520));
 sg13g2_a21oi_1 _2132_ (.A1(_0679_),
    .A2(net520),
    .Y(_0163_),
    .B1(_0430_));
 sg13g2_o21ai_1 _2133_ (.B1(net572),
    .Y(_0431_),
    .A1(net384),
    .A2(net523));
 sg13g2_a21oi_1 _2134_ (.A1(_0678_),
    .A2(net523),
    .Y(_0164_),
    .B1(_0431_));
 sg13g2_o21ai_1 _2135_ (.B1(net556),
    .Y(_0432_),
    .A1(\bitserial_cipher.datapath.shifter2[12] ),
    .A2(net517));
 sg13g2_a21oi_1 _2136_ (.A1(_0677_),
    .A2(net517),
    .Y(_0165_),
    .B1(_0432_));
 sg13g2_o21ai_1 _2137_ (.B1(net556),
    .Y(_0433_),
    .A1(net676),
    .A2(net514));
 sg13g2_a21oi_1 _2138_ (.A1(_0676_),
    .A2(net517),
    .Y(_0166_),
    .B1(_0433_));
 sg13g2_o21ai_1 _2139_ (.B1(net556),
    .Y(_0434_),
    .A1(\bitserial_cipher.datapath.shifter2[14] ),
    .A2(net514));
 sg13g2_a21oi_1 _2140_ (.A1(_0675_),
    .A2(net514),
    .Y(_0167_),
    .B1(_0434_));
 sg13g2_o21ai_1 _2141_ (.B1(net556),
    .Y(_0435_),
    .A1(net422),
    .A2(net514));
 sg13g2_a21oi_1 _2142_ (.A1(_0674_),
    .A2(net514),
    .Y(_0168_),
    .B1(_0435_));
 sg13g2_o21ai_1 _2143_ (.B1(net556),
    .Y(_0436_),
    .A1(\bitserial_cipher.datapath.shifter2[16] ),
    .A2(net514));
 sg13g2_a21oi_1 _2144_ (.A1(_0673_),
    .A2(net514),
    .Y(_0169_),
    .B1(_0436_));
 sg13g2_o21ai_1 _2145_ (.B1(net556),
    .Y(_0437_),
    .A1(net351),
    .A2(net514));
 sg13g2_a21oi_1 _2146_ (.A1(_0672_),
    .A2(net513),
    .Y(_0170_),
    .B1(_0437_));
 sg13g2_o21ai_1 _2147_ (.B1(net555),
    .Y(_0438_),
    .A1(\bitserial_cipher.datapath.shifter2[18] ),
    .A2(net513));
 sg13g2_a21oi_1 _2148_ (.A1(_0671_),
    .A2(net513),
    .Y(_0171_),
    .B1(_0438_));
 sg13g2_o21ai_1 _2149_ (.B1(net555),
    .Y(_0439_),
    .A1(net623),
    .A2(net513));
 sg13g2_a21oi_1 _2150_ (.A1(_0670_),
    .A2(net513),
    .Y(_0172_),
    .B1(_0439_));
 sg13g2_o21ai_1 _2151_ (.B1(net555),
    .Y(_0440_),
    .A1(\bitserial_cipher.datapath.shifter2[20] ),
    .A2(net513));
 sg13g2_a21oi_1 _2152_ (.A1(_0669_),
    .A2(net510),
    .Y(_0173_),
    .B1(_0440_));
 sg13g2_o21ai_1 _2153_ (.B1(net554),
    .Y(_0441_),
    .A1(\bitserial_cipher.datapath.shifter2[21] ),
    .A2(net509));
 sg13g2_a21oi_1 _2154_ (.A1(_0668_),
    .A2(net509),
    .Y(_0174_),
    .B1(_0441_));
 sg13g2_o21ai_1 _2155_ (.B1(net554),
    .Y(_0442_),
    .A1(net380),
    .A2(net509));
 sg13g2_a21oi_1 _2156_ (.A1(_0667_),
    .A2(net509),
    .Y(_0175_),
    .B1(_0442_));
 sg13g2_o21ai_1 _2157_ (.B1(net548),
    .Y(_0443_),
    .A1(\bitserial_cipher.datapath.shifter2[23] ),
    .A2(net496));
 sg13g2_a21oi_1 _2158_ (.A1(_0666_),
    .A2(net496),
    .Y(_0176_),
    .B1(_0443_));
 sg13g2_o21ai_1 _2159_ (.B1(net548),
    .Y(_0444_),
    .A1(\bitserial_cipher.datapath.shifter2[24] ),
    .A2(net497));
 sg13g2_a21oi_1 _2160_ (.A1(_0665_),
    .A2(net496),
    .Y(_0177_),
    .B1(_0444_));
 sg13g2_o21ai_1 _2161_ (.B1(net547),
    .Y(_0445_),
    .A1(net392),
    .A2(net495));
 sg13g2_a21oi_1 _2162_ (.A1(_0664_),
    .A2(net495),
    .Y(_0178_),
    .B1(_0445_));
 sg13g2_o21ai_1 _2163_ (.B1(net547),
    .Y(_0446_),
    .A1(net612),
    .A2(net495));
 sg13g2_a21oi_1 _2164_ (.A1(_0663_),
    .A2(net495),
    .Y(_0179_),
    .B1(_0446_));
 sg13g2_o21ai_1 _2165_ (.B1(net547),
    .Y(_0447_),
    .A1(\bitserial_cipher.datapath.shifter2[27] ),
    .A2(net495));
 sg13g2_a21oi_1 _2166_ (.A1(_0662_),
    .A2(net495),
    .Y(_0180_),
    .B1(_0447_));
 sg13g2_o21ai_1 _2167_ (.B1(net547),
    .Y(_0448_),
    .A1(net414),
    .A2(net495));
 sg13g2_a21oi_1 _2168_ (.A1(_0661_),
    .A2(net495),
    .Y(_0181_),
    .B1(_0448_));
 sg13g2_o21ai_1 _2169_ (.B1(net545),
    .Y(_0449_),
    .A1(net755),
    .A2(net492));
 sg13g2_a21oi_1 _2170_ (.A1(_0660_),
    .A2(net492),
    .Y(_0182_),
    .B1(_0449_));
 sg13g2_o21ai_1 _2171_ (.B1(net546),
    .Y(_0450_),
    .A1(\bitserial_cipher.datapath.shifter2[30] ),
    .A2(net492));
 sg13g2_a21oi_1 _2172_ (.A1(_0659_),
    .A2(net492),
    .Y(_0183_),
    .B1(_0450_));
 sg13g2_o21ai_1 _2173_ (.B1(net545),
    .Y(_0451_),
    .A1(net656),
    .A2(net491));
 sg13g2_a21oi_1 _2174_ (.A1(_0658_),
    .A2(net490),
    .Y(_0184_),
    .B1(_0451_));
 sg13g2_o21ai_1 _2175_ (.B1(net545),
    .Y(_0452_),
    .A1(\bitserial_cipher.datapath.shifter2[32] ),
    .A2(net490));
 sg13g2_a21oi_1 _2176_ (.A1(_0657_),
    .A2(net490),
    .Y(_0185_),
    .B1(_0452_));
 sg13g2_o21ai_1 _2177_ (.B1(net545),
    .Y(_0453_),
    .A1(\bitserial_cipher.datapath.shifter2[33] ),
    .A2(net490));
 sg13g2_a21oi_1 _2178_ (.A1(_0656_),
    .A2(net490),
    .Y(_0186_),
    .B1(_0453_));
 sg13g2_o21ai_1 _2179_ (.B1(net545),
    .Y(_0454_),
    .A1(net364),
    .A2(net490));
 sg13g2_a21oi_1 _2180_ (.A1(_0655_),
    .A2(net490),
    .Y(_0187_),
    .B1(_0454_));
 sg13g2_o21ai_1 _2181_ (.B1(net545),
    .Y(_0455_),
    .A1(net640),
    .A2(net490));
 sg13g2_a21oi_1 _2182_ (.A1(_0654_),
    .A2(net491),
    .Y(_0188_),
    .B1(_0455_));
 sg13g2_o21ai_1 _2183_ (.B1(net545),
    .Y(_0456_),
    .A1(\bitserial_cipher.datapath.shifter2[36] ),
    .A2(net491));
 sg13g2_a21oi_1 _2184_ (.A1(_0653_),
    .A2(net491),
    .Y(_0189_),
    .B1(_0456_));
 sg13g2_o21ai_1 _2185_ (.B1(net545),
    .Y(_0457_),
    .A1(net715),
    .A2(net491));
 sg13g2_a21oi_1 _2186_ (.A1(_0652_),
    .A2(net491),
    .Y(_0190_),
    .B1(_0457_));
 sg13g2_o21ai_1 _2187_ (.B1(net546),
    .Y(_0458_),
    .A1(\bitserial_cipher.datapath.shifter2[38] ),
    .A2(net493));
 sg13g2_a21oi_1 _2188_ (.A1(_0651_),
    .A2(net493),
    .Y(_0191_),
    .B1(_0458_));
 sg13g2_o21ai_1 _2189_ (.B1(net546),
    .Y(_0459_),
    .A1(net729),
    .A2(net493));
 sg13g2_a21oi_1 _2190_ (.A1(_0650_),
    .A2(net493),
    .Y(_0192_),
    .B1(_0459_));
 sg13g2_o21ai_1 _2191_ (.B1(net546),
    .Y(_0460_),
    .A1(\bitserial_cipher.datapath.shifter2[40] ),
    .A2(net494));
 sg13g2_a21oi_1 _2192_ (.A1(_0649_),
    .A2(net494),
    .Y(_0193_),
    .B1(_0460_));
 sg13g2_o21ai_1 _2193_ (.B1(net546),
    .Y(_0461_),
    .A1(\bitserial_cipher.datapath.shifter2[41] ),
    .A2(net493));
 sg13g2_a21oi_1 _2194_ (.A1(_0648_),
    .A2(net493),
    .Y(_0194_),
    .B1(_0461_));
 sg13g2_o21ai_1 _2195_ (.B1(net546),
    .Y(_0462_),
    .A1(net339),
    .A2(net493));
 sg13g2_a21oi_1 _2196_ (.A1(_0647_),
    .A2(net493),
    .Y(_0195_),
    .B1(_0462_));
 sg13g2_o21ai_1 _2197_ (.B1(net549),
    .Y(_0463_),
    .A1(\bitserial_cipher.datapath.shifter2[43] ),
    .A2(net498));
 sg13g2_a21oi_1 _2198_ (.A1(_0646_),
    .A2(net498),
    .Y(_0196_),
    .B1(_0463_));
 sg13g2_o21ai_1 _2199_ (.B1(net549),
    .Y(_0464_),
    .A1(net345),
    .A2(net498));
 sg13g2_a21oi_1 _2200_ (.A1(_0645_),
    .A2(net498),
    .Y(_0197_),
    .B1(_0464_));
 sg13g2_o21ai_1 _2201_ (.B1(net549),
    .Y(_0465_),
    .A1(net737),
    .A2(net498));
 sg13g2_a21oi_1 _2202_ (.A1(_0644_),
    .A2(net498),
    .Y(_0198_),
    .B1(_0465_));
 sg13g2_o21ai_1 _2203_ (.B1(net549),
    .Y(_0466_),
    .A1(\bitserial_cipher.datapath.shifter2[46] ),
    .A2(net499));
 sg13g2_a21oi_1 _2204_ (.A1(_0643_),
    .A2(net499),
    .Y(_0199_),
    .B1(_0466_));
 sg13g2_o21ai_1 _2205_ (.B1(net549),
    .Y(_0467_),
    .A1(\bitserial_cipher.datapath.shifter2[47] ),
    .A2(net499));
 sg13g2_a21oi_1 _2206_ (.A1(_0642_),
    .A2(net499),
    .Y(_0200_),
    .B1(_0467_));
 sg13g2_o21ai_1 _2207_ (.B1(net549),
    .Y(_0468_),
    .A1(net312),
    .A2(net498));
 sg13g2_a21oi_1 _2208_ (.A1(_0641_),
    .A2(net498),
    .Y(_0201_),
    .B1(_0468_));
 sg13g2_o21ai_1 _2209_ (.B1(net551),
    .Y(_0469_),
    .A1(net807),
    .A2(net502));
 sg13g2_a21oi_1 _2210_ (.A1(_0640_),
    .A2(net500),
    .Y(_0202_),
    .B1(_0469_));
 sg13g2_o21ai_1 _2211_ (.B1(net552),
    .Y(_0470_),
    .A1(\bitserial_cipher.datapath.shifter2[50] ),
    .A2(net504));
 sg13g2_a21oi_1 _2212_ (.A1(_0639_),
    .A2(net504),
    .Y(_0203_),
    .B1(_0470_));
 sg13g2_o21ai_1 _2213_ (.B1(net552),
    .Y(_0471_),
    .A1(\bitserial_cipher.datapath.shifter2[51] ),
    .A2(net505));
 sg13g2_a21oi_1 _2214_ (.A1(_0638_),
    .A2(net505),
    .Y(_0204_),
    .B1(_0471_));
 sg13g2_o21ai_1 _2215_ (.B1(net558),
    .Y(_0472_),
    .A1(\bitserial_cipher.datapath.shifter2[52] ),
    .A2(net511));
 sg13g2_a21oi_1 _2216_ (.A1(_0637_),
    .A2(net511),
    .Y(_0205_),
    .B1(_0472_));
 sg13g2_o21ai_1 _2217_ (.B1(net555),
    .Y(_0473_),
    .A1(net329),
    .A2(net512));
 sg13g2_a21oi_1 _2218_ (.A1(_0636_),
    .A2(net511),
    .Y(_0206_),
    .B1(_0473_));
 sg13g2_o21ai_1 _2219_ (.B1(net555),
    .Y(_0474_),
    .A1(net609),
    .A2(net511));
 sg13g2_a21oi_1 _2220_ (.A1(_0635_),
    .A2(net515),
    .Y(_0207_),
    .B1(_0474_));
 sg13g2_o21ai_1 _2221_ (.B1(net556),
    .Y(_0475_),
    .A1(\bitserial_cipher.datapath.shifter2[55] ),
    .A2(net515));
 sg13g2_a21oi_1 _2222_ (.A1(_0634_),
    .A2(net515),
    .Y(_0208_),
    .B1(_0475_));
 sg13g2_o21ai_1 _2223_ (.B1(net557),
    .Y(_0476_),
    .A1(net394),
    .A2(net516));
 sg13g2_a21oi_1 _2224_ (.A1(_0633_),
    .A2(net515),
    .Y(_0209_),
    .B1(_0476_));
 sg13g2_o21ai_1 _2225_ (.B1(net572),
    .Y(_0477_),
    .A1(\bitserial_cipher.datapath.shifter2[57] ),
    .A2(net522));
 sg13g2_a21oi_1 _2226_ (.A1(_0632_),
    .A2(net523),
    .Y(_0210_),
    .B1(_0477_));
 sg13g2_o21ai_1 _2227_ (.B1(net572),
    .Y(_0478_),
    .A1(\bitserial_cipher.datapath.shifter2[58] ),
    .A2(net523));
 sg13g2_a21oi_1 _2228_ (.A1(_0631_),
    .A2(net523),
    .Y(_0211_),
    .B1(_0478_));
 sg13g2_o21ai_1 _2229_ (.B1(net572),
    .Y(_0479_),
    .A1(net347),
    .A2(net523));
 sg13g2_a21oi_1 _2230_ (.A1(_0630_),
    .A2(net523),
    .Y(_0212_),
    .B1(_0479_));
 sg13g2_o21ai_1 _2231_ (.B1(net571),
    .Y(_0480_),
    .A1(\bitserial_cipher.datapath.shifter2[60] ),
    .A2(net524));
 sg13g2_a21oi_1 _2232_ (.A1(_0629_),
    .A2(net524),
    .Y(_0213_),
    .B1(_0480_));
 sg13g2_o21ai_1 _2233_ (.B1(net571),
    .Y(_0481_),
    .A1(\bitserial_cipher.datapath.shifter2[61] ),
    .A2(net524));
 sg13g2_a21oi_1 _2234_ (.A1(_0628_),
    .A2(net524),
    .Y(_0214_),
    .B1(_0481_));
 sg13g2_o21ai_1 _2235_ (.B1(net571),
    .Y(_0482_),
    .A1(\bitserial_cipher.datapath.shifter2[62] ),
    .A2(net526));
 sg13g2_a21oi_1 _2236_ (.A1(_0626_),
    .A2(net524),
    .Y(_0215_),
    .B1(_0482_));
 sg13g2_o21ai_1 _2237_ (.B1(net574),
    .Y(_0483_),
    .A1(net355),
    .A2(net528));
 sg13g2_a21oi_1 _2238_ (.A1(_0627_),
    .A2(net528),
    .Y(_0216_),
    .B1(_0483_));
 sg13g2_o21ai_1 _2239_ (.B1(net575),
    .Y(_0484_),
    .A1(\bitserial_cipher.datapath.fifo_ff56 ),
    .A2(net529));
 sg13g2_a21oi_1 _2240_ (.A1(_0625_),
    .A2(net529),
    .Y(_0217_),
    .B1(_0484_));
 sg13g2_nor2_1 _2241_ (.A(\bitserial_cipher.bit_counter[0] ),
    .B(_0297_),
    .Y(_0485_));
 sg13g2_o21ai_1 _2242_ (.B1(net574),
    .Y(_0486_),
    .A1(net528),
    .A2(net487));
 sg13g2_nor3_1 _2243_ (.A(net835),
    .B(net444),
    .C(_0833_),
    .Y(_0487_));
 sg13g2_nor3_1 _2244_ (.A(_0485_),
    .B(_0486_),
    .C(_0487_),
    .Y(_0218_));
 sg13g2_a21oi_1 _2245_ (.A1(\bitserial_cipher.bit_counter[0] ),
    .A2(_0297_),
    .Y(_0488_),
    .B1(net816));
 sg13g2_and3_1 _2246_ (.X(_0489_),
    .A(net816),
    .B(net846),
    .C(_0297_));
 sg13g2_nor3_1 _2247_ (.A(_0486_),
    .B(net817),
    .C(_0489_),
    .Y(_0219_));
 sg13g2_nor2_1 _2248_ (.A(net820),
    .B(_0489_),
    .Y(_0490_));
 sg13g2_and2_1 _2249_ (.A(net820),
    .B(_0489_),
    .X(_0491_));
 sg13g2_nor3_1 _2250_ (.A(_0486_),
    .B(_0490_),
    .C(_0491_),
    .Y(_0220_));
 sg13g2_nor2_1 _2251_ (.A(net848),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_and2_1 _2252_ (.A(net848),
    .B(_0491_),
    .X(_0493_));
 sg13g2_nor3_1 _2253_ (.A(_0486_),
    .B(_0492_),
    .C(_0493_),
    .Y(_0221_));
 sg13g2_and2_1 _2254_ (.A(net842),
    .B(_0493_),
    .X(_0494_));
 sg13g2_nor2_1 _2255_ (.A(net842),
    .B(_0493_),
    .Y(_0495_));
 sg13g2_nor3_1 _2256_ (.A(_0486_),
    .B(_0494_),
    .C(net843),
    .Y(_0222_));
 sg13g2_nor2_1 _2257_ (.A(net847),
    .B(_0494_),
    .Y(_0496_));
 sg13g2_and2_1 _2258_ (.A(net847),
    .B(_0494_),
    .X(_0497_));
 sg13g2_a21oi_2 _2259_ (.B1(net438),
    .Y(_0498_),
    .A2(_0833_),
    .A1(net444));
 sg13g2_nor3_1 _2260_ (.A(_0486_),
    .B(_0496_),
    .C(net438),
    .Y(_0223_));
 sg13g2_nand2_1 _2261_ (.Y(_0499_),
    .A(net442),
    .B(\bitserial_cipher.datapath.lut_ff62 ));
 sg13g2_o21ai_1 _2262_ (.B1(_0499_),
    .Y(_0500_),
    .A1(net442),
    .A2(_0623_));
 sg13g2_xor2_1 _2263_ (.B(\bitserial_cipher.cipher_data ),
    .A(\bitserial_cipher.datapath.key_in ),
    .X(_0501_));
 sg13g2_xnor2_1 _2264_ (.Y(_0502_),
    .A(_0500_),
    .B(_0501_));
 sg13g2_a21oi_1 _2265_ (.A1(\bitserial_cipher.datapath.fifo_ff63 ),
    .A2(\bitserial_cipher.datapath.fifo_ff56 ),
    .Y(_0503_),
    .B1(net442));
 sg13g2_nand2_1 _2266_ (.Y(_0504_),
    .A(\bitserial_cipher.datapath.lut_ff63 ),
    .B(\bitserial_cipher.datapath.lut_ff56 ));
 sg13g2_a21oi_1 _2267_ (.A1(net442),
    .A2(_0504_),
    .Y(_0505_),
    .B1(_0503_));
 sg13g2_xnor2_1 _2268_ (.Y(_0506_),
    .A(_0502_),
    .B(_0505_));
 sg13g2_o21ai_1 _2269_ (.B1(net574),
    .Y(_0507_),
    .A1(net442),
    .A2(_0506_));
 sg13g2_a21oi_1 _2270_ (.A1(net442),
    .A2(_0627_),
    .Y(_0224_),
    .B1(_0507_));
 sg13g2_and2_1 _2271_ (.A(net574),
    .B(net320),
    .X(_0225_));
 sg13g2_and2_1 _2272_ (.A(net574),
    .B(net359),
    .X(_0226_));
 sg13g2_and2_1 _2273_ (.A(net575),
    .B(net305),
    .X(_0227_));
 sg13g2_and2_1 _2274_ (.A(net575),
    .B(net307),
    .X(_0228_));
 sg13g2_and2_1 _2275_ (.A(net576),
    .B(net308),
    .X(_0229_));
 sg13g2_and2_1 _2276_ (.A(net575),
    .B(net309),
    .X(_0230_));
 sg13g2_o21ai_1 _2277_ (.B1(_0297_),
    .Y(_0508_),
    .A1(net855),
    .A2(_0506_));
 sg13g2_a21o_1 _2278_ (.A2(net855),
    .A1(_0627_),
    .B1(_0508_),
    .X(_0509_));
 sg13g2_a22oi_1 _2279_ (.Y(_0510_),
    .B1(net1),
    .B2(_0414_),
    .A2(_0832_),
    .A1(net823));
 sg13g2_a21oi_1 _2280_ (.A1(_0509_),
    .A2(_0510_),
    .Y(_0231_),
    .B1(_0834_));
 sg13g2_o21ai_1 _2281_ (.B1(net574),
    .Y(_0511_),
    .A1(\bitserial_cipher.datapath.fifo_ff62 ),
    .A2(net528));
 sg13g2_a21oi_1 _2282_ (.A1(_0624_),
    .A2(net528),
    .Y(_0232_),
    .B1(_0511_));
 sg13g2_o21ai_1 _2283_ (.B1(net575),
    .Y(_0512_),
    .A1(net611),
    .A2(net529));
 sg13g2_a21oi_1 _2284_ (.A1(_0623_),
    .A2(net532),
    .Y(_0233_),
    .B1(_0512_));
 sg13g2_and2_1 _2285_ (.A(net575),
    .B(net306),
    .X(_0234_));
 sg13g2_nor2_1 _2286_ (.A(net441),
    .B(net444),
    .Y(_0513_));
 sg13g2_a22oi_1 _2287_ (.Y(_0514_),
    .B1(_0513_),
    .B2(net438),
    .A2(_0498_),
    .A1(net441));
 sg13g2_nor2_1 _2288_ (.A(_0834_),
    .B(_0514_),
    .Y(_0235_));
 sg13g2_nand2_1 _2289_ (.Y(_0515_),
    .A(net440),
    .B(net441));
 sg13g2_xor2_1 _2290_ (.B(net441),
    .A(net440),
    .X(_0516_));
 sg13g2_a22oi_1 _2291_ (.Y(_0517_),
    .B1(_0516_),
    .B2(_0497_),
    .A2(_0498_),
    .A1(net440));
 sg13g2_nor2_1 _2292_ (.A(net443),
    .B(_0517_),
    .Y(_0236_));
 sg13g2_xor2_1 _2293_ (.B(_0515_),
    .A(net851),
    .X(_0518_));
 sg13g2_a22oi_1 _2294_ (.Y(_0519_),
    .B1(_0518_),
    .B2(net438),
    .A2(_0498_),
    .A1(net439));
 sg13g2_nor2_1 _2295_ (.A(net443),
    .B(net852),
    .Y(_0237_));
 sg13g2_nor2_2 _2296_ (.A(_0309_),
    .B(_0515_),
    .Y(_0520_));
 sg13g2_inv_1 _2297_ (.Y(_0521_),
    .A(_0520_));
 sg13g2_a22oi_1 _2298_ (.Y(_0522_),
    .B1(_0521_),
    .B2(net438),
    .A2(_0498_),
    .A1(net859));
 sg13g2_a21oi_1 _2299_ (.A1(net440),
    .A2(net441),
    .Y(_0523_),
    .B1(net859));
 sg13g2_nor4_1 _2300_ (.A(net443),
    .B(_0867_),
    .C(_0522_),
    .D(net860),
    .Y(_0238_));
 sg13g2_xnor2_1 _2301_ (.Y(_0524_),
    .A(_0002_),
    .B(_0520_));
 sg13g2_a22oi_1 _2302_ (.Y(_0525_),
    .B1(_0524_),
    .B2(net438),
    .A2(_0498_),
    .A1(net849));
 sg13g2_nor2_1 _2303_ (.A(net443),
    .B(net850),
    .Y(_0239_));
 sg13g2_nand3_1 _2304_ (.B(net849),
    .C(_0520_),
    .A(\bitserial_cipher.datapath.round_counter[5] ),
    .Y(_0526_));
 sg13g2_a21oi_1 _2305_ (.A1(net849),
    .A2(_0520_),
    .Y(_0527_),
    .B1(net858));
 sg13g2_a22oi_1 _2306_ (.Y(_0528_),
    .B1(_0526_),
    .B2(net438),
    .A2(_0498_),
    .A1(net858));
 sg13g2_nor3_1 _2307_ (.A(net443),
    .B(_0527_),
    .C(_0528_),
    .Y(_0240_));
 sg13g2_xnor2_1 _2308_ (.Y(_0529_),
    .A(_0836_),
    .B(_0526_));
 sg13g2_a22oi_1 _2309_ (.Y(_0530_),
    .B1(_0529_),
    .B2(net438),
    .A2(_0498_),
    .A1(net856));
 sg13g2_nor2_1 _2310_ (.A(net443),
    .B(net857),
    .Y(_0241_));
 sg13g2_o21ai_1 _2311_ (.B1(net567),
    .Y(_0531_),
    .A1(\bitserial_cipher.key_exp.lut_ff0 ),
    .A2(_0298_));
 sg13g2_a21oi_1 _2312_ (.A1(_0619_),
    .A2(_0298_),
    .Y(_0242_),
    .B1(_0531_));
 sg13g2_o21ai_1 _2313_ (.B1(net567),
    .Y(_0532_),
    .A1(\bitserial_cipher.key_exp.lut_ff1 ),
    .A2(_0298_));
 sg13g2_a21oi_1 _2314_ (.A1(_0618_),
    .A2(_0298_),
    .Y(_0243_),
    .B1(_0532_));
 sg13g2_o21ai_1 _2315_ (.B1(net567),
    .Y(_0533_),
    .A1(\bitserial_cipher.key_exp.lut_ff2 ),
    .A2(_0298_));
 sg13g2_a21oi_1 _2316_ (.A1(_0617_),
    .A2(_0298_),
    .Y(_0244_),
    .B1(_0533_));
 sg13g2_o21ai_1 _2317_ (.B1(net567),
    .Y(_0534_),
    .A1(_0299_),
    .A2(_0350_));
 sg13g2_a21oi_1 _2318_ (.A1(_0617_),
    .A2(_0299_),
    .Y(_0245_),
    .B1(_0534_));
 sg13g2_o21ai_1 _2319_ (.B1(net567),
    .Y(_0535_),
    .A1(\bitserial_cipher.key_exp.fifo_ff0 ),
    .A2(net486));
 sg13g2_a21oi_1 _2320_ (.A1(_0616_),
    .A2(net486),
    .Y(_0246_),
    .B1(_0535_));
 sg13g2_o21ai_1 _2321_ (.B1(net567),
    .Y(_0536_),
    .A1(net335),
    .A2(net486));
 sg13g2_a21oi_1 _2322_ (.A1(_0615_),
    .A2(net486),
    .Y(_0247_),
    .B1(_0536_));
 sg13g2_o21ai_1 _2323_ (.B1(net567),
    .Y(_0537_),
    .A1(net636),
    .A2(net486));
 sg13g2_a21oi_1 _2324_ (.A1(_0613_),
    .A2(net486),
    .Y(_0248_),
    .B1(_0537_));
 sg13g2_o21ai_1 _2325_ (.B1(net567),
    .Y(_0538_),
    .A1(net794),
    .A2(net488));
 sg13g2_a21oi_1 _2326_ (.A1(_0614_),
    .A2(net488),
    .Y(_0249_),
    .B1(_0538_));
 sg13g2_o21ai_1 _2327_ (.B1(net568),
    .Y(_0539_),
    .A1(\bitserial_cipher.datapath.key_in ),
    .A2(net488));
 sg13g2_a21oi_1 _2328_ (.A1(_0612_),
    .A2(net488),
    .Y(_0250_),
    .B1(_0539_));
 sg13g2_o21ai_1 _2329_ (.B1(net568),
    .Y(_0540_),
    .A1(net436),
    .A2(net489));
 sg13g2_a21oi_1 _2330_ (.A1(_0611_),
    .A2(net483),
    .Y(_0251_),
    .B1(_0540_));
 sg13g2_o21ai_1 _2331_ (.B1(net568),
    .Y(_0541_),
    .A1(\bitserial_cipher.key_exp.shifter2[2] ),
    .A2(net484));
 sg13g2_a21oi_1 _2332_ (.A1(_0610_),
    .A2(net484),
    .Y(_0252_),
    .B1(_0541_));
 sg13g2_o21ai_1 _2333_ (.B1(net565),
    .Y(_0542_),
    .A1(net627),
    .A2(net483));
 sg13g2_a21oi_1 _2334_ (.A1(_0609_),
    .A2(net483),
    .Y(_0253_),
    .B1(_0542_));
 sg13g2_o21ai_1 _2335_ (.B1(net565),
    .Y(_0543_),
    .A1(net671),
    .A2(net483));
 sg13g2_a21oi_1 _2336_ (.A1(_0608_),
    .A2(net483),
    .Y(_0254_),
    .B1(_0543_));
 sg13g2_o21ai_1 _2337_ (.B1(net565),
    .Y(_0544_),
    .A1(net763),
    .A2(net480));
 sg13g2_a21oi_1 _2338_ (.A1(_0607_),
    .A2(net480),
    .Y(_0255_),
    .B1(_0544_));
 sg13g2_o21ai_1 _2339_ (.B1(net564),
    .Y(_0545_),
    .A1(net768),
    .A2(net481));
 sg13g2_a21oi_1 _2340_ (.A1(_0606_),
    .A2(net480),
    .Y(_0256_),
    .B1(_0545_));
 sg13g2_o21ai_1 _2341_ (.B1(net564),
    .Y(_0546_),
    .A1(\bitserial_cipher.key_exp.shifter2[7] ),
    .A2(net481));
 sg13g2_a21oi_1 _2342_ (.A1(_0605_),
    .A2(net480),
    .Y(_0257_),
    .B1(_0546_));
 sg13g2_o21ai_1 _2343_ (.B1(net564),
    .Y(_0547_),
    .A1(net600),
    .A2(net481));
 sg13g2_a21oi_1 _2344_ (.A1(_0604_),
    .A2(net481),
    .Y(_0258_),
    .B1(_0547_));
 sg13g2_o21ai_1 _2345_ (.B1(net564),
    .Y(_0548_),
    .A1(net704),
    .A2(net482));
 sg13g2_a21oi_1 _2346_ (.A1(_0603_),
    .A2(net482),
    .Y(_0259_),
    .B1(_0548_));
 sg13g2_o21ai_1 _2347_ (.B1(net563),
    .Y(_0549_),
    .A1(\bitserial_cipher.key_exp.shifter2[10] ),
    .A2(net482));
 sg13g2_a21oi_1 _2348_ (.A1(_0602_),
    .A2(net478),
    .Y(_0260_),
    .B1(_0549_));
 sg13g2_o21ai_1 _2349_ (.B1(net563),
    .Y(_0550_),
    .A1(net310),
    .A2(net478));
 sg13g2_a21oi_1 _2350_ (.A1(_0601_),
    .A2(net478),
    .Y(_0261_),
    .B1(_0550_));
 sg13g2_o21ai_1 _2351_ (.B1(net563),
    .Y(_0551_),
    .A1(\bitserial_cipher.key_exp.shifter2[12] ),
    .A2(net477));
 sg13g2_a21oi_1 _2352_ (.A1(_0600_),
    .A2(net477),
    .Y(_0262_),
    .B1(_0551_));
 sg13g2_o21ai_1 _2353_ (.B1(net561),
    .Y(_0552_),
    .A1(\bitserial_cipher.key_exp.shifter2[13] ),
    .A2(net472));
 sg13g2_a21oi_1 _2354_ (.A1(_0599_),
    .A2(net472),
    .Y(_0263_),
    .B1(_0552_));
 sg13g2_o21ai_1 _2355_ (.B1(net560),
    .Y(_0553_),
    .A1(net654),
    .A2(net470));
 sg13g2_a21oi_1 _2356_ (.A1(_0598_),
    .A2(net470),
    .Y(_0264_),
    .B1(_0553_));
 sg13g2_o21ai_1 _2357_ (.B1(net560),
    .Y(_0554_),
    .A1(\bitserial_cipher.key_exp.shifter2[15] ),
    .A2(net461));
 sg13g2_a21oi_1 _2358_ (.A1(_0597_),
    .A2(net461),
    .Y(_0265_),
    .B1(_0554_));
 sg13g2_o21ai_1 _2359_ (.B1(net540),
    .Y(_0555_),
    .A1(net314),
    .A2(net462));
 sg13g2_a21oi_1 _2360_ (.A1(_0596_),
    .A2(net462),
    .Y(_0266_),
    .B1(_0555_));
 sg13g2_o21ai_1 _2361_ (.B1(net539),
    .Y(_0556_),
    .A1(\bitserial_cipher.key_exp.shifter2[17] ),
    .A2(net458));
 sg13g2_a21oi_1 _2362_ (.A1(_0595_),
    .A2(net457),
    .Y(_0267_),
    .B1(_0556_));
 sg13g2_o21ai_1 _2363_ (.B1(net539),
    .Y(_0557_),
    .A1(net663),
    .A2(net452));
 sg13g2_a21oi_1 _2364_ (.A1(_0594_),
    .A2(net452),
    .Y(_0268_),
    .B1(_0557_));
 sg13g2_o21ai_1 _2365_ (.B1(net535),
    .Y(_0558_),
    .A1(\bitserial_cipher.key_exp.shifter2[19] ),
    .A2(net451));
 sg13g2_a21oi_1 _2366_ (.A1(_0593_),
    .A2(net451),
    .Y(_0269_),
    .B1(_0558_));
 sg13g2_o21ai_1 _2367_ (.B1(net536),
    .Y(_0559_),
    .A1(net674),
    .A2(net450));
 sg13g2_a21oi_1 _2368_ (.A1(_0592_),
    .A2(net447),
    .Y(_0270_),
    .B1(_0559_));
 sg13g2_o21ai_1 _2369_ (.B1(net534),
    .Y(_0560_),
    .A1(\bitserial_cipher.key_exp.shifter2[21] ),
    .A2(net446));
 sg13g2_a21oi_1 _2370_ (.A1(_0591_),
    .A2(net446),
    .Y(_0271_),
    .B1(_0560_));
 sg13g2_o21ai_1 _2371_ (.B1(net534),
    .Y(_0561_),
    .A1(\bitserial_cipher.key_exp.shifter2[22] ),
    .A2(net446));
 sg13g2_a21oi_1 _2372_ (.A1(_0590_),
    .A2(net446),
    .Y(_0272_),
    .B1(_0561_));
 sg13g2_o21ai_1 _2373_ (.B1(net534),
    .Y(_0562_),
    .A1(net602),
    .A2(net445));
 sg13g2_a21oi_1 _2374_ (.A1(_0589_),
    .A2(net445),
    .Y(_0273_),
    .B1(_0562_));
 sg13g2_o21ai_1 _2375_ (.B1(net534),
    .Y(_0563_),
    .A1(\bitserial_cipher.key_exp.shifter2[24] ),
    .A2(net445));
 sg13g2_a21oi_1 _2376_ (.A1(_0588_),
    .A2(net445),
    .Y(_0274_),
    .B1(_0563_));
 sg13g2_o21ai_1 _2377_ (.B1(net534),
    .Y(_0564_),
    .A1(net587),
    .A2(net445));
 sg13g2_a21oi_1 _2378_ (.A1(_0587_),
    .A2(net445),
    .Y(_0275_),
    .B1(_0564_));
 sg13g2_o21ai_1 _2379_ (.B1(net534),
    .Y(_0565_),
    .A1(\bitserial_cipher.key_exp.shifter2[26] ),
    .A2(net445));
 sg13g2_a21oi_1 _2380_ (.A1(_0586_),
    .A2(net445),
    .Y(_0276_),
    .B1(_0565_));
 sg13g2_o21ai_1 _2381_ (.B1(net535),
    .Y(_0566_),
    .A1(net333),
    .A2(net447));
 sg13g2_a21oi_1 _2382_ (.A1(_0585_),
    .A2(net447),
    .Y(_0277_),
    .B1(_0566_));
 sg13g2_o21ai_1 _2383_ (.B1(net535),
    .Y(_0567_),
    .A1(\bitserial_cipher.key_exp.shifter2[28] ),
    .A2(net451));
 sg13g2_a21oi_1 _2384_ (.A1(_0584_),
    .A2(net451),
    .Y(_0278_),
    .B1(_0567_));
 sg13g2_o21ai_1 _2385_ (.B1(net535),
    .Y(_0568_),
    .A1(net727),
    .A2(net452));
 sg13g2_a21oi_1 _2386_ (.A1(_0583_),
    .A2(net452),
    .Y(_0279_),
    .B1(_0568_));
 sg13g2_o21ai_1 _2387_ (.B1(net539),
    .Y(_0569_),
    .A1(\bitserial_cipher.key_exp.shifter2[30] ),
    .A2(net457));
 sg13g2_a21oi_1 _2388_ (.A1(_0582_),
    .A2(net457),
    .Y(_0280_),
    .B1(_0569_));
 sg13g2_o21ai_1 _2389_ (.B1(net539),
    .Y(_0570_),
    .A1(net378),
    .A2(net457));
 sg13g2_a21oi_1 _2390_ (.A1(_0581_),
    .A2(net458),
    .Y(_0281_),
    .B1(_0570_));
 sg13g2_o21ai_1 _2391_ (.B1(net540),
    .Y(_0571_),
    .A1(\bitserial_cipher.key_exp.shifter2[32] ),
    .A2(net458));
 sg13g2_a21oi_1 _2392_ (.A1(_0580_),
    .A2(net462),
    .Y(_0282_),
    .B1(_0571_));
 sg13g2_o21ai_1 _2393_ (.B1(net540),
    .Y(_0572_),
    .A1(net368),
    .A2(net462));
 sg13g2_a21oi_1 _2394_ (.A1(_0579_),
    .A2(net462),
    .Y(_0283_),
    .B1(_0572_));
 sg13g2_o21ai_1 _2395_ (.B1(net540),
    .Y(_0573_),
    .A1(net608),
    .A2(net461));
 sg13g2_a21oi_1 _2396_ (.A1(_0578_),
    .A2(net461),
    .Y(_0284_),
    .B1(_0573_));
 sg13g2_o21ai_1 _2397_ (.B1(net540),
    .Y(_0574_),
    .A1(\bitserial_cipher.key_exp.shifter2[35] ),
    .A2(net461));
 sg13g2_a21oi_1 _2398_ (.A1(_0576_),
    .A2(net461),
    .Y(_0285_),
    .B1(_0574_));
 sg13g2_o21ai_1 _2399_ (.B1(net540),
    .Y(_0575_),
    .A1(net434),
    .A2(net461));
 sg13g2_a21oi_1 _2400_ (.A1(_0577_),
    .A2(net461),
    .Y(_0286_),
    .B1(_0575_));
 sg13g2_dfrbp_1 _2401_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net139),
    .D(net679),
    .Q_N(_1199_),
    .Q(\bitserial_cipher.key_exp.shifter2[37] ));
 sg13g2_dfrbp_1 _2402_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net131),
    .D(_0007_),
    .Q_N(_1198_),
    .Q(\bitserial_cipher.key_exp.shifter2[38] ));
 sg13g2_dfrbp_1 _2403_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net129),
    .D(net635),
    .Q_N(_1197_),
    .Q(\bitserial_cipher.key_exp.shifter2[39] ));
 sg13g2_dfrbp_1 _2404_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net127),
    .D(net405),
    .Q_N(_1196_),
    .Q(\bitserial_cipher.key_exp.shifter2[40] ));
 sg13g2_dfrbp_1 _2405_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net125),
    .D(_0010_),
    .Q_N(_1195_),
    .Q(\bitserial_cipher.key_exp.shifter2[41] ));
 sg13g2_dfrbp_1 _2406_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net123),
    .D(_0011_),
    .Q_N(_1194_),
    .Q(\bitserial_cipher.key_exp.shifter2[42] ));
 sg13g2_dfrbp_1 _2407_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net121),
    .D(_0012_),
    .Q_N(_1193_),
    .Q(\bitserial_cipher.key_exp.shifter2[43] ));
 sg13g2_dfrbp_1 _2408_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net119),
    .D(net649),
    .Q_N(_1192_),
    .Q(\bitserial_cipher.key_exp.shifter2[44] ));
 sg13g2_dfrbp_1 _2409_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net117),
    .D(_0014_),
    .Q_N(_1191_),
    .Q(\bitserial_cipher.key_exp.shifter2[45] ));
 sg13g2_dfrbp_1 _2410_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net115),
    .D(_0015_),
    .Q_N(_1190_),
    .Q(\bitserial_cipher.key_exp.shifter2[46] ));
 sg13g2_dfrbp_1 _2411_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net113),
    .D(net653),
    .Q_N(_1189_),
    .Q(\bitserial_cipher.key_exp.shifter2[47] ));
 sg13g2_dfrbp_1 _2412_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net111),
    .D(net399),
    .Q_N(_1188_),
    .Q(\bitserial_cipher.key_exp.shifter2[48] ));
 sg13g2_dfrbp_1 _2413_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net109),
    .D(_0018_),
    .Q_N(_1187_),
    .Q(\bitserial_cipher.key_exp.shifter2[49] ));
 sg13g2_dfrbp_1 _2414_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net107),
    .D(net668),
    .Q_N(_1186_),
    .Q(\bitserial_cipher.key_exp.shifter2[50] ));
 sg13g2_dfrbp_1 _2415_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net105),
    .D(_0020_),
    .Q_N(_1185_),
    .Q(\bitserial_cipher.key_exp.shifter2[51] ));
 sg13g2_dfrbp_1 _2416_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net103),
    .D(net586),
    .Q_N(_1184_),
    .Q(\bitserial_cipher.key_exp.shifter2[52] ));
 sg13g2_dfrbp_1 _2417_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net101),
    .D(_0022_),
    .Q_N(_1183_),
    .Q(\bitserial_cipher.key_exp.shifter2[53] ));
 sg13g2_dfrbp_1 _2418_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net99),
    .D(_0023_),
    .Q_N(_1182_),
    .Q(\bitserial_cipher.key_exp.shifter2[54] ));
 sg13g2_dfrbp_1 _2419_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net97),
    .D(net582),
    .Q_N(_1181_),
    .Q(\bitserial_cipher.key_exp.shifter2[55] ));
 sg13g2_dfrbp_1 _2420_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net95),
    .D(_0025_),
    .Q_N(_1180_),
    .Q(\bitserial_cipher.key_exp.shifter2[56] ));
 sg13g2_dfrbp_1 _2421_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net93),
    .D(_0026_),
    .Q_N(_1179_),
    .Q(\bitserial_cipher.key_exp.shifter2[57] ));
 sg13g2_dfrbp_1 _2422_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net91),
    .D(net614),
    .Q_N(_1178_),
    .Q(\bitserial_cipher.key_exp.shifter2[58] ));
 sg13g2_dfrbp_1 _2423_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net89),
    .D(net411),
    .Q_N(_1177_),
    .Q(\bitserial_cipher.key_exp.shifter2[59] ));
 sg13g2_dfrbp_1 _2424_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net87),
    .D(_0029_),
    .Q_N(_1176_),
    .Q(\bitserial_cipher.key_exp.shifter2[60] ));
 sg13g2_dfrbp_1 _2425_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net85),
    .D(_0030_),
    .Q_N(_1175_),
    .Q(\bitserial_cipher.key_exp.shifter2[61] ));
 sg13g2_dfrbp_1 _2426_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net83),
    .D(net373),
    .Q_N(_1174_),
    .Q(\bitserial_cipher.key_exp.shifter2[62] ));
 sg13g2_dfrbp_1 _2427_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net81),
    .D(_0032_),
    .Q_N(_1173_),
    .Q(\bitserial_cipher.key_exp.shifter2[63] ));
 sg13g2_dfrbp_1 _2428_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net79),
    .D(net673),
    .Q_N(_1172_),
    .Q(\bitserial_cipher.key_exp.shift_out1 ));
 sg13g2_dfrbp_1 _2429_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net77),
    .D(net344),
    .Q_N(_1171_),
    .Q(\bitserial_cipher.key_exp.shifter1[1] ));
 sg13g2_dfrbp_1 _2430_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net75),
    .D(_0035_),
    .Q_N(_1170_),
    .Q(\bitserial_cipher.key_exp.shifter1[2] ));
 sg13g2_dfrbp_1 _2431_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net73),
    .D(_0036_),
    .Q_N(_1169_),
    .Q(\bitserial_cipher.key_exp.shifter1[3] ));
 sg13g2_dfrbp_1 _2432_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net71),
    .D(net749),
    .Q_N(_1168_),
    .Q(\bitserial_cipher.key_exp.shifter1[4] ));
 sg13g2_dfrbp_1 _2433_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net69),
    .D(_0038_),
    .Q_N(_1167_),
    .Q(\bitserial_cipher.key_exp.shifter1[5] ));
 sg13g2_dfrbp_1 _2434_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net67),
    .D(net644),
    .Q_N(_1166_),
    .Q(\bitserial_cipher.key_exp.shifter1[6] ));
 sg13g2_dfrbp_1 _2435_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net65),
    .D(net622),
    .Q_N(_1165_),
    .Q(\bitserial_cipher.key_exp.shifter1[7] ));
 sg13g2_dfrbp_1 _2436_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net63),
    .D(_0041_),
    .Q_N(_1164_),
    .Q(\bitserial_cipher.key_exp.shifter1[8] ));
 sg13g2_dfrbp_1 _2437_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net61),
    .D(net651),
    .Q_N(_1163_),
    .Q(\bitserial_cipher.key_exp.shifter1[9] ));
 sg13g2_dfrbp_1 _2438_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net59),
    .D(net616),
    .Q_N(_1162_),
    .Q(\bitserial_cipher.key_exp.shifter1[10] ));
 sg13g2_dfrbp_1 _2439_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net57),
    .D(_0044_),
    .Q_N(_1161_),
    .Q(\bitserial_cipher.key_exp.shifter1[11] ));
 sg13g2_dfrbp_1 _2440_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net55),
    .D(net391),
    .Q_N(_1160_),
    .Q(\bitserial_cipher.key_exp.shifter1[12] ));
 sg13g2_dfrbp_1 _2441_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net53),
    .D(_0046_),
    .Q_N(_1159_),
    .Q(\bitserial_cipher.key_exp.shifter1[13] ));
 sg13g2_dfrbp_1 _2442_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net51),
    .D(net328),
    .Q_N(_1158_),
    .Q(\bitserial_cipher.key_exp.shifter1[14] ));
 sg13g2_dfrbp_1 _2443_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net49),
    .D(_0048_),
    .Q_N(_1157_),
    .Q(\bitserial_cipher.key_exp.shifter1[15] ));
 sg13g2_dfrbp_1 _2444_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net47),
    .D(net638),
    .Q_N(_1156_),
    .Q(\bitserial_cipher.key_exp.shifter1[16] ));
 sg13g2_dfrbp_1 _2445_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net45),
    .D(net596),
    .Q_N(_1155_),
    .Q(\bitserial_cipher.key_exp.shifter1[17] ));
 sg13g2_dfrbp_1 _2446_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net43),
    .D(net332),
    .Q_N(_1154_),
    .Q(\bitserial_cipher.key_exp.shifter1[18] ));
 sg13g2_dfrbp_1 _2447_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net41),
    .D(_0052_),
    .Q_N(_1153_),
    .Q(\bitserial_cipher.key_exp.shifter1[19] ));
 sg13g2_dfrbp_1 _2448_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net39),
    .D(_0053_),
    .Q_N(_1152_),
    .Q(\bitserial_cipher.key_exp.shifter1[20] ));
 sg13g2_dfrbp_1 _2449_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net37),
    .D(_0054_),
    .Q_N(_1151_),
    .Q(\bitserial_cipher.key_exp.shifter1[21] ));
 sg13g2_dfrbp_1 _2450_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net35),
    .D(_0055_),
    .Q_N(_1150_),
    .Q(\bitserial_cipher.key_exp.shifter1[22] ));
 sg13g2_dfrbp_1 _2451_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net33),
    .D(net594),
    .Q_N(_1149_),
    .Q(\bitserial_cipher.key_exp.shifter1[23] ));
 sg13g2_dfrbp_1 _2452_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net31),
    .D(_0057_),
    .Q_N(_1148_),
    .Q(\bitserial_cipher.key_exp.shifter1[24] ));
 sg13g2_dfrbp_1 _2453_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net29),
    .D(_0058_),
    .Q_N(_1147_),
    .Q(\bitserial_cipher.key_exp.shifter1[25] ));
 sg13g2_dfrbp_1 _2454_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net27),
    .D(net319),
    .Q_N(_1146_),
    .Q(\bitserial_cipher.key_exp.shifter1[26] ));
 sg13g2_dfrbp_1 _2455_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net25),
    .D(_0060_),
    .Q_N(_1145_),
    .Q(\bitserial_cipher.key_exp.shifter1[27] ));
 sg13g2_dfrbp_1 _2456_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net304),
    .D(_0061_),
    .Q_N(_1144_),
    .Q(\bitserial_cipher.key_exp.shifter1[28] ));
 sg13g2_dfrbp_1 _2457_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net302),
    .D(net687),
    .Q_N(_1143_),
    .Q(\bitserial_cipher.key_exp.shifter1[29] ));
 sg13g2_dfrbp_1 _2458_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net300),
    .D(_0063_),
    .Q_N(_1142_),
    .Q(\bitserial_cipher.key_exp.shifter1[30] ));
 sg13g2_dfrbp_1 _2459_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net298),
    .D(_0064_),
    .Q_N(_1141_),
    .Q(\bitserial_cipher.key_exp.shifter1[31] ));
 sg13g2_dfrbp_1 _2460_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net296),
    .D(_0065_),
    .Q_N(_1140_),
    .Q(\bitserial_cipher.key_exp.shifter1[32] ));
 sg13g2_dfrbp_1 _2461_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net294),
    .D(net361),
    .Q_N(_1139_),
    .Q(\bitserial_cipher.key_exp.shifter1[33] ));
 sg13g2_dfrbp_1 _2462_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net292),
    .D(_0067_),
    .Q_N(_1138_),
    .Q(\bitserial_cipher.key_exp.shifter1[34] ));
 sg13g2_dfrbp_1 _2463_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net290),
    .D(_0068_),
    .Q_N(_1137_),
    .Q(\bitserial_cipher.key_exp.shifter1[35] ));
 sg13g2_dfrbp_1 _2464_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net288),
    .D(net322),
    .Q_N(_1136_),
    .Q(\bitserial_cipher.key_exp.shifter1[36] ));
 sg13g2_dfrbp_1 _2465_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net286),
    .D(_0070_),
    .Q_N(_1135_),
    .Q(\bitserial_cipher.key_exp.shifter1[37] ));
 sg13g2_dfrbp_1 _2466_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net284),
    .D(_0071_),
    .Q_N(_1134_),
    .Q(\bitserial_cipher.key_exp.shifter1[38] ));
 sg13g2_dfrbp_1 _2467_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net282),
    .D(_0072_),
    .Q_N(_1133_),
    .Q(\bitserial_cipher.key_exp.shifter1[39] ));
 sg13g2_dfrbp_1 _2468_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net280),
    .D(net371),
    .Q_N(_1132_),
    .Q(\bitserial_cipher.key_exp.shifter1[40] ));
 sg13g2_dfrbp_1 _2469_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net278),
    .D(_0074_),
    .Q_N(_1131_),
    .Q(\bitserial_cipher.key_exp.shifter1[41] ));
 sg13g2_dfrbp_1 _2470_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net276),
    .D(_0075_),
    .Q_N(_1130_),
    .Q(\bitserial_cipher.key_exp.shifter1[42] ));
 sg13g2_dfrbp_1 _2471_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net274),
    .D(net403),
    .Q_N(_1129_),
    .Q(\bitserial_cipher.key_exp.shifter1[43] ));
 sg13g2_dfrbp_1 _2472_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net272),
    .D(_0077_),
    .Q_N(_1128_),
    .Q(\bitserial_cipher.key_exp.shifter1[44] ));
 sg13g2_dfrbp_1 _2473_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net270),
    .D(net590),
    .Q_N(_1127_),
    .Q(\bitserial_cipher.key_exp.shifter1[45] ));
 sg13g2_dfrbp_1 _2474_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net268),
    .D(_0079_),
    .Q_N(_1126_),
    .Q(\bitserial_cipher.key_exp.shifter1[46] ));
 sg13g2_dfrbp_1 _2475_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net266),
    .D(_0080_),
    .Q_N(_1125_),
    .Q(\bitserial_cipher.key_exp.shifter1[47] ));
 sg13g2_dfrbp_1 _2476_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net264),
    .D(net428),
    .Q_N(_1124_),
    .Q(\bitserial_cipher.key_exp.shifter1[48] ));
 sg13g2_dfrbp_1 _2477_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net262),
    .D(net383),
    .Q_N(_1123_),
    .Q(\bitserial_cipher.key_exp.shifter1[49] ));
 sg13g2_dfrbp_1 _2478_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net260),
    .D(_0083_),
    .Q_N(_1122_),
    .Q(\bitserial_cipher.key_exp.shifter1[50] ));
 sg13g2_dfrbp_1 _2479_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net258),
    .D(_0084_),
    .Q_N(_1121_),
    .Q(\bitserial_cipher.key_exp.shifter1[51] ));
 sg13g2_dfrbp_1 _2480_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net256),
    .D(net599),
    .Q_N(_1120_),
    .Q(\bitserial_cipher.key_exp.shifter1[52] ));
 sg13g2_dfrbp_1 _2481_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net254),
    .D(_0086_),
    .Q_N(_1119_),
    .Q(\bitserial_cipher.key_exp.shifter1[53] ));
 sg13g2_dfrbp_1 _2482_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net252),
    .D(net431),
    .Q_N(_1118_),
    .Q(\bitserial_cipher.key_exp.shifter1[54] ));
 sg13g2_dfrbp_1 _2483_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net250),
    .D(_0088_),
    .Q_N(_1117_),
    .Q(\bitserial_cipher.key_exp.shifter1[55] ));
 sg13g2_dfrbp_1 _2484_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net248),
    .D(net358),
    .Q_N(_1116_),
    .Q(\bitserial_cipher.key_exp.shifter1[56] ));
 sg13g2_dfrbp_1 _2485_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net246),
    .D(_0090_),
    .Q_N(_1115_),
    .Q(\bitserial_cipher.key_exp.shifter1[57] ));
 sg13g2_dfrbp_1 _2486_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net244),
    .D(_0091_),
    .Q_N(_1114_),
    .Q(\bitserial_cipher.key_exp.shifter1[58] ));
 sg13g2_dfrbp_1 _2487_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net242),
    .D(_0092_),
    .Q_N(_1113_),
    .Q(\bitserial_cipher.key_exp.shifter1[59] ));
 sg13g2_dfrbp_1 _2488_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net240),
    .D(net642),
    .Q_N(_1112_),
    .Q(\bitserial_cipher.datapath.fifo_ff57 ));
 sg13g2_dfrbp_1 _2489_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net238),
    .D(net389),
    .Q_N(_1111_),
    .Q(\bitserial_cipher.datapath.fifo_ff58 ));
 sg13g2_dfrbp_1 _2490_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net236),
    .D(net338),
    .Q_N(_1110_),
    .Q(\bitserial_cipher.datapath.fifo_ff59 ));
 sg13g2_dfrbp_1 _2491_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net234),
    .D(_0096_),
    .Q_N(_1109_),
    .Q(\bitserial_cipher.datapath.fifo_ff60 ));
 sg13g2_dfrbp_1 _2492_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net232),
    .D(net670),
    .Q_N(_1108_),
    .Q(\bitserial_cipher.datapath.shift_in2 ));
 sg13g2_dfrbp_1 _2493_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net230),
    .D(_0098_),
    .Q_N(_1107_),
    .Q(\bitserial_cipher.datapath.shifter1[1] ));
 sg13g2_dfrbp_1 _2494_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net228),
    .D(_0099_),
    .Q_N(_1106_),
    .Q(\bitserial_cipher.datapath.shifter1[2] ));
 sg13g2_dfrbp_1 _2495_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net226),
    .D(net811),
    .Q_N(_1105_),
    .Q(\bitserial_cipher.datapath.shifter1[3] ));
 sg13g2_dfrbp_1 _2496_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net224),
    .D(net719),
    .Q_N(_1104_),
    .Q(\bitserial_cipher.datapath.shifter1[4] ));
 sg13g2_dfrbp_1 _2497_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net222),
    .D(net607),
    .Q_N(_1103_),
    .Q(\bitserial_cipher.datapath.shifter1[5] ));
 sg13g2_dfrbp_1 _2498_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net220),
    .D(net377),
    .Q_N(_1102_),
    .Q(\bitserial_cipher.datapath.shifter1[6] ));
 sg13g2_dfrbp_1 _2499_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net218),
    .D(_0104_),
    .Q_N(_1101_),
    .Q(\bitserial_cipher.datapath.shifter1[7] ));
 sg13g2_dfrbp_1 _2500_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net216),
    .D(net363),
    .Q_N(_1100_),
    .Q(\bitserial_cipher.datapath.shifter1[8] ));
 sg13g2_dfrbp_1 _2501_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net214),
    .D(_0106_),
    .Q_N(_1099_),
    .Q(\bitserial_cipher.datapath.shifter1[9] ));
 sg13g2_dfrbp_1 _2502_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net212),
    .D(_0107_),
    .Q_N(_1098_),
    .Q(\bitserial_cipher.datapath.shifter1[10] ));
 sg13g2_dfrbp_1 _2503_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net210),
    .D(net631),
    .Q_N(_1097_),
    .Q(\bitserial_cipher.datapath.shifter1[11] ));
 sg13g2_dfrbp_1 _2504_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net208),
    .D(net605),
    .Q_N(_1096_),
    .Q(\bitserial_cipher.datapath.shifter1[12] ));
 sg13g2_dfrbp_1 _2505_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net206),
    .D(_0110_),
    .Q_N(_1095_),
    .Q(\bitserial_cipher.datapath.shifter1[13] ));
 sg13g2_dfrbp_1 _2506_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net204),
    .D(_0111_),
    .Q_N(_1094_),
    .Q(\bitserial_cipher.datapath.shifter1[14] ));
 sg13g2_dfrbp_1 _2507_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net202),
    .D(net659),
    .Q_N(_1093_),
    .Q(\bitserial_cipher.datapath.shifter1[15] ));
 sg13g2_dfrbp_1 _2508_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net200),
    .D(_0113_),
    .Q_N(_1092_),
    .Q(\bitserial_cipher.datapath.shifter1[16] ));
 sg13g2_dfrbp_1 _2509_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net198),
    .D(net317),
    .Q_N(_1091_),
    .Q(\bitserial_cipher.datapath.shifter1[17] ));
 sg13g2_dfrbp_1 _2510_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net196),
    .D(_0115_),
    .Q_N(_1090_),
    .Q(\bitserial_cipher.datapath.shifter1[18] ));
 sg13g2_dfrbp_1 _2511_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net194),
    .D(net413),
    .Q_N(_1089_),
    .Q(\bitserial_cipher.datapath.shifter1[19] ));
 sg13g2_dfrbp_1 _2512_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net192),
    .D(_0117_),
    .Q_N(_1088_),
    .Q(\bitserial_cipher.datapath.shifter1[20] ));
 sg13g2_dfrbp_1 _2513_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net190),
    .D(net683),
    .Q_N(_1087_),
    .Q(\bitserial_cipher.datapath.shifter1[21] ));
 sg13g2_dfrbp_1 _2514_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net188),
    .D(_0119_),
    .Q_N(_1086_),
    .Q(\bitserial_cipher.datapath.shifter1[22] ));
 sg13g2_dfrbp_1 _2515_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net186),
    .D(net342),
    .Q_N(_1085_),
    .Q(\bitserial_cipher.datapath.shifter1[23] ));
 sg13g2_dfrbp_1 _2516_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net184),
    .D(_0121_),
    .Q_N(_1084_),
    .Q(\bitserial_cipher.datapath.shifter1[24] ));
 sg13g2_dfrbp_1 _2517_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net182),
    .D(net699),
    .Q_N(_1083_),
    .Q(\bitserial_cipher.datapath.shifter1[25] ));
 sg13g2_dfrbp_1 _2518_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net180),
    .D(net433),
    .Q_N(_1082_),
    .Q(\bitserial_cipher.datapath.shifter1[26] ));
 sg13g2_dfrbp_1 _2519_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net178),
    .D(_0124_),
    .Q_N(_1081_),
    .Q(\bitserial_cipher.datapath.shifter1[27] ));
 sg13g2_dfrbp_1 _2520_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net176),
    .D(net354),
    .Q_N(_1080_),
    .Q(\bitserial_cipher.datapath.shifter1[28] ));
 sg13g2_dfrbp_1 _2521_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net174),
    .D(_0126_),
    .Q_N(_1079_),
    .Q(\bitserial_cipher.datapath.shifter1[29] ));
 sg13g2_dfrbp_1 _2522_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net172),
    .D(_0127_),
    .Q_N(_1078_),
    .Q(\bitserial_cipher.datapath.shifter1[30] ));
 sg13g2_dfrbp_1 _2523_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net170),
    .D(_0128_),
    .Q_N(_1077_),
    .Q(\bitserial_cipher.datapath.shifter1[31] ));
 sg13g2_dfrbp_1 _2524_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net168),
    .D(net592),
    .Q_N(_1076_),
    .Q(\bitserial_cipher.datapath.shifter1[32] ));
 sg13g2_dfrbp_1 _2525_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net166),
    .D(_0130_),
    .Q_N(_1075_),
    .Q(\bitserial_cipher.datapath.shifter1[33] ));
 sg13g2_dfrbp_1 _2526_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net164),
    .D(_0131_),
    .Q_N(_1074_),
    .Q(\bitserial_cipher.datapath.shifter1[34] ));
 sg13g2_dfrbp_1 _2527_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net162),
    .D(_0132_),
    .Q_N(_1073_),
    .Q(\bitserial_cipher.datapath.shifter1[35] ));
 sg13g2_dfrbp_1 _2528_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net160),
    .D(net796),
    .Q_N(_1072_),
    .Q(\bitserial_cipher.datapath.shifter1[36] ));
 sg13g2_dfrbp_1 _2529_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net158),
    .D(net781),
    .Q_N(_1071_),
    .Q(\bitserial_cipher.datapath.shifter1[37] ));
 sg13g2_dfrbp_1 _2530_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net156),
    .D(net419),
    .Q_N(_1070_),
    .Q(\bitserial_cipher.datapath.shifter1[38] ));
 sg13g2_dfrbp_1 _2531_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net154),
    .D(net326),
    .Q_N(_1069_),
    .Q(\bitserial_cipher.datapath.shifter1[39] ));
 sg13g2_dfrbp_1 _2532_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net152),
    .D(_0137_),
    .Q_N(_1068_),
    .Q(\bitserial_cipher.datapath.shifter1[40] ));
 sg13g2_dfrbp_1 _2533_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net150),
    .D(_0138_),
    .Q_N(_1067_),
    .Q(\bitserial_cipher.datapath.shifter1[41] ));
 sg13g2_dfrbp_1 _2534_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net148),
    .D(net350),
    .Q_N(_1066_),
    .Q(\bitserial_cipher.datapath.shifter1[42] ));
 sg13g2_dfrbp_1 _2535_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net146),
    .D(_0140_),
    .Q_N(_1065_),
    .Q(\bitserial_cipher.datapath.shifter1[43] ));
 sg13g2_dfrbp_1 _2536_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net144),
    .D(_0141_),
    .Q_N(_1064_),
    .Q(\bitserial_cipher.datapath.shifter1[44] ));
 sg13g2_dfrbp_1 _2537_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net142),
    .D(net791),
    .Q_N(_1063_),
    .Q(\bitserial_cipher.datapath.shifter1[45] ));
 sg13g2_dfrbp_1 _2538_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net140),
    .D(net735),
    .Q_N(_1062_),
    .Q(\bitserial_cipher.datapath.shifter1[46] ));
 sg13g2_dfrbp_1 _2539_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net138),
    .D(net694),
    .Q_N(_1061_),
    .Q(\bitserial_cipher.datapath.shifter1[47] ));
 sg13g2_dfrbp_1 _2540_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net136),
    .D(net619),
    .Q_N(_1060_),
    .Q(\bitserial_cipher.datapath.shifter1[48] ));
 sg13g2_dfrbp_1 _2541_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net134),
    .D(net397),
    .Q_N(_1059_),
    .Q(\bitserial_cipher.datapath.shifter1[49] ));
 sg13g2_dfrbp_1 _2542_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net132),
    .D(net375),
    .Q_N(_1058_),
    .Q(\bitserial_cipher.datapath.shifter1[50] ));
 sg13g2_dfrbp_1 _2543_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net128),
    .D(_0148_),
    .Q_N(_1057_),
    .Q(\bitserial_cipher.datapath.shifter1[51] ));
 sg13g2_dfrbp_1 _2544_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net124),
    .D(net324),
    .Q_N(_1056_),
    .Q(\bitserial_cipher.datapath.shifter1[52] ));
 sg13g2_dfrbp_1 _2545_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net120),
    .D(_0150_),
    .Q_N(_1055_),
    .Q(\bitserial_cipher.datapath.shifter1[53] ));
 sg13g2_dfrbp_1 _2546_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net116),
    .D(net709),
    .Q_N(_1054_),
    .Q(\bitserial_cipher.datapath.shifter1[54] ));
 sg13g2_dfrbp_1 _2547_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net112),
    .D(_0152_),
    .Q_N(_1053_),
    .Q(\bitserial_cipher.datapath.shifter1[55] ));
 sg13g2_dfrbp_1 _2548_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net108),
    .D(net580),
    .Q_N(_1052_),
    .Q(\bitserial_cipher.cipher_data ));
 sg13g2_dfrbp_1 _2549_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net104),
    .D(_0154_),
    .Q_N(_1051_),
    .Q(\bitserial_cipher.datapath.shifter2[1] ));
 sg13g2_dfrbp_1 _2550_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net100),
    .D(net421),
    .Q_N(_1050_),
    .Q(\bitserial_cipher.datapath.shifter2[2] ));
 sg13g2_dfrbp_1 _2551_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net96),
    .D(_0156_),
    .Q_N(_1049_),
    .Q(\bitserial_cipher.datapath.shifter2[3] ));
 sg13g2_dfrbp_1 _2552_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net92),
    .D(net401),
    .Q_N(_1048_),
    .Q(\bitserial_cipher.datapath.shifter2[4] ));
 sg13g2_dfrbp_1 _2553_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net88),
    .D(net367),
    .Q_N(_1047_),
    .Q(\bitserial_cipher.datapath.shifter2[5] ));
 sg13g2_dfrbp_1 _2554_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net84),
    .D(_0159_),
    .Q_N(_1046_),
    .Q(\bitserial_cipher.datapath.shifter2[6] ));
 sg13g2_dfrbp_1 _2555_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net80),
    .D(_0160_),
    .Q_N(_1045_),
    .Q(\bitserial_cipher.datapath.shifter2[7] ));
 sg13g2_dfrbp_1 _2556_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net76),
    .D(_0161_),
    .Q_N(_1044_),
    .Q(\bitserial_cipher.datapath.shifter2[8] ));
 sg13g2_dfrbp_1 _2557_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net72),
    .D(net696),
    .Q_N(_1043_),
    .Q(\bitserial_cipher.datapath.shifter2[9] ));
 sg13g2_dfrbp_1 _2558_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net68),
    .D(net385),
    .Q_N(_1042_),
    .Q(\bitserial_cipher.datapath.shifter2[10] ));
 sg13g2_dfrbp_1 _2559_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net64),
    .D(_0164_),
    .Q_N(_1041_),
    .Q(\bitserial_cipher.datapath.shifter2[11] ));
 sg13g2_dfrbp_1 _2560_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net60),
    .D(net677),
    .Q_N(_1040_),
    .Q(\bitserial_cipher.datapath.shifter2[12] ));
 sg13g2_dfrbp_1 _2561_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net56),
    .D(_0166_),
    .Q_N(_1039_),
    .Q(\bitserial_cipher.datapath.shifter2[13] ));
 sg13g2_dfrbp_1 _2562_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net52),
    .D(net423),
    .Q_N(_1038_),
    .Q(\bitserial_cipher.datapath.shifter2[14] ));
 sg13g2_dfrbp_1 _2563_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net48),
    .D(_0168_),
    .Q_N(_1037_),
    .Q(\bitserial_cipher.datapath.shifter2[15] ));
 sg13g2_dfrbp_1 _2564_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net44),
    .D(net352),
    .Q_N(_1036_),
    .Q(\bitserial_cipher.datapath.shifter2[16] ));
 sg13g2_dfrbp_1 _2565_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net40),
    .D(_0170_),
    .Q_N(_1035_),
    .Q(\bitserial_cipher.datapath.shifter2[17] ));
 sg13g2_dfrbp_1 _2566_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net36),
    .D(net624),
    .Q_N(_1034_),
    .Q(\bitserial_cipher.datapath.shifter2[18] ));
 sg13g2_dfrbp_1 _2567_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net32),
    .D(_0172_),
    .Q_N(_1033_),
    .Q(\bitserial_cipher.datapath.shifter2[19] ));
 sg13g2_dfrbp_1 _2568_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net28),
    .D(net409),
    .Q_N(_1032_),
    .Q(\bitserial_cipher.datapath.shifter2[20] ));
 sg13g2_dfrbp_1 _2569_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net24),
    .D(net381),
    .Q_N(_1031_),
    .Q(\bitserial_cipher.datapath.shifter2[21] ));
 sg13g2_dfrbp_1 _2570_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net301),
    .D(_0175_),
    .Q_N(_1030_),
    .Q(\bitserial_cipher.datapath.shifter2[22] ));
 sg13g2_dfrbp_1 _2571_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net297),
    .D(net707),
    .Q_N(_1029_),
    .Q(\bitserial_cipher.datapath.shifter2[23] ));
 sg13g2_dfrbp_1 _2572_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net293),
    .D(net393),
    .Q_N(_1028_),
    .Q(\bitserial_cipher.datapath.shifter2[24] ));
 sg13g2_dfrbp_1 _2573_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net289),
    .D(_0178_),
    .Q_N(_1027_),
    .Q(\bitserial_cipher.datapath.shifter2[25] ));
 sg13g2_dfrbp_1 _2574_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net285),
    .D(_0179_),
    .Q_N(_1026_),
    .Q(\bitserial_cipher.datapath.shifter2[26] ));
 sg13g2_dfrbp_1 _2575_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net281),
    .D(net415),
    .Q_N(_1025_),
    .Q(\bitserial_cipher.datapath.shifter2[27] ));
 sg13g2_dfrbp_1 _2576_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net277),
    .D(_0181_),
    .Q_N(_1024_),
    .Q(\bitserial_cipher.datapath.shifter2[28] ));
 sg13g2_dfrbp_1 _2577_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net273),
    .D(_0182_),
    .Q_N(_1023_),
    .Q(\bitserial_cipher.datapath.shifter2[29] ));
 sg13g2_dfrbp_1 _2578_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net269),
    .D(net657),
    .Q_N(_1022_),
    .Q(\bitserial_cipher.datapath.shifter2[30] ));
 sg13g2_dfrbp_1 _2579_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net265),
    .D(_0184_),
    .Q_N(_1021_),
    .Q(\bitserial_cipher.datapath.shifter2[31] ));
 sg13g2_dfrbp_1 _2580_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net261),
    .D(net426),
    .Q_N(_1020_),
    .Q(\bitserial_cipher.datapath.shifter2[32] ));
 sg13g2_dfrbp_1 _2581_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net257),
    .D(net365),
    .Q_N(_1019_),
    .Q(\bitserial_cipher.datapath.shifter2[33] ));
 sg13g2_dfrbp_1 _2582_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net253),
    .D(_0187_),
    .Q_N(_1018_),
    .Q(\bitserial_cipher.datapath.shifter2[34] ));
 sg13g2_dfrbp_1 _2583_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net249),
    .D(_0188_),
    .Q_N(_1017_),
    .Q(\bitserial_cipher.datapath.shifter2[35] ));
 sg13g2_dfrbp_1 _2584_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net245),
    .D(net716),
    .Q_N(_1016_),
    .Q(\bitserial_cipher.datapath.shifter2[36] ));
 sg13g2_dfrbp_1 _2585_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net241),
    .D(_0190_),
    .Q_N(_1015_),
    .Q(\bitserial_cipher.datapath.shifter2[37] ));
 sg13g2_dfrbp_1 _2586_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net237),
    .D(net730),
    .Q_N(_1014_),
    .Q(\bitserial_cipher.datapath.shifter2[38] ));
 sg13g2_dfrbp_1 _2587_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net233),
    .D(_0192_),
    .Q_N(_1013_),
    .Q(\bitserial_cipher.datapath.shifter2[39] ));
 sg13g2_dfrbp_1 _2588_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net229),
    .D(net407),
    .Q_N(_1012_),
    .Q(\bitserial_cipher.datapath.shifter2[40] ));
 sg13g2_dfrbp_1 _2589_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net225),
    .D(net340),
    .Q_N(_1011_),
    .Q(\bitserial_cipher.datapath.shifter2[41] ));
 sg13g2_dfrbp_1 _2590_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net221),
    .D(_0195_),
    .Q_N(_1010_),
    .Q(\bitserial_cipher.datapath.shifter2[42] ));
 sg13g2_dfrbp_1 _2591_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net217),
    .D(net346),
    .Q_N(_1009_),
    .Q(\bitserial_cipher.datapath.shifter2[43] ));
 sg13g2_dfrbp_1 _2592_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net213),
    .D(_0197_),
    .Q_N(_1008_),
    .Q(\bitserial_cipher.datapath.shifter2[44] ));
 sg13g2_dfrbp_1 _2593_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net209),
    .D(_0198_),
    .Q_N(_1007_),
    .Q(\bitserial_cipher.datapath.shifter2[45] ));
 sg13g2_dfrbp_1 _2594_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net205),
    .D(net777),
    .Q_N(_1006_),
    .Q(\bitserial_cipher.datapath.shifter2[46] ));
 sg13g2_dfrbp_1 _2595_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net201),
    .D(net313),
    .Q_N(_1005_),
    .Q(\bitserial_cipher.datapath.shifter2[47] ));
 sg13g2_dfrbp_1 _2596_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net197),
    .D(_0201_),
    .Q_N(_1004_),
    .Q(\bitserial_cipher.datapath.shifter2[48] ));
 sg13g2_dfrbp_1 _2597_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net193),
    .D(_0202_),
    .Q_N(_1003_),
    .Q(\bitserial_cipher.datapath.shifter2[49] ));
 sg13g2_dfrbp_1 _2598_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net189),
    .D(net765),
    .Q_N(_1002_),
    .Q(\bitserial_cipher.datapath.shifter2[50] ));
 sg13g2_dfrbp_1 _2599_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net185),
    .D(net584),
    .Q_N(_1001_),
    .Q(\bitserial_cipher.datapath.shifter2[51] ));
 sg13g2_dfrbp_1 _2600_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net181),
    .D(net330),
    .Q_N(_1000_),
    .Q(\bitserial_cipher.datapath.shifter2[52] ));
 sg13g2_dfrbp_1 _2601_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net177),
    .D(_0206_),
    .Q_N(_0999_),
    .Q(\bitserial_cipher.datapath.shifter2[53] ));
 sg13g2_dfrbp_1 _2602_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net173),
    .D(_0207_),
    .Q_N(_0998_),
    .Q(\bitserial_cipher.datapath.shifter2[54] ));
 sg13g2_dfrbp_1 _2603_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net169),
    .D(net395),
    .Q_N(_0997_),
    .Q(\bitserial_cipher.datapath.shifter2[55] ));
 sg13g2_dfrbp_1 _2604_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net165),
    .D(_0209_),
    .Q_N(_0996_),
    .Q(\bitserial_cipher.datapath.shifter2[56] ));
 sg13g2_dfrbp_1 _2605_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net161),
    .D(net681),
    .Q_N(_0995_),
    .Q(\bitserial_cipher.datapath.shifter2[57] ));
 sg13g2_dfrbp_1 _2606_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net157),
    .D(net348),
    .Q_N(_0994_),
    .Q(\bitserial_cipher.datapath.shifter2[58] ));
 sg13g2_dfrbp_1 _2607_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net153),
    .D(_0212_),
    .Q_N(_0993_),
    .Q(\bitserial_cipher.datapath.shifter2[59] ));
 sg13g2_dfrbp_1 _2608_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net149),
    .D(net762),
    .Q_N(_0992_),
    .Q(\bitserial_cipher.datapath.shifter2[60] ));
 sg13g2_dfrbp_1 _2609_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net145),
    .D(net417),
    .Q_N(_0991_),
    .Q(\bitserial_cipher.datapath.shifter2[61] ));
 sg13g2_dfrbp_1 _2610_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net141),
    .D(net356),
    .Q_N(_0990_),
    .Q(\bitserial_cipher.datapath.shifter2[62] ));
 sg13g2_dfrbp_1 _2611_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net137),
    .D(_0216_),
    .Q_N(_0989_),
    .Q(\bitserial_cipher.datapath.shifter2[63] ));
 sg13g2_dfrbp_1 _2612_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net133),
    .D(net647),
    .Q_N(_0988_),
    .Q(\bitserial_cipher.datapath.fifo_ff56 ));
 sg13g2_dfrbp_1 _2613_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net126),
    .D(net836),
    .Q_N(_0005_),
    .Q(\bitserial_cipher.bit_counter[0] ));
 sg13g2_dfrbp_1 _2614_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net118),
    .D(net818),
    .Q_N(_0987_),
    .Q(\bitserial_cipher.bit_counter[1] ));
 sg13g2_dfrbp_1 _2615_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net110),
    .D(_0220_),
    .Q_N(_0986_),
    .Q(\bitserial_cipher.bit_counter[2] ));
 sg13g2_dfrbp_1 _2616_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net102),
    .D(_0221_),
    .Q_N(_0985_),
    .Q(\bitserial_cipher.bit_counter[3] ));
 sg13g2_dfrbp_1 _2617_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net94),
    .D(_0222_),
    .Q_N(_0984_),
    .Q(\bitserial_cipher.bit_counter[4] ));
 sg13g2_dfrbp_1 _2618_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net86),
    .D(_0223_),
    .Q_N(_0983_),
    .Q(\bitserial_cipher.bit_counter[5] ));
 sg13g2_dfrbp_1 _2619_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net78),
    .D(_0224_),
    .Q_N(_0982_),
    .Q(\bitserial_cipher.datapath.lut_ff63 ));
 sg13g2_dfrbp_1 _2620_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net74),
    .D(_0225_),
    .Q_N(_0981_),
    .Q(\bitserial_cipher.datapath.lut_ff62 ));
 sg13g2_dfrbp_1 _2621_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net70),
    .D(_0226_),
    .Q_N(_0980_),
    .Q(\bitserial_cipher.datapath.lut_ff61 ));
 sg13g2_dfrbp_1 _2622_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net66),
    .D(_0227_),
    .Q_N(_0979_),
    .Q(\bitserial_cipher.datapath.lut_ff60 ));
 sg13g2_dfrbp_1 _2623_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net62),
    .D(_0228_),
    .Q_N(_0978_),
    .Q(\bitserial_cipher.datapath.lut_ff59 ));
 sg13g2_dfrbp_1 _2624_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net58),
    .D(_0229_),
    .Q_N(_0977_),
    .Q(\bitserial_cipher.datapath.lut_ff58 ));
 sg13g2_dfrbp_1 _2625_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net54),
    .D(_0230_),
    .Q_N(_0976_),
    .Q(\bitserial_cipher.datapath.lut_ff57 ));
 sg13g2_dfrbp_1 _2626_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net50),
    .D(_0231_),
    .Q_N(_0975_),
    .Q(\bitserial_cipher.datapath.fifo_ff63 ));
 sg13g2_dfrbp_1 _2627_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net42),
    .D(net824),
    .Q_N(_0974_),
    .Q(\bitserial_cipher.datapath.fifo_ff62 ));
 sg13g2_dfrbp_1 _2628_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net34),
    .D(_0233_),
    .Q_N(_0973_),
    .Q(\bitserial_cipher.datapath.fifo_ff61 ));
 sg13g2_dfrbp_1 _2629_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net26),
    .D(_0234_),
    .Q_N(_0972_),
    .Q(\bitserial_cipher.datapath.lut_ff56 ));
 sg13g2_dfrbp_1 _2630_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net303),
    .D(_0235_),
    .Q_N(_0000_),
    .Q(\bitserial_cipher.datapath.round_counter[0] ));
 sg13g2_dfrbp_1 _2631_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net295),
    .D(_0236_),
    .Q_N(_0004_),
    .Q(\bitserial_cipher.datapath.round_counter[1] ));
 sg13g2_dfrbp_1 _2632_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net287),
    .D(_0237_),
    .Q_N(_0001_),
    .Q(\bitserial_cipher.datapath.round_counter[2] ));
 sg13g2_dfrbp_1 _2633_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net279),
    .D(net861),
    .Q_N(_0971_),
    .Q(\bitserial_cipher.datapath.round_counter[3] ));
 sg13g2_dfrbp_1 _2634_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net271),
    .D(_0239_),
    .Q_N(_0002_),
    .Q(\bitserial_cipher.datapath.round_counter[4] ));
 sg13g2_dfrbp_1 _2635_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net263),
    .D(_0240_),
    .Q_N(_0970_),
    .Q(\bitserial_cipher.datapath.round_counter[5] ));
 sg13g2_dfrbp_1 _2636_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net255),
    .D(_0241_),
    .Q_N(_0003_),
    .Q(\bitserial_cipher.datapath.round_counter[6] ));
 sg13g2_dfrbp_1 _2637_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net247),
    .D(net787),
    .Q_N(_0969_),
    .Q(\bitserial_cipher.key_exp.lut_ff0 ));
 sg13g2_dfrbp_1 _2638_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net239),
    .D(net757),
    .Q_N(_0968_),
    .Q(\bitserial_cipher.key_exp.lut_ff1 ));
 sg13g2_dfrbp_1 _2639_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net231),
    .D(net747),
    .Q_N(_0967_),
    .Q(\bitserial_cipher.key_exp.lut_ff2 ));
 sg13g2_dfrbp_1 _2640_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net223),
    .D(_0245_),
    .Q_N(_0966_),
    .Q(\bitserial_cipher.key_exp.lut_ff3 ));
 sg13g2_dfrbp_1 _2641_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net215),
    .D(net336),
    .Q_N(_0965_),
    .Q(\bitserial_cipher.key_exp.fifo_ff0 ));
 sg13g2_dfrbp_1 _2642_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net207),
    .D(_0247_),
    .Q_N(_0964_),
    .Q(\bitserial_cipher.key_exp.fifo_ff1 ));
 sg13g2_dfrbp_1 _2643_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net199),
    .D(_0248_),
    .Q_N(_0963_),
    .Q(\bitserial_cipher.key_exp.fifo_ff2 ));
 sg13g2_dfrbp_1 _2644_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net191),
    .D(_0249_),
    .Q_N(_0962_),
    .Q(\bitserial_cipher.key_exp.fifo_ff3 ));
 sg13g2_dfrbp_1 _2645_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net183),
    .D(net437),
    .Q_N(_0961_),
    .Q(\bitserial_cipher.datapath.key_in ));
 sg13g2_dfrbp_1 _2646_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net175),
    .D(_0251_),
    .Q_N(_0960_),
    .Q(\bitserial_cipher.key_exp.shifter2[1] ));
 sg13g2_dfrbp_1 _2647_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net167),
    .D(net628),
    .Q_N(_0959_),
    .Q(\bitserial_cipher.key_exp.shifter2[2] ));
 sg13g2_dfrbp_1 _2648_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net159),
    .D(_0253_),
    .Q_N(_0958_),
    .Q(\bitserial_cipher.key_exp.shifter2[3] ));
 sg13g2_dfrbp_1 _2649_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net151),
    .D(_0254_),
    .Q_N(_0957_),
    .Q(\bitserial_cipher.key_exp.shifter2[4] ));
 sg13g2_dfrbp_1 _2650_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net143),
    .D(_0255_),
    .Q_N(_0956_),
    .Q(\bitserial_cipher.key_exp.shifter2[5] ));
 sg13g2_dfrbp_1 _2651_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net135),
    .D(_0256_),
    .Q_N(_0955_),
    .Q(\bitserial_cipher.key_exp.shifter2[6] ));
 sg13g2_dfrbp_1 _2652_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net122),
    .D(net601),
    .Q_N(_0954_),
    .Q(\bitserial_cipher.key_exp.shifter2[7] ));
 sg13g2_dfrbp_1 _2653_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net106),
    .D(_0258_),
    .Q_N(_0953_),
    .Q(\bitserial_cipher.key_exp.shifter2[8] ));
 sg13g2_dfrbp_1 _2654_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net90),
    .D(_0259_),
    .Q_N(_0952_),
    .Q(\bitserial_cipher.key_exp.shifter2[9] ));
 sg13g2_dfrbp_1 _2655_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net46),
    .D(net311),
    .Q_N(_0951_),
    .Q(\bitserial_cipher.key_exp.shifter2[10] ));
 sg13g2_dfrbp_1 _2656_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net30),
    .D(_0261_),
    .Q_N(_0950_),
    .Q(\bitserial_cipher.key_exp.shifter2[11] ));
 sg13g2_dfrbp_1 _2657_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net291),
    .D(net721),
    .Q_N(_0949_),
    .Q(\bitserial_cipher.key_exp.shifter2[12] ));
 sg13g2_dfrbp_1 _2658_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net275),
    .D(net655),
    .Q_N(_0948_),
    .Q(\bitserial_cipher.key_exp.shifter2[13] ));
 sg13g2_dfrbp_1 _2659_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net259),
    .D(_0264_),
    .Q_N(_0947_),
    .Q(\bitserial_cipher.key_exp.shifter2[14] ));
 sg13g2_dfrbp_1 _2660_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net243),
    .D(net315),
    .Q_N(_0946_),
    .Q(\bitserial_cipher.key_exp.shifter2[15] ));
 sg13g2_dfrbp_1 _2661_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net227),
    .D(_0266_),
    .Q_N(_0945_),
    .Q(\bitserial_cipher.key_exp.shifter2[16] ));
 sg13g2_dfrbp_1 _2662_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net211),
    .D(net664),
    .Q_N(_0944_),
    .Q(\bitserial_cipher.key_exp.shifter2[17] ));
 sg13g2_dfrbp_1 _2663_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net195),
    .D(_0268_),
    .Q_N(_0943_),
    .Q(\bitserial_cipher.key_exp.shifter2[18] ));
 sg13g2_dfrbp_1 _2664_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net179),
    .D(net675),
    .Q_N(_0942_),
    .Q(\bitserial_cipher.key_exp.shifter2[19] ));
 sg13g2_dfrbp_1 _2665_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net163),
    .D(_0270_),
    .Q_N(_0941_),
    .Q(\bitserial_cipher.key_exp.shifter2[20] ));
 sg13g2_dfrbp_1 _2666_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net147),
    .D(net685),
    .Q_N(_0940_),
    .Q(\bitserial_cipher.key_exp.shifter2[21] ));
 sg13g2_dfrbp_1 _2667_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net130),
    .D(net603),
    .Q_N(_0939_),
    .Q(\bitserial_cipher.key_exp.shifter2[22] ));
 sg13g2_dfrbp_1 _2668_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net98),
    .D(_0273_),
    .Q_N(_0938_),
    .Q(\bitserial_cipher.key_exp.shifter2[23] ));
 sg13g2_dfrbp_1 _2669_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net38),
    .D(net588),
    .Q_N(_0937_),
    .Q(\bitserial_cipher.key_exp.shifter2[24] ));
 sg13g2_dfrbp_1 _2670_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net283),
    .D(_0275_),
    .Q_N(_0936_),
    .Q(\bitserial_cipher.key_exp.shifter2[25] ));
 sg13g2_dfrbp_1 _2671_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net251),
    .D(net334),
    .Q_N(_0935_),
    .Q(\bitserial_cipher.key_exp.shifter2[26] ));
 sg13g2_dfrbp_1 _2672_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net219),
    .D(_0277_),
    .Q_N(_0934_),
    .Q(\bitserial_cipher.key_exp.shifter2[27] ));
 sg13g2_dfrbp_1 _2673_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net187),
    .D(net728),
    .Q_N(_0933_),
    .Q(\bitserial_cipher.key_exp.shifter2[28] ));
 sg13g2_dfrbp_1 _2674_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net155),
    .D(_0279_),
    .Q_N(_0932_),
    .Q(\bitserial_cipher.key_exp.shifter2[29] ));
 sg13g2_dfrbp_1 _2675_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net114),
    .D(net379),
    .Q_N(_0931_),
    .Q(\bitserial_cipher.key_exp.shifter2[30] ));
 sg13g2_dfrbp_1 _2676_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net299),
    .D(_0281_),
    .Q_N(_0930_),
    .Q(\bitserial_cipher.key_exp.shifter2[31] ));
 sg13g2_dfrbp_1 _2677_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net235),
    .D(net369),
    .Q_N(_0929_),
    .Q(\bitserial_cipher.key_exp.shifter2[32] ));
 sg13g2_dfrbp_1 _2678_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net171),
    .D(_0283_),
    .Q_N(_0928_),
    .Q(\bitserial_cipher.key_exp.shifter2[33] ));
 sg13g2_dfrbp_1 _2679_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net82),
    .D(_0284_),
    .Q_N(_0927_),
    .Q(\bitserial_cipher.key_exp.shifter2[34] ));
 sg13g2_dfrbp_1 _2680_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net203),
    .D(net435),
    .Q_N(_0926_),
    .Q(\bitserial_cipher.key_exp.shifter2[35] ));
 sg13g2_dfrbp_1 _2681_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net267),
    .D(_0286_),
    .Q_N(_0925_),
    .Q(\bitserial_cipher.key_exp.shifter2[36] ));
 sg13g2_tiehi _2455__25 (.L_HI(net25));
 sg13g2_tiehi _2629__26 (.L_HI(net26));
 sg13g2_tiehi _2454__27 (.L_HI(net27));
 sg13g2_tiehi _2568__28 (.L_HI(net28));
 sg13g2_tiehi _2453__29 (.L_HI(net29));
 sg13g2_tiehi _2656__30 (.L_HI(net30));
 sg13g2_tiehi _2452__31 (.L_HI(net31));
 sg13g2_tiehi _2567__32 (.L_HI(net32));
 sg13g2_tiehi _2451__33 (.L_HI(net33));
 sg13g2_tiehi _2628__34 (.L_HI(net34));
 sg13g2_tiehi _2450__35 (.L_HI(net35));
 sg13g2_tiehi _2566__36 (.L_HI(net36));
 sg13g2_tiehi _2449__37 (.L_HI(net37));
 sg13g2_tiehi _2669__38 (.L_HI(net38));
 sg13g2_tiehi _2448__39 (.L_HI(net39));
 sg13g2_tiehi _2565__40 (.L_HI(net40));
 sg13g2_tiehi _2447__41 (.L_HI(net41));
 sg13g2_tiehi _2627__42 (.L_HI(net42));
 sg13g2_tiehi _2446__43 (.L_HI(net43));
 sg13g2_tiehi _2564__44 (.L_HI(net44));
 sg13g2_tiehi _2445__45 (.L_HI(net45));
 sg13g2_tiehi _2655__46 (.L_HI(net46));
 sg13g2_tiehi _2444__47 (.L_HI(net47));
 sg13g2_tiehi _2563__48 (.L_HI(net48));
 sg13g2_tiehi _2443__49 (.L_HI(net49));
 sg13g2_tiehi _2626__50 (.L_HI(net50));
 sg13g2_tiehi _2442__51 (.L_HI(net51));
 sg13g2_tiehi _2562__52 (.L_HI(net52));
 sg13g2_tiehi _2441__53 (.L_HI(net53));
 sg13g2_tiehi _2625__54 (.L_HI(net54));
 sg13g2_tiehi _2440__55 (.L_HI(net55));
 sg13g2_tiehi _2561__56 (.L_HI(net56));
 sg13g2_tiehi _2439__57 (.L_HI(net57));
 sg13g2_tiehi _2624__58 (.L_HI(net58));
 sg13g2_tiehi _2438__59 (.L_HI(net59));
 sg13g2_tiehi _2560__60 (.L_HI(net60));
 sg13g2_tiehi _2437__61 (.L_HI(net61));
 sg13g2_tiehi _2623__62 (.L_HI(net62));
 sg13g2_tiehi _2436__63 (.L_HI(net63));
 sg13g2_tiehi _2559__64 (.L_HI(net64));
 sg13g2_tiehi _2435__65 (.L_HI(net65));
 sg13g2_tiehi _2622__66 (.L_HI(net66));
 sg13g2_tiehi _2434__67 (.L_HI(net67));
 sg13g2_tiehi _2558__68 (.L_HI(net68));
 sg13g2_tiehi _2433__69 (.L_HI(net69));
 sg13g2_tiehi _2621__70 (.L_HI(net70));
 sg13g2_tiehi _2432__71 (.L_HI(net71));
 sg13g2_tiehi _2557__72 (.L_HI(net72));
 sg13g2_tiehi _2431__73 (.L_HI(net73));
 sg13g2_tiehi _2620__74 (.L_HI(net74));
 sg13g2_tiehi _2430__75 (.L_HI(net75));
 sg13g2_tiehi _2556__76 (.L_HI(net76));
 sg13g2_tiehi _2429__77 (.L_HI(net77));
 sg13g2_tiehi _2619__78 (.L_HI(net78));
 sg13g2_tiehi _2428__79 (.L_HI(net79));
 sg13g2_tiehi _2555__80 (.L_HI(net80));
 sg13g2_tiehi _2427__81 (.L_HI(net81));
 sg13g2_tiehi _2679__82 (.L_HI(net82));
 sg13g2_tiehi _2426__83 (.L_HI(net83));
 sg13g2_tiehi _2554__84 (.L_HI(net84));
 sg13g2_tiehi _2425__85 (.L_HI(net85));
 sg13g2_tiehi _2618__86 (.L_HI(net86));
 sg13g2_tiehi _2424__87 (.L_HI(net87));
 sg13g2_tiehi _2553__88 (.L_HI(net88));
 sg13g2_tiehi _2423__89 (.L_HI(net89));
 sg13g2_tiehi _2654__90 (.L_HI(net90));
 sg13g2_tiehi _2422__91 (.L_HI(net91));
 sg13g2_tiehi _2552__92 (.L_HI(net92));
 sg13g2_tiehi _2421__93 (.L_HI(net93));
 sg13g2_tiehi _2617__94 (.L_HI(net94));
 sg13g2_tiehi _2420__95 (.L_HI(net95));
 sg13g2_tiehi _2551__96 (.L_HI(net96));
 sg13g2_tiehi _2419__97 (.L_HI(net97));
 sg13g2_tiehi _2668__98 (.L_HI(net98));
 sg13g2_tiehi _2418__99 (.L_HI(net99));
 sg13g2_tiehi _2550__100 (.L_HI(net100));
 sg13g2_tiehi _2417__101 (.L_HI(net101));
 sg13g2_tiehi _2616__102 (.L_HI(net102));
 sg13g2_tiehi _2416__103 (.L_HI(net103));
 sg13g2_tiehi _2549__104 (.L_HI(net104));
 sg13g2_tiehi _2415__105 (.L_HI(net105));
 sg13g2_tiehi _2653__106 (.L_HI(net106));
 sg13g2_tiehi _2414__107 (.L_HI(net107));
 sg13g2_tiehi _2548__108 (.L_HI(net108));
 sg13g2_tiehi _2413__109 (.L_HI(net109));
 sg13g2_tiehi _2615__110 (.L_HI(net110));
 sg13g2_tiehi _2412__111 (.L_HI(net111));
 sg13g2_tiehi _2547__112 (.L_HI(net112));
 sg13g2_tiehi _2411__113 (.L_HI(net113));
 sg13g2_tiehi _2675__114 (.L_HI(net114));
 sg13g2_tiehi _2410__115 (.L_HI(net115));
 sg13g2_tiehi _2546__116 (.L_HI(net116));
 sg13g2_tiehi _2409__117 (.L_HI(net117));
 sg13g2_tiehi _2614__118 (.L_HI(net118));
 sg13g2_tiehi _2408__119 (.L_HI(net119));
 sg13g2_tiehi _2545__120 (.L_HI(net120));
 sg13g2_tiehi _2407__121 (.L_HI(net121));
 sg13g2_tiehi _2652__122 (.L_HI(net122));
 sg13g2_tiehi _2406__123 (.L_HI(net123));
 sg13g2_tiehi _2544__124 (.L_HI(net124));
 sg13g2_tiehi _2405__125 (.L_HI(net125));
 sg13g2_tiehi _2613__126 (.L_HI(net126));
 sg13g2_tiehi _2404__127 (.L_HI(net127));
 sg13g2_tiehi _2543__128 (.L_HI(net128));
 sg13g2_tiehi _2403__129 (.L_HI(net129));
 sg13g2_tiehi _2667__130 (.L_HI(net130));
 sg13g2_tiehi _2402__131 (.L_HI(net131));
 sg13g2_tiehi _2542__132 (.L_HI(net132));
 sg13g2_tiehi _2612__133 (.L_HI(net133));
 sg13g2_tiehi _2541__134 (.L_HI(net134));
 sg13g2_tiehi _2651__135 (.L_HI(net135));
 sg13g2_tiehi _2540__136 (.L_HI(net136));
 sg13g2_tiehi _2611__137 (.L_HI(net137));
 sg13g2_tiehi _2539__138 (.L_HI(net138));
 sg13g2_tiehi _2401__139 (.L_HI(net139));
 sg13g2_tiehi _2538__140 (.L_HI(net140));
 sg13g2_tiehi _2610__141 (.L_HI(net141));
 sg13g2_tiehi _2537__142 (.L_HI(net142));
 sg13g2_tiehi _2650__143 (.L_HI(net143));
 sg13g2_tiehi _2536__144 (.L_HI(net144));
 sg13g2_tiehi _2609__145 (.L_HI(net145));
 sg13g2_tiehi _2535__146 (.L_HI(net146));
 sg13g2_tiehi _2666__147 (.L_HI(net147));
 sg13g2_tiehi _2534__148 (.L_HI(net148));
 sg13g2_tiehi _2608__149 (.L_HI(net149));
 sg13g2_tiehi _2533__150 (.L_HI(net150));
 sg13g2_tiehi _2649__151 (.L_HI(net151));
 sg13g2_tiehi _2532__152 (.L_HI(net152));
 sg13g2_tiehi _2607__153 (.L_HI(net153));
 sg13g2_tiehi _2531__154 (.L_HI(net154));
 sg13g2_tiehi _2674__155 (.L_HI(net155));
 sg13g2_tiehi _2530__156 (.L_HI(net156));
 sg13g2_tiehi _2606__157 (.L_HI(net157));
 sg13g2_tiehi _2529__158 (.L_HI(net158));
 sg13g2_tiehi _2648__159 (.L_HI(net159));
 sg13g2_tiehi _2528__160 (.L_HI(net160));
 sg13g2_tiehi _2605__161 (.L_HI(net161));
 sg13g2_tiehi _2527__162 (.L_HI(net162));
 sg13g2_tiehi _2665__163 (.L_HI(net163));
 sg13g2_tiehi _2526__164 (.L_HI(net164));
 sg13g2_tiehi _2604__165 (.L_HI(net165));
 sg13g2_tiehi _2525__166 (.L_HI(net166));
 sg13g2_tiehi _2647__167 (.L_HI(net167));
 sg13g2_tiehi _2524__168 (.L_HI(net168));
 sg13g2_tiehi _2603__169 (.L_HI(net169));
 sg13g2_tiehi _2523__170 (.L_HI(net170));
 sg13g2_tiehi _2678__171 (.L_HI(net171));
 sg13g2_tiehi _2522__172 (.L_HI(net172));
 sg13g2_tiehi _2602__173 (.L_HI(net173));
 sg13g2_tiehi _2521__174 (.L_HI(net174));
 sg13g2_tiehi _2646__175 (.L_HI(net175));
 sg13g2_tiehi _2520__176 (.L_HI(net176));
 sg13g2_tiehi _2601__177 (.L_HI(net177));
 sg13g2_tiehi _2519__178 (.L_HI(net178));
 sg13g2_tiehi _2664__179 (.L_HI(net179));
 sg13g2_tiehi _2518__180 (.L_HI(net180));
 sg13g2_tiehi _2600__181 (.L_HI(net181));
 sg13g2_tiehi _2517__182 (.L_HI(net182));
 sg13g2_tiehi _2645__183 (.L_HI(net183));
 sg13g2_tiehi _2516__184 (.L_HI(net184));
 sg13g2_tiehi _2599__185 (.L_HI(net185));
 sg13g2_tiehi _2515__186 (.L_HI(net186));
 sg13g2_tiehi _2673__187 (.L_HI(net187));
 sg13g2_tiehi _2514__188 (.L_HI(net188));
 sg13g2_tiehi _2598__189 (.L_HI(net189));
 sg13g2_tiehi _2513__190 (.L_HI(net190));
 sg13g2_tiehi _2644__191 (.L_HI(net191));
 sg13g2_tiehi _2512__192 (.L_HI(net192));
 sg13g2_tiehi _2597__193 (.L_HI(net193));
 sg13g2_tiehi _2511__194 (.L_HI(net194));
 sg13g2_tiehi _2663__195 (.L_HI(net195));
 sg13g2_tiehi _2510__196 (.L_HI(net196));
 sg13g2_tiehi _2596__197 (.L_HI(net197));
 sg13g2_tiehi _2509__198 (.L_HI(net198));
 sg13g2_tiehi _2643__199 (.L_HI(net199));
 sg13g2_tiehi _2508__200 (.L_HI(net200));
 sg13g2_tiehi _2595__201 (.L_HI(net201));
 sg13g2_tiehi _2507__202 (.L_HI(net202));
 sg13g2_tiehi _2680__203 (.L_HI(net203));
 sg13g2_tiehi _2506__204 (.L_HI(net204));
 sg13g2_tiehi _2594__205 (.L_HI(net205));
 sg13g2_tiehi _2505__206 (.L_HI(net206));
 sg13g2_tiehi _2642__207 (.L_HI(net207));
 sg13g2_tiehi _2504__208 (.L_HI(net208));
 sg13g2_tiehi _2593__209 (.L_HI(net209));
 sg13g2_tiehi _2503__210 (.L_HI(net210));
 sg13g2_tiehi _2662__211 (.L_HI(net211));
 sg13g2_tiehi _2502__212 (.L_HI(net212));
 sg13g2_tiehi _2592__213 (.L_HI(net213));
 sg13g2_tiehi _2501__214 (.L_HI(net214));
 sg13g2_tiehi _2641__215 (.L_HI(net215));
 sg13g2_tiehi _2500__216 (.L_HI(net216));
 sg13g2_tiehi _2591__217 (.L_HI(net217));
 sg13g2_tiehi _2499__218 (.L_HI(net218));
 sg13g2_tiehi _2672__219 (.L_HI(net219));
 sg13g2_tiehi _2498__220 (.L_HI(net220));
 sg13g2_tiehi _2590__221 (.L_HI(net221));
 sg13g2_tiehi _2497__222 (.L_HI(net222));
 sg13g2_tiehi _2640__223 (.L_HI(net223));
 sg13g2_tiehi _2496__224 (.L_HI(net224));
 sg13g2_tiehi _2589__225 (.L_HI(net225));
 sg13g2_tiehi _2495__226 (.L_HI(net226));
 sg13g2_tiehi _2661__227 (.L_HI(net227));
 sg13g2_tiehi _2494__228 (.L_HI(net228));
 sg13g2_tiehi _2588__229 (.L_HI(net229));
 sg13g2_tiehi _2493__230 (.L_HI(net230));
 sg13g2_tiehi _2639__231 (.L_HI(net231));
 sg13g2_tiehi _2492__232 (.L_HI(net232));
 sg13g2_tiehi _2587__233 (.L_HI(net233));
 sg13g2_tiehi _2491__234 (.L_HI(net234));
 sg13g2_tiehi _2677__235 (.L_HI(net235));
 sg13g2_tiehi _2490__236 (.L_HI(net236));
 sg13g2_tiehi _2586__237 (.L_HI(net237));
 sg13g2_tiehi _2489__238 (.L_HI(net238));
 sg13g2_tiehi _2638__239 (.L_HI(net239));
 sg13g2_tiehi _2488__240 (.L_HI(net240));
 sg13g2_tiehi _2585__241 (.L_HI(net241));
 sg13g2_tiehi _2487__242 (.L_HI(net242));
 sg13g2_tiehi _2660__243 (.L_HI(net243));
 sg13g2_tiehi _2486__244 (.L_HI(net244));
 sg13g2_tiehi _2584__245 (.L_HI(net245));
 sg13g2_tiehi _2485__246 (.L_HI(net246));
 sg13g2_tiehi _2637__247 (.L_HI(net247));
 sg13g2_tiehi _2484__248 (.L_HI(net248));
 sg13g2_tiehi _2583__249 (.L_HI(net249));
 sg13g2_tiehi _2483__250 (.L_HI(net250));
 sg13g2_tiehi _2671__251 (.L_HI(net251));
 sg13g2_tiehi _2482__252 (.L_HI(net252));
 sg13g2_tiehi _2582__253 (.L_HI(net253));
 sg13g2_tiehi _2481__254 (.L_HI(net254));
 sg13g2_tiehi _2636__255 (.L_HI(net255));
 sg13g2_tiehi _2480__256 (.L_HI(net256));
 sg13g2_tiehi _2581__257 (.L_HI(net257));
 sg13g2_tiehi _2479__258 (.L_HI(net258));
 sg13g2_tiehi _2659__259 (.L_HI(net259));
 sg13g2_tiehi _2478__260 (.L_HI(net260));
 sg13g2_tiehi _2580__261 (.L_HI(net261));
 sg13g2_tiehi _2477__262 (.L_HI(net262));
 sg13g2_tiehi _2635__263 (.L_HI(net263));
 sg13g2_tiehi _2476__264 (.L_HI(net264));
 sg13g2_tiehi _2579__265 (.L_HI(net265));
 sg13g2_tiehi _2475__266 (.L_HI(net266));
 sg13g2_tiehi _2681__267 (.L_HI(net267));
 sg13g2_tiehi _2474__268 (.L_HI(net268));
 sg13g2_tiehi _2578__269 (.L_HI(net269));
 sg13g2_tiehi _2473__270 (.L_HI(net270));
 sg13g2_tiehi _2634__271 (.L_HI(net271));
 sg13g2_tiehi _2472__272 (.L_HI(net272));
 sg13g2_tiehi _2577__273 (.L_HI(net273));
 sg13g2_tiehi _2471__274 (.L_HI(net274));
 sg13g2_tiehi _2658__275 (.L_HI(net275));
 sg13g2_tiehi _2470__276 (.L_HI(net276));
 sg13g2_tiehi _2576__277 (.L_HI(net277));
 sg13g2_tiehi _2469__278 (.L_HI(net278));
 sg13g2_tiehi _2633__279 (.L_HI(net279));
 sg13g2_tiehi _2468__280 (.L_HI(net280));
 sg13g2_tiehi _2575__281 (.L_HI(net281));
 sg13g2_tiehi _2467__282 (.L_HI(net282));
 sg13g2_tiehi _2670__283 (.L_HI(net283));
 sg13g2_tiehi _2466__284 (.L_HI(net284));
 sg13g2_tiehi _2574__285 (.L_HI(net285));
 sg13g2_tiehi _2465__286 (.L_HI(net286));
 sg13g2_tiehi _2632__287 (.L_HI(net287));
 sg13g2_tiehi _2464__288 (.L_HI(net288));
 sg13g2_tiehi _2573__289 (.L_HI(net289));
 sg13g2_tiehi _2463__290 (.L_HI(net290));
 sg13g2_tiehi _2657__291 (.L_HI(net291));
 sg13g2_tiehi _2462__292 (.L_HI(net292));
 sg13g2_tiehi _2572__293 (.L_HI(net293));
 sg13g2_tiehi _2461__294 (.L_HI(net294));
 sg13g2_tiehi _2631__295 (.L_HI(net295));
 sg13g2_tiehi _2460__296 (.L_HI(net296));
 sg13g2_tiehi _2571__297 (.L_HI(net297));
 sg13g2_tiehi _2459__298 (.L_HI(net298));
 sg13g2_tiehi _2676__299 (.L_HI(net299));
 sg13g2_tiehi _2458__300 (.L_HI(net300));
 sg13g2_tiehi _2570__301 (.L_HI(net301));
 sg13g2_tiehi _2457__302 (.L_HI(net302));
 sg13g2_tiehi _2630__303 (.L_HI(net303));
 sg13g2_tiehi _2456__304 (.L_HI(net304));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_simon_cipher_2 (.L_LO(net2));
 sg13g2_tielo tt_um_simon_cipher_3 (.L_LO(net3));
 sg13g2_tielo tt_um_simon_cipher_4 (.L_LO(net4));
 sg13g2_tielo tt_um_simon_cipher_5 (.L_LO(net5));
 sg13g2_tielo tt_um_simon_cipher_6 (.L_LO(net6));
 sg13g2_tielo tt_um_simon_cipher_7 (.L_LO(net7));
 sg13g2_tielo tt_um_simon_cipher_8 (.L_LO(net8));
 sg13g2_tielo tt_um_simon_cipher_9 (.L_LO(net9));
 sg13g2_tielo tt_um_simon_cipher_10 (.L_LO(net10));
 sg13g2_tielo tt_um_simon_cipher_11 (.L_LO(net11));
 sg13g2_tielo tt_um_simon_cipher_12 (.L_LO(net12));
 sg13g2_tielo tt_um_simon_cipher_13 (.L_LO(net13));
 sg13g2_tielo tt_um_simon_cipher_14 (.L_LO(net14));
 sg13g2_tielo tt_um_simon_cipher_15 (.L_LO(net15));
 sg13g2_tielo tt_um_simon_cipher_16 (.L_LO(net16));
 sg13g2_tielo tt_um_simon_cipher_17 (.L_LO(net17));
 sg13g2_tielo tt_um_simon_cipher_18 (.L_LO(net18));
 sg13g2_tielo tt_um_simon_cipher_19 (.L_LO(net19));
 sg13g2_tielo tt_um_simon_cipher_20 (.L_LO(net20));
 sg13g2_tielo tt_um_simon_cipher_21 (.L_LO(net21));
 sg13g2_tielo tt_um_simon_cipher_22 (.L_LO(net22));
 sg13g2_tielo tt_um_simon_cipher_23 (.L_LO(net23));
 sg13g2_tiehi _2569__24 (.L_HI(net24));
 sg13g2_buf_2 _2986_ (.A(\bitserial_cipher.cipher_data ),
    .X(uo_out[0]));
 sg13g2_buf_1 _2987_ (.A(\bitserial_cipher.datapath.valid ),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout438 (.X(net438),
    .A(_0497_));
 sg13g2_buf_2 fanout439 (.A(\bitserial_cipher.datapath.round_counter[2] ),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(net862),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(net854),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(net854),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_0834_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_0832_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(net447),
    .X(net445));
 sg13g2_buf_1 fanout446 (.A(net447),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(net450),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(net449),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(net450),
    .X(net449));
 sg13g2_buf_1 fanout450 (.A(net456),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(net453),
    .X(net451));
 sg13g2_buf_1 fanout452 (.A(net453),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(net456),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(net455),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(net456),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(ui_in[7]),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(net460),
    .X(net457));
 sg13g2_buf_1 fanout458 (.A(net460),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(net460),
    .X(net459));
 sg13g2_buf_1 fanout460 (.A(net469),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(net462),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(net465),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(net465),
    .X(net463));
 sg13g2_buf_1 fanout464 (.A(net465),
    .X(net464));
 sg13g2_buf_1 fanout465 (.A(net469),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(net467),
    .X(net466));
 sg13g2_buf_1 fanout467 (.A(net469),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(net469),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(ui_in[7]),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(net474),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(net474),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(net474),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(net474),
    .X(net473));
 sg13g2_buf_1 fanout474 (.A(net489),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(net489),
    .X(net475));
 sg13g2_buf_1 fanout476 (.A(net489),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(net479),
    .X(net477));
 sg13g2_buf_1 fanout478 (.A(net479),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(net485),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(net485),
    .X(net480));
 sg13g2_buf_1 fanout481 (.A(net482),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(net485),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(net484),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(net485),
    .X(net484));
 sg13g2_buf_1 fanout485 (.A(net489),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(net488),
    .X(net486));
 sg13g2_buf_1 fanout487 (.A(net488),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(net489),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(ui_in[7]),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(net491),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(net492),
    .X(net491));
 sg13g2_buf_1 fanout492 (.A(net494),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(net494),
    .X(net493));
 sg13g2_buf_1 fanout494 (.A(net507),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(net497),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(net497),
    .X(net496));
 sg13g2_buf_1 fanout497 (.A(net507),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(net500),
    .X(net498));
 sg13g2_buf_1 fanout499 (.A(net500),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(net507),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(net503),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(net503),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(net507),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(net506),
    .X(net504));
 sg13g2_buf_1 fanout505 (.A(net506),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(net507),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(net533),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net510),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(net518),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(net513),
    .X(net511));
 sg13g2_buf_1 fanout512 (.A(net513),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(net518),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(net517),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(net517),
    .X(net515));
 sg13g2_buf_1 fanout516 (.A(net517),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(net518),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(net533),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(net521),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(net521),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(net527),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(net523),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(net527),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(net526),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(net526),
    .X(net525));
 sg13g2_buf_1 fanout526 (.A(net527),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(net533),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(net532),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(net531),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(net532),
    .X(net530));
 sg13g2_buf_1 fanout531 (.A(net532),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(net533),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(ui_in[6]),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net536),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(net536),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(net544),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(net544),
    .X(net537));
 sg13g2_buf_1 fanout538 (.A(net544),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(net541),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(net541),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(net544),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(net543),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(net544),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(net578),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net546),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(net548),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(net548),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net559),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(net551),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(net551),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(net559),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_1 fanout554 (.A(net559),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(net558),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(net558),
    .X(net556));
 sg13g2_buf_1 fanout557 (.A(net558),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(net578),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(net561),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net562),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(net569),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(net566),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(net566),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(net566),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(net569),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(net569),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(net569),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(net578),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(net573),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(net573),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(net577),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net577),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(net577),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(rst_n),
    .X(net578));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_35_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_12_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_17_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\bitserial_cipher.datapath.lut_ff61 ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold2 (.A(\bitserial_cipher.datapath.lut_ff57 ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold3 (.A(\bitserial_cipher.datapath.lut_ff60 ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold4 (.A(\bitserial_cipher.datapath.lut_ff59 ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold5 (.A(\bitserial_cipher.datapath.lut_ff58 ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold6 (.A(\bitserial_cipher.key_exp.shifter2[11] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0260_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold8 (.A(\bitserial_cipher.datapath.shifter2[48] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0200_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold10 (.A(\bitserial_cipher.key_exp.shifter2[16] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0265_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold12 (.A(\bitserial_cipher.datapath.shifter1[18] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0114_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold14 (.A(\bitserial_cipher.key_exp.shifter1[27] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0059_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold16 (.A(\bitserial_cipher.datapath.lut_ff63 ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold17 (.A(\bitserial_cipher.key_exp.shifter1[37] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0069_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold19 (.A(\bitserial_cipher.datapath.shifter1[53] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0149_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold21 (.A(\bitserial_cipher.datapath.shifter1[40] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0136_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold23 (.A(\bitserial_cipher.key_exp.shifter1[15] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0047_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold25 (.A(\bitserial_cipher.datapath.shifter2[53] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0205_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold27 (.A(\bitserial_cipher.key_exp.shifter1[19] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0051_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold29 (.A(\bitserial_cipher.key_exp.shifter2[27] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0276_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold31 (.A(\bitserial_cipher.key_exp.fifo_ff1 ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0246_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold33 (.A(\bitserial_cipher.datapath.fifo_ff60 ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0095_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold35 (.A(\bitserial_cipher.datapath.shifter2[42] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0194_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold37 (.A(\bitserial_cipher.datapath.shifter1[24] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0120_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold39 (.A(\bitserial_cipher.key_exp.shifter1[2] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0034_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold41 (.A(\bitserial_cipher.datapath.shifter2[44] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0196_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold43 (.A(\bitserial_cipher.datapath.shifter2[59] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0211_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold45 (.A(\bitserial_cipher.datapath.shifter1[43] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0139_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold47 (.A(\bitserial_cipher.datapath.shifter2[17] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0169_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold49 (.A(\bitserial_cipher.datapath.shifter1[29] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0125_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold51 (.A(\bitserial_cipher.datapath.shifter2[63] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0215_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold53 (.A(\bitserial_cipher.key_exp.shifter1[57] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0089_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold55 (.A(\bitserial_cipher.datapath.lut_ff62 ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold56 (.A(\bitserial_cipher.key_exp.shifter1[34] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0066_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold58 (.A(\bitserial_cipher.datapath.shifter1[9] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0105_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold60 (.A(\bitserial_cipher.datapath.shifter2[34] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0186_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold62 (.A(\bitserial_cipher.datapath.shifter2[6] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0158_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold64 (.A(\bitserial_cipher.key_exp.shifter2[33] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0282_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold66 (.A(\bitserial_cipher.key_exp.shifter1[41] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0073_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold68 (.A(\bitserial_cipher.key_exp.shifter2[63] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0031_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold70 (.A(\bitserial_cipher.datapath.shifter1[51] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0147_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold72 (.A(\bitserial_cipher.datapath.shifter1[7] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0103_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold74 (.A(\bitserial_cipher.key_exp.shifter2[31] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0280_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold76 (.A(\bitserial_cipher.datapath.shifter2[22] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0174_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold78 (.A(\bitserial_cipher.key_exp.shifter1[50] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0082_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold80 (.A(\bitserial_cipher.datapath.shifter2[11] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0163_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold82 (.A(\bitserial_cipher.datapath.shifter2[7] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold83 (.A(\bitserial_cipher.key_exp.shifter1[20] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold84 (.A(\bitserial_cipher.datapath.fifo_ff59 ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0094_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold86 (.A(\bitserial_cipher.key_exp.shifter1[13] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0045_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold88 (.A(\bitserial_cipher.datapath.shifter2[25] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0177_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold90 (.A(\bitserial_cipher.datapath.shifter2[56] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0208_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold92 (.A(\bitserial_cipher.datapath.shifter1[50] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0146_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold94 (.A(\bitserial_cipher.key_exp.shifter2[49] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0017_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold96 (.A(\bitserial_cipher.datapath.shifter2[5] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0157_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold98 (.A(\bitserial_cipher.key_exp.shifter1[44] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0076_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold100 (.A(\bitserial_cipher.key_exp.shifter2[41] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0009_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold102 (.A(\bitserial_cipher.datapath.shifter2[41] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0193_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold104 (.A(\bitserial_cipher.datapath.shifter2[21] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0173_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold106 (.A(\bitserial_cipher.key_exp.shifter2[60] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0028_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold108 (.A(\bitserial_cipher.datapath.shifter1[20] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0116_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold110 (.A(\bitserial_cipher.datapath.shifter2[28] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0180_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold112 (.A(\bitserial_cipher.datapath.shifter2[62] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0214_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold114 (.A(\bitserial_cipher.datapath.shifter1[39] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0135_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold116 (.A(\bitserial_cipher.datapath.shifter2[3] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0155_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold118 (.A(\bitserial_cipher.datapath.shifter2[15] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0167_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold120 (.A(\bitserial_cipher.key_exp.shifter1[58] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold121 (.A(\bitserial_cipher.datapath.shifter2[33] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0185_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold123 (.A(\bitserial_cipher.key_exp.shifter1[49] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0081_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold125 (.A(\bitserial_cipher.key_exp.shifter2[42] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold126 (.A(\bitserial_cipher.key_exp.shifter1[55] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0087_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold128 (.A(\bitserial_cipher.datapath.shifter1[27] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0123_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold130 (.A(\bitserial_cipher.key_exp.shifter2[36] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0285_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold132 (.A(\bitserial_cipher.key_exp.shifter2[1] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0250_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold134 (.A(\bitserial_cipher.datapath.shifter2[1] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0153_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold136 (.A(\bitserial_cipher.key_exp.shifter2[56] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0024_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold138 (.A(\bitserial_cipher.datapath.shifter2[52] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0204_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold140 (.A(\bitserial_cipher.key_exp.shifter2[53] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0021_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold142 (.A(\bitserial_cipher.key_exp.shifter2[25] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0274_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold144 (.A(\bitserial_cipher.key_exp.shifter1[46] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0078_),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold146 (.A(\bitserial_cipher.datapath.shifter1[33] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0129_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold148 (.A(\bitserial_cipher.key_exp.shifter1[24] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0056_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold150 (.A(\bitserial_cipher.key_exp.shifter1[18] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0050_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold152 (.A(\bitserial_cipher.key_exp.shifter2[43] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold153 (.A(\bitserial_cipher.key_exp.shifter1[53] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0085_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold155 (.A(\bitserial_cipher.key_exp.shifter2[8] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0257_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold157 (.A(\bitserial_cipher.key_exp.shifter2[23] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0272_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold159 (.A(\bitserial_cipher.datapath.shifter1[13] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0109_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold161 (.A(\bitserial_cipher.datapath.shifter1[6] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0102_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold163 (.A(\bitserial_cipher.key_exp.shifter2[34] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold164 (.A(\bitserial_cipher.datapath.shifter2[54] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold165 (.A(\bitserial_cipher.key_exp.shifter1[25] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold166 (.A(\bitserial_cipher.datapath.fifo_ff61 ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold167 (.A(\bitserial_cipher.datapath.shifter2[26] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold168 (.A(\bitserial_cipher.key_exp.shifter2[59] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0027_),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold170 (.A(\bitserial_cipher.key_exp.shifter1[11] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0043_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold172 (.A(\bitserial_cipher.key_exp.shifter2[61] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold173 (.A(\bitserial_cipher.datapath.shifter1[49] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0145_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold175 (.A(\bitserial_cipher.key_exp.shifter2[24] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold176 (.A(\bitserial_cipher.key_exp.shifter1[8] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0040_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold178 (.A(\bitserial_cipher.datapath.shifter2[19] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0171_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold180 (.A(\bitserial_cipher.key_exp.shifter2[35] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold181 (.A(\bitserial_cipher.datapath.shifter1[34] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold182 (.A(\bitserial_cipher.key_exp.shifter2[3] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0252_),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold184 (.A(\bitserial_cipher.datapath.shifter1[14] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold185 (.A(\bitserial_cipher.datapath.shifter1[12] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0108_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold187 (.A(\bitserial_cipher.key_exp.shifter1[28] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold188 (.A(\bitserial_cipher.datapath.shifter2[18] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold189 (.A(\bitserial_cipher.key_exp.shifter2[40] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0008_),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold191 (.A(\bitserial_cipher.key_exp.fifo_ff2 ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold192 (.A(\bitserial_cipher.key_exp.shifter1[17] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0049_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold194 (.A(\bitserial_cipher.datapath.shifter1[41] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold195 (.A(\bitserial_cipher.datapath.shifter2[35] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold196 (.A(\bitserial_cipher.datapath.fifo_ff58 ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0093_),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold198 (.A(\bitserial_cipher.key_exp.shifter1[7] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0039_),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold200 (.A(\bitserial_cipher.datapath.shifter1[10] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold201 (.A(\bitserial_cipher.datapath.fifo_ff57 ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0217_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold203 (.A(\bitserial_cipher.key_exp.shifter2[45] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0013_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold205 (.A(\bitserial_cipher.key_exp.shifter1[10] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0042_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold207 (.A(\bitserial_cipher.key_exp.shifter2[48] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0016_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold209 (.A(\bitserial_cipher.key_exp.shifter2[14] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0263_),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold211 (.A(\bitserial_cipher.datapath.shifter2[31] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0183_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold213 (.A(\bitserial_cipher.datapath.shifter1[16] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0112_),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold215 (.A(\bitserial_cipher.datapath.shifter1[19] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold216 (.A(\bitserial_cipher.datapath.shifter2[8] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold217 (.A(\bitserial_cipher.key_exp.shifter1[56] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold218 (.A(\bitserial_cipher.key_exp.shifter2[18] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0267_),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold220 (.A(\bitserial_cipher.datapath.shifter1[11] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold221 (.A(\bitserial_cipher.datapath.shifter2[16] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold222 (.A(\bitserial_cipher.key_exp.shifter2[51] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0019_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold224 (.A(\bitserial_cipher.datapath.shifter1[1] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0097_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold226 (.A(\bitserial_cipher.key_exp.shifter2[4] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold227 (.A(\bitserial_cipher.key_exp.shifter1[1] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0033_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold229 (.A(\bitserial_cipher.key_exp.shifter2[20] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0269_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold231 (.A(\bitserial_cipher.datapath.shifter2[13] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0165_),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold233 (.A(\bitserial_cipher.key_exp.shifter2[38] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0006_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold235 (.A(\bitserial_cipher.datapath.shifter2[58] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0210_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold237 (.A(\bitserial_cipher.datapath.shifter1[22] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0118_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold239 (.A(\bitserial_cipher.key_exp.shifter2[22] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0271_),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold241 (.A(\bitserial_cipher.key_exp.shifter1[30] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0062_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold243 (.A(\bitserial_cipher.key_exp.shifter1[31] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold244 (.A(\bitserial_cipher.key_exp.shifter2[32] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold245 (.A(\bitserial_cipher.key_exp.shifter1[42] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold246 (.A(\bitserial_cipher.key_exp.shifter1[38] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold247 (.A(\bitserial_cipher.key_exp.shifter2[26] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold248 (.A(\bitserial_cipher.datapath.shifter1[48] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0144_),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold250 (.A(\bitserial_cipher.datapath.shifter2[10] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0162_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold252 (.A(\bitserial_cipher.key_exp.shifter1[45] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold253 (.A(\bitserial_cipher.datapath.shifter1[26] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0122_),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold255 (.A(\bitserial_cipher.key_exp.shifter1[47] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold256 (.A(\bitserial_cipher.datapath.shifter2[4] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold257 (.A(\bitserial_cipher.key_exp.shifter1[29] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold258 (.A(\bitserial_cipher.key_exp.shifter1[51] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold259 (.A(\bitserial_cipher.key_exp.shifter2[9] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold260 (.A(\bitserial_cipher.key_exp.shifter2[54] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold261 (.A(\bitserial_cipher.datapath.shifter2[24] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0176_),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold263 (.A(\bitserial_cipher.datapath.shifter1[54] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0151_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold265 (.A(\bitserial_cipher.datapath.shifter2[23] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold266 (.A(\bitserial_cipher.key_exp.shifter2[2] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold267 (.A(\bitserial_cipher.datapath.shifter2[12] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold268 (.A(\bitserial_cipher.key_exp.shifter1[52] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold269 (.A(\bitserial_cipher.key_exp.shifter2[21] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold270 (.A(\bitserial_cipher.datapath.shifter2[37] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0189_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold272 (.A(\bitserial_cipher.datapath.shifter1[44] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold273 (.A(\bitserial_cipher.datapath.shifter1[5] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0101_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold275 (.A(\bitserial_cipher.key_exp.shifter2[13] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0262_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold277 (.A(\bitserial_cipher.datapath.shifter1[42] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold278 (.A(\bitserial_cipher.key_exp.shifter1[3] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold279 (.A(\bitserial_cipher.datapath.shifter1[15] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold280 (.A(\bitserial_cipher.datapath.shifter2[36] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold281 (.A(\bitserial_cipher.key_exp.shifter1[35] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold282 (.A(\bitserial_cipher.key_exp.shifter2[29] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0278_),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold284 (.A(\bitserial_cipher.datapath.shifter2[39] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0191_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold286 (.A(\bitserial_cipher.datapath.shifter2[20] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold287 (.A(\bitserial_cipher.datapath.shifter2[43] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold288 (.A(\bitserial_cipher.datapath.shifter2[32] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold289 (.A(\bitserial_cipher.datapath.shifter1[47] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0143_),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold291 (.A(\bitserial_cipher.key_exp.shifter2[50] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold292 (.A(\bitserial_cipher.datapath.shifter2[45] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold293 (.A(\bitserial_cipher.key_exp.shifter1[14] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold294 (.A(\bitserial_cipher.key_exp.shifter2[46] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold295 (.A(\bitserial_cipher.key_exp.shifter1[21] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold296 (.A(\bitserial_cipher.datapath.shifter2[9] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold297 (.A(\bitserial_cipher.key_exp.shifter1[16] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold298 (.A(\bitserial_cipher.key_exp.shifter1[48] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold299 (.A(\bitserial_cipher.key_exp.shifter2[44] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold300 (.A(\bitserial_cipher.datapath.shifter1[30] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold301 (.A(\bitserial_cipher.key_exp.lut_ff3 ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0244_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold303 (.A(\bitserial_cipher.key_exp.shifter1[5] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0037_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold305 (.A(\bitserial_cipher.key_exp.shifter2[57] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold306 (.A(\bitserial_cipher.key_exp.shifter1[39] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold307 (.A(\bitserial_cipher.datapath.shifter2[2] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold308 (.A(\bitserial_cipher.datapath.shifter1[17] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold309 (.A(\bitserial_cipher.datapath.shifter1[8] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold310 (.A(\bitserial_cipher.datapath.shifter2[29] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold311 (.A(\bitserial_cipher.key_exp.lut_ff2 ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0243_),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold313 (.A(\bitserial_cipher.datapath.shifter2[14] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold314 (.A(\bitserial_cipher.key_exp.shifter1[22] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold315 (.A(\bitserial_cipher.datapath.shifter1[31] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold316 (.A(\bitserial_cipher.datapath.shifter2[61] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0213_),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold318 (.A(\bitserial_cipher.key_exp.shifter2[5] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold319 (.A(\bitserial_cipher.datapath.shifter2[51] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0203_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold321 (.A(\bitserial_cipher.key_exp.shifter2[30] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold322 (.A(\bitserial_cipher.key_exp.shifter1[9] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold323 (.A(\bitserial_cipher.key_exp.shifter2[6] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold324 (.A(\bitserial_cipher.datapath.shifter2[40] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold325 (.A(\bitserial_cipher.key_exp.shifter1[12] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold326 (.A(\bitserial_cipher.datapath.shifter2[27] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold327 (.A(\bitserial_cipher.datapath.shifter1[32] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold328 (.A(\bitserial_cipher.key_exp.shifter2[15] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold329 (.A(\bitserial_cipher.key_exp.shifter2[47] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold330 (.A(\bitserial_cipher.datapath.shifter1[28] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold331 (.A(\bitserial_cipher.datapath.shifter2[47] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0199_),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold333 (.A(\bitserial_cipher.datapath.shifter1[2] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold334 (.A(\bitserial_cipher.datapath.shifter1[21] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold335 (.A(\bitserial_cipher.datapath.shifter1[38] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0134_),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold337 (.A(\bitserial_cipher.key_exp.shifter2[28] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold338 (.A(\bitserial_cipher.datapath.shifter1[25] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold339 (.A(\bitserial_cipher.key_exp.shifter1[6] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold340 (.A(\bitserial_cipher.datapath.shifter2[57] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold341 (.A(\bitserial_cipher.key_exp.lut_ff1 ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0242_),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold343 (.A(\bitserial_cipher.datapath.shifter1[55] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0419_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold345 (.A(\bitserial_cipher.datapath.shifter1[46] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0142_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold347 (.A(\bitserial_cipher.key_exp.shifter2[39] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold348 (.A(\bitserial_cipher.datapath.shifter2[60] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold349 (.A(\bitserial_cipher.key_exp.fifo_ff3 ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold350 (.A(\bitserial_cipher.datapath.shifter1[37] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0133_),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold352 (.A(\bitserial_cipher.key_exp.shifter1[26] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold353 (.A(\bitserial_cipher.datapath.shifter1[45] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold354 (.A(\bitserial_cipher.key_exp.shifter2[62] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold355 (.A(\bitserial_cipher.datapath.shifter1[35] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold356 (.A(\bitserial_cipher.datapath.shifter2[55] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold357 (.A(\bitserial_cipher.key_exp.shifter2[52] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold358 (.A(\bitserial_cipher.key_exp.shifter1[32] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold359 (.A(\bitserial_cipher.key_exp.shifter1[36] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold360 (.A(\bitserial_cipher.key_exp.shifter2[19] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold361 (.A(\bitserial_cipher.datapath.shifter2[30] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold362 (.A(\bitserial_cipher.datapath.shifter2[49] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold363 (.A(\bitserial_cipher.key_exp.shifter2[37] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold364 (.A(\bitserial_cipher.key_exp.shifter1[23] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold365 (.A(\bitserial_cipher.datapath.shifter1[4] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0100_),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold367 (.A(\bitserial_cipher.key_exp.shifter1[43] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold368 (.A(\bitserial_cipher.key_exp.shifter2[17] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold369 (.A(\bitserial_cipher.datapath.shifter2[38] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold370 (.A(\bitserial_cipher.datapath.shifter1[52] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold371 (.A(\bitserial_cipher.bit_counter[1] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0488_),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0219_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold374 (.A(\bitserial_cipher.key_exp.shifter1[4] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold375 (.A(\bitserial_cipher.bit_counter[2] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold376 (.A(\bitserial_cipher.key_exp.shifter1[59] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold377 (.A(\bitserial_cipher.datapath.shifter1[36] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold378 (.A(\bitserial_cipher.datapath.fifo_ff63 ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0232_),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold380 (.A(\bitserial_cipher.datapath.shifter1[3] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold381 (.A(\bitserial_cipher.datapath.shifter2[50] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold382 (.A(\bitserial_cipher.key_exp.shifter2[58] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold383 (.A(\bitserial_cipher.key_exp.shifter2[55] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold384 (.A(\bitserial_cipher.key_exp.shifter1[54] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold385 (.A(\bitserial_cipher.key_exp.shifter1[40] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold386 (.A(\bitserial_cipher.key_exp.shifter1[33] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold387 (.A(\bitserial_cipher.key_exp.shifter2[7] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold388 (.A(\bitserial_cipher.key_exp.shifter2[10] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold389 (.A(\bitserial_cipher.datapath.fifo_ff62 ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0005_),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0218_),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold392 (.A(\bitserial_cipher.datapath.shifter2[46] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold393 (.A(\bitserial_cipher.key_exp.lut_ff0 ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0874_),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold395 (.A(\bitserial_cipher.datapath.shifter1[23] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold396 (.A(\bitserial_cipher.key_exp.shift_out1 ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold397 (.A(\bitserial_cipher.bit_counter[4] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold398 (.A(_0495_),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold399 (.A(\bitserial_cipher.key_exp.shifter2[12] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold400 (.A(\bitserial_cipher.datapath.shift_in2 ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold401 (.A(\bitserial_cipher.bit_counter[0] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold402 (.A(\bitserial_cipher.bit_counter[5] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold403 (.A(\bitserial_cipher.bit_counter[3] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold404 (.A(\bitserial_cipher.datapath.round_counter[4] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0525_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0001_),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0519_),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold408 (.A(\bitserial_cipher.key_exp.fifo_ff0 ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold409 (.A(\bitserial_cipher.datapath.round_counter[0] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0000_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold411 (.A(\bitserial_cipher.datapath.round_counter[6] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0530_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold413 (.A(\bitserial_cipher.datapath.round_counter[5] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold414 (.A(\bitserial_cipher.datapath.round_counter[3] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0523_),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0238_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold417 (.A(\bitserial_cipher.datapath.round_counter[1] ),
    .X(net862));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_4 FILLER_11_322 ();
 sg13g2_fill_2 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_331 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_decap_8 FILLER_11_345 ();
 sg13g2_decap_8 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_fill_1 FILLER_12_140 ();
 sg13g2_fill_2 FILLER_12_152 ();
 sg13g2_fill_1 FILLER_12_154 ();
 sg13g2_fill_2 FILLER_12_159 ();
 sg13g2_fill_1 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_165 ();
 sg13g2_decap_8 FILLER_12_172 ();
 sg13g2_decap_8 FILLER_12_179 ();
 sg13g2_decap_8 FILLER_12_186 ();
 sg13g2_decap_8 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_214 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_4 FILLER_12_245 ();
 sg13g2_fill_1 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_4 FILLER_12_301 ();
 sg13g2_fill_1 FILLER_12_305 ();
 sg13g2_decap_4 FILLER_12_314 ();
 sg13g2_fill_1 FILLER_12_318 ();
 sg13g2_fill_2 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_decap_8 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_4 FILLER_13_119 ();
 sg13g2_fill_2 FILLER_13_123 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_fill_1 FILLER_13_166 ();
 sg13g2_decap_8 FILLER_13_180 ();
 sg13g2_decap_8 FILLER_13_187 ();
 sg13g2_decap_8 FILLER_13_194 ();
 sg13g2_decap_8 FILLER_13_201 ();
 sg13g2_decap_8 FILLER_13_208 ();
 sg13g2_decap_8 FILLER_13_215 ();
 sg13g2_decap_4 FILLER_13_222 ();
 sg13g2_fill_1 FILLER_13_226 ();
 sg13g2_fill_2 FILLER_13_243 ();
 sg13g2_decap_8 FILLER_13_271 ();
 sg13g2_fill_2 FILLER_13_278 ();
 sg13g2_fill_1 FILLER_13_280 ();
 sg13g2_fill_2 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_289 ();
 sg13g2_decap_4 FILLER_13_296 ();
 sg13g2_fill_2 FILLER_13_300 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_decap_8 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_fill_2 FILLER_14_112 ();
 sg13g2_fill_1 FILLER_14_203 ();
 sg13g2_decap_4 FILLER_14_213 ();
 sg13g2_fill_2 FILLER_14_291 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_1 FILLER_14_330 ();
 sg13g2_decap_8 FILLER_14_366 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_fill_2 FILLER_15_105 ();
 sg13g2_fill_1 FILLER_15_213 ();
 sg13g2_fill_1 FILLER_15_250 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_4 FILLER_16_105 ();
 sg13g2_fill_2 FILLER_16_109 ();
 sg13g2_fill_2 FILLER_16_151 ();
 sg13g2_fill_2 FILLER_16_162 ();
 sg13g2_fill_2 FILLER_16_218 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_fill_1 FILLER_17_137 ();
 sg13g2_fill_2 FILLER_17_148 ();
 sg13g2_fill_1 FILLER_17_211 ();
 sg13g2_fill_2 FILLER_17_253 ();
 sg13g2_fill_2 FILLER_17_263 ();
 sg13g2_fill_1 FILLER_17_356 ();
 sg13g2_fill_2 FILLER_17_363 ();
 sg13g2_fill_1 FILLER_17_365 ();
 sg13g2_fill_2 FILLER_17_373 ();
 sg13g2_fill_1 FILLER_17_375 ();
 sg13g2_fill_2 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_fill_1 FILLER_18_162 ();
 sg13g2_decap_4 FILLER_18_177 ();
 sg13g2_fill_2 FILLER_18_267 ();
 sg13g2_fill_1 FILLER_18_274 ();
 sg13g2_fill_2 FILLER_18_283 ();
 sg13g2_fill_1 FILLER_18_322 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_4 FILLER_19_119 ();
 sg13g2_fill_1 FILLER_19_123 ();
 sg13g2_fill_1 FILLER_19_158 ();
 sg13g2_fill_2 FILLER_19_198 ();
 sg13g2_fill_2 FILLER_19_205 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_fill_1 FILLER_19_258 ();
 sg13g2_fill_2 FILLER_19_278 ();
 sg13g2_fill_2 FILLER_19_317 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_fill_2 FILLER_20_119 ();
 sg13g2_fill_1 FILLER_20_187 ();
 sg13g2_decap_4 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_227 ();
 sg13g2_fill_2 FILLER_20_232 ();
 sg13g2_fill_2 FILLER_20_376 ();
 sg13g2_fill_1 FILLER_20_392 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_fill_1 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_160 ();
 sg13g2_decap_4 FILLER_21_187 ();
 sg13g2_fill_2 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_fill_2 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_223 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_fill_2 FILLER_21_237 ();
 sg13g2_fill_2 FILLER_21_299 ();
 sg13g2_fill_2 FILLER_21_349 ();
 sg13g2_fill_2 FILLER_21_379 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_4 FILLER_22_112 ();
 sg13g2_fill_2 FILLER_22_116 ();
 sg13g2_fill_1 FILLER_22_138 ();
 sg13g2_fill_2 FILLER_22_153 ();
 sg13g2_fill_2 FILLER_22_160 ();
 sg13g2_fill_1 FILLER_22_177 ();
 sg13g2_fill_2 FILLER_22_187 ();
 sg13g2_fill_1 FILLER_22_221 ();
 sg13g2_decap_4 FILLER_22_239 ();
 sg13g2_fill_2 FILLER_22_243 ();
 sg13g2_fill_2 FILLER_22_275 ();
 sg13g2_fill_1 FILLER_22_286 ();
 sg13g2_fill_2 FILLER_22_327 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_119 ();
 sg13g2_fill_1 FILLER_23_173 ();
 sg13g2_fill_2 FILLER_23_204 ();
 sg13g2_decap_4 FILLER_23_246 ();
 sg13g2_fill_1 FILLER_23_250 ();
 sg13g2_fill_2 FILLER_23_283 ();
 sg13g2_fill_1 FILLER_23_290 ();
 sg13g2_fill_2 FILLER_23_303 ();
 sg13g2_fill_1 FILLER_23_322 ();
 sg13g2_fill_1 FILLER_23_352 ();
 sg13g2_fill_1 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_fill_2 FILLER_24_145 ();
 sg13g2_decap_4 FILLER_24_165 ();
 sg13g2_fill_1 FILLER_24_174 ();
 sg13g2_decap_4 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_267 ();
 sg13g2_decap_8 FILLER_24_274 ();
 sg13g2_fill_2 FILLER_24_347 ();
 sg13g2_fill_1 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_fill_1 FILLER_25_139 ();
 sg13g2_fill_1 FILLER_25_150 ();
 sg13g2_fill_1 FILLER_25_217 ();
 sg13g2_fill_1 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_250 ();
 sg13g2_fill_1 FILLER_25_252 ();
 sg13g2_fill_2 FILLER_25_257 ();
 sg13g2_fill_2 FILLER_25_269 ();
 sg13g2_fill_1 FILLER_25_340 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_126 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_306 ();
 sg13g2_fill_1 FILLER_26_344 ();
 sg13g2_fill_2 FILLER_26_350 ();
 sg13g2_fill_2 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_178 ();
 sg13g2_fill_1 FILLER_27_188 ();
 sg13g2_fill_1 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_fill_2 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_321 ();
 sg13g2_fill_1 FILLER_27_356 ();
 sg13g2_fill_1 FILLER_27_376 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_4 FILLER_28_126 ();
 sg13g2_fill_2 FILLER_28_130 ();
 sg13g2_decap_4 FILLER_28_149 ();
 sg13g2_decap_8 FILLER_28_167 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_206 ();
 sg13g2_fill_2 FILLER_28_280 ();
 sg13g2_fill_1 FILLER_28_301 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_143 ();
 sg13g2_fill_1 FILLER_29_162 ();
 sg13g2_fill_2 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_191 ();
 sg13g2_fill_2 FILLER_29_252 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_fill_2 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_4 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_116 ();
 sg13g2_fill_2 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_180 ();
 sg13g2_fill_1 FILLER_31_196 ();
 sg13g2_fill_1 FILLER_31_207 ();
 sg13g2_decap_8 FILLER_31_240 ();
 sg13g2_fill_2 FILLER_31_247 ();
 sg13g2_fill_1 FILLER_31_256 ();
 sg13g2_fill_1 FILLER_31_279 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_fill_2 FILLER_31_385 ();
 sg13g2_fill_1 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_4 FILLER_32_112 ();
 sg13g2_fill_2 FILLER_32_116 ();
 sg13g2_decap_8 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_242 ();
 sg13g2_decap_8 FILLER_32_249 ();
 sg13g2_decap_8 FILLER_32_256 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_fill_1 FILLER_32_279 ();
 sg13g2_fill_1 FILLER_32_283 ();
 sg13g2_fill_1 FILLER_32_288 ();
 sg13g2_fill_2 FILLER_32_321 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_4 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_128 ();
 sg13g2_fill_2 FILLER_33_160 ();
 sg13g2_fill_1 FILLER_33_166 ();
 sg13g2_decap_8 FILLER_33_180 ();
 sg13g2_fill_2 FILLER_33_187 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_fill_2 FILLER_33_211 ();
 sg13g2_fill_1 FILLER_33_223 ();
 sg13g2_decap_8 FILLER_33_250 ();
 sg13g2_decap_8 FILLER_33_257 ();
 sg13g2_decap_8 FILLER_33_264 ();
 sg13g2_fill_1 FILLER_33_271 ();
 sg13g2_fill_1 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_353 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_4 FILLER_34_112 ();
 sg13g2_fill_2 FILLER_34_116 ();
 sg13g2_decap_4 FILLER_34_166 ();
 sg13g2_fill_2 FILLER_34_173 ();
 sg13g2_decap_8 FILLER_34_178 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_fill_2 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_215 ();
 sg13g2_decap_8 FILLER_34_244 ();
 sg13g2_decap_4 FILLER_34_251 ();
 sg13g2_fill_1 FILLER_34_255 ();
 sg13g2_decap_4 FILLER_34_259 ();
 sg13g2_fill_1 FILLER_34_263 ();
 sg13g2_fill_1 FILLER_34_290 ();
 sg13g2_fill_2 FILLER_34_339 ();
 sg13g2_fill_1 FILLER_34_357 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_fill_2 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_fill_2 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_202 ();
 sg13g2_fill_1 FILLER_35_365 ();
 sg13g2_fill_1 FILLER_35_380 ();
 sg13g2_fill_2 FILLER_35_395 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_fill_1 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_fill_2 FILLER_36_292 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_4 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_116 ();
 sg13g2_fill_2 FILLER_37_121 ();
 sg13g2_fill_1 FILLER_37_205 ();
 sg13g2_fill_2 FILLER_37_222 ();
 sg13g2_fill_1 FILLER_37_234 ();
 sg13g2_fill_1 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_4 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_113 ();
 sg13g2_fill_2 FILLER_38_151 ();
 sg13g2_fill_2 FILLER_38_162 ();
 sg13g2_fill_2 FILLER_38_245 ();
 sg13g2_fill_2 FILLER_38_273 ();
 sg13g2_fill_1 FILLER_38_313 ();
 sg13g2_fill_1 FILLER_38_352 ();
 sg13g2_fill_1 FILLER_38_376 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_fill_1 FILLER_39_124 ();
 sg13g2_fill_2 FILLER_39_153 ();
 sg13g2_fill_2 FILLER_39_190 ();
 sg13g2_fill_1 FILLER_39_257 ();
 sg13g2_fill_2 FILLER_39_323 ();
 sg13g2_fill_1 FILLER_39_339 ();
 sg13g2_fill_2 FILLER_39_354 ();
 sg13g2_fill_2 FILLER_39_360 ();
 sg13g2_fill_1 FILLER_39_375 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_4 FILLER_40_105 ();
 sg13g2_fill_2 FILLER_40_152 ();
 sg13g2_fill_1 FILLER_40_154 ();
 sg13g2_fill_1 FILLER_40_165 ();
 sg13g2_fill_1 FILLER_40_175 ();
 sg13g2_fill_1 FILLER_40_248 ();
 sg13g2_fill_1 FILLER_40_274 ();
 sg13g2_fill_2 FILLER_40_298 ();
 sg13g2_fill_1 FILLER_40_329 ();
 sg13g2_fill_2 FILLER_40_385 ();
 sg13g2_fill_1 FILLER_40_387 ();
 sg13g2_decap_8 FILLER_40_397 ();
 sg13g2_decap_4 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_4 FILLER_41_98 ();
 sg13g2_fill_2 FILLER_41_119 ();
 sg13g2_fill_1 FILLER_41_130 ();
 sg13g2_fill_2 FILLER_41_136 ();
 sg13g2_fill_2 FILLER_41_164 ();
 sg13g2_fill_1 FILLER_41_176 ();
 sg13g2_fill_1 FILLER_41_191 ();
 sg13g2_fill_2 FILLER_41_211 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_fill_2 FILLER_41_231 ();
 sg13g2_decap_4 FILLER_41_238 ();
 sg13g2_fill_1 FILLER_41_249 ();
 sg13g2_fill_2 FILLER_41_276 ();
 sg13g2_fill_1 FILLER_41_309 ();
 sg13g2_fill_2 FILLER_41_381 ();
 sg13g2_decap_8 FILLER_41_389 ();
 sg13g2_decap_4 FILLER_41_405 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_4 FILLER_42_91 ();
 sg13g2_fill_2 FILLER_42_95 ();
 sg13g2_fill_1 FILLER_42_153 ();
 sg13g2_fill_1 FILLER_42_180 ();
 sg13g2_fill_2 FILLER_42_201 ();
 sg13g2_decap_4 FILLER_42_207 ();
 sg13g2_fill_1 FILLER_42_211 ();
 sg13g2_fill_2 FILLER_42_225 ();
 sg13g2_fill_1 FILLER_42_227 ();
 sg13g2_fill_2 FILLER_42_285 ();
 sg13g2_fill_1 FILLER_42_352 ();
 sg13g2_fill_1 FILLER_42_379 ();
 sg13g2_decap_8 FILLER_42_397 ();
 sg13g2_decap_4 FILLER_42_404 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_4 FILLER_43_91 ();
 sg13g2_fill_1 FILLER_43_95 ();
 sg13g2_fill_2 FILLER_43_126 ();
 sg13g2_fill_2 FILLER_43_172 ();
 sg13g2_fill_1 FILLER_43_200 ();
 sg13g2_decap_4 FILLER_43_255 ();
 sg13g2_fill_1 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_271 ();
 sg13g2_fill_2 FILLER_43_278 ();
 sg13g2_fill_2 FILLER_43_289 ();
 sg13g2_fill_1 FILLER_43_291 ();
 sg13g2_fill_2 FILLER_43_324 ();
 sg13g2_fill_1 FILLER_43_335 ();
 sg13g2_decap_4 FILLER_43_405 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_4 FILLER_44_84 ();
 sg13g2_fill_2 FILLER_44_141 ();
 sg13g2_fill_1 FILLER_44_160 ();
 sg13g2_decap_8 FILLER_44_170 ();
 sg13g2_fill_2 FILLER_44_177 ();
 sg13g2_fill_1 FILLER_44_179 ();
 sg13g2_fill_1 FILLER_44_206 ();
 sg13g2_fill_1 FILLER_44_212 ();
 sg13g2_fill_1 FILLER_44_245 ();
 sg13g2_decap_8 FILLER_44_260 ();
 sg13g2_decap_8 FILLER_44_267 ();
 sg13g2_decap_8 FILLER_44_274 ();
 sg13g2_decap_8 FILLER_44_281 ();
 sg13g2_fill_1 FILLER_44_288 ();
 sg13g2_decap_4 FILLER_44_296 ();
 sg13g2_fill_1 FILLER_44_320 ();
 sg13g2_fill_2 FILLER_44_359 ();
 sg13g2_fill_1 FILLER_44_369 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_4 FILLER_45_91 ();
 sg13g2_fill_2 FILLER_45_95 ();
 sg13g2_fill_2 FILLER_45_161 ();
 sg13g2_fill_2 FILLER_45_179 ();
 sg13g2_fill_1 FILLER_45_181 ();
 sg13g2_fill_1 FILLER_45_187 ();
 sg13g2_decap_8 FILLER_45_262 ();
 sg13g2_decap_8 FILLER_45_269 ();
 sg13g2_decap_4 FILLER_45_276 ();
 sg13g2_decap_4 FILLER_45_305 ();
 sg13g2_fill_1 FILLER_45_309 ();
 sg13g2_fill_2 FILLER_45_315 ();
 sg13g2_fill_1 FILLER_45_317 ();
 sg13g2_fill_1 FILLER_45_371 ();
 sg13g2_fill_2 FILLER_45_386 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_fill_2 FILLER_46_114 ();
 sg13g2_fill_1 FILLER_46_130 ();
 sg13g2_fill_2 FILLER_46_141 ();
 sg13g2_decap_8 FILLER_46_200 ();
 sg13g2_fill_1 FILLER_46_211 ();
 sg13g2_fill_2 FILLER_46_217 ();
 sg13g2_decap_4 FILLER_46_255 ();
 sg13g2_decap_4 FILLER_46_311 ();
 sg13g2_fill_1 FILLER_46_315 ();
 sg13g2_fill_2 FILLER_46_320 ();
 sg13g2_fill_2 FILLER_46_379 ();
 sg13g2_decap_4 FILLER_46_405 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_fill_1 FILLER_47_112 ();
 sg13g2_decap_4 FILLER_47_155 ();
 sg13g2_fill_1 FILLER_47_159 ();
 sg13g2_decap_4 FILLER_47_174 ();
 sg13g2_fill_2 FILLER_47_178 ();
 sg13g2_fill_2 FILLER_47_193 ();
 sg13g2_fill_1 FILLER_47_195 ();
 sg13g2_decap_4 FILLER_47_205 ();
 sg13g2_fill_2 FILLER_47_209 ();
 sg13g2_fill_1 FILLER_47_214 ();
 sg13g2_decap_4 FILLER_47_220 ();
 sg13g2_fill_2 FILLER_47_246 ();
 sg13g2_fill_1 FILLER_47_248 ();
 sg13g2_fill_2 FILLER_47_303 ();
 sg13g2_fill_1 FILLER_47_393 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_4 FILLER_48_119 ();
 sg13g2_fill_1 FILLER_48_139 ();
 sg13g2_decap_4 FILLER_48_152 ();
 sg13g2_fill_2 FILLER_48_156 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_fill_1 FILLER_48_194 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_fill_2 FILLER_48_245 ();
 sg13g2_fill_2 FILLER_48_267 ();
 sg13g2_fill_1 FILLER_48_278 ();
 sg13g2_fill_2 FILLER_48_328 ();
 sg13g2_fill_2 FILLER_48_341 ();
 sg13g2_fill_1 FILLER_48_343 ();
 sg13g2_fill_2 FILLER_48_349 ();
 sg13g2_fill_1 FILLER_48_351 ();
 sg13g2_fill_2 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_401 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_fill_1 FILLER_49_126 ();
 sg13g2_fill_2 FILLER_49_146 ();
 sg13g2_decap_8 FILLER_49_153 ();
 sg13g2_fill_1 FILLER_49_160 ();
 sg13g2_fill_1 FILLER_49_170 ();
 sg13g2_fill_2 FILLER_49_219 ();
 sg13g2_fill_2 FILLER_49_283 ();
 sg13g2_fill_1 FILLER_49_304 ();
 sg13g2_fill_1 FILLER_49_331 ();
 sg13g2_fill_2 FILLER_49_341 ();
 sg13g2_fill_2 FILLER_49_352 ();
 sg13g2_fill_1 FILLER_49_354 ();
 sg13g2_decap_4 FILLER_49_376 ();
 sg13g2_fill_1 FILLER_49_380 ();
 sg13g2_decap_8 FILLER_49_394 ();
 sg13g2_decap_8 FILLER_49_401 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_4 FILLER_50_105 ();
 sg13g2_fill_2 FILLER_50_109 ();
 sg13g2_fill_1 FILLER_50_137 ();
 sg13g2_fill_2 FILLER_50_167 ();
 sg13g2_fill_1 FILLER_50_169 ();
 sg13g2_decap_4 FILLER_50_175 ();
 sg13g2_fill_2 FILLER_50_250 ();
 sg13g2_fill_2 FILLER_50_265 ();
 sg13g2_fill_1 FILLER_50_272 ();
 sg13g2_fill_1 FILLER_50_377 ();
 sg13g2_decap_8 FILLER_50_381 ();
 sg13g2_decap_8 FILLER_50_388 ();
 sg13g2_decap_8 FILLER_50_395 ();
 sg13g2_decap_8 FILLER_50_402 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_4 FILLER_51_105 ();
 sg13g2_fill_1 FILLER_51_109 ();
 sg13g2_decap_4 FILLER_51_186 ();
 sg13g2_fill_2 FILLER_51_190 ();
 sg13g2_fill_1 FILLER_51_201 ();
 sg13g2_fill_2 FILLER_51_228 ();
 sg13g2_fill_2 FILLER_51_247 ();
 sg13g2_fill_1 FILLER_51_298 ();
 sg13g2_fill_1 FILLER_51_366 ();
 sg13g2_decap_8 FILLER_51_402 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_fill_2 FILLER_52_105 ();
 sg13g2_fill_2 FILLER_52_256 ();
 sg13g2_fill_1 FILLER_52_322 ();
 sg13g2_decap_8 FILLER_52_394 ();
 sg13g2_decap_8 FILLER_52_401 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_4 FILLER_53_98 ();
 sg13g2_fill_1 FILLER_53_102 ();
 sg13g2_fill_1 FILLER_53_207 ();
 sg13g2_decap_8 FILLER_53_250 ();
 sg13g2_decap_8 FILLER_53_257 ();
 sg13g2_decap_4 FILLER_53_264 ();
 sg13g2_decap_8 FILLER_53_401 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_fill_2 FILLER_54_112 ();
 sg13g2_fill_1 FILLER_54_114 ();
 sg13g2_fill_1 FILLER_54_180 ();
 sg13g2_fill_2 FILLER_54_186 ();
 sg13g2_fill_1 FILLER_54_188 ();
 sg13g2_fill_2 FILLER_54_198 ();
 sg13g2_decap_4 FILLER_54_257 ();
 sg13g2_fill_2 FILLER_54_261 ();
 sg13g2_decap_8 FILLER_54_268 ();
 sg13g2_fill_1 FILLER_54_323 ();
 sg13g2_decap_8 FILLER_54_331 ();
 sg13g2_fill_2 FILLER_54_338 ();
 sg13g2_decap_8 FILLER_54_401 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_fill_2 FILLER_55_112 ();
 sg13g2_decap_4 FILLER_55_197 ();
 sg13g2_decap_8 FILLER_55_204 ();
 sg13g2_fill_2 FILLER_55_211 ();
 sg13g2_fill_2 FILLER_55_282 ();
 sg13g2_fill_1 FILLER_55_284 ();
 sg13g2_fill_2 FILLER_55_329 ();
 sg13g2_decap_8 FILLER_55_393 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_fill_2 FILLER_56_171 ();
 sg13g2_decap_4 FILLER_56_204 ();
 sg13g2_decap_4 FILLER_56_220 ();
 sg13g2_fill_1 FILLER_56_228 ();
 sg13g2_fill_1 FILLER_56_289 ();
 sg13g2_fill_2 FILLER_56_344 ();
 sg13g2_fill_1 FILLER_56_378 ();
 sg13g2_decap_8 FILLER_56_388 ();
 sg13g2_decap_8 FILLER_56_395 ();
 sg13g2_decap_8 FILLER_56_402 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_fill_2 FILLER_57_105 ();
 sg13g2_fill_1 FILLER_57_147 ();
 sg13g2_decap_4 FILLER_57_155 ();
 sg13g2_fill_1 FILLER_57_159 ();
 sg13g2_fill_1 FILLER_57_186 ();
 sg13g2_fill_1 FILLER_57_213 ();
 sg13g2_fill_2 FILLER_57_240 ();
 sg13g2_fill_1 FILLER_57_242 ();
 sg13g2_fill_2 FILLER_57_248 ();
 sg13g2_fill_1 FILLER_57_283 ();
 sg13g2_fill_2 FILLER_57_293 ();
 sg13g2_fill_1 FILLER_57_295 ();
 sg13g2_decap_8 FILLER_57_391 ();
 sg13g2_decap_8 FILLER_57_398 ();
 sg13g2_decap_4 FILLER_57_405 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_4 FILLER_58_112 ();
 sg13g2_fill_1 FILLER_58_116 ();
 sg13g2_fill_2 FILLER_58_130 ();
 sg13g2_fill_1 FILLER_58_141 ();
 sg13g2_decap_8 FILLER_58_146 ();
 sg13g2_fill_2 FILLER_58_153 ();
 sg13g2_fill_1 FILLER_58_203 ();
 sg13g2_fill_2 FILLER_58_230 ();
 sg13g2_fill_1 FILLER_58_232 ();
 sg13g2_fill_1 FILLER_58_248 ();
 sg13g2_fill_2 FILLER_58_343 ();
 sg13g2_fill_1 FILLER_58_345 ();
 sg13g2_fill_2 FILLER_58_356 ();
 sg13g2_decap_8 FILLER_58_380 ();
 sg13g2_decap_8 FILLER_58_387 ();
 sg13g2_decap_8 FILLER_58_394 ();
 sg13g2_decap_8 FILLER_58_401 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_4 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_139 ();
 sg13g2_decap_4 FILLER_59_146 ();
 sg13g2_fill_2 FILLER_59_150 ();
 sg13g2_fill_1 FILLER_59_318 ();
 sg13g2_decap_8 FILLER_59_375 ();
 sg13g2_decap_8 FILLER_59_382 ();
 sg13g2_decap_8 FILLER_59_389 ();
 sg13g2_decap_8 FILLER_59_396 ();
 sg13g2_decap_4 FILLER_59_403 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_4 FILLER_60_98 ();
 sg13g2_fill_1 FILLER_60_137 ();
 sg13g2_fill_1 FILLER_60_177 ();
 sg13g2_fill_2 FILLER_60_225 ();
 sg13g2_fill_2 FILLER_60_251 ();
 sg13g2_fill_2 FILLER_60_262 ();
 sg13g2_fill_2 FILLER_60_290 ();
 sg13g2_fill_2 FILLER_60_309 ();
 sg13g2_fill_2 FILLER_60_351 ();
 sg13g2_fill_1 FILLER_60_353 ();
 sg13g2_decap_8 FILLER_60_385 ();
 sg13g2_decap_8 FILLER_60_392 ();
 sg13g2_decap_8 FILLER_60_399 ();
 sg13g2_fill_2 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_4 FILLER_61_98 ();
 sg13g2_fill_1 FILLER_61_102 ();
 sg13g2_fill_1 FILLER_61_159 ();
 sg13g2_fill_1 FILLER_61_185 ();
 sg13g2_fill_1 FILLER_61_229 ();
 sg13g2_fill_2 FILLER_61_335 ();
 sg13g2_decap_8 FILLER_61_391 ();
 sg13g2_decap_8 FILLER_61_398 ();
 sg13g2_decap_4 FILLER_61_405 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_fill_1 FILLER_62_143 ();
 sg13g2_decap_8 FILLER_62_174 ();
 sg13g2_fill_1 FILLER_62_181 ();
 sg13g2_fill_1 FILLER_62_208 ();
 sg13g2_fill_2 FILLER_62_232 ();
 sg13g2_fill_2 FILLER_62_247 ();
 sg13g2_fill_2 FILLER_62_284 ();
 sg13g2_fill_1 FILLER_62_346 ();
 sg13g2_decap_8 FILLER_62_386 ();
 sg13g2_decap_8 FILLER_62_393 ();
 sg13g2_decap_8 FILLER_62_400 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_fill_1 FILLER_63_98 ();
 sg13g2_fill_2 FILLER_63_247 ();
 sg13g2_fill_1 FILLER_63_249 ();
 sg13g2_fill_2 FILLER_63_255 ();
 sg13g2_fill_2 FILLER_63_262 ();
 sg13g2_fill_1 FILLER_63_264 ();
 sg13g2_fill_1 FILLER_63_283 ();
 sg13g2_fill_1 FILLER_63_288 ();
 sg13g2_fill_2 FILLER_63_307 ();
 sg13g2_decap_8 FILLER_63_371 ();
 sg13g2_decap_8 FILLER_63_378 ();
 sg13g2_decap_8 FILLER_63_385 ();
 sg13g2_decap_8 FILLER_63_392 ();
 sg13g2_decap_8 FILLER_63_399 ();
 sg13g2_fill_2 FILLER_63_406 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_fill_1 FILLER_64_98 ();
 sg13g2_fill_2 FILLER_64_137 ();
 sg13g2_fill_1 FILLER_64_149 ();
 sg13g2_fill_2 FILLER_64_197 ();
 sg13g2_fill_1 FILLER_64_217 ();
 sg13g2_fill_1 FILLER_64_226 ();
 sg13g2_fill_2 FILLER_64_236 ();
 sg13g2_fill_1 FILLER_64_238 ();
 sg13g2_fill_2 FILLER_64_249 ();
 sg13g2_fill_2 FILLER_64_271 ();
 sg13g2_fill_1 FILLER_64_303 ();
 sg13g2_fill_2 FILLER_64_353 ();
 sg13g2_decap_8 FILLER_64_365 ();
 sg13g2_decap_8 FILLER_64_372 ();
 sg13g2_decap_8 FILLER_64_379 ();
 sg13g2_decap_8 FILLER_64_386 ();
 sg13g2_decap_8 FILLER_64_393 ();
 sg13g2_decap_8 FILLER_64_400 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_fill_1 FILLER_65_105 ();
 sg13g2_fill_2 FILLER_65_136 ();
 sg13g2_fill_2 FILLER_65_260 ();
 sg13g2_fill_1 FILLER_65_266 ();
 sg13g2_fill_1 FILLER_65_280 ();
 sg13g2_fill_1 FILLER_65_300 ();
 sg13g2_fill_2 FILLER_65_359 ();
 sg13g2_decap_8 FILLER_65_373 ();
 sg13g2_decap_8 FILLER_65_380 ();
 sg13g2_decap_8 FILLER_65_387 ();
 sg13g2_decap_8 FILLER_65_394 ();
 sg13g2_decap_8 FILLER_65_401 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_fill_1 FILLER_66_112 ();
 sg13g2_fill_1 FILLER_66_147 ();
 sg13g2_fill_1 FILLER_66_188 ();
 sg13g2_fill_1 FILLER_66_250 ();
 sg13g2_fill_2 FILLER_66_334 ();
 sg13g2_decap_8 FILLER_66_371 ();
 sg13g2_decap_8 FILLER_66_378 ();
 sg13g2_decap_8 FILLER_66_385 ();
 sg13g2_decap_8 FILLER_66_392 ();
 sg13g2_decap_8 FILLER_66_399 ();
 sg13g2_fill_2 FILLER_66_406 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_4 FILLER_67_112 ();
 sg13g2_fill_1 FILLER_67_116 ();
 sg13g2_fill_2 FILLER_67_150 ();
 sg13g2_fill_1 FILLER_67_183 ();
 sg13g2_fill_2 FILLER_67_230 ();
 sg13g2_fill_1 FILLER_67_232 ();
 sg13g2_decap_4 FILLER_67_237 ();
 sg13g2_fill_1 FILLER_67_241 ();
 sg13g2_fill_2 FILLER_67_260 ();
 sg13g2_fill_1 FILLER_67_262 ();
 sg13g2_decap_8 FILLER_67_374 ();
 sg13g2_decap_8 FILLER_67_381 ();
 sg13g2_decap_8 FILLER_67_388 ();
 sg13g2_decap_8 FILLER_67_395 ();
 sg13g2_decap_8 FILLER_67_402 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_fill_2 FILLER_68_112 ();
 sg13g2_fill_1 FILLER_68_174 ();
 sg13g2_fill_1 FILLER_68_201 ();
 sg13g2_decap_8 FILLER_68_228 ();
 sg13g2_decap_8 FILLER_68_235 ();
 sg13g2_fill_2 FILLER_68_246 ();
 sg13g2_fill_1 FILLER_68_248 ();
 sg13g2_fill_2 FILLER_68_258 ();
 sg13g2_fill_1 FILLER_68_335 ();
 sg13g2_decap_8 FILLER_68_365 ();
 sg13g2_decap_8 FILLER_68_372 ();
 sg13g2_decap_8 FILLER_68_379 ();
 sg13g2_decap_8 FILLER_68_386 ();
 sg13g2_decap_8 FILLER_68_393 ();
 sg13g2_decap_8 FILLER_68_400 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_4 FILLER_69_98 ();
 sg13g2_fill_2 FILLER_69_128 ();
 sg13g2_fill_1 FILLER_69_152 ();
 sg13g2_fill_2 FILLER_69_181 ();
 sg13g2_decap_8 FILLER_69_230 ();
 sg13g2_fill_1 FILLER_69_237 ();
 sg13g2_fill_2 FILLER_69_281 ();
 sg13g2_fill_1 FILLER_69_297 ();
 sg13g2_decap_8 FILLER_69_325 ();
 sg13g2_decap_4 FILLER_69_332 ();
 sg13g2_fill_1 FILLER_69_336 ();
 sg13g2_fill_2 FILLER_69_351 ();
 sg13g2_decap_8 FILLER_69_370 ();
 sg13g2_decap_8 FILLER_69_377 ();
 sg13g2_decap_8 FILLER_69_384 ();
 sg13g2_decap_8 FILLER_69_391 ();
 sg13g2_decap_8 FILLER_69_398 ();
 sg13g2_decap_4 FILLER_69_405 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_fill_1 FILLER_70_124 ();
 sg13g2_fill_1 FILLER_70_141 ();
 sg13g2_fill_2 FILLER_70_157 ();
 sg13g2_fill_1 FILLER_70_159 ();
 sg13g2_fill_1 FILLER_70_173 ();
 sg13g2_fill_2 FILLER_70_182 ();
 sg13g2_fill_2 FILLER_70_224 ();
 sg13g2_decap_8 FILLER_70_265 ();
 sg13g2_fill_2 FILLER_70_272 ();
 sg13g2_fill_1 FILLER_70_274 ();
 sg13g2_fill_1 FILLER_70_301 ();
 sg13g2_fill_1 FILLER_70_307 ();
 sg13g2_decap_4 FILLER_70_334 ();
 sg13g2_fill_2 FILLER_70_338 ();
 sg13g2_decap_8 FILLER_70_363 ();
 sg13g2_decap_8 FILLER_70_370 ();
 sg13g2_decap_8 FILLER_70_377 ();
 sg13g2_decap_8 FILLER_70_384 ();
 sg13g2_decap_8 FILLER_70_391 ();
 sg13g2_decap_8 FILLER_70_398 ();
 sg13g2_decap_4 FILLER_70_405 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_4 FILLER_71_91 ();
 sg13g2_fill_2 FILLER_71_95 ();
 sg13g2_fill_1 FILLER_71_155 ();
 sg13g2_fill_1 FILLER_71_179 ();
 sg13g2_fill_2 FILLER_71_213 ();
 sg13g2_fill_2 FILLER_71_257 ();
 sg13g2_fill_1 FILLER_71_259 ();
 sg13g2_decap_8 FILLER_71_269 ();
 sg13g2_decap_8 FILLER_71_276 ();
 sg13g2_decap_4 FILLER_71_283 ();
 sg13g2_fill_1 FILLER_71_292 ();
 sg13g2_fill_1 FILLER_71_327 ();
 sg13g2_decap_8 FILLER_71_357 ();
 sg13g2_decap_8 FILLER_71_364 ();
 sg13g2_decap_8 FILLER_71_371 ();
 sg13g2_decap_8 FILLER_71_378 ();
 sg13g2_decap_8 FILLER_71_385 ();
 sg13g2_decap_8 FILLER_71_392 ();
 sg13g2_decap_8 FILLER_71_399 ();
 sg13g2_fill_2 FILLER_71_406 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_fill_2 FILLER_72_98 ();
 sg13g2_fill_2 FILLER_72_126 ();
 sg13g2_fill_2 FILLER_72_221 ();
 sg13g2_fill_1 FILLER_72_230 ();
 sg13g2_fill_1 FILLER_72_253 ();
 sg13g2_decap_8 FILLER_72_276 ();
 sg13g2_fill_2 FILLER_72_283 ();
 sg13g2_fill_1 FILLER_72_285 ();
 sg13g2_decap_8 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_371 ();
 sg13g2_decap_8 FILLER_72_378 ();
 sg13g2_decap_8 FILLER_72_385 ();
 sg13g2_decap_8 FILLER_72_392 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_fill_2 FILLER_72_406 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_fill_2 FILLER_73_98 ();
 sg13g2_fill_1 FILLER_73_100 ();
 sg13g2_fill_2 FILLER_73_132 ();
 sg13g2_fill_2 FILLER_73_210 ();
 sg13g2_decap_8 FILLER_73_221 ();
 sg13g2_fill_1 FILLER_73_228 ();
 sg13g2_fill_1 FILLER_73_277 ();
 sg13g2_fill_1 FILLER_73_330 ();
 sg13g2_fill_2 FILLER_73_336 ();
 sg13g2_decap_8 FILLER_73_373 ();
 sg13g2_decap_8 FILLER_73_380 ();
 sg13g2_decap_8 FILLER_73_387 ();
 sg13g2_decap_8 FILLER_73_394 ();
 sg13g2_decap_8 FILLER_73_401 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_4 FILLER_74_98 ();
 sg13g2_fill_1 FILLER_74_102 ();
 sg13g2_fill_2 FILLER_74_138 ();
 sg13g2_fill_2 FILLER_74_205 ();
 sg13g2_fill_1 FILLER_74_310 ();
 sg13g2_fill_2 FILLER_74_338 ();
 sg13g2_decap_8 FILLER_74_374 ();
 sg13g2_decap_8 FILLER_74_381 ();
 sg13g2_decap_8 FILLER_74_388 ();
 sg13g2_decap_8 FILLER_74_395 ();
 sg13g2_decap_8 FILLER_74_402 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_fill_1 FILLER_75_112 ();
 sg13g2_fill_1 FILLER_75_120 ();
 sg13g2_fill_2 FILLER_75_126 ();
 sg13g2_fill_1 FILLER_75_135 ();
 sg13g2_fill_1 FILLER_75_146 ();
 sg13g2_fill_1 FILLER_75_161 ();
 sg13g2_fill_2 FILLER_75_166 ();
 sg13g2_fill_2 FILLER_75_183 ();
 sg13g2_fill_2 FILLER_75_194 ();
 sg13g2_decap_8 FILLER_75_200 ();
 sg13g2_fill_2 FILLER_75_207 ();
 sg13g2_fill_1 FILLER_75_209 ();
 sg13g2_fill_2 FILLER_75_236 ();
 sg13g2_fill_1 FILLER_75_238 ();
 sg13g2_decap_8 FILLER_75_368 ();
 sg13g2_decap_8 FILLER_75_375 ();
 sg13g2_decap_8 FILLER_75_382 ();
 sg13g2_decap_8 FILLER_75_389 ();
 sg13g2_decap_8 FILLER_75_396 ();
 sg13g2_decap_4 FILLER_75_403 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_4 FILLER_76_112 ();
 sg13g2_fill_2 FILLER_76_116 ();
 sg13g2_decap_8 FILLER_76_193 ();
 sg13g2_decap_8 FILLER_76_200 ();
 sg13g2_fill_2 FILLER_76_207 ();
 sg13g2_fill_1 FILLER_76_209 ();
 sg13g2_fill_1 FILLER_76_251 ();
 sg13g2_fill_2 FILLER_76_301 ();
 sg13g2_fill_1 FILLER_76_303 ();
 sg13g2_decap_4 FILLER_76_313 ();
 sg13g2_fill_1 FILLER_76_317 ();
 sg13g2_fill_2 FILLER_76_332 ();
 sg13g2_decap_8 FILLER_76_356 ();
 sg13g2_decap_8 FILLER_76_363 ();
 sg13g2_decap_8 FILLER_76_370 ();
 sg13g2_decap_8 FILLER_76_377 ();
 sg13g2_decap_8 FILLER_76_384 ();
 sg13g2_decap_8 FILLER_76_391 ();
 sg13g2_decap_8 FILLER_76_398 ();
 sg13g2_decap_4 FILLER_76_405 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_fill_1 FILLER_77_112 ();
 sg13g2_fill_1 FILLER_77_132 ();
 sg13g2_fill_1 FILLER_77_159 ();
 sg13g2_fill_1 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_199 ();
 sg13g2_decap_4 FILLER_77_206 ();
 sg13g2_fill_2 FILLER_77_222 ();
 sg13g2_fill_1 FILLER_77_275 ();
 sg13g2_decap_4 FILLER_77_302 ();
 sg13g2_fill_2 FILLER_77_320 ();
 sg13g2_fill_1 FILLER_77_330 ();
 sg13g2_decap_8 FILLER_77_345 ();
 sg13g2_decap_8 FILLER_77_352 ();
 sg13g2_decap_8 FILLER_77_359 ();
 sg13g2_decap_8 FILLER_77_366 ();
 sg13g2_decap_8 FILLER_77_373 ();
 sg13g2_decap_8 FILLER_77_380 ();
 sg13g2_decap_8 FILLER_77_387 ();
 sg13g2_decap_8 FILLER_77_394 ();
 sg13g2_decap_8 FILLER_77_401 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_4 FILLER_78_112 ();
 sg13g2_fill_2 FILLER_78_116 ();
 sg13g2_decap_8 FILLER_78_205 ();
 sg13g2_decap_4 FILLER_78_212 ();
 sg13g2_fill_2 FILLER_78_216 ();
 sg13g2_fill_1 FILLER_78_280 ();
 sg13g2_decap_8 FILLER_78_359 ();
 sg13g2_decap_8 FILLER_78_366 ();
 sg13g2_decap_8 FILLER_78_373 ();
 sg13g2_decap_8 FILLER_78_380 ();
 sg13g2_decap_8 FILLER_78_387 ();
 sg13g2_decap_8 FILLER_78_394 ();
 sg13g2_decap_8 FILLER_78_401 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_fill_1 FILLER_79_133 ();
 sg13g2_fill_1 FILLER_79_138 ();
 sg13g2_fill_2 FILLER_79_148 ();
 sg13g2_fill_1 FILLER_79_164 ();
 sg13g2_fill_1 FILLER_79_174 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_4 FILLER_79_224 ();
 sg13g2_fill_1 FILLER_79_228 ();
 sg13g2_fill_2 FILLER_79_233 ();
 sg13g2_fill_1 FILLER_79_235 ();
 sg13g2_fill_1 FILLER_79_276 ();
 sg13g2_fill_1 FILLER_79_281 ();
 sg13g2_decap_8 FILLER_79_356 ();
 sg13g2_decap_8 FILLER_79_363 ();
 sg13g2_decap_8 FILLER_79_370 ();
 sg13g2_decap_8 FILLER_79_377 ();
 sg13g2_decap_8 FILLER_79_384 ();
 sg13g2_decap_8 FILLER_79_391 ();
 sg13g2_decap_8 FILLER_79_398 ();
 sg13g2_decap_4 FILLER_79_405 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_fill_2 FILLER_80_156 ();
 sg13g2_fill_1 FILLER_80_158 ();
 sg13g2_fill_1 FILLER_80_167 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_4 FILLER_80_187 ();
 sg13g2_fill_1 FILLER_80_191 ();
 sg13g2_decap_4 FILLER_80_196 ();
 sg13g2_decap_4 FILLER_80_204 ();
 sg13g2_decap_4 FILLER_80_212 ();
 sg13g2_decap_4 FILLER_80_220 ();
 sg13g2_decap_4 FILLER_80_228 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_decap_8 FILLER_80_243 ();
 sg13g2_decap_8 FILLER_80_267 ();
 sg13g2_decap_8 FILLER_80_274 ();
 sg13g2_decap_8 FILLER_80_281 ();
 sg13g2_decap_8 FILLER_80_288 ();
 sg13g2_decap_4 FILLER_80_308 ();
 sg13g2_decap_8 FILLER_80_316 ();
 sg13g2_fill_1 FILLER_80_323 ();
 sg13g2_decap_8 FILLER_80_337 ();
 sg13g2_decap_8 FILLER_80_344 ();
 sg13g2_decap_8 FILLER_80_351 ();
 sg13g2_decap_8 FILLER_80_358 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_372 ();
 sg13g2_decap_8 FILLER_80_379 ();
 sg13g2_decap_8 FILLER_80_386 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_8 FILLER_80_400 ();
 sg13g2_fill_2 FILLER_80_407 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
 assign uo_out[1] = net18;
 assign uo_out[2] = net19;
 assign uo_out[3] = net20;
 assign uo_out[4] = net21;
 assign uo_out[5] = net22;
 assign uo_out[6] = net23;
endmodule

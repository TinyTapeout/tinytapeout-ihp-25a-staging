module tt_um_wokwi_412635532198550529 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire \and1.b ;
 wire \and10.a ;
 wire \and100.a ;
 wire \and101.a ;
 wire \and102.a ;
 wire \and104.b ;
 wire \and106.a ;
 wire \and107.b ;
 wire \and108.b ;
 wire \and11.b ;
 wire \and110.b ;
 wire \and112.a ;
 wire \and113.a ;
 wire \and115.b ;
 wire \and116.a ;
 wire \and118.a ;
 wire \and119.a ;
 wire \and122.a ;
 wire \and125.a ;
 wire \and126.a ;
 wire \and127.a ;
 wire \and128.b ;
 wire \and129.a ;
 wire \and131.b ;
 wire \and73.a ;
 wire \and74.a ;
 wire \and74.b ;
 wire \and75.a ;
 wire \and76.a ;
 wire \and81.b ;
 wire \and82.a ;
 wire \and83.a ;
 wire \and83.b ;
 wire \and84.a ;
 wire \and85.a ;
 wire \and86.a ;
 wire \and92.a ;
 wire \and93.a ;
 wire \and94.a ;
 wire \flop10.d ;
 wire \flop10.q ;
 wire \flop11.q ;
 wire \flop12.d ;
 wire \flop12.q ;
 wire \flop13.d ;
 wire \flop13.q ;
 wire \flop14.d ;
 wire \flop14.q ;
 wire \flop15.d ;
 wire \flop15.q ;
 wire \flop16.d ;
 wire \flop16.q ;
 wire \flop17.d ;
 wire \flop17.q ;
 wire \flop18.d ;
 wire \flop18.q ;
 wire \flop19.d ;
 wire \flop20.notq ;
 wire \flop21.notq ;
 wire \flop22.notq ;
 wire \flop23.notq ;
 wire \flop24.notq ;
 wire \flop25.q ;
 wire \flop26.q ;
 wire \flop27.d ;
 wire \flop28.notq ;
 wire \flop29.notq ;
 wire \flop30.notq ;
 wire \flop31.notq ;
 wire \flop32.notq ;
 wire \flop33.notq ;
 wire \flop34.notq ;
 wire \flop35.notq ;
 wire \flop36.notq ;
 wire \flop37.notq ;
 wire \flop38.notq ;
 wire \flop39.notq ;
 wire \flop40.notq ;
 wire \flop42.notq ;
 wire \flop43.q ;
 wire \flop44.q ;
 wire \flop45.q ;
 wire \flop46.q ;
 wire \flop47.q ;
 wire \flop48.q ;
 wire \flop49.q ;
 wire \flop50.q ;
 wire \flop51.q ;
 wire \flop52.q ;
 wire \flop53.q ;
 wire \flop54.q ;
 wire \flop55.q ;
 wire \flop56.q ;
 wire \flop57.q ;
 wire \flop58.q ;
 wire \flop59.q ;
 wire \flop60.q ;
 wire \flop61.q ;
 wire \flop62.q ;
 wire \flop63.q ;
 wire \flop64.q ;
 wire \flop65.q ;
 wire \flop66.q ;
 wire \flop67.q ;
 wire \flop68.q ;
 wire \flop69.q ;
 wire \flop70.q ;
 wire \flop71.q ;
 wire \flop72.q ;
 wire \flop73.q ;
 wire \flop74.q ;
 wire \flop83.d ;
 wire \flop83.q ;
 wire \flop84.q ;
 wire \flop85.q ;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net26;
 wire clknet_0_clk;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net216;

 sg13g2_inv_1 _0559_ (.Y(_0092_),
    .A(net48));
 sg13g2_inv_1 _0560_ (.Y(_0093_),
    .A(net50));
 sg13g2_inv_1 _0561_ (.Y(_0094_),
    .A(net184));
 sg13g2_inv_1 _0562_ (.Y(_0095_),
    .A(net188));
 sg13g2_inv_1 _0563_ (.Y(_0096_),
    .A(net191));
 sg13g2_inv_1 _0564_ (.Y(_0097_),
    .A(_0000_));
 sg13g2_inv_1 _0565_ (.Y(_0098_),
    .A(\and128.b ));
 sg13g2_inv_2 _0566_ (.Y(_0099_),
    .A(net156));
 sg13g2_inv_1 _0567_ (.Y(_0100_),
    .A(\flop66.q ));
 sg13g2_inv_1 _0568_ (.Y(_0101_),
    .A(\flop74.q ));
 sg13g2_inv_1 _0569_ (.Y(_0102_),
    .A(\flop50.q ));
 sg13g2_inv_1 _0570_ (.Y(_0103_),
    .A(\flop58.q ));
 sg13g2_inv_1 _0571_ (.Y(_0104_),
    .A(net135));
 sg13g2_inv_1 _0572_ (.Y(_0105_),
    .A(\and126.a ));
 sg13g2_inv_1 _0573_ (.Y(_0106_),
    .A(_0003_));
 sg13g2_inv_1 _0574_ (.Y(_0107_),
    .A(_0004_));
 sg13g2_inv_1 _0575_ (.Y(_0108_),
    .A(_0005_));
 sg13g2_inv_1 _0576_ (.Y(_0109_),
    .A(net5));
 sg13g2_inv_1 _0577_ (.Y(_0110_),
    .A(net144));
 sg13g2_inv_2 _0578_ (.Y(_0111_),
    .A(_0006_));
 sg13g2_inv_1 _0579_ (.Y(_0112_),
    .A(net4));
 sg13g2_inv_1 _0580_ (.Y(_0113_),
    .A(net146));
 sg13g2_inv_2 _0581_ (.Y(_0114_),
    .A(net133));
 sg13g2_inv_1 _0582_ (.Y(_0115_),
    .A(_0008_));
 sg13g2_inv_1 _0583_ (.Y(_0116_),
    .A(net3));
 sg13g2_inv_1 _0584_ (.Y(_0117_),
    .A(_0009_));
 sg13g2_inv_1 _0585_ (.Y(_0118_),
    .A(_0011_));
 sg13g2_inv_1 _0586_ (.Y(_0119_),
    .A(_0010_));
 sg13g2_inv_1 _0587_ (.Y(_0120_),
    .A(_0013_));
 sg13g2_inv_1 _0588_ (.Y(_0121_),
    .A(_0012_));
 sg13g2_inv_1 _0589_ (.Y(_0122_),
    .A(net1));
 sg13g2_inv_1 _0590_ (.Y(_0123_),
    .A(net46));
 sg13g2_inv_1 _0591_ (.Y(_0124_),
    .A(net39));
 sg13g2_inv_1 _0592_ (.Y(_0125_),
    .A(\flop31.notq ));
 sg13g2_inv_2 _0593_ (.Y(_0126_),
    .A(net31));
 sg13g2_nand3b_1 _0594_ (.B(\and74.a ),
    .C(\and74.b ),
    .Y(_0127_),
    .A_N(\flop21.notq ));
 sg13g2_nor2_1 _0595_ (.A(\flop22.notq ),
    .B(_0127_),
    .Y(_0128_));
 sg13g2_nor3_2 _0596_ (.A(\flop23.notq ),
    .B(\flop22.notq ),
    .C(_0127_),
    .Y(_0129_));
 sg13g2_nor2b_1 _0597_ (.A(net93),
    .B_N(_0129_),
    .Y(_0130_));
 sg13g2_nor2_1 _0598_ (.A(net70),
    .B(_0129_),
    .Y(_0131_));
 sg13g2_nor2_1 _0599_ (.A(_0130_),
    .B(net71),
    .Y(_0080_));
 sg13g2_nor2_1 _0600_ (.A(net67),
    .B(_0128_),
    .Y(_0132_));
 sg13g2_nor2_1 _0601_ (.A(_0129_),
    .B(net68),
    .Y(_0079_));
 sg13g2_a21oi_1 _0602_ (.A1(_0092_),
    .A2(_0127_),
    .Y(_0078_),
    .B1(_0128_));
 sg13g2_a21o_1 _0603_ (.A2(\and74.b ),
    .A1(\and74.a ),
    .B1(net140),
    .X(_0133_));
 sg13g2_and2_1 _0604_ (.A(_0127_),
    .B(net141),
    .X(_0077_));
 sg13g2_mux2_1 _0605_ (.A0(\and74.a ),
    .A1(net34),
    .S(\and74.b ),
    .X(_0076_));
 sg13g2_nor2_1 _0606_ (.A(net154),
    .B(net197),
    .Y(_0134_));
 sg13g2_nand2_2 _0607_ (.Y(_0135_),
    .A(net186),
    .B(net189));
 sg13g2_nor4_2 _0608_ (.A(net182),
    .B(net184),
    .C(_0001_),
    .Y(_0136_),
    .D(_0135_));
 sg13g2_or4_1 _0609_ (.A(net182),
    .B(net185),
    .C(_0001_),
    .D(_0135_),
    .X(_0137_));
 sg13g2_nand2_1 _0610_ (.Y(_0138_),
    .A(net185),
    .B(net189));
 sg13g2_mux2_2 _0611_ (.A0(\and128.b ),
    .A1(net193),
    .S(_0138_),
    .X(_0139_));
 sg13g2_mux2_2 _0612_ (.A0(\and131.b ),
    .A1(\and115.b ),
    .S(_0138_),
    .X(_0140_));
 sg13g2_mux4_1 _0613_ (.S0(net176),
    .A0(_0120_),
    .A1(_0121_),
    .A2(_0118_),
    .A3(_0119_),
    .S1(net175),
    .X(_0141_));
 sg13g2_mux4_1 _0614_ (.S0(net176),
    .A0(_0013_),
    .A1(_0012_),
    .A2(_0011_),
    .A3(_0010_),
    .S1(net175),
    .X(_0142_));
 sg13g2_a21oi_1 _0615_ (.A1(_0117_),
    .A2(_0141_),
    .Y(_0143_),
    .B1(_0137_));
 sg13g2_nor4_2 _0616_ (.A(net182),
    .B(net184),
    .C(_0000_),
    .Y(_0144_),
    .D(_0135_));
 sg13g2_or4_2 _0617_ (.A(net182),
    .B(net184),
    .C(_0000_),
    .D(_0135_),
    .X(_0145_));
 sg13g2_mux4_1 _0618_ (.S0(net176),
    .A0(\flop43.q ),
    .A1(\flop51.q ),
    .A2(\flop59.q ),
    .A3(\flop67.q ),
    .S1(net175),
    .X(_0146_));
 sg13g2_o21ai_1 _0619_ (.B1(_0144_),
    .Y(_0147_),
    .A1(_0117_),
    .A2(_0146_));
 sg13g2_or2_1 _0620_ (.X(_0148_),
    .B(_0147_),
    .A(_0143_));
 sg13g2_nand2_1 _0621_ (.Y(_0149_),
    .A(\and116.a ),
    .B(_0136_));
 sg13g2_xnor2_1 _0622_ (.Y(_0150_),
    .A(_0141_),
    .B(_0149_));
 sg13g2_nand2_1 _0623_ (.Y(_0151_),
    .A(\and129.a ),
    .B(\and112.a ));
 sg13g2_nor2_1 _0624_ (.A(net184),
    .B(_0151_),
    .Y(_0152_));
 sg13g2_nand2b_1 _0625_ (.Y(_0153_),
    .B(_0094_),
    .A_N(_0151_));
 sg13g2_nor2_2 _0626_ (.A(_0095_),
    .B(_0152_),
    .Y(_0154_));
 sg13g2_inv_1 _0627_ (.Y(_0155_),
    .A(_0154_));
 sg13g2_a21oi_1 _0628_ (.A1(_0145_),
    .A2(_0150_),
    .Y(_0156_),
    .B1(_0155_));
 sg13g2_nand2_1 _0629_ (.Y(_0157_),
    .A(net181),
    .B(_0122_));
 sg13g2_nor2b_2 _0630_ (.A(\and128.b ),
    .B_N(net194),
    .Y(_0158_));
 sg13g2_nand2b_1 _0631_ (.Y(_0159_),
    .B(_0158_),
    .A_N(net183));
 sg13g2_o21ai_1 _0632_ (.B1(_0159_),
    .Y(_0160_),
    .A1(net178),
    .A2(_0146_));
 sg13g2_nand3_1 _0633_ (.B(net182),
    .C(net188),
    .A(net186),
    .Y(_0161_));
 sg13g2_nor2_2 _0634_ (.A(net184),
    .B(_0161_),
    .Y(_0162_));
 sg13g2_nand2_1 _0635_ (.Y(_0163_),
    .A(net188),
    .B(_0152_));
 sg13g2_nand2_1 _0636_ (.Y(_0164_),
    .A(_0098_),
    .B(\flop84.q ));
 sg13g2_o21ai_1 _0637_ (.B1(\and131.b ),
    .Y(_0165_),
    .A1(net194),
    .A2(_0115_));
 sg13g2_a21oi_1 _0638_ (.A1(net193),
    .A2(_0164_),
    .Y(_0166_),
    .B1(_0165_));
 sg13g2_nand2b_1 _0639_ (.Y(_0167_),
    .B(_0162_),
    .A_N(_0166_));
 sg13g2_a21oi_1 _0640_ (.A1(net180),
    .A2(_0160_),
    .Y(_0168_),
    .B1(_0167_));
 sg13g2_a221oi_1 _0641_ (.B2(_0156_),
    .C1(_0168_),
    .B1(_0148_),
    .A1(net181),
    .Y(_0169_),
    .A2(_0122_));
 sg13g2_nor2_1 _0642_ (.A(net184),
    .B(net180),
    .Y(_0170_));
 sg13g2_nor3_2 _0643_ (.A(net184),
    .B(net179),
    .C(_0104_),
    .Y(_0171_));
 sg13g2_a21oi_1 _0644_ (.A1(net183),
    .A2(_0171_),
    .Y(_0172_),
    .B1(net186));
 sg13g2_o21ai_1 _0645_ (.B1(_0172_),
    .Y(_0173_),
    .A1(net183),
    .A2(_0171_));
 sg13g2_xnor2_1 _0646_ (.Y(_0174_),
    .A(_0169_),
    .B(_0173_));
 sg13g2_a21oi_2 _0647_ (.B1(_0134_),
    .Y(_0175_),
    .A2(_0174_),
    .A1(net197));
 sg13g2_nor2_1 _0648_ (.A(\and106.a ),
    .B(net11),
    .Y(_0176_));
 sg13g2_a21oi_2 _0649_ (.B1(_0176_),
    .Y(_0177_),
    .A2(net11),
    .A1(net10));
 sg13g2_nand2b_2 _0650_ (.Y(_0178_),
    .B(net182),
    .A_N(net186));
 sg13g2_a21oi_1 _0651_ (.A1(_0000_),
    .A2(_0160_),
    .Y(_0179_),
    .B1(_0167_));
 sg13g2_a21oi_1 _0652_ (.A1(_0009_),
    .A2(_0142_),
    .Y(_0180_),
    .B1(_0144_));
 sg13g2_nand2b_1 _0653_ (.Y(_0181_),
    .B(_0142_),
    .A_N(_0001_));
 sg13g2_and2_1 _0654_ (.A(net183),
    .B(_0144_),
    .X(_0182_));
 sg13g2_a21o_1 _0655_ (.A2(_0146_),
    .A1(net177),
    .B1(_0162_),
    .X(_0183_));
 sg13g2_a221oi_1 _0656_ (.B2(_0182_),
    .C1(_0183_),
    .B1(_0181_),
    .A1(_0143_),
    .Y(_0184_),
    .A2(_0180_));
 sg13g2_o21ai_1 _0657_ (.B1(net189),
    .Y(_0185_),
    .A1(_0179_),
    .A2(_0184_));
 sg13g2_mux4_1 _0658_ (.S0(_0139_),
    .A0(\flop44.q ),
    .A1(\flop52.q ),
    .A2(\flop60.q ),
    .A3(\flop68.q ),
    .S1(_0140_),
    .X(_0186_));
 sg13g2_a21o_1 _0659_ (.A2(_0186_),
    .A1(_0115_),
    .B1(_0144_),
    .X(_0187_));
 sg13g2_nor2_1 _0660_ (.A(_0114_),
    .B(_0145_),
    .Y(_0188_));
 sg13g2_a21oi_1 _0661_ (.A1(_0186_),
    .A2(_0188_),
    .Y(_0189_),
    .B1(net177));
 sg13g2_nand2_2 _0662_ (.Y(_0190_),
    .A(net177),
    .B(_0145_));
 sg13g2_a21oi_1 _0663_ (.A1(net177),
    .A2(_0145_),
    .Y(_0191_),
    .B1(_0008_));
 sg13g2_o21ai_1 _0664_ (.B1(_0154_),
    .Y(_0192_),
    .A1(_0186_),
    .A2(_0191_));
 sg13g2_a21oi_1 _0665_ (.A1(_0187_),
    .A2(_0189_),
    .Y(_0193_),
    .B1(_0192_));
 sg13g2_a21oi_1 _0666_ (.A1(_0114_),
    .A2(_0158_),
    .Y(_0194_),
    .B1(net191));
 sg13g2_o21ai_1 _0667_ (.B1(_0194_),
    .Y(_0195_),
    .A1(_0098_),
    .A2(_0186_));
 sg13g2_nor2_1 _0668_ (.A(net194),
    .B(_0007_),
    .Y(_0196_));
 sg13g2_a21oi_1 _0669_ (.A1(net194),
    .A2(_0117_),
    .Y(_0197_),
    .B1(_0196_));
 sg13g2_a21oi_1 _0670_ (.A1(net191),
    .A2(_0197_),
    .Y(_0198_),
    .B1(_0163_));
 sg13g2_a22oi_1 _0671_ (.Y(_0199_),
    .B1(_0195_),
    .B2(_0198_),
    .A2(net2),
    .A1(net181));
 sg13g2_nand2b_1 _0672_ (.Y(_0200_),
    .B(_0199_),
    .A_N(_0193_));
 sg13g2_a21oi_1 _0673_ (.A1(_0157_),
    .A2(_0185_),
    .Y(_0201_),
    .B1(_0200_));
 sg13g2_mux4_1 _0674_ (.S0(_0139_),
    .A0(\flop45.q ),
    .A1(\flop53.q ),
    .A2(\flop61.q ),
    .A3(\flop69.q ),
    .S1(_0140_),
    .X(_0202_));
 sg13g2_a21oi_1 _0675_ (.A1(\and122.a ),
    .A2(_0190_),
    .Y(_0203_),
    .B1(_0202_));
 sg13g2_nand2_1 _0676_ (.Y(_0204_),
    .A(\and122.a ),
    .B(_0202_));
 sg13g2_nor2_1 _0677_ (.A(_0007_),
    .B(_0145_),
    .Y(_0205_));
 sg13g2_a221oi_1 _0678_ (.B2(_0202_),
    .C1(net177),
    .B1(_0205_),
    .A1(_0145_),
    .Y(_0206_),
    .A2(_0204_));
 sg13g2_o21ai_1 _0679_ (.B1(_0154_),
    .Y(_0207_),
    .A1(_0203_),
    .A2(_0206_));
 sg13g2_nand2_1 _0680_ (.Y(_0208_),
    .A(_0113_),
    .B(_0158_));
 sg13g2_o21ai_1 _0681_ (.B1(net191),
    .Y(_0209_),
    .A1(net195),
    .A2(_0111_));
 sg13g2_a21o_1 _0682_ (.A2(_0008_),
    .A1(net194),
    .B1(_0209_),
    .X(_0210_));
 sg13g2_o21ai_1 _0683_ (.B1(_0208_),
    .Y(_0211_),
    .A1(net178),
    .A2(_0202_));
 sg13g2_a21oi_1 _0684_ (.A1(net180),
    .A2(_0211_),
    .Y(_0212_),
    .B1(_0163_));
 sg13g2_a22oi_1 _0685_ (.Y(_0213_),
    .B1(_0210_),
    .B2(_0212_),
    .A2(_0116_),
    .A1(net181));
 sg13g2_nand2_1 _0686_ (.Y(_0214_),
    .A(_0207_),
    .B(_0213_));
 sg13g2_a221oi_1 _0687_ (.B2(_0213_),
    .C1(_0200_),
    .B1(_0207_),
    .A1(_0157_),
    .Y(_0215_),
    .A2(_0185_));
 sg13g2_nor2_1 _0688_ (.A(_0178_),
    .B(_0215_),
    .Y(_0216_));
 sg13g2_mux4_1 _0689_ (.S0(net176),
    .A0(\flop46.q ),
    .A1(\flop54.q ),
    .A2(\flop62.q ),
    .A3(\flop70.q ),
    .S1(net175),
    .X(_0217_));
 sg13g2_a21oi_1 _0690_ (.A1(_0111_),
    .A2(_0190_),
    .Y(_0218_),
    .B1(_0217_));
 sg13g2_a21oi_1 _0691_ (.A1(_0111_),
    .A2(_0217_),
    .Y(_0219_),
    .B1(_0097_));
 sg13g2_and3_1 _0692_ (.X(_0220_),
    .A(_0111_),
    .B(_0144_),
    .C(_0217_));
 sg13g2_nor3_1 _0693_ (.A(net177),
    .B(_0219_),
    .C(_0220_),
    .Y(_0221_));
 sg13g2_o21ai_1 _0694_ (.B1(_0154_),
    .Y(_0222_),
    .A1(_0218_),
    .A2(_0221_));
 sg13g2_nand2_1 _0695_ (.Y(_0223_),
    .A(_0110_),
    .B(_0158_));
 sg13g2_o21ai_1 _0696_ (.B1(_0223_),
    .Y(_0224_),
    .A1(net178),
    .A2(_0217_));
 sg13g2_nand2_1 _0697_ (.Y(_0225_),
    .A(net179),
    .B(_0224_));
 sg13g2_o21ai_1 _0698_ (.B1(net191),
    .Y(_0226_),
    .A1(net195),
    .A2(_0108_));
 sg13g2_a21oi_1 _0699_ (.A1(net195),
    .A2(_0007_),
    .Y(_0227_),
    .B1(_0226_));
 sg13g2_nor2_1 _0700_ (.A(_0163_),
    .B(_0227_),
    .Y(_0228_));
 sg13g2_a22oi_1 _0701_ (.Y(_0229_),
    .B1(_0225_),
    .B2(_0228_),
    .A2(_0112_),
    .A1(net181));
 sg13g2_nand2_1 _0702_ (.Y(_0230_),
    .A(_0222_),
    .B(_0229_));
 sg13g2_a21oi_1 _0703_ (.A1(_0215_),
    .A2(_0230_),
    .Y(_0231_),
    .B1(_0178_));
 sg13g2_mux4_1 _0704_ (.S0(net176),
    .A0(\flop47.q ),
    .A1(\flop55.q ),
    .A2(\flop63.q ),
    .A3(\flop71.q ),
    .S1(net175),
    .X(_0232_));
 sg13g2_a21oi_1 _0705_ (.A1(_0108_),
    .A2(_0190_),
    .Y(_0233_),
    .B1(_0232_));
 sg13g2_and2_1 _0706_ (.A(_0108_),
    .B(_0232_),
    .X(_0234_));
 sg13g2_xnor2_1 _0707_ (.Y(_0235_),
    .A(_0000_),
    .B(_0234_));
 sg13g2_a21oi_1 _0708_ (.A1(_0136_),
    .A2(_0235_),
    .Y(_0236_),
    .B1(_0233_));
 sg13g2_nand2b_1 _0709_ (.Y(_0237_),
    .B(_0158_),
    .A_N(\and11.b ));
 sg13g2_nand2b_1 _0710_ (.Y(_0238_),
    .B(_0004_),
    .A_N(net192));
 sg13g2_a21oi_1 _0711_ (.A1(net192),
    .A2(_0006_),
    .Y(_0239_),
    .B1(net179));
 sg13g2_o21ai_1 _0712_ (.B1(_0237_),
    .Y(_0240_),
    .A1(net178),
    .A2(_0232_));
 sg13g2_a22oi_1 _0713_ (.Y(_0241_),
    .B1(_0240_),
    .B2(net179),
    .A2(_0239_),
    .A1(_0238_));
 sg13g2_a22oi_1 _0714_ (.Y(_0242_),
    .B1(_0162_),
    .B2(_0241_),
    .A2(_0109_),
    .A1(net181));
 sg13g2_o21ai_1 _0715_ (.B1(_0242_),
    .Y(_0243_),
    .A1(_0155_),
    .A2(_0236_));
 sg13g2_nor2_1 _0716_ (.A(_0178_),
    .B(_0243_),
    .Y(_0244_));
 sg13g2_nor2_1 _0717_ (.A(_0231_),
    .B(_0244_),
    .Y(_0245_));
 sg13g2_mux4_1 _0718_ (.S0(net176),
    .A0(\flop48.q ),
    .A1(\flop56.q ),
    .A2(\flop64.q ),
    .A3(\flop72.q ),
    .S1(net175),
    .X(_0246_));
 sg13g2_nand2b_1 _0719_ (.Y(_0247_),
    .B(_0158_),
    .A_N(\and125.a ));
 sg13g2_nand2b_1 _0720_ (.Y(_0248_),
    .B(_0003_),
    .A_N(net192));
 sg13g2_o21ai_1 _0721_ (.B1(_0247_),
    .Y(_0249_),
    .A1(net178),
    .A2(_0246_));
 sg13g2_a21oi_1 _0722_ (.A1(net192),
    .A2(_0005_),
    .Y(_0250_),
    .B1(net179));
 sg13g2_a221oi_1 _0723_ (.B2(_0248_),
    .C1(net181),
    .B1(_0250_),
    .A1(net179),
    .Y(_0251_),
    .A2(_0249_));
 sg13g2_nand2_1 _0724_ (.Y(_0252_),
    .A(_0107_),
    .B(_0246_));
 sg13g2_o21ai_1 _0725_ (.B1(_0136_),
    .Y(_0253_),
    .A1(_0000_),
    .A2(_0252_));
 sg13g2_a21oi_1 _0726_ (.A1(_0000_),
    .A2(_0252_),
    .Y(_0254_),
    .B1(_0253_));
 sg13g2_a21oi_1 _0727_ (.A1(_0107_),
    .A2(_0190_),
    .Y(_0255_),
    .B1(_0246_));
 sg13g2_or3_1 _0728_ (.A(_0162_),
    .B(_0254_),
    .C(_0255_),
    .X(_0256_));
 sg13g2_o21ai_1 _0729_ (.B1(_0256_),
    .Y(_0257_),
    .A1(_0154_),
    .A2(_0251_));
 sg13g2_o21ai_1 _0730_ (.B1(_0257_),
    .Y(_0258_),
    .A1(net188),
    .A2(net6));
 sg13g2_xor2_1 _0731_ (.B(_0258_),
    .A(_0245_),
    .X(_0259_));
 sg13g2_xor2_1 _0732_ (.B(_0243_),
    .A(_0231_),
    .X(_0260_));
 sg13g2_nor2_1 _0733_ (.A(_0005_),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_xor2_1 _0734_ (.B(_0230_),
    .A(_0216_),
    .X(_0262_));
 sg13g2_nor2_1 _0735_ (.A(_0006_),
    .B(_0262_),
    .Y(_0263_));
 sg13g2_o21ai_1 _0736_ (.B1(_0214_),
    .Y(_0264_),
    .A1(_0178_),
    .A2(_0201_));
 sg13g2_or3_1 _0737_ (.A(_0178_),
    .B(_0201_),
    .C(_0214_),
    .X(_0265_));
 sg13g2_nand2_1 _0738_ (.Y(_0266_),
    .A(_0264_),
    .B(_0265_));
 sg13g2_nand3b_1 _0739_ (.B(_0264_),
    .C(_0265_),
    .Y(_0267_),
    .A_N(_0007_));
 sg13g2_a21oi_1 _0740_ (.A1(_0264_),
    .A2(_0265_),
    .Y(_0268_),
    .B1(\and122.a ));
 sg13g2_nand3_1 _0741_ (.B(_0171_),
    .C(_0185_),
    .A(_0157_),
    .Y(_0269_));
 sg13g2_a22oi_1 _0742_ (.Y(_0270_),
    .B1(_0171_),
    .B2(net183),
    .A2(_0169_),
    .A1(_0117_));
 sg13g2_nand3_1 _0743_ (.B(_0269_),
    .C(_0270_),
    .A(_0008_),
    .Y(_0271_));
 sg13g2_a21oi_1 _0744_ (.A1(_0269_),
    .A2(_0270_),
    .Y(_0272_),
    .B1(_0114_));
 sg13g2_nand3b_1 _0745_ (.B(net182),
    .C(_0169_),
    .Y(_0273_),
    .A_N(net186));
 sg13g2_xnor2_1 _0746_ (.Y(_0274_),
    .A(_0200_),
    .B(_0273_));
 sg13g2_a21oi_2 _0747_ (.B1(_0272_),
    .Y(_0275_),
    .A2(_0274_),
    .A1(_0271_));
 sg13g2_a21oi_1 _0748_ (.A1(_0267_),
    .A2(_0275_),
    .Y(_0276_),
    .B1(_0268_));
 sg13g2_a221oi_1 _0749_ (.B2(_0275_),
    .C1(_0268_),
    .B1(_0267_),
    .A1(_0110_),
    .Y(_0277_),
    .A2(_0262_));
 sg13g2_nor2_1 _0750_ (.A(_0263_),
    .B(_0277_),
    .Y(_0278_));
 sg13g2_nand2b_1 _0751_ (.Y(_0279_),
    .B(_0260_),
    .A_N(\and11.b ));
 sg13g2_or3_1 _0752_ (.A(_0261_),
    .B(_0263_),
    .C(_0277_),
    .X(_0280_));
 sg13g2_and3_1 _0753_ (.X(_0281_),
    .A(\and125.a ),
    .B(_0279_),
    .C(_0280_));
 sg13g2_a21oi_1 _0754_ (.A1(_0279_),
    .A2(_0280_),
    .Y(_0282_),
    .B1(\and125.a ));
 sg13g2_nor3_1 _0755_ (.A(net187),
    .B(_0281_),
    .C(_0282_),
    .Y(_0283_));
 sg13g2_xnor2_1 _0756_ (.Y(_0284_),
    .A(_0259_),
    .B(_0283_));
 sg13g2_mux2_1 _0757_ (.A0(net147),
    .A1(_0284_),
    .S(net196),
    .X(_0285_));
 sg13g2_nor2_1 _0758_ (.A(net157),
    .B(net197),
    .Y(_0286_));
 sg13g2_and3_1 _0759_ (.X(_0287_),
    .A(_0114_),
    .B(_0269_),
    .C(_0270_));
 sg13g2_nor3_1 _0760_ (.A(net186),
    .B(_0272_),
    .C(_0287_),
    .Y(_0288_));
 sg13g2_xor2_1 _0761_ (.B(_0288_),
    .A(_0274_),
    .X(_0289_));
 sg13g2_a21oi_2 _0762_ (.B1(_0286_),
    .Y(_0290_),
    .A2(_0289_),
    .A1(net197));
 sg13g2_mux2_2 _0763_ (.A0(_0285_),
    .A1(_0290_),
    .S(_0177_),
    .X(_0291_));
 sg13g2_inv_1 _0764_ (.Y(_0292_),
    .A(_0291_));
 sg13g2_xor2_1 _0765_ (.B(_0278_),
    .A(\and11.b ),
    .X(_0293_));
 sg13g2_nor2_1 _0766_ (.A(net187),
    .B(_0293_),
    .Y(_0294_));
 sg13g2_xor2_1 _0767_ (.B(_0294_),
    .A(_0260_),
    .X(_0295_));
 sg13g2_mux2_1 _0768_ (.A0(net153),
    .A1(_0295_),
    .S(net196),
    .X(_0296_));
 sg13g2_mux2_2 _0769_ (.A0(_0296_),
    .A1(_0175_),
    .S(_0177_),
    .X(_0297_));
 sg13g2_inv_1 _0770_ (.Y(_0298_),
    .A(_0297_));
 sg13g2_mux4_1 _0771_ (.S0(net176),
    .A0(\flop49.q ),
    .A1(\flop57.q ),
    .A2(\flop65.q ),
    .A3(\flop73.q ),
    .S1(net175),
    .X(_0299_));
 sg13g2_nand2_1 _0772_ (.Y(_0300_),
    .A(_0106_),
    .B(_0299_));
 sg13g2_xnor2_1 _0773_ (.Y(_0301_),
    .A(_0000_),
    .B(_0300_));
 sg13g2_a21oi_1 _0774_ (.A1(_0106_),
    .A2(_0190_),
    .Y(_0302_),
    .B1(_0299_));
 sg13g2_nor2_1 _0775_ (.A(_0162_),
    .B(_0302_),
    .Y(_0303_));
 sg13g2_o21ai_1 _0776_ (.B1(_0303_),
    .Y(_0304_),
    .A1(net177),
    .A2(_0301_));
 sg13g2_nand2_1 _0777_ (.Y(_0305_),
    .A(net192),
    .B(_0105_));
 sg13g2_nor2_1 _0778_ (.A(net192),
    .B(_0002_),
    .Y(_0306_));
 sg13g2_a21oi_1 _0779_ (.A1(net192),
    .A2(_0107_),
    .Y(_0307_),
    .B1(_0306_));
 sg13g2_a21oi_1 _0780_ (.A1(net191),
    .A2(_0307_),
    .Y(_0308_),
    .B1(_0153_));
 sg13g2_nor2_1 _0781_ (.A(net178),
    .B(_0299_),
    .Y(_0309_));
 sg13g2_o21ai_1 _0782_ (.B1(net179),
    .Y(_0310_),
    .A1(\and128.b ),
    .A2(_0305_));
 sg13g2_o21ai_1 _0783_ (.B1(_0308_),
    .Y(_0311_),
    .A1(_0309_),
    .A2(_0310_));
 sg13g2_nand3_1 _0784_ (.B(_0304_),
    .C(_0311_),
    .A(net188),
    .Y(_0312_));
 sg13g2_o21ai_1 _0785_ (.B1(_0312_),
    .Y(_0313_),
    .A1(net188),
    .A2(net7));
 sg13g2_a21oi_1 _0786_ (.A1(_0245_),
    .A2(_0258_),
    .Y(_0314_),
    .B1(_0178_));
 sg13g2_xnor2_1 _0787_ (.Y(_0315_),
    .A(_0313_),
    .B(_0314_));
 sg13g2_nor2_1 _0788_ (.A(\and126.a ),
    .B(_0315_),
    .Y(_0316_));
 sg13g2_nand2_1 _0789_ (.Y(_0317_),
    .A(\and126.a ),
    .B(_0315_));
 sg13g2_nand2b_1 _0790_ (.Y(_0318_),
    .B(_0317_),
    .A_N(_0316_));
 sg13g2_nor2_1 _0791_ (.A(\and125.a ),
    .B(_0259_),
    .Y(_0319_));
 sg13g2_a22oi_1 _0792_ (.Y(_0320_),
    .B1(_0279_),
    .B2(_0280_),
    .A2(_0259_),
    .A1(_0107_));
 sg13g2_or2_1 _0793_ (.X(_0321_),
    .B(_0320_),
    .A(_0319_));
 sg13g2_xnor2_1 _0794_ (.Y(_0322_),
    .A(_0318_),
    .B(_0321_));
 sg13g2_mux2_2 _0795_ (.A0(_0322_),
    .A1(_0313_),
    .S(net187),
    .X(_0323_));
 sg13g2_nand2_1 _0796_ (.Y(_0324_),
    .A(net197),
    .B(_0323_));
 sg13g2_o21ai_1 _0797_ (.B1(_0324_),
    .Y(_0325_),
    .A1(net145),
    .A2(net197));
 sg13g2_nor2_1 _0798_ (.A(net158),
    .B(net12),
    .Y(_0326_));
 sg13g2_xnor2_1 _0799_ (.Y(_0327_),
    .A(_0113_),
    .B(_0275_));
 sg13g2_nor2_1 _0800_ (.A(net187),
    .B(_0327_),
    .Y(_0328_));
 sg13g2_xnor2_1 _0801_ (.Y(_0329_),
    .A(_0266_),
    .B(_0328_));
 sg13g2_inv_1 _0802_ (.Y(_0330_),
    .A(_0329_));
 sg13g2_a21oi_1 _0803_ (.A1(net12),
    .A2(_0329_),
    .Y(_0331_),
    .B1(_0326_));
 sg13g2_mux4_1 _0804_ (.S0(_0177_),
    .A0(_0105_),
    .A1(_0007_),
    .A2(_0323_),
    .A3(_0330_),
    .S1(net197),
    .X(_0332_));
 sg13g2_inv_1 _0805_ (.Y(_0333_),
    .A(net162));
 sg13g2_nand2_1 _0806_ (.Y(_0334_),
    .A(_0298_),
    .B(_0333_));
 sg13g2_o21ai_1 _0807_ (.B1(_0291_),
    .Y(_0335_),
    .A1(_0297_),
    .A2(net162));
 sg13g2_nor2_1 _0808_ (.A(net155),
    .B(net196),
    .Y(_0336_));
 sg13g2_xnor2_1 _0809_ (.Y(_0337_),
    .A(\and10.a ),
    .B(_0276_));
 sg13g2_nor2_1 _0810_ (.A(net187),
    .B(_0337_),
    .Y(_0338_));
 sg13g2_xnor2_1 _0811_ (.Y(_0339_),
    .A(_0262_),
    .B(_0338_));
 sg13g2_inv_1 _0812_ (.Y(_0340_),
    .A(_0339_));
 sg13g2_a21oi_1 _0813_ (.A1(net196),
    .A2(_0339_),
    .Y(_0341_),
    .B1(_0336_));
 sg13g2_mux4_1 _0814_ (.S0(net176),
    .A0(_0102_),
    .A1(_0103_),
    .A2(_0100_),
    .A3(_0101_),
    .S1(net175),
    .X(_0342_));
 sg13g2_nor2_1 _0815_ (.A(_0002_),
    .B(_0342_),
    .Y(_0343_));
 sg13g2_xnor2_1 _0816_ (.Y(_0344_),
    .A(_0097_),
    .B(_0343_));
 sg13g2_nand2b_1 _0817_ (.Y(_0345_),
    .B(_0190_),
    .A_N(_0002_));
 sg13g2_a21oi_1 _0818_ (.A1(_0342_),
    .A2(_0345_),
    .Y(_0346_),
    .B1(_0162_));
 sg13g2_o21ai_1 _0819_ (.B1(_0346_),
    .Y(_0347_),
    .A1(net177),
    .A2(_0344_));
 sg13g2_nand2_1 _0820_ (.Y(_0348_),
    .A(\and128.b ),
    .B(_0342_));
 sg13g2_nand2b_1 _0821_ (.Y(_0349_),
    .B(net192),
    .A_N(\and127.a ));
 sg13g2_o21ai_1 _0822_ (.B1(_0348_),
    .Y(_0350_),
    .A1(\and128.b ),
    .A2(_0349_));
 sg13g2_nand3_1 _0823_ (.B(\and115.b ),
    .C(net190),
    .A(\and128.b ),
    .Y(_0351_));
 sg13g2_nand2_1 _0824_ (.Y(_0352_),
    .A(_0164_),
    .B(_0351_));
 sg13g2_o21ai_1 _0825_ (.B1(_0305_),
    .Y(_0353_),
    .A1(net194),
    .A2(_0352_));
 sg13g2_a21oi_1 _0826_ (.A1(net191),
    .A2(_0353_),
    .Y(_0354_),
    .B1(_0153_));
 sg13g2_o21ai_1 _0827_ (.B1(_0354_),
    .Y(_0355_),
    .A1(net191),
    .A2(_0350_));
 sg13g2_nand3_1 _0828_ (.B(_0347_),
    .C(_0355_),
    .A(net188),
    .Y(_0356_));
 sg13g2_o21ai_1 _0829_ (.B1(_0356_),
    .Y(_0357_),
    .A1(net8),
    .A2(net188));
 sg13g2_nor2_1 _0830_ (.A(_0178_),
    .B(_0313_),
    .Y(_0358_));
 sg13g2_nor2_1 _0831_ (.A(_0314_),
    .B(_0358_),
    .Y(_0359_));
 sg13g2_xnor2_1 _0832_ (.Y(_0360_),
    .A(_0357_),
    .B(_0359_));
 sg13g2_inv_1 _0833_ (.Y(_0361_),
    .A(_0360_));
 sg13g2_nand2_1 _0834_ (.Y(_0362_),
    .A(net187),
    .B(_0361_));
 sg13g2_xnor2_1 _0835_ (.Y(_0363_),
    .A(net190),
    .B(_0360_));
 sg13g2_a21oi_1 _0836_ (.A1(_0317_),
    .A2(_0321_),
    .Y(_0364_),
    .B1(_0316_));
 sg13g2_xnor2_1 _0837_ (.Y(_0365_),
    .A(_0363_),
    .B(_0364_));
 sg13g2_mux2_1 _0838_ (.A0(_0365_),
    .A1(_0360_),
    .S(net187),
    .X(_0366_));
 sg13g2_o21ai_1 _0839_ (.B1(_0362_),
    .Y(_0367_),
    .A1(net187),
    .A2(_0365_));
 sg13g2_mux4_1 _0840_ (.S0(_0177_),
    .A0(_0002_),
    .A1(_0006_),
    .A2(_0366_),
    .A3(_0340_),
    .S1(net196),
    .X(_0368_));
 sg13g2_nand2_1 _0841_ (.Y(_0369_),
    .A(_0291_),
    .B(net162));
 sg13g2_nand2_1 _0842_ (.Y(_0370_),
    .A(_0298_),
    .B(_0369_));
 sg13g2_nor2_1 _0843_ (.A(net190),
    .B(net196),
    .Y(_0371_));
 sg13g2_a21oi_1 _0844_ (.A1(net196),
    .A2(_0366_),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_mux4_1 _0845_ (.S0(_0177_),
    .A0(net190),
    .A1(_0111_),
    .A2(_0367_),
    .A3(_0339_),
    .S1(net196),
    .X(_0373_));
 sg13g2_nand2_1 _0846_ (.Y(_0374_),
    .A(_0297_),
    .B(net162));
 sg13g2_inv_1 _0847_ (.Y(_0375_),
    .A(_0374_));
 sg13g2_o21ai_1 _0848_ (.B1(_0370_),
    .Y(_0376_),
    .A1(_0373_),
    .A2(_0375_));
 sg13g2_a221oi_1 _0849_ (.B2(_0368_),
    .C1(net198),
    .B1(_0335_),
    .A1(_0292_),
    .Y(_0377_),
    .A2(_0333_));
 sg13g2_a22oi_1 _0850_ (.Y(\flop12.d ),
    .B1(_0376_),
    .B2(_0377_),
    .A2(_0175_),
    .A1(net198));
 sg13g2_o21ai_1 _0851_ (.B1(_0298_),
    .Y(_0378_),
    .A1(_0291_),
    .A2(_0368_));
 sg13g2_nor2_1 _0852_ (.A(_0292_),
    .B(_0373_),
    .Y(_0379_));
 sg13g2_or2_1 _0853_ (.X(_0380_),
    .B(_0379_),
    .A(_0378_));
 sg13g2_or2_1 _0854_ (.X(_0381_),
    .B(_0368_),
    .A(net162));
 sg13g2_nand2_1 _0855_ (.Y(_0382_),
    .A(_0335_),
    .B(_0374_));
 sg13g2_a21oi_1 _0856_ (.A1(_0381_),
    .A2(_0382_),
    .Y(_0383_),
    .B1(net198));
 sg13g2_a22oi_1 _0857_ (.Y(\flop13.d ),
    .B1(_0380_),
    .B2(_0383_),
    .A2(_0290_),
    .A1(net199));
 sg13g2_nand2_1 _0858_ (.Y(_0384_),
    .A(_0292_),
    .B(net162));
 sg13g2_a221oi_1 _0859_ (.B2(_0368_),
    .C1(net198),
    .B1(_0384_),
    .A1(net162),
    .Y(_0385_),
    .A2(_0373_));
 sg13g2_a22oi_1 _0860_ (.Y(\flop14.d ),
    .B1(_0378_),
    .B2(_0385_),
    .A2(_0331_),
    .A1(net198));
 sg13g2_nor3_1 _0861_ (.A(_0291_),
    .B(_0297_),
    .C(_0332_),
    .Y(_0386_));
 sg13g2_or2_1 _0862_ (.X(_0387_),
    .B(_0386_),
    .A(_0382_));
 sg13g2_a221oi_1 _0863_ (.B2(_0368_),
    .C1(net198),
    .B1(_0375_),
    .A1(_0291_),
    .Y(_0388_),
    .A2(_0373_));
 sg13g2_a22oi_1 _0864_ (.Y(\flop15.d ),
    .B1(_0387_),
    .B2(_0388_),
    .A2(_0341_),
    .A1(net198));
 sg13g2_nor2_1 _0865_ (.A(_0292_),
    .B(net162),
    .Y(_0389_));
 sg13g2_nand2_1 _0866_ (.Y(_0390_),
    .A(_0291_),
    .B(_0333_));
 sg13g2_a221oi_1 _0867_ (.B2(_0297_),
    .C1(net198),
    .B1(_0390_),
    .A1(_0369_),
    .Y(_0391_),
    .A2(_0373_));
 sg13g2_a21oi_1 _0868_ (.A1(net199),
    .A2(_0296_),
    .Y(\flop16.d ),
    .B1(_0391_));
 sg13g2_a21oi_1 _0869_ (.A1(_0368_),
    .A2(_0389_),
    .Y(_0392_),
    .B1(net199));
 sg13g2_a22oi_1 _0870_ (.Y(_0393_),
    .B1(_0390_),
    .B2(_0373_),
    .A2(_0384_),
    .A1(_0297_));
 sg13g2_a22oi_1 _0871_ (.Y(\flop17.d ),
    .B1(_0392_),
    .B2(_0393_),
    .A2(_0285_),
    .A1(net199));
 sg13g2_nand2_1 _0872_ (.Y(_0394_),
    .A(_0297_),
    .B(_0333_));
 sg13g2_a22oi_1 _0873_ (.Y(_0395_),
    .B1(_0373_),
    .B2(_0394_),
    .A2(_0334_),
    .A1(_0292_));
 sg13g2_a22oi_1 _0874_ (.Y(\flop18.d ),
    .B1(_0392_),
    .B2(_0395_),
    .A2(_0325_),
    .A1(net199));
 sg13g2_mux2_1 _0875_ (.A0(_0177_),
    .A1(_0372_),
    .S(net199),
    .X(\flop83.d ));
 sg13g2_nand3b_1 _0876_ (.B(\and83.a ),
    .C(\and83.b ),
    .Y(_0396_),
    .A_N(\flop29.notq ));
 sg13g2_nor2_1 _0877_ (.A(\flop30.notq ),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_nor4_2 _0878_ (.A(\flop30.notq ),
    .B(\flop31.notq ),
    .C(\flop32.notq ),
    .Y(_0398_),
    .D(_0396_));
 sg13g2_nor2b_1 _0879_ (.A(\flop33.notq ),
    .B_N(_0398_),
    .Y(_0399_));
 sg13g2_nor2b_1 _0880_ (.A(\flop34.notq ),
    .B_N(_0399_),
    .Y(_0400_));
 sg13g2_nor2b_1 _0881_ (.A(\flop35.notq ),
    .B_N(_0400_),
    .Y(_0401_));
 sg13g2_nand2b_1 _0882_ (.Y(_0402_),
    .B(_0401_),
    .A_N(net44));
 sg13g2_nor2_1 _0883_ (.A(\flop37.notq ),
    .B(_0402_),
    .Y(_0403_));
 sg13g2_nor3_2 _0884_ (.A(\flop37.notq ),
    .B(\flop38.notq ),
    .C(_0402_),
    .Y(_0404_));
 sg13g2_nor2_1 _0885_ (.A(net54),
    .B(_0403_),
    .Y(_0405_));
 sg13g2_nor2_1 _0886_ (.A(_0404_),
    .B(net55),
    .Y(_0021_));
 sg13g2_nor3_1 _0887_ (.A(net180),
    .B(\and128.b ),
    .C(_0161_),
    .Y(_0406_));
 sg13g2_nor2b_2 _0888_ (.A(\flop26.q ),
    .B_N(net30),
    .Y(_0407_));
 sg13g2_nand2_1 _0889_ (.Y(_0408_),
    .A(_0094_),
    .B(_0407_));
 sg13g2_a21oi_2 _0890_ (.B1(_0408_),
    .Y(_0409_),
    .A2(_0406_),
    .A1(_0099_));
 sg13g2_nand2_1 _0891_ (.Y(_0410_),
    .A(_0339_),
    .B(net172));
 sg13g2_o21ai_1 _0892_ (.B1(_0410_),
    .Y(_0022_),
    .A1(_0110_),
    .A2(net172));
 sg13g2_nor2b_1 _0893_ (.A(\flop39.notq ),
    .B_N(_0404_),
    .Y(_0411_));
 sg13g2_nand2b_1 _0894_ (.Y(_0412_),
    .B(_0404_),
    .A_N(\flop39.notq ));
 sg13g2_nor2_1 _0895_ (.A(\flop40.notq ),
    .B(_0412_),
    .Y(_0413_));
 sg13g2_a21oi_1 _0896_ (.A1(_0093_),
    .A2(_0412_),
    .Y(_0023_),
    .B1(_0413_));
 sg13g2_a21oi_1 _0897_ (.A1(net41),
    .A2(_0411_),
    .Y(_0414_),
    .B1(\and106.a ));
 sg13g2_nor4_1 _0898_ (.A(\flop40.notq ),
    .B(\flop42.notq ),
    .C(net41),
    .D(_0412_),
    .Y(_0415_));
 sg13g2_nor2_1 _0899_ (.A(net42),
    .B(_0415_),
    .Y(_0024_));
 sg13g2_mux2_1 _0900_ (.A0(\and110.b ),
    .A1(net52),
    .S(_0413_),
    .X(_0025_));
 sg13g2_nand2_1 _0901_ (.Y(_0416_),
    .A(net185),
    .B(_0407_));
 sg13g2_nor3_1 _0902_ (.A(\and115.b ),
    .B(net193),
    .C(_0416_),
    .Y(_0417_));
 sg13g2_nor3_2 _0903_ (.A(_0094_),
    .B(net189),
    .C(_0151_),
    .Y(_0418_));
 sg13g2_nand2b_1 _0904_ (.Y(_0419_),
    .B(net174),
    .A_N(net183));
 sg13g2_o21ai_1 _0905_ (.B1(_0419_),
    .Y(_0420_),
    .A1(_0174_),
    .A2(net174));
 sg13g2_nor2_1 _0906_ (.A(net111),
    .B(net170),
    .Y(_0421_));
 sg13g2_a21oi_1 _0907_ (.A1(net170),
    .A2(_0420_),
    .Y(_0026_),
    .B1(_0421_));
 sg13g2_nor2_1 _0908_ (.A(net117),
    .B(net170),
    .Y(_0422_));
 sg13g2_nand2_1 _0909_ (.Y(_0423_),
    .A(_0114_),
    .B(net174));
 sg13g2_o21ai_1 _0910_ (.B1(_0423_),
    .Y(_0424_),
    .A1(_0289_),
    .A2(net174));
 sg13g2_a21oi_1 _0911_ (.A1(net170),
    .A2(_0424_),
    .Y(_0027_),
    .B1(_0422_));
 sg13g2_nand2_1 _0912_ (.Y(_0425_),
    .A(_0113_),
    .B(net174));
 sg13g2_o21ai_1 _0913_ (.B1(_0425_),
    .Y(_0426_),
    .A1(_0329_),
    .A2(_0418_));
 sg13g2_nor2_1 _0914_ (.A(net91),
    .B(net170),
    .Y(_0427_));
 sg13g2_a21oi_1 _0915_ (.A1(_0417_),
    .A2(_0426_),
    .Y(_0028_),
    .B1(_0427_));
 sg13g2_nand2_1 _0916_ (.Y(_0428_),
    .A(_0110_),
    .B(net174));
 sg13g2_o21ai_1 _0917_ (.B1(_0428_),
    .Y(_0429_),
    .A1(_0339_),
    .A2(net174));
 sg13g2_nor2_1 _0918_ (.A(net123),
    .B(net169),
    .Y(_0430_));
 sg13g2_a21oi_1 _0919_ (.A1(net170),
    .A2(_0429_),
    .Y(_0029_),
    .B1(_0430_));
 sg13g2_nor2_1 _0920_ (.A(net103),
    .B(net170),
    .Y(_0431_));
 sg13g2_nor2_1 _0921_ (.A(_0295_),
    .B(net173),
    .Y(_0432_));
 sg13g2_a21oi_2 _0922_ (.B1(_0432_),
    .Y(_0433_),
    .A2(net173),
    .A1(\and11.b ));
 sg13g2_a21oi_1 _0923_ (.A1(net169),
    .A2(_0433_),
    .Y(_0030_),
    .B1(_0431_));
 sg13g2_nor2_1 _0924_ (.A(_0284_),
    .B(net173),
    .Y(_0434_));
 sg13g2_a21oi_2 _0925_ (.B1(_0434_),
    .Y(_0435_),
    .A2(net173),
    .A1(\and125.a ));
 sg13g2_nor2_1 _0926_ (.A(net131),
    .B(net169),
    .Y(_0436_));
 sg13g2_a21oi_1 _0927_ (.A1(net169),
    .A2(_0435_),
    .Y(_0031_),
    .B1(_0436_));
 sg13g2_nor2_1 _0928_ (.A(net134),
    .B(net172),
    .Y(_0437_));
 sg13g2_a21oi_1 _0929_ (.A1(_0295_),
    .A2(net171),
    .Y(_0032_),
    .B1(_0437_));
 sg13g2_nor2_1 _0930_ (.A(net101),
    .B(net169),
    .Y(_0438_));
 sg13g2_nor2_1 _0931_ (.A(_0366_),
    .B(net173),
    .Y(_0439_));
 sg13g2_a21oi_2 _0932_ (.B1(_0439_),
    .Y(_0440_),
    .A2(net173),
    .A1(net190));
 sg13g2_a21oi_1 _0933_ (.A1(net169),
    .A2(_0440_),
    .Y(_0033_),
    .B1(_0438_));
 sg13g2_nand3_1 _0934_ (.B(net193),
    .C(_0407_),
    .A(net185),
    .Y(_0441_));
 sg13g2_nor2_1 _0935_ (.A(\and115.b ),
    .B(_0441_),
    .Y(_0442_));
 sg13g2_nor2_1 _0936_ (.A(net85),
    .B(net168),
    .Y(_0443_));
 sg13g2_a21oi_1 _0937_ (.A1(_0420_),
    .A2(net168),
    .Y(_0034_),
    .B1(_0443_));
 sg13g2_nor2_1 _0938_ (.A(net82),
    .B(net168),
    .Y(_0444_));
 sg13g2_a21oi_1 _0939_ (.A1(_0424_),
    .A2(net168),
    .Y(_0035_),
    .B1(_0444_));
 sg13g2_nor2_1 _0940_ (.A(net96),
    .B(net168),
    .Y(_0445_));
 sg13g2_a21oi_1 _0941_ (.A1(_0426_),
    .A2(_0442_),
    .Y(_0036_),
    .B1(_0445_));
 sg13g2_nor2_1 _0942_ (.A(net95),
    .B(net167),
    .Y(_0446_));
 sg13g2_a21oi_1 _0943_ (.A1(_0429_),
    .A2(net168),
    .Y(_0037_),
    .B1(_0446_));
 sg13g2_nor2_1 _0944_ (.A(net89),
    .B(net168),
    .Y(_0447_));
 sg13g2_a21oi_1 _0945_ (.A1(_0433_),
    .A2(net167),
    .Y(_0038_),
    .B1(_0447_));
 sg13g2_nor2_1 _0946_ (.A(net119),
    .B(net167),
    .Y(_0448_));
 sg13g2_a21oi_1 _0947_ (.A1(_0435_),
    .A2(net167),
    .Y(_0039_),
    .B1(_0448_));
 sg13g2_nor2_1 _0948_ (.A(_0323_),
    .B(net173),
    .Y(_0449_));
 sg13g2_a21oi_2 _0949_ (.B1(_0449_),
    .Y(_0450_),
    .A2(net173),
    .A1(\and126.a ));
 sg13g2_nor2_1 _0950_ (.A(net124),
    .B(net167),
    .Y(_0451_));
 sg13g2_a21oi_1 _0951_ (.A1(net167),
    .A2(_0450_),
    .Y(_0040_),
    .B1(_0451_));
 sg13g2_nor2_1 _0952_ (.A(net76),
    .B(net167),
    .Y(_0452_));
 sg13g2_a21oi_1 _0953_ (.A1(_0440_),
    .A2(net167),
    .Y(_0041_),
    .B1(_0452_));
 sg13g2_nor2_1 _0954_ (.A(net143),
    .B(net171),
    .Y(_0453_));
 sg13g2_a21oi_1 _0955_ (.A1(_0284_),
    .A2(net171),
    .Y(_0042_),
    .B1(_0453_));
 sg13g2_nor3_1 _0956_ (.A(_0099_),
    .B(net193),
    .C(_0416_),
    .Y(_0454_));
 sg13g2_nor2_1 _0957_ (.A(net99),
    .B(net166),
    .Y(_0455_));
 sg13g2_a21oi_1 _0958_ (.A1(_0424_),
    .A2(net166),
    .Y(_0043_),
    .B1(_0455_));
 sg13g2_nor2_1 _0959_ (.A(net129),
    .B(net166),
    .Y(_0456_));
 sg13g2_a21oi_1 _0960_ (.A1(_0426_),
    .A2(_0454_),
    .Y(_0044_),
    .B1(_0456_));
 sg13g2_nor2_1 _0961_ (.A(net98),
    .B(net165),
    .Y(_0457_));
 sg13g2_a21oi_1 _0962_ (.A1(_0429_),
    .A2(net166),
    .Y(_0045_),
    .B1(_0457_));
 sg13g2_nor2_1 _0963_ (.A(net109),
    .B(net166),
    .Y(_0458_));
 sg13g2_a21oi_1 _0964_ (.A1(_0433_),
    .A2(net165),
    .Y(_0046_),
    .B1(_0458_));
 sg13g2_nor2_1 _0965_ (.A(net107),
    .B(net165),
    .Y(_0459_));
 sg13g2_a21oi_1 _0966_ (.A1(_0435_),
    .A2(net165),
    .Y(_0047_),
    .B1(_0459_));
 sg13g2_nor2_1 _0967_ (.A(net105),
    .B(net165),
    .Y(_0460_));
 sg13g2_a21oi_1 _0968_ (.A1(_0450_),
    .A2(net165),
    .Y(_0048_),
    .B1(_0460_));
 sg13g2_nor2_1 _0969_ (.A(net84),
    .B(net165),
    .Y(_0461_));
 sg13g2_a21oi_1 _0970_ (.A1(_0440_),
    .A2(net165),
    .Y(_0049_),
    .B1(_0461_));
 sg13g2_nor2_1 _0971_ (.A(_0099_),
    .B(_0441_),
    .Y(_0462_));
 sg13g2_nor2_1 _0972_ (.A(net102),
    .B(net164),
    .Y(_0463_));
 sg13g2_a21oi_1 _0973_ (.A1(_0420_),
    .A2(net164),
    .Y(_0050_),
    .B1(_0463_));
 sg13g2_nor2_1 _0974_ (.A(net86),
    .B(_0462_),
    .Y(_0464_));
 sg13g2_a21oi_1 _0975_ (.A1(_0424_),
    .A2(net164),
    .Y(_0051_),
    .B1(net87));
 sg13g2_nor2_1 _0976_ (.A(net145),
    .B(net171),
    .Y(_0465_));
 sg13g2_a21oi_1 _0977_ (.A1(_0323_),
    .A2(net171),
    .Y(_0052_),
    .B1(_0465_));
 sg13g2_nor2_1 _0978_ (.A(net126),
    .B(net164),
    .Y(_0466_));
 sg13g2_a21oi_1 _0979_ (.A1(_0429_),
    .A2(net164),
    .Y(_0053_),
    .B1(_0466_));
 sg13g2_nor2_1 _0980_ (.A(net121),
    .B(net163),
    .Y(_0467_));
 sg13g2_a21oi_1 _0981_ (.A1(_0433_),
    .A2(net163),
    .Y(_0054_),
    .B1(_0467_));
 sg13g2_nor2_1 _0982_ (.A(net115),
    .B(net163),
    .Y(_0468_));
 sg13g2_a21oi_1 _0983_ (.A1(_0435_),
    .A2(net163),
    .Y(_0055_),
    .B1(_0468_));
 sg13g2_nor2_1 _0984_ (.A(net127),
    .B(net163),
    .Y(_0469_));
 sg13g2_a21oi_1 _0985_ (.A1(_0450_),
    .A2(net163),
    .Y(_0056_),
    .B1(_0469_));
 sg13g2_nor2_1 _0986_ (.A(net77),
    .B(net163),
    .Y(_0470_));
 sg13g2_a21oi_1 _0987_ (.A1(_0440_),
    .A2(net163),
    .Y(_0057_),
    .B1(_0470_));
 sg13g2_nor2_1 _0988_ (.A(net193),
    .B(net201),
    .Y(_0471_));
 sg13g2_a21oi_1 _0989_ (.A1(_0122_),
    .A2(net201),
    .Y(_0058_),
    .B1(_0471_));
 sg13g2_nand2_1 _0990_ (.Y(_0472_),
    .A(net2),
    .B(net200));
 sg13g2_o21ai_1 _0991_ (.B1(_0472_),
    .Y(_0059_),
    .A1(_0099_),
    .A2(net201));
 sg13g2_nand2_1 _0992_ (.Y(_0473_),
    .A(net3),
    .B(net201));
 sg13g2_o21ai_1 _0993_ (.B1(_0473_),
    .Y(_0060_),
    .A1(net178),
    .A2(net200));
 sg13g2_nand2_1 _0994_ (.Y(_0474_),
    .A(net4),
    .B(net201));
 sg13g2_o21ai_1 _0995_ (.B1(_0474_),
    .Y(_0061_),
    .A1(net179),
    .A2(net201));
 sg13g2_nor2_1 _0996_ (.A(net190),
    .B(net171),
    .Y(_0475_));
 sg13g2_a21oi_1 _0997_ (.A1(_0366_),
    .A2(net171),
    .Y(_0062_),
    .B1(_0475_));
 sg13g2_nand2_1 _0998_ (.Y(_0476_),
    .A(net6),
    .B(net200));
 sg13g2_o21ai_1 _0999_ (.B1(_0476_),
    .Y(_0063_),
    .A1(net181),
    .A2(net200));
 sg13g2_mux2_1 _1000_ (.A0(net186),
    .A1(net7),
    .S(net200),
    .X(_0064_));
 sg13g2_nand2_1 _1001_ (.Y(_0477_),
    .A(net8),
    .B(net200));
 sg13g2_o21ai_1 _1002_ (.B1(_0477_),
    .Y(_0065_),
    .A1(_0094_),
    .A2(net200));
 sg13g2_nand3b_1 _1003_ (.B(_0170_),
    .C(net178),
    .Y(_0478_),
    .A_N(_0161_));
 sg13g2_inv_1 _1004_ (.Y(_0479_),
    .A(_0478_));
 sg13g2_nand3b_1 _1005_ (.B(_0170_),
    .C(\and115.b ),
    .Y(_0480_),
    .A_N(net193));
 sg13g2_o21ai_1 _1006_ (.B1(net186),
    .Y(_0481_),
    .A1(_0161_),
    .A2(_0480_));
 sg13g2_o21ai_1 _1007_ (.B1(_0407_),
    .Y(_0482_),
    .A1(_0479_),
    .A2(_0481_));
 sg13g2_o21ai_1 _1008_ (.B1(_0364_),
    .Y(_0483_),
    .A1(net190),
    .A2(_0361_));
 sg13g2_o21ai_1 _1009_ (.B1(_0483_),
    .Y(_0484_),
    .A1(_0002_),
    .A2(_0360_));
 sg13g2_o21ai_1 _1010_ (.B1(_0478_),
    .Y(_0485_),
    .A1(_0014_),
    .A2(_0484_));
 sg13g2_a21o_1 _1011_ (.A2(_0484_),
    .A1(_0014_),
    .B1(_0485_),
    .X(_0486_));
 sg13g2_a21oi_1 _1012_ (.A1(net194),
    .A2(_0104_),
    .Y(_0487_),
    .B1(_0478_));
 sg13g2_nor2_1 _1013_ (.A(\and115.b ),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_mux2_1 _1014_ (.A0(net183),
    .A1(net190),
    .S(net193),
    .X(_0489_));
 sg13g2_a221oi_1 _1015_ (.B2(\and115.b ),
    .C1(_0482_),
    .B1(_0489_),
    .A1(_0486_),
    .Y(_0490_),
    .A2(_0488_));
 sg13g2_a21oi_1 _1016_ (.A1(_0104_),
    .A2(_0482_),
    .Y(_0066_),
    .B1(_0490_));
 sg13g2_nor2b_1 _1017_ (.A(_0174_),
    .B_N(_0409_),
    .Y(_0491_));
 sg13g2_inv_1 _1018_ (.Y(_0492_),
    .A(_0491_));
 sg13g2_nor2_1 _1019_ (.A(net183),
    .B(_0409_),
    .Y(_0493_));
 sg13g2_nor2_1 _1020_ (.A(_0491_),
    .B(net149),
    .Y(_0067_));
 sg13g2_a21o_1 _1021_ (.A2(\and83.a ),
    .A1(\and83.b ),
    .B1(net137),
    .X(_0494_));
 sg13g2_and2_1 _1022_ (.A(_0396_),
    .B(net138),
    .X(_0068_));
 sg13g2_nor2_1 _1023_ (.A(net57),
    .B(_0404_),
    .Y(_0495_));
 sg13g2_nor2_1 _1024_ (.A(_0411_),
    .B(net58),
    .Y(_0069_));
 sg13g2_nor2_1 _1025_ (.A(net113),
    .B(net169),
    .Y(_0496_));
 sg13g2_a21oi_1 _1026_ (.A1(net169),
    .A2(_0450_),
    .Y(_0070_),
    .B1(_0496_));
 sg13g2_nor2_1 _1027_ (.A(net112),
    .B(net166),
    .Y(_0497_));
 sg13g2_a21oi_1 _1028_ (.A1(_0420_),
    .A2(net166),
    .Y(_0071_),
    .B1(_0497_));
 sg13g2_nor2_1 _1029_ (.A(net78),
    .B(net164),
    .Y(_0498_));
 sg13g2_a21oi_1 _1030_ (.A1(_0426_),
    .A2(net164),
    .Y(_0072_),
    .B1(_0498_));
 sg13g2_mux2_1 _1031_ (.A0(net182),
    .A1(net5),
    .S(net200),
    .X(_0073_));
 sg13g2_nand2b_1 _1032_ (.Y(_0499_),
    .B(net66),
    .A_N(net171));
 sg13g2_nor4_1 _1033_ (.A(_0289_),
    .B(_0329_),
    .C(_0339_),
    .D(_0492_),
    .Y(_0500_));
 sg13g2_nand4_1 _1034_ (.B(_0295_),
    .C(_0323_),
    .A(_0284_),
    .Y(_0501_),
    .D(_0500_));
 sg13g2_o21ai_1 _1035_ (.B1(_0499_),
    .Y(_0074_),
    .A1(_0367_),
    .A2(_0501_));
 sg13g2_a21oi_2 _1036_ (.B1(net211),
    .Y(_0502_),
    .A2(net161),
    .A1(_0126_));
 sg13g2_o21ai_1 _1037_ (.B1(_0502_),
    .Y(_0015_),
    .A1(_0126_),
    .A2(net159));
 sg13g2_nand2_1 _1038_ (.Y(_0503_),
    .A(_0289_),
    .B(net172));
 sg13g2_o21ai_1 _1039_ (.B1(_0503_),
    .Y(_0075_),
    .A1(_0114_),
    .A2(net172));
 sg13g2_nor2_1 _1040_ (.A(net30),
    .B(net94),
    .Y(_0504_));
 sg13g2_a21oi_1 _1041_ (.A1(_0126_),
    .A2(net94),
    .Y(_0081_),
    .B1(_0504_));
 sg13g2_mux2_1 _1042_ (.A0(\and83.a ),
    .A1(net32),
    .S(\and83.b ),
    .X(_0082_));
 sg13g2_nand2_1 _1043_ (.Y(_0505_),
    .A(_0329_),
    .B(net172));
 sg13g2_o21ai_1 _1044_ (.B1(_0505_),
    .Y(_0083_),
    .A1(_0113_),
    .A2(net172));
 sg13g2_a21oi_1 _1045_ (.A1(_0123_),
    .A2(_0396_),
    .Y(_0084_),
    .B1(_0397_));
 sg13g2_nor2_1 _1046_ (.A(net73),
    .B(_0397_),
    .Y(_0506_));
 sg13g2_a21oi_1 _1047_ (.A1(_0125_),
    .A2(_0397_),
    .Y(_0085_),
    .B1(net74));
 sg13g2_a21oi_1 _1048_ (.A1(_0125_),
    .A2(_0397_),
    .Y(_0507_),
    .B1(net36));
 sg13g2_nor2_1 _1049_ (.A(_0398_),
    .B(net37),
    .Y(_0086_));
 sg13g2_nor2_1 _1050_ (.A(net60),
    .B(_0398_),
    .Y(_0508_));
 sg13g2_nor2_1 _1051_ (.A(_0399_),
    .B(net61),
    .Y(_0087_));
 sg13g2_nor2_1 _1052_ (.A(net63),
    .B(_0399_),
    .Y(_0509_));
 sg13g2_nor2_1 _1053_ (.A(_0400_),
    .B(net64),
    .Y(_0088_));
 sg13g2_nor2_1 _1054_ (.A(net79),
    .B(_0400_),
    .Y(_0510_));
 sg13g2_nor2_1 _1055_ (.A(_0401_),
    .B(net80),
    .Y(_0089_));
 sg13g2_mux2_1 _1056_ (.A0(\and94.a ),
    .A1(net44),
    .S(_0401_),
    .X(_0090_));
 sg13g2_a21oi_1 _1057_ (.A1(_0124_),
    .A2(_0402_),
    .Y(_0091_),
    .B1(_0403_));
 sg13g2_o21ai_1 _1058_ (.B1(_0502_),
    .Y(_0016_),
    .A1(_0126_),
    .A2(net159));
 sg13g2_o21ai_1 _1059_ (.B1(_0502_),
    .Y(_0017_),
    .A1(_0126_),
    .A2(net159));
 sg13g2_o21ai_1 _1060_ (.B1(_0502_),
    .Y(_0018_),
    .A1(_0126_),
    .A2(net159));
 sg13g2_o21ai_1 _1061_ (.B1(_0502_),
    .Y(_0019_),
    .A1(_0126_),
    .A2(net159));
 sg13g2_o21ai_1 _1062_ (.B1(_0502_),
    .Y(_0020_),
    .A1(_0126_),
    .A2(net159));
 sg13g2_dfrbp_1 _1063_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net208),
    .D(net56),
    .Q_N(\flop38.notq ),
    .Q(\and102.a ));
 sg13g2_dfrbp_1 _1064_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net205),
    .D(_0022_),
    .Q_N(_0006_),
    .Q(\and10.a ));
 sg13g2_dfrbp_1 _1065_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net208),
    .D(net51),
    .Q_N(\flop40.notq ),
    .Q(\and107.b ));
 sg13g2_dfrbp_1 _1066_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net208),
    .D(net43),
    .Q_N(\and108.b ),
    .Q(\and106.a ));
 sg13g2_dfrbp_1 _1067_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net208),
    .D(net53),
    .Q_N(\flop42.notq ),
    .Q(\and110.b ));
 sg13g2_dfrbp_1 _1068_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net212),
    .D(_0026_),
    .Q_N(_0013_),
    .Q(\flop43.q ));
 sg13g2_dfrbp_1 _1069_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net210),
    .D(net118),
    .Q_N(_0546_),
    .Q(\flop44.q ));
 sg13g2_dfrbp_1 _1070_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net210),
    .D(net92),
    .Q_N(_0545_),
    .Q(\flop45.q ));
 sg13g2_dfrbp_1 _1071_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net204),
    .D(_0029_),
    .Q_N(_0544_),
    .Q(\flop46.q ));
 sg13g2_dfrbp_1 _1072_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net204),
    .D(net104),
    .Q_N(_0543_),
    .Q(\flop47.q ));
 sg13g2_dfrbp_1 _1073_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net203),
    .D(net132),
    .Q_N(_0542_),
    .Q(\flop48.q ));
 sg13g2_dfrbp_1 _1074_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net205),
    .D(_0032_),
    .Q_N(_0005_),
    .Q(\and11.b ));
 sg13g2_dfrbp_1 _1075_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net202),
    .D(_0033_),
    .Q_N(_0541_),
    .Q(\flop50.q ));
 sg13g2_dfrbp_1 _1076_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net211),
    .D(_0034_),
    .Q_N(_0012_),
    .Q(\flop51.q ));
 sg13g2_dfrbp_1 _1077_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net210),
    .D(net83),
    .Q_N(_0540_),
    .Q(\flop52.q ));
 sg13g2_dfrbp_1 _1078_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net210),
    .D(net97),
    .Q_N(_0539_),
    .Q(\flop53.q ));
 sg13g2_dfrbp_1 _1079_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net204),
    .D(_0037_),
    .Q_N(_0538_),
    .Q(\flop54.q ));
 sg13g2_dfrbp_1 _1080_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net205),
    .D(net90),
    .Q_N(_0537_),
    .Q(\flop55.q ));
 sg13g2_dfrbp_1 _1081_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net203),
    .D(net120),
    .Q_N(_0536_),
    .Q(\flop56.q ));
 sg13g2_dfrbp_1 _1082_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net203),
    .D(net125),
    .Q_N(_0535_),
    .Q(\flop57.q ));
 sg13g2_dfrbp_1 _1083_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net202),
    .D(_0041_),
    .Q_N(_0534_),
    .Q(\flop58.q ));
 sg13g2_dfrbp_1 _1084_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net209),
    .D(_0042_),
    .Q_N(_0004_),
    .Q(\and125.a ));
 sg13g2_dfrbp_1 _1085_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net211),
    .D(net100),
    .Q_N(_0533_),
    .Q(\flop60.q ));
 sg13g2_dfrbp_1 _1086_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net210),
    .D(net130),
    .Q_N(_0532_),
    .Q(\flop61.q ));
 sg13g2_dfrbp_1 _1087_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net204),
    .D(_0045_),
    .Q_N(_0531_),
    .Q(\flop62.q ));
 sg13g2_dfrbp_1 _1088_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net204),
    .D(net110),
    .Q_N(_0530_),
    .Q(\flop63.q ));
 sg13g2_dfrbp_1 _1089_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net203),
    .D(net108),
    .Q_N(_0529_),
    .Q(\flop64.q ));
 sg13g2_dfrbp_1 _1090_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net207),
    .D(net106),
    .Q_N(_0528_),
    .Q(\flop65.q ));
 sg13g2_dfrbp_1 _1091_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net202),
    .D(_0049_),
    .Q_N(_0527_),
    .Q(\flop66.q ));
 sg13g2_dfrbp_1 _1092_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net212),
    .D(_0050_),
    .Q_N(_0010_),
    .Q(\flop67.q ));
 sg13g2_dfrbp_1 _1093_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net211),
    .D(net88),
    .Q_N(_0526_),
    .Q(\flop68.q ));
 sg13g2_dfrbp_1 _1094_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net209),
    .D(_0052_),
    .Q_N(_0003_),
    .Q(\and126.a ));
 sg13g2_dfrbp_1 _1095_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net204),
    .D(_0053_),
    .Q_N(_0525_),
    .Q(\flop70.q ));
 sg13g2_dfrbp_1 _1096_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net204),
    .D(net122),
    .Q_N(_0524_),
    .Q(\flop71.q ));
 sg13g2_dfrbp_1 _1097_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net205),
    .D(net116),
    .Q_N(_0523_),
    .Q(\flop72.q ));
 sg13g2_dfrbp_1 _1098_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net202),
    .D(net128),
    .Q_N(_0522_),
    .Q(\flop73.q ));
 sg13g2_dfrbp_1 _1099_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net204),
    .D(_0057_),
    .Q_N(_0521_),
    .Q(\flop74.q ));
 sg13g2_dfrbp_1 _1100_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net214),
    .D(_0058_),
    .Q_N(_0014_),
    .Q(\and113.a ));
 sg13g2_dfrbp_1 _1101_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net214),
    .D(_0059_),
    .Q_N(_0520_),
    .Q(\and115.b ));
 sg13g2_dfrbp_1 _1102_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net213),
    .D(_0060_),
    .Q_N(_0001_),
    .Q(\and128.b ));
 sg13g2_dfrbp_1 _1103_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net213),
    .D(_0061_),
    .Q_N(_0000_),
    .Q(\and131.b ));
 sg13g2_dfrbp_1 _1104_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net207),
    .D(_0062_),
    .Q_N(_0002_),
    .Q(\and127.a ));
 sg13g2_dfrbp_1 _1105_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net214),
    .D(_0063_),
    .Q_N(_0519_),
    .Q(\and119.a ));
 sg13g2_dfrbp_1 _1106_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net213),
    .D(_0064_),
    .Q_N(_0547_),
    .Q(\and129.a ));
 sg13g2_dfrbp_1 _1107_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net208),
    .D(\flop83.d ),
    .Q_N(_0518_),
    .Q(\flop83.q ));
 sg13g2_dfrbp_1 _1108_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net213),
    .D(_0065_),
    .Q_N(_0517_),
    .Q(\and118.a ));
 sg13g2_dfrbp_1 _1109_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net213),
    .D(net136),
    .Q_N(_0516_),
    .Q(\flop84.q ));
 sg13g2_dfrbp_1 _1110_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net212),
    .D(_0067_),
    .Q_N(_0009_),
    .Q(\and116.a ));
 sg13g2_dfrbp_1 _1111_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net202),
    .D(net139),
    .Q_N(\flop29.notq ),
    .Q(\and84.a ));
 sg13g2_dfrbp_1 _1112_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net208),
    .D(net59),
    .Q_N(\flop39.notq ),
    .Q(\and104.b ));
 sg13g2_dfrbp_1 _1113_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net207),
    .D(net114),
    .Q_N(_0515_),
    .Q(\flop49.q ));
 sg13g2_dfrbp_1 _1114_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net211),
    .D(_0071_),
    .Q_N(_0011_),
    .Q(\flop59.q ));
 sg13g2_dfrbp_1 _1115_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net210),
    .D(_0072_),
    .Q_N(_0514_),
    .Q(\flop69.q ));
 sg13g2_dfrbp_1 _1116_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net213),
    .D(_0073_),
    .Q_N(_0548_),
    .Q(\and112.a ));
 sg13g2_dfrbp_1 _1117_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net213),
    .D(net9),
    .Q_N(_0549_),
    .Q(\flop10.d ));
 sg13g2_dfrbp_1 _1118_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net213),
    .D(net29),
    .Q_N(_0550_),
    .Q(\flop10.q ));
 sg13g2_dfrbp_1 _1119_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net211),
    .D(net31),
    .Q_N(_0513_),
    .Q(\flop11.q ));
 sg13g2_dfrbp_1 _1120_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net207),
    .D(_0074_),
    .Q_N(_0551_),
    .Q(\flop85.q ));
 sg13g2_dfrbp_1 _1121_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net214),
    .D(\flop12.d ),
    .Q_N(_0552_),
    .Q(\flop12.q ));
 sg13g2_dfrbp_1 _1122_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net209),
    .D(\flop13.d ),
    .Q_N(_0553_),
    .Q(\flop13.q ));
 sg13g2_dfrbp_1 _1123_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net214),
    .D(\flop14.d ),
    .Q_N(_0554_),
    .Q(\flop14.q ));
 sg13g2_dfrbp_1 _1124_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net209),
    .D(\flop15.d ),
    .Q_N(_0555_),
    .Q(\flop15.q ));
 sg13g2_dfrbp_1 _1125_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net209),
    .D(\flop16.d ),
    .Q_N(_0556_),
    .Q(\flop16.q ));
 sg13g2_dfrbp_1 _1126_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net209),
    .D(\flop17.d ),
    .Q_N(_0557_),
    .Q(\flop17.q ));
 sg13g2_dfrbp_1 _1127_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net208),
    .D(\flop18.d ),
    .Q_N(_0512_),
    .Q(\flop18.q ));
 sg13g2_dfrbp_1 _1128_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(_0015_),
    .D(net28),
    .Q_N(\flop19.d ),
    .Q(\and74.b ));
 sg13g2_dfrbp_1 _1129_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net210),
    .D(_0075_),
    .Q_N(_0008_),
    .Q(\and1.b ));
 sg13g2_dfrbp_1 _1130_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(_0016_),
    .D(net35),
    .Q_N(\flop20.notq ),
    .Q(\and74.a ));
 sg13g2_dfrbp_1 _1131_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(_0017_),
    .D(net142),
    .Q_N(\flop21.notq ),
    .Q(\and73.a ));
 sg13g2_dfrbp_1 _1132_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net160),
    .D(net49),
    .Q_N(\flop22.notq ),
    .Q(\and75.a ));
 sg13g2_dfrbp_1 _1133_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(_0019_),
    .D(net69),
    .Q_N(\flop23.notq ),
    .Q(\and76.a ));
 sg13g2_dfrbp_1 _1134_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(_0020_),
    .D(net72),
    .Q_N(\flop24.notq ),
    .Q(\and81.b ));
 sg13g2_dfrbp_1 _1135_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net211),
    .D(net30),
    .Q_N(_0558_),
    .Q(\flop26.q ));
 sg13g2_dfrbp_1 _1136_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net202),
    .D(net27),
    .Q_N(\flop27.d ),
    .Q(\and83.b ));
 sg13g2_dfrbp_1 _1137_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net211),
    .D(_0081_),
    .Q_N(_0511_),
    .Q(\flop25.q ));
 sg13g2_dfrbp_1 _1138_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net202),
    .D(net33),
    .Q_N(\flop28.notq ),
    .Q(\and83.a ));
 sg13g2_dfrbp_1 _1139_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net210),
    .D(_0083_),
    .Q_N(_0007_),
    .Q(\and122.a ));
 sg13g2_dfrbp_1 _1140_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net202),
    .D(net47),
    .Q_N(\flop30.notq ),
    .Q(\and85.a ));
 sg13g2_dfrbp_1 _1141_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net203),
    .D(net75),
    .Q_N(\flop31.notq ),
    .Q(\and86.a ));
 sg13g2_dfrbp_1 _1142_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net203),
    .D(net38),
    .Q_N(\flop32.notq ),
    .Q(\and100.a ));
 sg13g2_dfrbp_1 _1143_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net203),
    .D(net62),
    .Q_N(\flop33.notq ),
    .Q(\and82.a ));
 sg13g2_dfrbp_1 _1144_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net207),
    .D(net65),
    .Q_N(\flop34.notq ),
    .Q(\and92.a ));
 sg13g2_dfrbp_1 _1145_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net207),
    .D(net81),
    .Q_N(\flop35.notq ),
    .Q(\and93.a ));
 sg13g2_dfrbp_1 _1146_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net207),
    .D(net45),
    .Q_N(\flop36.notq ),
    .Q(\and94.a ));
 sg13g2_dfrbp_1 _1147_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net207),
    .D(net40),
    .Q_N(\flop37.notq ),
    .Q(\and101.a ));
 sg13g2_tiehi tt_um_wokwi_412635532198550529_26 (.L_HI(net26));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_wokwi_412635532198550529_14 (.L_LO(net14));
 sg13g2_tielo tt_um_wokwi_412635532198550529_15 (.L_LO(net15));
 sg13g2_tielo tt_um_wokwi_412635532198550529_16 (.L_LO(net16));
 sg13g2_tielo tt_um_wokwi_412635532198550529_17 (.L_LO(net17));
 sg13g2_tielo tt_um_wokwi_412635532198550529_18 (.L_LO(net18));
 sg13g2_tielo tt_um_wokwi_412635532198550529_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wokwi_412635532198550529_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wokwi_412635532198550529_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wokwi_412635532198550529_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wokwi_412635532198550529_23 (.L_LO(net23));
 sg13g2_tielo tt_um_wokwi_412635532198550529_24 (.L_LO(net24));
 sg13g2_tiehi tt_um_wokwi_412635532198550529_25 (.L_HI(net25));
 sg13g2_buf_2 _1162_ (.A(\flop84.q ),
    .X(uio_out[6]));
 sg13g2_buf_1 _1163_ (.A(\flop85.q ),
    .X(uio_out[7]));
 sg13g2_buf_1 _1164_ (.A(\flop12.q ),
    .X(uo_out[0]));
 sg13g2_buf_1 _1165_ (.A(\flop13.q ),
    .X(uo_out[1]));
 sg13g2_buf_1 _1166_ (.A(\flop14.q ),
    .X(uo_out[2]));
 sg13g2_buf_1 _1167_ (.A(\flop15.q ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1168_ (.A(\flop16.q ),
    .X(uo_out[4]));
 sg13g2_buf_1 _1169_ (.A(\flop17.q ),
    .X(uo_out[5]));
 sg13g2_buf_1 _1170_ (.A(\flop18.q ),
    .X(uo_out[6]));
 sg13g2_buf_1 _1171_ (.A(\flop83.q ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout162 (.A(_0332_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_0462_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(net166),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_0454_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(net168),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_0442_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(net170),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_0417_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_0409_),
    .X(net172));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(net174));
 sg13g2_buf_2 fanout174 (.A(_0418_),
    .X(net174));
 sg13g2_buf_4 fanout175 (.X(net175),
    .A(_0140_));
 sg13g2_buf_8 fanout176 (.A(_0139_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_0137_),
    .X(net177));
 sg13g2_buf_4 fanout178 (.X(net178),
    .A(_0098_));
 sg13g2_buf_2 fanout179 (.A(_0096_),
    .X(net179));
 sg13g2_buf_1 fanout180 (.A(_0096_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_0095_),
    .X(net181));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(net151));
 sg13g2_buf_2 fanout183 (.A(net148),
    .X(net183));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(net216));
 sg13g2_buf_2 fanout185 (.A(\and118.a ),
    .X(net185));
 sg13g2_buf_4 fanout186 (.X(net186),
    .A(net150));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(\and129.a ));
 sg13g2_buf_2 fanout188 (.A(\and119.a ),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(\and119.a ),
    .X(net189));
 sg13g2_buf_4 fanout190 (.X(net190),
    .A(net152));
 sg13g2_buf_2 fanout191 (.A(\and131.b ),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(net195),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(net194),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(\and113.a ),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(net197),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(net12),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(net199),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(uio_in[2]),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(uio_in[0]),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(uio_in[0]),
    .X(net201));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(net206));
 sg13g2_buf_4 fanout203 (.X(net203),
    .A(net206));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(net206));
 sg13g2_buf_2 fanout205 (.A(net206),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(net215),
    .X(net206));
 sg13g2_buf_4 fanout207 (.X(net207),
    .A(net209));
 sg13g2_buf_4 fanout208 (.X(net208),
    .A(net209));
 sg13g2_buf_4 fanout209 (.X(net209),
    .A(net215));
 sg13g2_buf_4 fanout210 (.X(net210),
    .A(net212));
 sg13g2_buf_4 fanout211 (.X(net211),
    .A(net212));
 sg13g2_buf_2 fanout212 (.A(net215),
    .X(net212));
 sg13g2_buf_4 fanout213 (.X(net213),
    .A(net214));
 sg13g2_buf_4 fanout214 (.X(net214),
    .A(net215));
 sg13g2_buf_2 fanout215 (.A(rst_n),
    .X(net215));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_tielo tt_um_wokwi_412635532198550529_13 (.L_LO(net13));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\flop27.d ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold2 (.A(\flop19.d ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold3 (.A(\flop10.d ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold4 (.A(\flop25.q ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold5 (.A(\flop10.q ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold6 (.A(\flop28.notq ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0082_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold8 (.A(\flop20.notq ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0076_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold10 (.A(\and100.a ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0507_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0086_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold13 (.A(\and101.a ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0091_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold15 (.A(\and108.b ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0414_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0024_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold18 (.A(\flop36.notq ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0090_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold20 (.A(\and85.a ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0084_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold22 (.A(\and75.a ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0078_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold24 (.A(\and107.b ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0023_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold26 (.A(\flop42.notq ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0025_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold28 (.A(\and102.a ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0405_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0021_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold31 (.A(\and104.b ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0495_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0069_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold34 (.A(\and82.a ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0508_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0087_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold37 (.A(\and92.a ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0509_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0088_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold40 (.A(\flop85.q ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold41 (.A(\and76.a ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0132_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0079_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold44 (.A(\and81.b ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0131_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0080_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold47 (.A(\and86.a ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0506_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0085_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold50 (.A(\flop58.q ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold51 (.A(\flop74.q ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold52 (.A(\flop69.q ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold53 (.A(\and93.a ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0510_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0089_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold56 (.A(\flop52.q ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0035_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold58 (.A(\flop66.q ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold59 (.A(\flop51.q ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold60 (.A(\flop68.q ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0464_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0051_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold63 (.A(\flop55.q ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0038_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold65 (.A(\flop45.q ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0028_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold67 (.A(\flop24.notq ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0130_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold69 (.A(\flop54.q ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold70 (.A(\flop53.q ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0036_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold72 (.A(\flop62.q ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold73 (.A(\flop60.q ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0043_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold75 (.A(\flop50.q ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold76 (.A(\flop67.q ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold77 (.A(\flop47.q ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0030_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold79 (.A(\flop65.q ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0048_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold81 (.A(\flop64.q ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0047_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold83 (.A(\flop63.q ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0046_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold85 (.A(\flop43.q ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold86 (.A(\flop59.q ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold87 (.A(\flop49.q ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0070_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold89 (.A(\flop72.q ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0055_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold91 (.A(\flop44.q ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0027_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold93 (.A(\flop56.q ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0039_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold95 (.A(\flop71.q ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0054_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold97 (.A(\flop46.q ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold98 (.A(\flop57.q ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0040_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold100 (.A(\flop70.q ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold101 (.A(\flop73.q ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0056_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold103 (.A(\flop61.q ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0044_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold105 (.A(\flop48.q ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0031_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold107 (.A(\and1.b ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold108 (.A(\and11.b ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold109 (.A(\flop84.q ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0066_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold111 (.A(\and84.a ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0494_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0068_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold114 (.A(\and73.a ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0133_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0077_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold117 (.A(\and125.a ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold118 (.A(\and10.a ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold119 (.A(\and126.a ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold120 (.A(\and122.a ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0004_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold122 (.A(\and116.a ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0493_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold124 (.A(\and129.a ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold125 (.A(\and112.a ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold126 (.A(\and127.a ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0005_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0009_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0006_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold130 (.A(\and115.b ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0008_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0007_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold133 (.A(\flop11.q ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0018_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold135 (.A(\flop11.q ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold136 (.A(\and118.a ),
    .X(net216));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_4 FILLER_12_371 ();
 sg13g2_fill_2 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_4 FILLER_13_364 ();
 sg13g2_fill_2 FILLER_13_373 ();
 sg13g2_fill_1 FILLER_13_375 ();
 sg13g2_fill_2 FILLER_13_385 ();
 sg13g2_fill_2 FILLER_13_394 ();
 sg13g2_fill_1 FILLER_13_396 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_4 FILLER_14_350 ();
 sg13g2_fill_2 FILLER_14_354 ();
 sg13g2_fill_1 FILLER_14_361 ();
 sg13g2_fill_2 FILLER_14_367 ();
 sg13g2_fill_1 FILLER_14_397 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_fill_1 FILLER_15_343 ();
 sg13g2_fill_2 FILLER_15_379 ();
 sg13g2_fill_1 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_fill_1 FILLER_16_329 ();
 sg13g2_fill_1 FILLER_16_334 ();
 sg13g2_fill_2 FILLER_16_339 ();
 sg13g2_fill_1 FILLER_16_341 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_4 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_121 ();
 sg13g2_decap_8 FILLER_17_128 ();
 sg13g2_decap_8 FILLER_17_135 ();
 sg13g2_decap_8 FILLER_17_142 ();
 sg13g2_decap_8 FILLER_17_149 ();
 sg13g2_decap_8 FILLER_17_156 ();
 sg13g2_decap_8 FILLER_17_163 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_177 ();
 sg13g2_decap_8 FILLER_17_184 ();
 sg13g2_decap_8 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_205 ();
 sg13g2_decap_8 FILLER_17_212 ();
 sg13g2_decap_8 FILLER_17_219 ();
 sg13g2_decap_8 FILLER_17_226 ();
 sg13g2_decap_8 FILLER_17_233 ();
 sg13g2_decap_8 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_247 ();
 sg13g2_decap_8 FILLER_17_254 ();
 sg13g2_decap_8 FILLER_17_261 ();
 sg13g2_decap_8 FILLER_17_268 ();
 sg13g2_decap_8 FILLER_17_275 ();
 sg13g2_decap_8 FILLER_17_282 ();
 sg13g2_decap_8 FILLER_17_289 ();
 sg13g2_decap_8 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_17_310 ();
 sg13g2_fill_2 FILLER_17_317 ();
 sg13g2_fill_1 FILLER_17_319 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_fill_2 FILLER_18_70 ();
 sg13g2_decap_4 FILLER_18_115 ();
 sg13g2_fill_2 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_147 ();
 sg13g2_fill_2 FILLER_18_153 ();
 sg13g2_fill_2 FILLER_18_159 ();
 sg13g2_decap_8 FILLER_18_170 ();
 sg13g2_decap_8 FILLER_18_177 ();
 sg13g2_decap_4 FILLER_18_184 ();
 sg13g2_fill_2 FILLER_18_188 ();
 sg13g2_decap_8 FILLER_18_204 ();
 sg13g2_fill_2 FILLER_18_224 ();
 sg13g2_fill_2 FILLER_18_231 ();
 sg13g2_fill_1 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_260 ();
 sg13g2_decap_8 FILLER_18_267 ();
 sg13g2_decap_8 FILLER_18_274 ();
 sg13g2_decap_8 FILLER_18_281 ();
 sg13g2_decap_8 FILLER_18_288 ();
 sg13g2_decap_8 FILLER_18_295 ();
 sg13g2_fill_1 FILLER_18_302 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_fill_1 FILLER_18_323 ();
 sg13g2_fill_1 FILLER_18_338 ();
 sg13g2_fill_2 FILLER_18_353 ();
 sg13g2_fill_1 FILLER_18_355 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_4 FILLER_19_70 ();
 sg13g2_fill_2 FILLER_19_74 ();
 sg13g2_fill_2 FILLER_19_114 ();
 sg13g2_fill_1 FILLER_19_116 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_133 ();
 sg13g2_fill_1 FILLER_19_217 ();
 sg13g2_fill_2 FILLER_19_223 ();
 sg13g2_decap_8 FILLER_19_260 ();
 sg13g2_decap_4 FILLER_19_267 ();
 sg13g2_fill_2 FILLER_19_271 ();
 sg13g2_decap_8 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_333 ();
 sg13g2_fill_2 FILLER_19_391 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_fill_2 FILLER_20_70 ();
 sg13g2_decap_4 FILLER_20_118 ();
 sg13g2_fill_2 FILLER_20_122 ();
 sg13g2_decap_4 FILLER_20_132 ();
 sg13g2_fill_2 FILLER_20_159 ();
 sg13g2_fill_1 FILLER_20_161 ();
 sg13g2_fill_2 FILLER_20_165 ();
 sg13g2_fill_1 FILLER_20_167 ();
 sg13g2_fill_2 FILLER_20_180 ();
 sg13g2_fill_1 FILLER_20_182 ();
 sg13g2_fill_2 FILLER_20_192 ();
 sg13g2_fill_1 FILLER_20_194 ();
 sg13g2_decap_4 FILLER_20_209 ();
 sg13g2_fill_2 FILLER_20_230 ();
 sg13g2_fill_2 FILLER_20_237 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_fill_2 FILLER_20_259 ();
 sg13g2_fill_1 FILLER_20_261 ();
 sg13g2_fill_2 FILLER_20_301 ();
 sg13g2_fill_1 FILLER_20_303 ();
 sg13g2_fill_2 FILLER_20_313 ();
 sg13g2_fill_1 FILLER_20_315 ();
 sg13g2_fill_1 FILLER_20_364 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_4 FILLER_21_63 ();
 sg13g2_fill_1 FILLER_21_67 ();
 sg13g2_fill_1 FILLER_21_117 ();
 sg13g2_decap_4 FILLER_21_182 ();
 sg13g2_fill_1 FILLER_21_186 ();
 sg13g2_fill_2 FILLER_21_226 ();
 sg13g2_fill_1 FILLER_21_228 ();
 sg13g2_decap_4 FILLER_21_281 ();
 sg13g2_fill_1 FILLER_21_325 ();
 sg13g2_fill_2 FILLER_21_335 ();
 sg13g2_fill_2 FILLER_21_375 ();
 sg13g2_fill_1 FILLER_21_377 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_fill_2 FILLER_22_56 ();
 sg13g2_fill_1 FILLER_22_58 ();
 sg13g2_fill_1 FILLER_22_85 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_fill_2 FILLER_22_238 ();
 sg13g2_fill_1 FILLER_22_240 ();
 sg13g2_fill_1 FILLER_22_254 ();
 sg13g2_fill_1 FILLER_22_359 ();
 sg13g2_fill_1 FILLER_22_377 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_fill_2 FILLER_23_109 ();
 sg13g2_fill_2 FILLER_23_145 ();
 sg13g2_fill_1 FILLER_23_147 ();
 sg13g2_fill_2 FILLER_23_218 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_fill_1 FILLER_23_231 ();
 sg13g2_fill_2 FILLER_23_267 ();
 sg13g2_fill_1 FILLER_23_269 ();
 sg13g2_fill_2 FILLER_23_279 ();
 sg13g2_fill_2 FILLER_23_310 ();
 sg13g2_fill_1 FILLER_23_312 ();
 sg13g2_fill_1 FILLER_23_322 ();
 sg13g2_fill_2 FILLER_23_362 ();
 sg13g2_fill_1 FILLER_23_369 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_4 FILLER_24_49 ();
 sg13g2_fill_2 FILLER_24_53 ();
 sg13g2_fill_2 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_139 ();
 sg13g2_fill_1 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_4 FILLER_24_252 ();
 sg13g2_fill_2 FILLER_24_328 ();
 sg13g2_fill_1 FILLER_24_349 ();
 sg13g2_fill_1 FILLER_24_368 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_4 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_121 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_fill_2 FILLER_25_180 ();
 sg13g2_fill_1 FILLER_25_182 ();
 sg13g2_fill_1 FILLER_25_192 ();
 sg13g2_decap_4 FILLER_25_206 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_247 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_decap_8 FILLER_25_265 ();
 sg13g2_decap_4 FILLER_25_272 ();
 sg13g2_fill_1 FILLER_25_276 ();
 sg13g2_fill_2 FILLER_25_318 ();
 sg13g2_fill_1 FILLER_25_320 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_95 ();
 sg13g2_fill_2 FILLER_26_148 ();
 sg13g2_fill_1 FILLER_26_150 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_fill_2 FILLER_26_208 ();
 sg13g2_decap_4 FILLER_26_223 ();
 sg13g2_fill_1 FILLER_26_227 ();
 sg13g2_fill_2 FILLER_26_252 ();
 sg13g2_fill_2 FILLER_26_280 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_fill_1 FILLER_26_352 ();
 sg13g2_fill_2 FILLER_26_358 ();
 sg13g2_fill_1 FILLER_26_360 ();
 sg13g2_fill_2 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_88 ();
 sg13g2_fill_1 FILLER_27_98 ();
 sg13g2_fill_2 FILLER_27_125 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_fill_2 FILLER_27_137 ();
 sg13g2_fill_1 FILLER_27_139 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_fill_1 FILLER_27_170 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_fill_2 FILLER_27_201 ();
 sg13g2_fill_2 FILLER_27_226 ();
 sg13g2_decap_4 FILLER_27_232 ();
 sg13g2_decap_8 FILLER_27_248 ();
 sg13g2_fill_2 FILLER_27_255 ();
 sg13g2_fill_1 FILLER_27_270 ();
 sg13g2_decap_8 FILLER_27_313 ();
 sg13g2_decap_4 FILLER_27_320 ();
 sg13g2_fill_1 FILLER_27_324 ();
 sg13g2_fill_2 FILLER_27_337 ();
 sg13g2_fill_1 FILLER_27_355 ();
 sg13g2_decap_8 FILLER_27_374 ();
 sg13g2_fill_1 FILLER_27_381 ();
 sg13g2_fill_2 FILLER_27_385 ();
 sg13g2_fill_1 FILLER_27_387 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_4 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_53 ();
 sg13g2_fill_2 FILLER_28_150 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_fill_2 FILLER_28_173 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_fill_1 FILLER_28_195 ();
 sg13g2_decap_8 FILLER_28_205 ();
 sg13g2_fill_1 FILLER_28_212 ();
 sg13g2_decap_8 FILLER_28_226 ();
 sg13g2_fill_2 FILLER_28_258 ();
 sg13g2_decap_8 FILLER_28_272 ();
 sg13g2_fill_2 FILLER_28_308 ();
 sg13g2_fill_1 FILLER_28_310 ();
 sg13g2_fill_1 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_347 ();
 sg13g2_fill_2 FILLER_28_366 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_4 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_53 ();
 sg13g2_fill_1 FILLER_29_170 ();
 sg13g2_fill_2 FILLER_29_186 ();
 sg13g2_decap_4 FILLER_29_236 ();
 sg13g2_fill_2 FILLER_29_240 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_decap_4 FILLER_29_275 ();
 sg13g2_fill_1 FILLER_29_279 ();
 sg13g2_fill_1 FILLER_29_285 ();
 sg13g2_fill_1 FILLER_29_299 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_decap_4 FILLER_29_336 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_fill_2 FILLER_29_365 ();
 sg13g2_fill_1 FILLER_29_367 ();
 sg13g2_decap_8 FILLER_29_377 ();
 sg13g2_fill_1 FILLER_29_394 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_89 ();
 sg13g2_fill_1 FILLER_30_91 ();
 sg13g2_fill_2 FILLER_30_115 ();
 sg13g2_fill_2 FILLER_30_140 ();
 sg13g2_fill_2 FILLER_30_156 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_fill_2 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_202 ();
 sg13g2_fill_2 FILLER_30_208 ();
 sg13g2_fill_2 FILLER_30_228 ();
 sg13g2_decap_4 FILLER_30_256 ();
 sg13g2_decap_4 FILLER_30_282 ();
 sg13g2_fill_1 FILLER_30_310 ();
 sg13g2_fill_2 FILLER_30_326 ();
 sg13g2_fill_1 FILLER_30_338 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_1 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_fill_2 FILLER_31_42 ();
 sg13g2_fill_1 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_123 ();
 sg13g2_fill_2 FILLER_31_161 ();
 sg13g2_fill_2 FILLER_31_185 ();
 sg13g2_decap_4 FILLER_31_204 ();
 sg13g2_fill_2 FILLER_31_213 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_fill_2 FILLER_31_254 ();
 sg13g2_fill_2 FILLER_31_259 ();
 sg13g2_decap_4 FILLER_31_279 ();
 sg13g2_fill_1 FILLER_31_283 ();
 sg13g2_fill_1 FILLER_31_296 ();
 sg13g2_decap_4 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_decap_8 FILLER_31_311 ();
 sg13g2_fill_2 FILLER_31_318 ();
 sg13g2_fill_2 FILLER_31_359 ();
 sg13g2_fill_1 FILLER_31_366 ();
 sg13g2_decap_4 FILLER_31_376 ();
 sg13g2_fill_1 FILLER_31_380 ();
 sg13g2_fill_2 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_403 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_fill_2 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_63 ();
 sg13g2_fill_1 FILLER_32_112 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_fill_1 FILLER_32_183 ();
 sg13g2_decap_8 FILLER_32_194 ();
 sg13g2_decap_8 FILLER_32_201 ();
 sg13g2_fill_2 FILLER_32_208 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_fill_1 FILLER_32_229 ();
 sg13g2_fill_2 FILLER_32_247 ();
 sg13g2_fill_2 FILLER_32_273 ();
 sg13g2_decap_4 FILLER_32_378 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_4 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_107 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_fill_1 FILLER_33_167 ();
 sg13g2_decap_8 FILLER_33_179 ();
 sg13g2_decap_8 FILLER_33_200 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_fill_1 FILLER_33_235 ();
 sg13g2_decap_8 FILLER_33_271 ();
 sg13g2_fill_2 FILLER_33_278 ();
 sg13g2_fill_1 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_289 ();
 sg13g2_decap_4 FILLER_33_296 ();
 sg13g2_fill_1 FILLER_33_300 ();
 sg13g2_decap_8 FILLER_33_305 ();
 sg13g2_decap_4 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_329 ();
 sg13g2_fill_2 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_353 ();
 sg13g2_fill_1 FILLER_33_359 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_96 ();
 sg13g2_fill_2 FILLER_34_131 ();
 sg13g2_fill_1 FILLER_34_160 ();
 sg13g2_fill_1 FILLER_34_187 ();
 sg13g2_decap_4 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_209 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_226 ();
 sg13g2_decap_8 FILLER_34_248 ();
 sg13g2_fill_1 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_311 ();
 sg13g2_fill_2 FILLER_34_318 ();
 sg13g2_fill_1 FILLER_34_320 ();
 sg13g2_fill_2 FILLER_34_343 ();
 sg13g2_fill_1 FILLER_34_350 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_decap_8 FILLER_34_383 ();
 sg13g2_fill_2 FILLER_34_390 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_4 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_32 ();
 sg13g2_fill_1 FILLER_35_60 ();
 sg13g2_fill_2 FILLER_35_94 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_fill_2 FILLER_35_131 ();
 sg13g2_fill_2 FILLER_35_160 ();
 sg13g2_decap_8 FILLER_35_173 ();
 sg13g2_decap_8 FILLER_35_190 ();
 sg13g2_decap_8 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_decap_8 FILLER_35_214 ();
 sg13g2_decap_8 FILLER_35_221 ();
 sg13g2_decap_8 FILLER_35_228 ();
 sg13g2_decap_4 FILLER_35_235 ();
 sg13g2_fill_2 FILLER_35_239 ();
 sg13g2_fill_2 FILLER_35_246 ();
 sg13g2_decap_8 FILLER_35_263 ();
 sg13g2_fill_2 FILLER_35_270 ();
 sg13g2_fill_1 FILLER_35_272 ();
 sg13g2_decap_4 FILLER_35_277 ();
 sg13g2_fill_1 FILLER_35_281 ();
 sg13g2_decap_8 FILLER_35_311 ();
 sg13g2_fill_1 FILLER_35_318 ();
 sg13g2_fill_2 FILLER_35_344 ();
 sg13g2_fill_1 FILLER_35_346 ();
 sg13g2_fill_2 FILLER_35_375 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_fill_1 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_79 ();
 sg13g2_decap_8 FILLER_36_111 ();
 sg13g2_decap_4 FILLER_36_123 ();
 sg13g2_fill_1 FILLER_36_127 ();
 sg13g2_decap_4 FILLER_36_133 ();
 sg13g2_decap_4 FILLER_36_161 ();
 sg13g2_decap_4 FILLER_36_192 ();
 sg13g2_fill_2 FILLER_36_226 ();
 sg13g2_decap_4 FILLER_36_233 ();
 sg13g2_decap_4 FILLER_36_245 ();
 sg13g2_fill_2 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_341 ();
 sg13g2_fill_1 FILLER_36_343 ();
 sg13g2_fill_2 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_51 ();
 sg13g2_decap_8 FILLER_37_87 ();
 sg13g2_decap_8 FILLER_37_94 ();
 sg13g2_fill_1 FILLER_37_101 ();
 sg13g2_fill_2 FILLER_37_128 ();
 sg13g2_fill_2 FILLER_37_135 ();
 sg13g2_fill_1 FILLER_37_145 ();
 sg13g2_fill_2 FILLER_37_185 ();
 sg13g2_decap_8 FILLER_37_199 ();
 sg13g2_decap_8 FILLER_37_206 ();
 sg13g2_fill_2 FILLER_37_213 ();
 sg13g2_fill_1 FILLER_37_215 ();
 sg13g2_decap_8 FILLER_37_246 ();
 sg13g2_decap_4 FILLER_37_253 ();
 sg13g2_fill_1 FILLER_37_271 ();
 sg13g2_decap_4 FILLER_37_276 ();
 sg13g2_decap_8 FILLER_37_284 ();
 sg13g2_fill_1 FILLER_37_351 ();
 sg13g2_fill_2 FILLER_37_364 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_fill_2 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_51 ();
 sg13g2_fill_1 FILLER_38_64 ();
 sg13g2_fill_2 FILLER_38_78 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_fill_1 FILLER_38_153 ();
 sg13g2_fill_1 FILLER_38_193 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_231 ();
 sg13g2_fill_1 FILLER_38_233 ();
 sg13g2_fill_2 FILLER_38_264 ();
 sg13g2_fill_1 FILLER_38_266 ();
 sg13g2_fill_1 FILLER_38_293 ();
 sg13g2_fill_2 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_329 ();
 sg13g2_fill_1 FILLER_38_360 ();
 sg13g2_fill_1 FILLER_38_387 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net13;
 assign uio_oe[1] = net14;
 assign uio_oe[2] = net15;
 assign uio_oe[3] = net16;
 assign uio_oe[4] = net17;
 assign uio_oe[5] = net18;
 assign uio_oe[6] = net25;
 assign uio_oe[7] = net26;
 assign uio_out[0] = net19;
 assign uio_out[1] = net20;
 assign uio_out[2] = net21;
 assign uio_out[3] = net22;
 assign uio_out[4] = net23;
 assign uio_out[5] = net24;
endmodule

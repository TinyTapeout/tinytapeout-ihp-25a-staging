module tt_um_htfab_bouncy_capsule (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire bitmap_pixel;
 wire \capsule_color[0] ;
 wire \capsule_color[1] ;
 wire \capsule_color[2] ;
 wire \capsule_color[3] ;
 wire \center_x[0] ;
 wire \center_x[1] ;
 wire \center_x[2] ;
 wire \center_x[3] ;
 wire \center_x[4] ;
 wire \center_x[5] ;
 wire \center_x[6] ;
 wire \center_x[7] ;
 wire \center_x[8] ;
 wire \center_x[9] ;
 wire \center_y[0] ;
 wire \center_y[1] ;
 wire \center_y[2] ;
 wire \center_y[3] ;
 wire \center_y[4] ;
 wire \center_y[5] ;
 wire \center_y[6] ;
 wire \center_y[7] ;
 wire \center_y[8] ;
 wire \center_y[9] ;
 wire \collision_impact[0] ;
 wire \collision_impact[1] ;
 wire \color_entropy[0] ;
 wire \color_entropy[1] ;
 wire handle_impact;
 wire hsync;
 wire \i_bitmap.in[0] ;
 wire \i_bitmap.in[10] ;
 wire \i_bitmap.in[11] ;
 wire \i_bitmap.in[12] ;
 wire \i_bitmap.in[1] ;
 wire \i_bitmap.in[2] ;
 wire \i_bitmap.in[3] ;
 wire \i_bitmap.in[4] ;
 wire \i_bitmap.in[5] ;
 wire \i_bitmap.in[6] ;
 wire \i_bitmap.in[7] ;
 wire \i_bitmap.in[8] ;
 wire \i_bitmap.in[9] ;
 wire \i_capsule.tf_x[0] ;
 wire \i_capsule.tf_x[8] ;
 wire \i_capsule.tf_x[9] ;
 wire \i_capsule.tf_y[0] ;
 wire \i_capsule.tf_y[7] ;
 wire \i_capsule.tf_y[8] ;
 wire \i_capsule.tf_y[9] ;
 wire \i_collision.i_coll_table.in[0] ;
 wire \i_collision.i_coll_table.in[1] ;
 wire \i_collision.i_coll_table.in[3] ;
 wire \i_collision.i_coll_table.in[4] ;
 wire \i_collision.i_coll_table.in[5] ;
 wire \i_collision.mirror ;
 wire \i_collision.phi[1] ;
 wire \i_collision.rotate ;
 wire \i_collision.update ;
 wire \i_collision.vx[0] ;
 wire \i_collision.vx[1] ;
 wire \i_collision.vx[2] ;
 wire \i_collision.vy[0] ;
 wire \i_collision.vy[1] ;
 wire \i_collision.vy[2] ;
 wire \i_colors.capsule_color[4] ;
 wire \i_colors.capsule_color[5] ;
 wire \i_colors.channel[0] ;
 wire \i_colors.channel[1] ;
 wire \i_colors.channel[2] ;
 wire \i_delta_sigma.acc[0] ;
 wire \i_delta_sigma.acc[10] ;
 wire \i_delta_sigma.acc[11] ;
 wire \i_delta_sigma.acc[12] ;
 wire \i_delta_sigma.acc[13] ;
 wire \i_delta_sigma.acc[1] ;
 wire \i_delta_sigma.acc[2] ;
 wire \i_delta_sigma.acc[3] ;
 wire \i_delta_sigma.acc[4] ;
 wire \i_delta_sigma.acc[5] ;
 wire \i_delta_sigma.acc[6] ;
 wire \i_delta_sigma.acc[7] ;
 wire \i_delta_sigma.acc[8] ;
 wire \i_delta_sigma.acc[9] ;
 wire \i_delta_sigma.sample[0] ;
 wire \i_delta_sigma.sample[10] ;
 wire \i_delta_sigma.sample[11] ;
 wire \i_delta_sigma.sample[1] ;
 wire \i_delta_sigma.sample[2] ;
 wire \i_delta_sigma.sample[3] ;
 wire \i_delta_sigma.sample[4] ;
 wire \i_delta_sigma.sample[5] ;
 wire \i_delta_sigma.sample[6] ;
 wire \i_delta_sigma.sample[7] ;
 wire \i_delta_sigma.sample[8] ;
 wire \i_delta_sigma.sample[9] ;
 wire \i_kinematics.center_x_lo[0] ;
 wire \i_kinematics.center_x_lo[1] ;
 wire \i_kinematics.center_y_lo[0] ;
 wire \i_kinematics.center_y_lo[1] ;
 wire \i_kinematics.phi[0] ;
 wire \i_kinematics.phi[10] ;
 wire \i_kinematics.phi[1] ;
 wire \i_kinematics.phi[2] ;
 wire \i_kinematics.phi[3] ;
 wire \i_kinematics.phi[4] ;
 wire \i_kinematics.phi[5] ;
 wire \i_kinematics.phi[6] ;
 wire \i_kinematics.phi[7] ;
 wire \i_kinematics.update ;
 wire \i_orchestrator.hit_bottom ;
 wire \i_orchestrator.hit_left ;
 wire \i_orchestrator.hit_priority[0] ;
 wire \i_orchestrator.hit_priority[1] ;
 wire \i_orchestrator.hit_right ;
 wire \i_orchestrator.hit_top ;
 wire \i_orchestrator.lfsr[1] ;
 wire \i_orchestrator.lfsr[2] ;
 wire \i_orchestrator.lfsr[3] ;
 wire \i_orchestrator.lfsr[4] ;
 wire \i_orchestrator.lfsr[5] ;
 wire \i_orchestrator.lfsr[6] ;
 wire \i_orchestrator.lfsr[7] ;
 wire \i_orchestrator.sample_counter[0] ;
 wire \i_orchestrator.sample_counter[1] ;
 wire \i_orchestrator.sample_counter[2] ;
 wire \i_orchestrator.sample_counter[3] ;
 wire \i_orchestrator.sample_counter[4] ;
 wire \i_orchestrator.sample_counter[5] ;
 wire \i_orchestrator.sample_counter[6] ;
 wire \i_orchestrator.sample_counter[7] ;
 wire \i_orchestrator.sample_counter[8] ;
 wire \i_orchestrator.sample_counter[9] ;
 wire \i_orchestrator.tension[1] ;
 wire \i_orchestrator.tension[2] ;
 wire \i_orchestrator.tension[3] ;
 wire \i_orchestrator.trigger_debounce ;
 wire \i_orchestrator.trigger_resonator[0] ;
 wire \i_orchestrator.trigger_resonator[1] ;
 wire \i_orchestrator.update_resonator ;
 wire \i_orchestrator.update_transform ;
 wire \i_orchestrator.vga_x[0] ;
 wire \i_orchestrator.vga_x[1] ;
 wire \i_orchestrator.vga_x[2] ;
 wire \i_orchestrator.vga_x[3] ;
 wire \i_orchestrator.vga_x[4] ;
 wire \i_orchestrator.vga_x[5] ;
 wire \i_orchestrator.vga_x[6] ;
 wire \i_orchestrator.vga_x[7] ;
 wire \i_orchestrator.vga_x[8] ;
 wire \i_orchestrator.vga_x[9] ;
 wire \i_orchestrator.vga_y[0] ;
 wire \i_orchestrator.vga_y[1] ;
 wire \i_orchestrator.vga_y[2] ;
 wire \i_orchestrator.vga_y[3] ;
 wire \i_orchestrator.vga_y[4] ;
 wire \i_orchestrator.vga_y[5] ;
 wire \i_orchestrator.vga_y[6] ;
 wire \i_orchestrator.vga_y[7] ;
 wire \i_orchestrator.vga_y[8] ;
 wire \i_orchestrator.vga_y[9] ;
 wire \i_resonator.counter[0] ;
 wire \i_resonator.counter[1] ;
 wire \i_resonator.counter[2] ;
 wire \i_resonator.counter[3] ;
 wire \i_resonator.v[0] ;
 wire \i_resonator.v[10] ;
 wire \i_resonator.v[11] ;
 wire \i_resonator.v[12] ;
 wire \i_resonator.v[13] ;
 wire \i_resonator.v[14] ;
 wire \i_resonator.v[15] ;
 wire \i_resonator.v[1] ;
 wire \i_resonator.v[2] ;
 wire \i_resonator.v[3] ;
 wire \i_resonator.v[4] ;
 wire \i_resonator.v[5] ;
 wire \i_resonator.v[6] ;
 wire \i_resonator.v[7] ;
 wire \i_resonator.v[8] ;
 wire \i_resonator.v[9] ;
 wire \i_transform.image_x[0] ;
 wire \i_transform.image_x[1] ;
 wire \i_transform.image_x[2] ;
 wire \i_transform.image_x[3] ;
 wire \i_transform.image_x[4] ;
 wire \i_transform.image_x[5] ;
 wire \i_transform.image_y[0] ;
 wire \i_transform.image_y[1] ;
 wire \i_transform.image_y[2] ;
 wire \i_transform.image_y[3] ;
 wire \i_transform.image_y[4] ;
 wire \i_transform.image_y[5] ;
 wire \i_transform.track_x[0] ;
 wire \i_transform.track_x[1] ;
 wire \i_transform.track_x[2] ;
 wire \i_transform.track_x[3] ;
 wire \i_transform.track_x[4] ;
 wire \i_transform.track_x[5] ;
 wire \i_transform.track_x[6] ;
 wire \i_transform.track_x[7] ;
 wire \i_transform.track_x[8] ;
 wire \i_transform.track_x[9] ;
 wire \i_transform.track_y[0] ;
 wire \i_transform.track_y[1] ;
 wire \i_transform.track_y[2] ;
 wire \i_transform.track_y[3] ;
 wire \i_transform.track_y[4] ;
 wire \i_transform.track_y[5] ;
 wire \i_transform.track_y[6] ;
 wire \i_transform.track_y[7] ;
 wire \i_transform.track_y[8] ;
 wire \i_transform.track_y[9] ;
 wire \i_vga_beam.vsync ;
 wire orient;
 wire pdm_out;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire clknet_leaf_0_clk;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;

 sg13g2_inv_2 _3226_ (.Y(_2373_),
    .A(net996));
 sg13g2_inv_4 _3227_ (.A(net998),
    .Y(_2374_));
 sg13g2_inv_1 _3228_ (.Y(_2375_),
    .A(net1010));
 sg13g2_inv_1 _3229_ (.Y(_2376_),
    .A(net550));
 sg13g2_inv_2 _3230_ (.Y(_2377_),
    .A(net546));
 sg13g2_inv_1 _3231_ (.Y(_2378_),
    .A(\i_resonator.v[9] ));
 sg13g2_inv_1 _3232_ (.Y(_2379_),
    .A(\i_resonator.v[8] ));
 sg13g2_inv_1 _3233_ (.Y(_2380_),
    .A(net1013));
 sg13g2_inv_1 _3234_ (.Y(_2381_),
    .A(\i_delta_sigma.sample[8] ));
 sg13g2_inv_1 _3235_ (.Y(_2382_),
    .A(\i_delta_sigma.sample[7] ));
 sg13g2_inv_1 _3236_ (.Y(_2383_),
    .A(\i_delta_sigma.sample[6] ));
 sg13g2_inv_1 _3237_ (.Y(_2384_),
    .A(net356));
 sg13g2_inv_2 _3238_ (.Y(_2385_),
    .A(net1016));
 sg13g2_inv_1 _3239_ (.Y(_2386_),
    .A(\capsule_color[3] ));
 sg13g2_inv_1 _3240_ (.Y(_2387_),
    .A(net1019));
 sg13g2_inv_1 _3241_ (.Y(_2388_),
    .A(net247));
 sg13g2_inv_1 _3242_ (.Y(_2389_),
    .A(\i_transform.image_x[3] ));
 sg13g2_inv_1 _3243_ (.Y(_2390_),
    .A(\i_transform.image_y[3] ));
 sg13g2_inv_1 _3244_ (.Y(_2391_),
    .A(net1039));
 sg13g2_inv_1 _3245_ (.Y(_2392_),
    .A(net1020));
 sg13g2_inv_1 _3246_ (.Y(_2393_),
    .A(\i_kinematics.phi[5] ));
 sg13g2_inv_1 _3247_ (.Y(_2394_),
    .A(\i_kinematics.phi[1] ));
 sg13g2_inv_1 _3248_ (.Y(_2395_),
    .A(\center_x[3] ));
 sg13g2_inv_2 _3249_ (.Y(_2396_),
    .A(net1027));
 sg13g2_inv_1 _3250_ (.Y(_2397_),
    .A(net385));
 sg13g2_inv_1 _3251_ (.Y(_2398_),
    .A(net372));
 sg13g2_inv_2 _3252_ (.Y(_2399_),
    .A(\i_capsule.tf_x[9] ));
 sg13g2_inv_1 _3253_ (.Y(_2400_),
    .A(\i_capsule.tf_x[8] ));
 sg13g2_inv_1 _3254_ (.Y(_2401_),
    .A(\i_bitmap.in[6] ));
 sg13g2_inv_1 _3255_ (.Y(_2402_),
    .A(\i_bitmap.in[4] ));
 sg13g2_inv_1 _3256_ (.Y(_2403_),
    .A(net1032));
 sg13g2_inv_1 _3257_ (.Y(_2404_),
    .A(net365));
 sg13g2_inv_1 _3258_ (.Y(_2405_),
    .A(net381));
 sg13g2_inv_1 _3259_ (.Y(_2406_),
    .A(net338));
 sg13g2_inv_1 _3260_ (.Y(_2407_),
    .A(net295));
 sg13g2_inv_1 _3261_ (.Y(_2408_),
    .A(net279));
 sg13g2_inv_1 _3262_ (.Y(_2409_),
    .A(net292));
 sg13g2_inv_1 _3263_ (.Y(_2410_),
    .A(net268));
 sg13g2_inv_1 _3264_ (.Y(_2411_),
    .A(\i_orchestrator.lfsr[4] ));
 sg13g2_inv_1 _3265_ (.Y(_2412_),
    .A(net266));
 sg13g2_inv_1 _3266_ (.Y(_2413_),
    .A(net270));
 sg13g2_inv_4 _3267_ (.A(net1049),
    .Y(_2414_));
 sg13g2_inv_1 _3268_ (.Y(_2415_),
    .A(net240));
 sg13g2_inv_1 _3269_ (.Y(_2416_),
    .A(\i_capsule.tf_y[8] ));
 sg13g2_inv_1 _3270_ (.Y(_2417_),
    .A(\i_capsule.tf_y[7] ));
 sg13g2_inv_1 _3271_ (.Y(_2418_),
    .A(\i_bitmap.in[11] ));
 sg13g2_inv_1 _3272_ (.Y(_2419_),
    .A(\i_delta_sigma.acc[10] ));
 sg13g2_inv_1 _3273_ (.Y(_2420_),
    .A(\i_delta_sigma.acc[8] ));
 sg13g2_inv_1 _3274_ (.Y(_2421_),
    .A(net346));
 sg13g2_inv_1 _3275_ (.Y(_2422_),
    .A(net1053));
 sg13g2_inv_1 _3276_ (.Y(_2423_),
    .A(net325));
 sg13g2_inv_1 _3277_ (.Y(_2424_),
    .A(\i_transform.track_y[6] ));
 sg13g2_inv_2 _3278_ (.Y(_2425_),
    .A(net370));
 sg13g2_inv_1 _3279_ (.Y(_2426_),
    .A(\i_transform.track_y[4] ));
 sg13g2_inv_1 _3280_ (.Y(_2427_),
    .A(\i_transform.track_y[9] ));
 sg13g2_inv_1 _3281_ (.Y(_2428_),
    .A(_0062_));
 sg13g2_inv_1 _3282_ (.Y(_2429_),
    .A(net264));
 sg13g2_inv_1 _3283_ (.Y(_2430_),
    .A(\i_transform.track_x[2] ));
 sg13g2_inv_2 _3284_ (.Y(_2431_),
    .A(net1072));
 sg13g2_inv_1 _3285_ (.Y(_2432_),
    .A(\i_orchestrator.trigger_resonator[0] ));
 sg13g2_inv_2 _3286_ (.Y(_2433_),
    .A(net1047));
 sg13g2_inv_1 _3287_ (.Y(_2434_),
    .A(_0009_));
 sg13g2_inv_1 _3288_ (.Y(_2435_),
    .A(net272));
 sg13g2_inv_1 _3289_ (.Y(_2436_),
    .A(net376));
 sg13g2_inv_1 _3290_ (.Y(_2437_),
    .A(net281));
 sg13g2_inv_1 _3291_ (.Y(_2438_),
    .A(_0019_));
 sg13g2_inv_1 _3292_ (.Y(_2439_),
    .A(_0029_));
 sg13g2_inv_1 _3293_ (.Y(_2440_),
    .A(_0034_));
 sg13g2_inv_1 _3294_ (.Y(_2441_),
    .A(_0036_));
 sg13g2_inv_1 _3295_ (.Y(_2442_),
    .A(_0037_));
 sg13g2_inv_1 _3296_ (.Y(_2443_),
    .A(_0038_));
 sg13g2_inv_1 _3297_ (.Y(_2444_),
    .A(_0050_));
 sg13g2_nor2b_1 _3298_ (.A(net7),
    .B_N(net450),
    .Y(_2445_));
 sg13g2_nand2b_2 _3299_ (.Y(_2446_),
    .B(net450),
    .A_N(net7));
 sg13g2_nand4_1 _3300_ (.B(net1075),
    .C(net423),
    .A(net306),
    .Y(_2447_),
    .D(_2445_));
 sg13g2_nand3_1 _3301_ (.B(\i_colors.channel[2] ),
    .C(_2446_),
    .A(net1075),
    .Y(_2448_));
 sg13g2_nand2b_1 _3302_ (.Y(_2449_),
    .B(net1075),
    .A_N(net306));
 sg13g2_nor2_1 _3303_ (.A(_2446_),
    .B(_2449_),
    .Y(_2450_));
 sg13g2_nand2_1 _3304_ (.Y(_2451_),
    .A(net432),
    .B(_2450_));
 sg13g2_nand3_1 _3305_ (.B(_2448_),
    .C(_2451_),
    .A(_2447_),
    .Y(_0003_));
 sg13g2_nand3_1 _3306_ (.B(net449),
    .C(_2445_),
    .A(net306),
    .Y(_2452_));
 sg13g2_nand3_1 _3307_ (.B(net432),
    .C(_2446_),
    .A(net1075),
    .Y(_2453_));
 sg13g2_a21oi_1 _3308_ (.A1(net423),
    .A2(_2450_),
    .Y(_2454_),
    .B1(net1066));
 sg13g2_nand3_1 _3309_ (.B(_2453_),
    .C(_2454_),
    .A(_2452_),
    .Y(_0001_));
 sg13g2_nand4_1 _3310_ (.B(net1075),
    .C(\i_colors.channel[0] ),
    .A(net306),
    .Y(_2455_),
    .D(_2445_));
 sg13g2_nand3_1 _3311_ (.B(net423),
    .C(_2446_),
    .A(net1075),
    .Y(_2456_));
 sg13g2_nand2_1 _3312_ (.Y(_2457_),
    .A(\i_colors.channel[2] ),
    .B(_2450_));
 sg13g2_nand3_1 _3313_ (.B(_2456_),
    .C(_2457_),
    .A(_2455_),
    .Y(_0002_));
 sg13g2_nor2_2 _3314_ (.A(net4),
    .B(\i_delta_sigma.acc[13] ),
    .Y(pdm_out));
 sg13g2_nand2_1 _3315_ (.Y(_2458_),
    .A(\i_orchestrator.vga_y[7] ),
    .B(\i_orchestrator.vga_y[6] ));
 sg13g2_and3_2 _3316_ (.X(_2459_),
    .A(\i_orchestrator.vga_y[7] ),
    .B(\i_orchestrator.vga_y[6] ),
    .C(\i_orchestrator.vga_y[5] ));
 sg13g2_nor2b_2 _3317_ (.A(net382),
    .B_N(\i_orchestrator.vga_y[8] ),
    .Y(_2460_));
 sg13g2_nand2_2 _3318_ (.Y(_2461_),
    .A(_2459_),
    .B(_2460_));
 sg13g2_nand3b_1 _3319_ (.B(net1057),
    .C(net1055),
    .Y(_2462_),
    .A_N(net1059));
 sg13g2_or4_1 _3320_ (.A(net1053),
    .B(net533),
    .C(_2461_),
    .D(_2462_),
    .X(_2463_));
 sg13g2_nor2_1 _3321_ (.A(\i_orchestrator.vga_y[9] ),
    .B(\i_orchestrator.vga_y[8] ),
    .Y(_2464_));
 sg13g2_or2_1 _3322_ (.X(_2465_),
    .B(\i_orchestrator.vga_y[8] ),
    .A(\i_orchestrator.vga_y[9] ));
 sg13g2_a21o_1 _3323_ (.A2(net1057),
    .A1(net1059),
    .B1(net1056),
    .X(_2466_));
 sg13g2_nand4_1 _3324_ (.B(_2459_),
    .C(_2465_),
    .A(net1055),
    .Y(_2467_),
    .D(_2466_));
 sg13g2_nor2_1 _3325_ (.A(net1059),
    .B(net1057),
    .Y(_2468_));
 sg13g2_nand2_1 _3326_ (.Y(_2469_),
    .A(net1056),
    .B(net1055));
 sg13g2_o21ai_1 _3327_ (.B1(_2422_),
    .Y(_2470_),
    .A1(_2468_),
    .A2(_2469_));
 sg13g2_nand2_1 _3328_ (.Y(_2471_),
    .A(net1057),
    .B(_2460_));
 sg13g2_a221oi_1 _3329_ (.B2(_2459_),
    .C1(_2471_),
    .B1(_2470_),
    .A1(_2463_),
    .Y(_0007_),
    .A2(_2467_));
 sg13g2_and3_1 _3330_ (.X(_2472_),
    .A(net538),
    .B(net1062),
    .C(net307));
 sg13g2_nor3_1 _3331_ (.A(\i_orchestrator.vga_x[4] ),
    .B(net1062),
    .C(\i_orchestrator.vga_x[6] ),
    .Y(_2473_));
 sg13g2_nand2_1 _3332_ (.Y(_2474_),
    .A(net1061),
    .B(net1060));
 sg13g2_nor4_1 _3333_ (.A(net417),
    .B(_2472_),
    .C(_2473_),
    .D(_2474_),
    .Y(_0006_));
 sg13g2_nor2_2 _3334_ (.A(net1069),
    .B(net535),
    .Y(_2475_));
 sg13g2_nand2b_1 _3335_ (.Y(_2476_),
    .B(net1073),
    .A_N(\i_orchestrator.update_transform ));
 sg13g2_xnor2_1 _3336_ (.Y(_2477_),
    .A(\i_kinematics.phi[10] ),
    .B(orient));
 sg13g2_xor2_1 _3337_ (.B(orient),
    .A(\i_kinematics.phi[10] ),
    .X(_2478_));
 sg13g2_xnor2_1 _3338_ (.Y(_2479_),
    .A(_0031_),
    .B(net971));
 sg13g2_inv_1 _3339_ (.Y(_2480_),
    .A(_2479_));
 sg13g2_xor2_1 _3340_ (.B(net1022),
    .A(net1020),
    .X(_2481_));
 sg13g2_xnor2_1 _3341_ (.Y(_2482_),
    .A(net1020),
    .B(net1022));
 sg13g2_xor2_1 _3342_ (.B(\i_kinematics.phi[7] ),
    .A(net1022),
    .X(_2483_));
 sg13g2_xnor2_1 _3343_ (.Y(_2484_),
    .A(net1022),
    .B(\i_kinematics.phi[7] ));
 sg13g2_xor2_1 _3344_ (.B(\i_kinematics.phi[6] ),
    .A(net1021),
    .X(_2485_));
 sg13g2_xnor2_1 _3345_ (.Y(_2486_),
    .A(net1021),
    .B(\i_kinematics.phi[6] ));
 sg13g2_xor2_1 _3346_ (.B(\i_kinematics.phi[5] ),
    .A(net1021),
    .X(_2487_));
 sg13g2_xnor2_1 _3347_ (.Y(_2488_),
    .A(net1021),
    .B(\i_kinematics.phi[5] ));
 sg13g2_xor2_1 _3348_ (.B(\i_kinematics.phi[4] ),
    .A(net1021),
    .X(_2489_));
 sg13g2_xnor2_1 _3349_ (.Y(_2490_),
    .A(net1021),
    .B(\i_kinematics.phi[4] ));
 sg13g2_xor2_1 _3350_ (.B(\i_kinematics.phi[3] ),
    .A(net1021),
    .X(_2491_));
 sg13g2_xnor2_1 _3351_ (.Y(_2492_),
    .A(net1021),
    .B(\i_kinematics.phi[3] ));
 sg13g2_o21ai_1 _3352_ (.B1(net957),
    .Y(_2493_),
    .A1(net955),
    .A2(_2491_));
 sg13g2_and2_1 _3353_ (.A(net959),
    .B(_2493_),
    .X(_2494_));
 sg13g2_nor2_2 _3354_ (.A(net963),
    .B(_2494_),
    .Y(_2495_));
 sg13g2_nor2_1 _3355_ (.A(net965),
    .B(_2495_),
    .Y(_2496_));
 sg13g2_nand2_1 _3356_ (.Y(_2497_),
    .A(net957),
    .B(_2489_));
 sg13g2_nand4_1 _3357_ (.B(net961),
    .C(_2487_),
    .A(_2483_),
    .Y(_2498_),
    .D(_2489_));
 sg13g2_nor2_1 _3358_ (.A(net957),
    .B(net955),
    .Y(_2499_));
 sg13g2_nand2_1 _3359_ (.Y(_2500_),
    .A(_2488_),
    .B(_2490_));
 sg13g2_o21ai_1 _3360_ (.B1(net963),
    .Y(_2501_),
    .A1(net959),
    .A2(_2499_));
 sg13g2_a22oi_1 _3361_ (.Y(_2502_),
    .B1(_2501_),
    .B2(_2496_),
    .A2(_2498_),
    .A1(net965));
 sg13g2_nand2_1 _3362_ (.Y(_2503_),
    .A(net956),
    .B(_2491_));
 sg13g2_nor3_1 _3363_ (.A(net960),
    .B(net957),
    .C(net954),
    .Y(_2504_));
 sg13g2_xnor2_1 _3364_ (.Y(_2505_),
    .A(_2490_),
    .B(_2504_));
 sg13g2_nor2_1 _3365_ (.A(net956),
    .B(_2491_),
    .Y(_2506_));
 sg13g2_nor3_1 _3366_ (.A(net957),
    .B(net955),
    .C(net954),
    .Y(_2507_));
 sg13g2_nand3_1 _3367_ (.B(_2490_),
    .C(_2491_),
    .A(net956),
    .Y(_2508_));
 sg13g2_o21ai_1 _3368_ (.B1(net960),
    .Y(_2509_),
    .A1(_2506_),
    .A2(_2507_));
 sg13g2_nand2_1 _3369_ (.Y(_2510_),
    .A(net955),
    .B(_2491_));
 sg13g2_nand2_1 _3370_ (.Y(_2511_),
    .A(net955),
    .B(net954));
 sg13g2_nand3_1 _3371_ (.B(net955),
    .C(net954),
    .A(net956),
    .Y(_2512_));
 sg13g2_a21oi_1 _3372_ (.A1(_2490_),
    .A2(_2491_),
    .Y(_2513_),
    .B1(net961));
 sg13g2_a21oi_1 _3373_ (.A1(_2512_),
    .A2(_2513_),
    .Y(_2514_),
    .B1(net962));
 sg13g2_a22oi_1 _3374_ (.Y(_2515_),
    .B1(_2509_),
    .B2(_2514_),
    .A2(_2505_),
    .A1(net962));
 sg13g2_xor2_1 _3375_ (.B(\i_kinematics.phi[3] ),
    .A(\i_kinematics.phi[4] ),
    .X(_2516_));
 sg13g2_nor2_1 _3376_ (.A(net956),
    .B(_2516_),
    .Y(_2517_));
 sg13g2_mux2_1 _3377_ (.A0(_2490_),
    .A1(_2516_),
    .S(net957),
    .X(_2518_));
 sg13g2_nand2_1 _3378_ (.Y(_2519_),
    .A(net960),
    .B(_2518_));
 sg13g2_nor3_2 _3379_ (.A(net956),
    .B(_2490_),
    .C(net954),
    .Y(_2520_));
 sg13g2_a21oi_1 _3380_ (.A1(net958),
    .A2(_2520_),
    .Y(_2521_),
    .B1(_2483_));
 sg13g2_nand2_1 _3381_ (.Y(_2522_),
    .A(_2519_),
    .B(_2521_));
 sg13g2_nor3_1 _3382_ (.A(net958),
    .B(net955),
    .C(net954),
    .Y(_2523_));
 sg13g2_a221oi_1 _3383_ (.B2(net956),
    .C1(_2523_),
    .B1(_2511_),
    .A1(net958),
    .Y(_2524_),
    .A2(_2506_));
 sg13g2_nor2_1 _3384_ (.A(net958),
    .B(net957),
    .Y(_2525_));
 sg13g2_and2_1 _3385_ (.A(net956),
    .B(_2523_),
    .X(_2526_));
 sg13g2_o21ai_1 _3386_ (.B1(_2483_),
    .Y(_2527_),
    .A1(_2524_),
    .A2(_2526_));
 sg13g2_nand3_1 _3387_ (.B(_2522_),
    .C(_2527_),
    .A(net964),
    .Y(_2528_));
 sg13g2_or2_1 _3388_ (.X(_2529_),
    .B(_2515_),
    .A(net964));
 sg13g2_and2_1 _3389_ (.A(_2528_),
    .B(_2529_),
    .X(_2530_));
 sg13g2_and3_1 _3390_ (.X(_2531_),
    .A(net967),
    .B(_2528_),
    .C(_2529_));
 sg13g2_nor3_1 _3391_ (.A(net958),
    .B(net957),
    .C(net954),
    .Y(_2532_));
 sg13g2_nor3_1 _3392_ (.A(_2506_),
    .B(_2507_),
    .C(_2532_),
    .Y(_2533_));
 sg13g2_o21ai_1 _3393_ (.B1(net958),
    .Y(_2534_),
    .A1(_2507_),
    .A2(_2517_));
 sg13g2_and2_1 _3394_ (.A(net961),
    .B(_2516_),
    .X(_2535_));
 sg13g2_a21oi_1 _3395_ (.A1(_2508_),
    .A2(_2535_),
    .Y(_2536_),
    .B1(net962));
 sg13g2_a22oi_1 _3396_ (.Y(_2537_),
    .B1(_2534_),
    .B2(_2536_),
    .A2(_2533_),
    .A1(net962));
 sg13g2_nor2_1 _3397_ (.A(net964),
    .B(_2537_),
    .Y(_2538_));
 sg13g2_nand3b_1 _3398_ (.B(net960),
    .C(_2500_),
    .Y(_2539_),
    .A_N(_2520_));
 sg13g2_nand2_1 _3399_ (.Y(_2540_),
    .A(net962),
    .B(_2539_));
 sg13g2_or2_1 _3400_ (.X(_2541_),
    .B(_2518_),
    .A(net960));
 sg13g2_a21oi_1 _3401_ (.A1(net955),
    .A2(net954),
    .Y(_2542_),
    .B1(net958));
 sg13g2_a21oi_1 _3402_ (.A1(_2503_),
    .A2(_2542_),
    .Y(_2543_),
    .B1(net962));
 sg13g2_a22oi_1 _3403_ (.Y(_2544_),
    .B1(_2541_),
    .B2(_2543_),
    .A2(_2539_),
    .A1(net963));
 sg13g2_a21oi_2 _3404_ (.B1(_2538_),
    .Y(_2545_),
    .A2(_2544_),
    .A1(net964));
 sg13g2_a21oi_1 _3405_ (.A1(net960),
    .A2(_2518_),
    .Y(_2546_),
    .B1(_2483_));
 sg13g2_nand3_1 _3406_ (.B(_2493_),
    .C(_2500_),
    .A(net958),
    .Y(_2547_));
 sg13g2_a21oi_1 _3407_ (.A1(_2510_),
    .A2(_2525_),
    .Y(_2548_),
    .B1(net962));
 sg13g2_nand2_1 _3408_ (.Y(_2549_),
    .A(net961),
    .B(_2520_));
 sg13g2_a221oi_1 _3409_ (.B2(_2510_),
    .C1(net962),
    .B1(_2525_),
    .A1(net960),
    .Y(_2550_),
    .A2(_2520_));
 sg13g2_a22oi_1 _3410_ (.Y(_2551_),
    .B1(_2547_),
    .B2(_2550_),
    .A2(_2546_),
    .A1(_2541_));
 sg13g2_nor2_1 _3411_ (.A(net965),
    .B(_2551_),
    .Y(_2552_));
 sg13g2_a21oi_1 _3412_ (.A1(_2492_),
    .A2(_2499_),
    .Y(_2553_),
    .B1(net959));
 sg13g2_nand2_1 _3413_ (.Y(_2554_),
    .A(_2497_),
    .B(_2553_));
 sg13g2_a22oi_1 _3414_ (.Y(_2555_),
    .B1(_2554_),
    .B2(_2495_),
    .A2(_2549_),
    .A1(net963));
 sg13g2_a21oi_2 _3415_ (.B1(_2552_),
    .Y(_2556_),
    .A2(_2555_),
    .A1(net964));
 sg13g2_nor3_1 _3416_ (.A(_2531_),
    .B(_2545_),
    .C(_2556_),
    .Y(_2557_));
 sg13g2_nor2_1 _3417_ (.A(net971),
    .B(_2557_),
    .Y(_2558_));
 sg13g2_o21ai_1 _3418_ (.B1(_2495_),
    .Y(_2559_),
    .A1(net959),
    .A2(_2497_));
 sg13g2_o21ai_1 _3419_ (.B1(_2548_),
    .Y(_2560_),
    .A1(net960),
    .A2(_2493_));
 sg13g2_o21ai_1 _3420_ (.B1(_2560_),
    .Y(_2561_),
    .A1(_2494_),
    .A2(_2540_));
 sg13g2_mux2_1 _3421_ (.A0(_2559_),
    .A1(_2561_),
    .S(_2482_),
    .X(_2562_));
 sg13g2_nor4_1 _3422_ (.A(_2531_),
    .B(_2545_),
    .C(_2556_),
    .D(_2562_),
    .Y(_2563_));
 sg13g2_nor2_1 _3423_ (.A(net971),
    .B(_2563_),
    .Y(_2564_));
 sg13g2_a21oi_1 _3424_ (.A1(_2502_),
    .A2(_2563_),
    .Y(_2565_),
    .B1(net971));
 sg13g2_xnor2_1 _3425_ (.Y(_2566_),
    .A(_2496_),
    .B(_2565_));
 sg13g2_nand2_1 _3426_ (.Y(_2567_),
    .A(\i_transform.image_y[5] ),
    .B(net899));
 sg13g2_xnor2_1 _3427_ (.Y(_2568_),
    .A(\i_transform.image_y[5] ),
    .B(net899));
 sg13g2_xnor2_1 _3428_ (.Y(_2569_),
    .A(_2558_),
    .B(_2562_));
 sg13g2_nor2_1 _3429_ (.A(_2390_),
    .B(net898),
    .Y(_2570_));
 sg13g2_xnor2_1 _3430_ (.Y(_2571_),
    .A(_2390_),
    .B(net898));
 sg13g2_and2_1 _3431_ (.A(\i_transform.image_y[0] ),
    .B(net909),
    .X(_2572_));
 sg13g2_xor2_1 _3432_ (.B(_2545_),
    .A(_2531_),
    .X(_2573_));
 sg13g2_inv_1 _3433_ (.Y(_2574_),
    .A(_2573_));
 sg13g2_xnor2_1 _3434_ (.Y(_2575_),
    .A(_0013_),
    .B(_2573_));
 sg13g2_and2_1 _3435_ (.A(\i_transform.image_y[1] ),
    .B(_2573_),
    .X(_2576_));
 sg13g2_a21o_1 _3436_ (.A2(_2575_),
    .A1(_2572_),
    .B1(_2576_),
    .X(_2577_));
 sg13g2_o21ai_1 _3437_ (.B1(net967),
    .Y(_2578_),
    .A1(net909),
    .A2(_2545_));
 sg13g2_xor2_1 _3438_ (.B(_2578_),
    .A(_2556_),
    .X(_2579_));
 sg13g2_xnor2_1 _3439_ (.Y(_2580_),
    .A(\i_transform.image_y[2] ),
    .B(_2579_));
 sg13g2_nand2_1 _3440_ (.Y(_2581_),
    .A(_2577_),
    .B(_2580_));
 sg13g2_nor2_1 _3441_ (.A(_0014_),
    .B(_2579_),
    .Y(_2582_));
 sg13g2_a21oi_1 _3442_ (.A1(_2577_),
    .A2(_2580_),
    .Y(_2583_),
    .B1(_2582_));
 sg13g2_nor2_1 _3443_ (.A(_2571_),
    .B(_2583_),
    .Y(_2584_));
 sg13g2_xor2_1 _3444_ (.B(_2564_),
    .A(_2502_),
    .X(_2585_));
 sg13g2_xnor2_1 _3445_ (.Y(_2586_),
    .A(\i_transform.image_y[4] ),
    .B(_2585_));
 sg13g2_o21ai_1 _3446_ (.B1(_2586_),
    .Y(_2587_),
    .A1(_2570_),
    .A2(_2584_));
 sg13g2_or2_1 _3447_ (.X(_2588_),
    .B(_2585_),
    .A(_0016_));
 sg13g2_a21o_1 _3448_ (.A2(_2588_),
    .A1(_2587_),
    .B1(_2568_),
    .X(_2589_));
 sg13g2_xnor2_1 _3449_ (.Y(_2590_),
    .A(_0032_),
    .B(net967));
 sg13g2_inv_1 _3450_ (.Y(_2591_),
    .A(_2590_));
 sg13g2_a21oi_1 _3451_ (.A1(_2567_),
    .A2(_2589_),
    .Y(_2592_),
    .B1(_2591_));
 sg13g2_a21o_1 _3452_ (.A2(_0031_),
    .A1(\i_capsule.tf_y[0] ),
    .B1(\i_bitmap.in[7] ),
    .X(_2593_));
 sg13g2_a22oi_1 _3453_ (.Y(_2594_),
    .B1(_2593_),
    .B2(net966),
    .A2(_2592_),
    .A1(_2480_));
 sg13g2_xnor2_1 _3454_ (.Y(_2595_),
    .A(_2440_),
    .B(net970));
 sg13g2_inv_1 _3455_ (.Y(_2596_),
    .A(_2595_));
 sg13g2_nand2b_2 _3456_ (.Y(_2597_),
    .B(_2460_),
    .A_N(_2459_));
 sg13g2_nand2_1 _3457_ (.Y(_2598_),
    .A(_2465_),
    .B(_2597_));
 sg13g2_o21ai_1 _3458_ (.B1(net1060),
    .Y(_2599_),
    .A1(net1061),
    .A2(\i_orchestrator.vga_x[8] ));
 sg13g2_and2_1 _3459_ (.A(net928),
    .B(_2599_),
    .X(_2600_));
 sg13g2_nand2_1 _3460_ (.Y(_2601_),
    .A(net928),
    .B(_2599_));
 sg13g2_a21oi_1 _3461_ (.A1(net1060),
    .A2(net918),
    .Y(_2602_),
    .B1(_0068_));
 sg13g2_nand2_1 _3462_ (.Y(_2603_),
    .A(\i_orchestrator.vga_x[8] ),
    .B(net918));
 sg13g2_a21oi_1 _3463_ (.A1(\i_transform.track_x[8] ),
    .A2(_2603_),
    .Y(_2604_),
    .B1(_2602_));
 sg13g2_or2_1 _3464_ (.X(_2605_),
    .B(_2603_),
    .A(\i_transform.track_x[8] ));
 sg13g2_nand2_1 _3465_ (.Y(_2606_),
    .A(\i_orchestrator.vga_x[6] ),
    .B(net917));
 sg13g2_xor2_1 _3466_ (.B(_2606_),
    .A(\i_transform.track_x[6] ),
    .X(_2607_));
 sg13g2_nand3_1 _3467_ (.B(_0065_),
    .C(net920),
    .A(\i_orchestrator.vga_x[7] ),
    .Y(_2608_));
 sg13g2_a21o_1 _3468_ (.A2(net918),
    .A1(net1061),
    .B1(_0065_),
    .X(_2609_));
 sg13g2_nand3_1 _3469_ (.B(_0066_),
    .C(net918),
    .A(net1062),
    .Y(_2610_));
 sg13g2_nand4_1 _3470_ (.B(_2608_),
    .C(_2609_),
    .A(_2607_),
    .Y(_2611_),
    .D(_2610_));
 sg13g2_nand3_1 _3471_ (.B(_0067_),
    .C(net917),
    .A(\i_orchestrator.vga_x[4] ),
    .Y(_2612_));
 sg13g2_a21oi_1 _3472_ (.A1(\i_orchestrator.vga_x[3] ),
    .A2(net917),
    .Y(_2613_),
    .B1(_0064_));
 sg13g2_nand2_1 _3473_ (.Y(_2614_),
    .A(\i_orchestrator.vga_x[2] ),
    .B(net919));
 sg13g2_a21oi_1 _3474_ (.A1(\i_transform.track_x[2] ),
    .A2(_2614_),
    .Y(_2615_),
    .B1(_2613_));
 sg13g2_nand3_1 _3475_ (.B(_2430_),
    .C(net917),
    .A(\i_orchestrator.vga_x[2] ),
    .Y(_2616_));
 sg13g2_nand3_1 _3476_ (.B(_0064_),
    .C(net917),
    .A(\i_orchestrator.vga_x[3] ),
    .Y(_2617_));
 sg13g2_nand3_1 _3477_ (.B(_2616_),
    .C(_2617_),
    .A(_2615_),
    .Y(_2618_));
 sg13g2_nor2_1 _3478_ (.A(_0074_),
    .B(_2601_),
    .Y(_2619_));
 sg13g2_nand2_1 _3479_ (.Y(_2620_),
    .A(_0063_),
    .B(_2619_));
 sg13g2_nand2_1 _3480_ (.Y(_2621_),
    .A(\i_orchestrator.vga_x[1] ),
    .B(net919));
 sg13g2_o21ai_1 _3481_ (.B1(_2620_),
    .Y(_2622_),
    .A1(\i_transform.track_x[1] ),
    .A2(_2621_));
 sg13g2_nand2_1 _3482_ (.Y(_2623_),
    .A(\i_transform.track_x[1] ),
    .B(_2621_));
 sg13g2_a21oi_1 _3483_ (.A1(_2622_),
    .A2(_2623_),
    .Y(_2624_),
    .B1(_2618_));
 sg13g2_nor2b_1 _3484_ (.A(_2615_),
    .B_N(_2617_),
    .Y(_2625_));
 sg13g2_o21ai_1 _3485_ (.B1(_2612_),
    .Y(_2626_),
    .A1(_2624_),
    .A2(_2625_));
 sg13g2_a21oi_1 _3486_ (.A1(net1062),
    .A2(net917),
    .Y(_2627_),
    .B1(_0066_));
 sg13g2_a21oi_1 _3487_ (.A1(\i_orchestrator.vga_x[4] ),
    .A2(net917),
    .Y(_2628_),
    .B1(_0067_));
 sg13g2_nor2_1 _3488_ (.A(_2627_),
    .B(_2628_),
    .Y(_2629_));
 sg13g2_a21o_1 _3489_ (.A2(_2629_),
    .A1(_2626_),
    .B1(_2611_),
    .X(_2630_));
 sg13g2_nand3_1 _3490_ (.B(_2606_),
    .C(_2608_),
    .A(\i_transform.track_x[6] ),
    .Y(_2631_));
 sg13g2_nand3_1 _3491_ (.B(_2630_),
    .C(_2631_),
    .A(_2609_),
    .Y(_2632_));
 sg13g2_and2_1 _3492_ (.A(_2605_),
    .B(_2632_),
    .X(_2633_));
 sg13g2_nor2b_1 _3493_ (.A(_2633_),
    .B_N(_2604_),
    .Y(_2634_));
 sg13g2_nand3_1 _3494_ (.B(_0068_),
    .C(net917),
    .A(net1060),
    .Y(_2635_));
 sg13g2_nand3_1 _3495_ (.B(_2430_),
    .C(\i_transform.track_x[5] ),
    .A(_2429_),
    .Y(_2636_));
 sg13g2_nor4_1 _3496_ (.A(\i_transform.track_x[0] ),
    .B(\i_transform.track_x[1] ),
    .C(\i_transform.track_x[4] ),
    .D(_2636_),
    .Y(_2637_));
 sg13g2_nand2b_1 _3497_ (.Y(_2638_),
    .B(_0066_),
    .A_N(\i_transform.track_x[8] ));
 sg13g2_or4_1 _3498_ (.A(\i_transform.track_x[7] ),
    .B(\i_transform.track_x[6] ),
    .C(\i_transform.track_x[9] ),
    .D(_2638_),
    .X(_2639_));
 sg13g2_o21ai_1 _3499_ (.B1(_2635_),
    .Y(_2640_),
    .A1(_2637_),
    .A2(_2639_));
 sg13g2_or2_1 _3500_ (.X(_2641_),
    .B(_2619_),
    .A(_0063_));
 sg13g2_nor3_1 _3501_ (.A(_2622_),
    .B(_2627_),
    .C(_2628_),
    .Y(_2642_));
 sg13g2_nand4_1 _3502_ (.B(_2623_),
    .C(_2635_),
    .A(_2604_),
    .Y(_2643_),
    .D(_2642_));
 sg13g2_nand3_1 _3503_ (.B(_2612_),
    .C(_2641_),
    .A(_2605_),
    .Y(_2644_));
 sg13g2_nor4_2 _3504_ (.A(_2611_),
    .B(_2618_),
    .C(_2643_),
    .Y(_2645_),
    .D(_2644_));
 sg13g2_or2_1 _3505_ (.X(_2646_),
    .B(_2644_),
    .A(_2611_));
 sg13g2_nor3_1 _3506_ (.A(_2634_),
    .B(_2640_),
    .C(_2645_),
    .Y(_2647_));
 sg13g2_or3_2 _3507_ (.A(_2634_),
    .B(_2640_),
    .C(_2645_),
    .X(_2648_));
 sg13g2_xnor2_1 _3508_ (.Y(_2649_),
    .A(_2594_),
    .B(_2596_));
 sg13g2_a21oi_1 _3509_ (.A1(net1053),
    .A2(net926),
    .Y(_2650_),
    .B1(_0061_));
 sg13g2_a21oi_1 _3510_ (.A1(net1052),
    .A2(net926),
    .Y(_2651_),
    .B1(_0060_));
 sg13g2_nor2_1 _3511_ (.A(_2650_),
    .B(_2651_),
    .Y(_2652_));
 sg13g2_nand3_1 _3512_ (.B(_0061_),
    .C(net926),
    .A(net1053),
    .Y(_2653_));
 sg13g2_nand3_1 _3513_ (.B(_0058_),
    .C(net926),
    .A(net1055),
    .Y(_2654_));
 sg13g2_and2_1 _3514_ (.A(_2653_),
    .B(_2654_),
    .X(_2655_));
 sg13g2_nand2_1 _3515_ (.Y(_2656_),
    .A(_2652_),
    .B(_2655_));
 sg13g2_nand3_1 _3516_ (.B(_0060_),
    .C(net926),
    .A(net1052),
    .Y(_2657_));
 sg13g2_nand2_1 _3517_ (.Y(_2658_),
    .A(\i_orchestrator.vga_y[6] ),
    .B(net927));
 sg13g2_o21ai_1 _3518_ (.B1(_2657_),
    .Y(_2659_),
    .A1(\i_transform.track_y[6] ),
    .A2(_2658_));
 sg13g2_a21oi_1 _3519_ (.A1(net1055),
    .A2(net927),
    .Y(_2660_),
    .B1(_0058_));
 sg13g2_nand2_1 _3520_ (.Y(_2661_),
    .A(net1056),
    .B(net926));
 sg13g2_a21o_1 _3521_ (.A2(_2661_),
    .A1(\i_transform.track_y[2] ),
    .B1(_2660_),
    .X(_2662_));
 sg13g2_nand2_1 _3522_ (.Y(_2663_),
    .A(net1058),
    .B(net927));
 sg13g2_nand2_1 _3523_ (.Y(_2664_),
    .A(\i_transform.track_y[1] ),
    .B(_2663_));
 sg13g2_a21oi_1 _3524_ (.A1(_2465_),
    .A2(_2597_),
    .Y(_2665_),
    .B1(_0073_));
 sg13g2_nand2_1 _3525_ (.Y(_2666_),
    .A(_0057_),
    .B(_2665_));
 sg13g2_o21ai_1 _3526_ (.B1(_2666_),
    .Y(_2667_),
    .A1(\i_transform.track_y[1] ),
    .A2(_2663_));
 sg13g2_nor2b_1 _3527_ (.A(_2667_),
    .B_N(_2664_),
    .Y(_2668_));
 sg13g2_nor2_1 _3528_ (.A(\i_transform.track_y[2] ),
    .B(_2661_),
    .Y(_2669_));
 sg13g2_a21oi_1 _3529_ (.A1(\i_transform.track_y[8] ),
    .A2(_2597_),
    .Y(_2670_),
    .B1(_2428_));
 sg13g2_o21ai_1 _3530_ (.B1(_2670_),
    .Y(_2671_),
    .A1(_0057_),
    .A2(_2665_));
 sg13g2_nor2_1 _3531_ (.A(_2669_),
    .B(_2671_),
    .Y(_2672_));
 sg13g2_a21oi_1 _3532_ (.A1(\i_orchestrator.vga_y[7] ),
    .A2(net926),
    .Y(_2673_),
    .B1(_0059_));
 sg13g2_a21o_1 _3533_ (.A2(_2658_),
    .A1(\i_transform.track_y[6] ),
    .B1(_2673_),
    .X(_2674_));
 sg13g2_nand3_1 _3534_ (.B(_0059_),
    .C(net926),
    .A(\i_orchestrator.vga_y[7] ),
    .Y(_2675_));
 sg13g2_o21ai_1 _3535_ (.B1(_2675_),
    .Y(_2676_),
    .A1(\i_transform.track_y[8] ),
    .A2(_2597_));
 sg13g2_inv_1 _3536_ (.Y(_2677_),
    .A(_2676_));
 sg13g2_nor3_1 _3537_ (.A(_2656_),
    .B(_2659_),
    .C(_2674_),
    .Y(_2678_));
 sg13g2_nor2_1 _3538_ (.A(_2662_),
    .B(_2676_),
    .Y(_2679_));
 sg13g2_and4_1 _3539_ (.A(_2668_),
    .B(_2672_),
    .C(_2678_),
    .D(_2679_),
    .X(_2680_));
 sg13g2_nand4_1 _3540_ (.B(_2672_),
    .C(_2678_),
    .A(_2668_),
    .Y(_2681_),
    .D(_2679_));
 sg13g2_nand2_1 _3541_ (.Y(_2682_),
    .A(_0033_),
    .B(_2530_));
 sg13g2_xnor2_1 _3542_ (.Y(_2683_),
    .A(_0032_),
    .B(_2573_));
 sg13g2_nor2b_1 _3543_ (.A(_2683_),
    .B_N(_2682_),
    .Y(_2684_));
 sg13g2_a21oi_1 _3544_ (.A1(\i_capsule.tf_y[0] ),
    .A2(_2574_),
    .Y(_2685_),
    .B1(_2684_));
 sg13g2_xnor2_1 _3545_ (.Y(_2686_),
    .A(_0031_),
    .B(_2579_));
 sg13g2_nor2b_1 _3546_ (.A(_2685_),
    .B_N(_2686_),
    .Y(_2687_));
 sg13g2_a21o_1 _3547_ (.A2(_2579_),
    .A1(\i_bitmap.in[7] ),
    .B1(_2687_),
    .X(_2688_));
 sg13g2_xnor2_1 _3548_ (.Y(_2689_),
    .A(_2440_),
    .B(_2569_));
 sg13g2_nor2b_1 _3549_ (.A(_2688_),
    .B_N(_2689_),
    .Y(_2690_));
 sg13g2_nor2b_1 _3550_ (.A(_2689_),
    .B_N(_2688_),
    .Y(_2691_));
 sg13g2_nor3_1 _3551_ (.A(net874),
    .B(_2690_),
    .C(_2691_),
    .Y(_2692_));
 sg13g2_nor2_1 _3552_ (.A(net902),
    .B(_2692_),
    .Y(_2693_));
 sg13g2_o21ai_1 _3553_ (.B1(_2693_),
    .Y(_2694_),
    .A1(net877),
    .A2(_2649_));
 sg13g2_and2_2 _3554_ (.A(_2645_),
    .B(_2680_),
    .X(_2695_));
 sg13g2_nand2_1 _3555_ (.Y(_2696_),
    .A(_2645_),
    .B(net906));
 sg13g2_xnor2_1 _3556_ (.Y(_2697_),
    .A(net1020),
    .B(net971));
 sg13g2_xnor2_1 _3557_ (.Y(_2698_),
    .A(_2392_),
    .B(net971));
 sg13g2_xnor2_1 _3558_ (.Y(_2699_),
    .A(\i_bitmap.in[7] ),
    .B(net939));
 sg13g2_nor2_1 _3559_ (.A(_2482_),
    .B(_2495_),
    .Y(_2700_));
 sg13g2_mux2_1 _3560_ (.A0(_2559_),
    .A1(_2561_),
    .S(net965),
    .X(_2701_));
 sg13g2_nand2b_1 _3561_ (.Y(_2702_),
    .B(net964),
    .A_N(_2515_));
 sg13g2_nand3_1 _3562_ (.B(_2522_),
    .C(_2527_),
    .A(_2482_),
    .Y(_2703_));
 sg13g2_nand2_2 _3563_ (.Y(_2704_),
    .A(_2702_),
    .B(_2703_));
 sg13g2_and2_2 _3564_ (.A(_2702_),
    .B(_2703_),
    .X(_2705_));
 sg13g2_nor2_1 _3565_ (.A(net964),
    .B(_2544_),
    .Y(_2706_));
 sg13g2_a21oi_2 _3566_ (.B1(_2706_),
    .Y(_2707_),
    .A2(_2537_),
    .A1(net964));
 sg13g2_nor2_1 _3567_ (.A(_2482_),
    .B(_2551_),
    .Y(_2708_));
 sg13g2_a21oi_1 _3568_ (.A1(_2482_),
    .A2(_2555_),
    .Y(_2709_),
    .B1(_2708_));
 sg13g2_a21oi_2 _3569_ (.B1(net936),
    .Y(_2710_),
    .A2(_2707_),
    .A1(_2704_));
 sg13g2_and2_1 _3570_ (.A(net939),
    .B(_2709_),
    .X(_2711_));
 sg13g2_nor2_1 _3571_ (.A(_2710_),
    .B(_2711_),
    .Y(_2712_));
 sg13g2_and2_1 _3572_ (.A(net939),
    .B(_2701_),
    .X(_2713_));
 sg13g2_nor3_1 _3573_ (.A(_2710_),
    .B(_2711_),
    .C(_2713_),
    .Y(_2714_));
 sg13g2_a22oi_1 _3574_ (.Y(_2715_),
    .B1(_2501_),
    .B2(_2700_),
    .A2(_2498_),
    .A1(_2482_));
 sg13g2_o21ai_1 _3575_ (.B1(_2714_),
    .Y(_2716_),
    .A1(net936),
    .A2(_2715_));
 sg13g2_xnor2_1 _3576_ (.Y(_2717_),
    .A(_2700_),
    .B(_2716_));
 sg13g2_or2_1 _3577_ (.X(_2718_),
    .B(_2717_),
    .A(_0033_));
 sg13g2_xnor2_1 _3578_ (.Y(_2719_),
    .A(_0033_),
    .B(_2717_));
 sg13g2_inv_1 _3579_ (.Y(_2720_),
    .A(_2719_));
 sg13g2_xor2_1 _3580_ (.B(_2712_),
    .A(_2701_),
    .X(_2721_));
 sg13g2_nand2b_1 _3581_ (.Y(_2722_),
    .B(_2721_),
    .A_N(_0015_));
 sg13g2_nand3_1 _3582_ (.B(_2702_),
    .C(_2703_),
    .A(net939),
    .Y(_2723_));
 sg13g2_xor2_1 _3583_ (.B(_2723_),
    .A(_2707_),
    .X(_2724_));
 sg13g2_inv_1 _3584_ (.Y(_2725_),
    .A(_2724_));
 sg13g2_or2_1 _3585_ (.X(_2726_),
    .B(_2724_),
    .A(_0013_));
 sg13g2_xnor2_1 _3586_ (.Y(_2727_),
    .A(_0013_),
    .B(_2724_));
 sg13g2_a21o_1 _3587_ (.A2(_2705_),
    .A1(_0012_),
    .B1(_2727_),
    .X(_2728_));
 sg13g2_xnor2_1 _3588_ (.Y(_2729_),
    .A(_2709_),
    .B(_2710_));
 sg13g2_xor2_1 _3589_ (.B(_2729_),
    .A(_0014_),
    .X(_2730_));
 sg13g2_a21o_1 _3590_ (.A2(_2728_),
    .A1(_2726_),
    .B1(_2730_),
    .X(_2731_));
 sg13g2_nand2_1 _3591_ (.Y(_2732_),
    .A(\i_transform.image_y[2] ),
    .B(_2729_));
 sg13g2_xor2_1 _3592_ (.B(_2721_),
    .A(_0015_),
    .X(_2733_));
 sg13g2_a21o_1 _3593_ (.A2(_2732_),
    .A1(_2731_),
    .B1(_2733_),
    .X(_2734_));
 sg13g2_xnor2_1 _3594_ (.Y(_2735_),
    .A(_2714_),
    .B(_2715_));
 sg13g2_xor2_1 _3595_ (.B(_2735_),
    .A(_0016_),
    .X(_2736_));
 sg13g2_a21oi_1 _3596_ (.A1(_2722_),
    .A2(_2734_),
    .Y(_2737_),
    .B1(_2736_));
 sg13g2_and2_1 _3597_ (.A(\i_transform.image_y[4] ),
    .B(_2735_),
    .X(_2738_));
 sg13g2_o21ai_1 _3598_ (.B1(_2720_),
    .Y(_2739_),
    .A1(_2737_),
    .A2(_2738_));
 sg13g2_xnor2_1 _3599_ (.Y(_2740_),
    .A(\i_capsule.tf_y[0] ),
    .B(net936));
 sg13g2_a21oi_2 _3600_ (.B1(_2740_),
    .Y(_2741_),
    .A2(_2739_),
    .A1(_2718_));
 sg13g2_o21ai_1 _3601_ (.B1(_0031_),
    .Y(_2742_),
    .A1(\i_bitmap.in[7] ),
    .A2(_0032_));
 sg13g2_nor2_1 _3602_ (.A(_0032_),
    .B(net939),
    .Y(_2743_));
 sg13g2_a22oi_1 _3603_ (.Y(_2744_),
    .B1(_2742_),
    .B2(net936),
    .A2(_2741_),
    .A1(_2699_));
 sg13g2_xnor2_1 _3604_ (.Y(_2745_),
    .A(\i_bitmap.in[8] ),
    .B(net936));
 sg13g2_and2_1 _3605_ (.A(_2744_),
    .B(_2745_),
    .X(_2746_));
 sg13g2_a21oi_1 _3606_ (.A1(_2664_),
    .A2(_2667_),
    .Y(_2747_),
    .B1(_2669_));
 sg13g2_o21ai_1 _3607_ (.B1(_2655_),
    .Y(_2748_),
    .A1(_2662_),
    .A2(_2747_));
 sg13g2_a21oi_1 _3608_ (.A1(_2652_),
    .A2(_2748_),
    .Y(_2749_),
    .B1(_2659_));
 sg13g2_o21ai_1 _3609_ (.B1(_2677_),
    .Y(_2750_),
    .A1(_2674_),
    .A2(_2749_));
 sg13g2_a21oi_1 _3610_ (.A1(_2670_),
    .A2(_2750_),
    .Y(_2751_),
    .B1(net906));
 sg13g2_nor2_1 _3611_ (.A(\i_transform.track_y[0] ),
    .B(\i_transform.track_y[1] ),
    .Y(_2752_));
 sg13g2_nor3_1 _3612_ (.A(\i_transform.track_y[3] ),
    .B(\i_transform.track_y[2] ),
    .C(_2425_),
    .Y(_2753_));
 sg13g2_nand3_1 _3613_ (.B(_2752_),
    .C(_2753_),
    .A(_2426_),
    .Y(_2754_));
 sg13g2_nor3_1 _3614_ (.A(\i_transform.track_y[7] ),
    .B(\i_transform.track_y[6] ),
    .C(\i_transform.track_y[8] ),
    .Y(_2755_));
 sg13g2_nand4_1 _3615_ (.B(_2427_),
    .C(_2754_),
    .A(_0060_),
    .Y(_2756_),
    .D(_2755_));
 sg13g2_and2_1 _3616_ (.A(_2751_),
    .B(_2756_),
    .X(_2757_));
 sg13g2_nand2_1 _3617_ (.Y(_2758_),
    .A(_2751_),
    .B(_2756_));
 sg13g2_nor2_1 _3618_ (.A(_2744_),
    .B(_2745_),
    .Y(_2759_));
 sg13g2_o21ai_1 _3619_ (.B1(net886),
    .Y(_2760_),
    .A1(_2744_),
    .A2(_2745_));
 sg13g2_nor2_1 _3620_ (.A(_0032_),
    .B(_2725_),
    .Y(_2761_));
 sg13g2_nand2_1 _3621_ (.Y(_2762_),
    .A(\i_transform.image_y[5] ),
    .B(_2705_));
 sg13g2_xnor2_1 _3622_ (.Y(_2763_),
    .A(_0032_),
    .B(_2724_));
 sg13g2_nor2b_1 _3623_ (.A(_2762_),
    .B_N(_2763_),
    .Y(_2764_));
 sg13g2_xnor2_1 _3624_ (.Y(_2765_),
    .A(\i_bitmap.in[7] ),
    .B(_2729_));
 sg13g2_o21ai_1 _3625_ (.B1(_2765_),
    .Y(_2766_),
    .A1(_2761_),
    .A2(_2764_));
 sg13g2_or2_1 _3626_ (.X(_2767_),
    .B(_2729_),
    .A(_0031_));
 sg13g2_and2_1 _3627_ (.A(_2766_),
    .B(_2767_),
    .X(_2768_));
 sg13g2_xor2_1 _3628_ (.B(_2721_),
    .A(\i_bitmap.in[8] ),
    .X(_2769_));
 sg13g2_or2_1 _3629_ (.X(_2770_),
    .B(_2769_),
    .A(_2768_));
 sg13g2_a21oi_1 _3630_ (.A1(_2768_),
    .A2(_2769_),
    .Y(_2771_),
    .B1(net886));
 sg13g2_a21oi_1 _3631_ (.A1(_2770_),
    .A2(_2771_),
    .Y(_2772_),
    .B1(net905));
 sg13g2_o21ai_1 _3632_ (.B1(_2772_),
    .Y(_2773_),
    .A1(_2746_),
    .A2(_2760_));
 sg13g2_nor4_1 _3633_ (.A(_2618_),
    .B(_2643_),
    .C(_2646_),
    .D(net902),
    .Y(_2774_));
 sg13g2_nand3_1 _3634_ (.B(net894),
    .C(_2773_),
    .A(_2694_),
    .Y(_2775_));
 sg13g2_o21ai_1 _3635_ (.B1(_2775_),
    .Y(_2776_),
    .A1(_0034_),
    .A2(net894));
 sg13g2_and2_2 _3636_ (.A(net987),
    .B(_2776_),
    .X(_2777_));
 sg13g2_nand2_1 _3637_ (.Y(_2778_),
    .A(net987),
    .B(_2776_));
 sg13g2_xnor2_1 _3638_ (.Y(_2779_),
    .A(_0029_),
    .B(net974));
 sg13g2_a21oi_1 _3639_ (.A1(\i_bitmap.in[3] ),
    .A2(_0028_),
    .Y(_2780_),
    .B1(\i_bitmap.in[4] ));
 sg13g2_or2_1 _3640_ (.X(_2781_),
    .B(_2780_),
    .A(net973));
 sg13g2_and2_1 _3641_ (.A(_0026_),
    .B(net971),
    .X(_2782_));
 sg13g2_nor2_1 _3642_ (.A(_0026_),
    .B(net970),
    .Y(_2783_));
 sg13g2_a21o_1 _3643_ (.A2(_0018_),
    .A1(\i_capsule.tf_x[0] ),
    .B1(\i_bitmap.in[0] ),
    .X(_2784_));
 sg13g2_and2_1 _3644_ (.A(net967),
    .B(_2784_),
    .X(_2785_));
 sg13g2_xor2_1 _3645_ (.B(net899),
    .A(\i_transform.image_x[5] ),
    .X(_2786_));
 sg13g2_nor2b_1 _3646_ (.A(_0024_),
    .B_N(_2573_),
    .Y(_2787_));
 sg13g2_xnor2_1 _3647_ (.Y(_2788_),
    .A(_0024_),
    .B(_2573_));
 sg13g2_nand2b_1 _3648_ (.Y(_2789_),
    .B(net909),
    .A_N(_0025_));
 sg13g2_inv_1 _3649_ (.Y(_2790_),
    .A(_2789_));
 sg13g2_a21oi_2 _3650_ (.B1(_2787_),
    .Y(_2791_),
    .A2(_2790_),
    .A1(_2788_));
 sg13g2_xor2_1 _3651_ (.B(_2579_),
    .A(\i_transform.image_x[2] ),
    .X(_2792_));
 sg13g2_nor2_1 _3652_ (.A(_2791_),
    .B(_2792_),
    .Y(_2793_));
 sg13g2_or2_1 _3653_ (.X(_2794_),
    .B(_2579_),
    .A(_0023_));
 sg13g2_o21ai_1 _3654_ (.B1(_2794_),
    .Y(_2795_),
    .A1(_2791_),
    .A2(_2792_));
 sg13g2_xor2_1 _3655_ (.B(net898),
    .A(_0022_),
    .X(_2796_));
 sg13g2_nand2_1 _3656_ (.Y(_2797_),
    .A(_2795_),
    .B(_2796_));
 sg13g2_nor2_1 _3657_ (.A(_2389_),
    .B(net898),
    .Y(_2798_));
 sg13g2_a21oi_1 _3658_ (.A1(_2795_),
    .A2(_2796_),
    .Y(_2799_),
    .B1(_2798_));
 sg13g2_o21ai_1 _3659_ (.B1(_2797_),
    .Y(_2800_),
    .A1(_2389_),
    .A2(net898));
 sg13g2_xnor2_1 _3660_ (.Y(_2801_),
    .A(\i_transform.image_x[4] ),
    .B(_2585_));
 sg13g2_nand2_1 _3661_ (.Y(_2802_),
    .A(_2786_),
    .B(_2801_));
 sg13g2_nor2_1 _3662_ (.A(_0020_),
    .B(_2585_),
    .Y(_2803_));
 sg13g2_a22oi_1 _3663_ (.Y(_2804_),
    .B1(_2786_),
    .B2(_2803_),
    .A2(net899),
    .A1(_2438_));
 sg13g2_o21ai_1 _3664_ (.B1(_2804_),
    .Y(_2805_),
    .A1(_2799_),
    .A2(_2802_));
 sg13g2_xnor2_1 _3665_ (.Y(_2806_),
    .A(_0018_),
    .B(net970));
 sg13g2_xnor2_1 _3666_ (.Y(_2807_),
    .A(_0021_),
    .B(net970));
 sg13g2_inv_1 _3667_ (.Y(_2808_),
    .A(_2807_));
 sg13g2_nor2_1 _3668_ (.A(_2806_),
    .B(_2807_),
    .Y(_2809_));
 sg13g2_a21o_1 _3669_ (.A2(_2809_),
    .A1(_2805_),
    .B1(_2785_),
    .X(_2810_));
 sg13g2_xnor2_1 _3670_ (.Y(_2811_),
    .A(_0017_),
    .B(net966));
 sg13g2_a22oi_1 _3671_ (.Y(_2812_),
    .B1(_2810_),
    .B2(_2811_),
    .A2(net966),
    .A1(net1032));
 sg13g2_a221oi_1 _3672_ (.B2(_2811_),
    .C1(_2783_),
    .B1(_2810_),
    .A1(net1032),
    .Y(_2813_),
    .A2(net966));
 sg13g2_xnor2_1 _3673_ (.Y(_2814_),
    .A(_0027_),
    .B(net972));
 sg13g2_nor3_1 _3674_ (.A(_2782_),
    .B(_2813_),
    .C(_2814_),
    .Y(_2815_));
 sg13g2_xnor2_1 _3675_ (.Y(_2816_),
    .A(_0028_),
    .B(net972));
 sg13g2_or4_2 _3676_ (.A(_2782_),
    .B(_2813_),
    .C(_2814_),
    .D(_2816_),
    .X(_2817_));
 sg13g2_a21o_1 _3677_ (.A2(_2817_),
    .A1(_2781_),
    .B1(_2779_),
    .X(_2818_));
 sg13g2_o21ai_1 _3678_ (.B1(_2818_),
    .Y(_2819_),
    .A1(_0029_),
    .A2(net975));
 sg13g2_xnor2_1 _3679_ (.Y(_2820_),
    .A(_0030_),
    .B(net975));
 sg13g2_xor2_1 _3680_ (.B(_2820_),
    .A(_2819_),
    .X(_2821_));
 sg13g2_nor2_2 _3681_ (.A(net906),
    .B(net893),
    .Y(_2822_));
 sg13g2_xnor2_1 _3682_ (.Y(_2823_),
    .A(\i_bitmap.in[6] ),
    .B(net975));
 sg13g2_o21ai_1 _3683_ (.B1(_0029_),
    .Y(_2824_),
    .A1(\i_bitmap.in[5] ),
    .A2(_2402_));
 sg13g2_nand2_1 _3684_ (.Y(_2825_),
    .A(net974),
    .B(_2824_));
 sg13g2_xnor2_1 _3685_ (.Y(_2826_),
    .A(\i_bitmap.in[5] ),
    .B(net969));
 sg13g2_nor2_1 _3686_ (.A(_0027_),
    .B(_2566_),
    .Y(_2827_));
 sg13g2_xnor2_1 _3687_ (.Y(_2828_),
    .A(_0027_),
    .B(net899));
 sg13g2_and2_1 _3688_ (.A(net1032),
    .B(net898),
    .X(_2829_));
 sg13g2_nand2_1 _3689_ (.Y(_2830_),
    .A(_0019_),
    .B(net909));
 sg13g2_xnor2_1 _3690_ (.Y(_2831_),
    .A(_0021_),
    .B(_2573_));
 sg13g2_nor2b_1 _3691_ (.A(_2831_),
    .B_N(_2830_),
    .Y(_2832_));
 sg13g2_nor2b_1 _3692_ (.A(_2573_),
    .B_N(\i_capsule.tf_x[0] ),
    .Y(_2833_));
 sg13g2_xnor2_1 _3693_ (.Y(_2834_),
    .A(_0018_),
    .B(_2579_));
 sg13g2_o21ai_1 _3694_ (.B1(_2834_),
    .Y(_2835_),
    .A1(_2832_),
    .A2(_2833_));
 sg13g2_nand2_1 _3695_ (.Y(_2836_),
    .A(\i_bitmap.in[0] ),
    .B(_2579_));
 sg13g2_xnor2_1 _3696_ (.Y(_2837_),
    .A(net1032),
    .B(net898));
 sg13g2_a21oi_1 _3697_ (.A1(_2835_),
    .A2(_2836_),
    .Y(_2838_),
    .B1(_2837_));
 sg13g2_xnor2_1 _3698_ (.Y(_2839_),
    .A(_0026_),
    .B(_2585_));
 sg13g2_o21ai_1 _3699_ (.B1(_2839_),
    .Y(_2840_),
    .A1(_2829_),
    .A2(_2838_));
 sg13g2_nand2_1 _3700_ (.Y(_2841_),
    .A(\i_bitmap.in[2] ),
    .B(_2585_));
 sg13g2_a21oi_2 _3701_ (.B1(_2828_),
    .Y(_2842_),
    .A2(_2841_),
    .A1(_2840_));
 sg13g2_nand2_1 _3702_ (.Y(_2843_),
    .A(\i_bitmap.in[4] ),
    .B(net974));
 sg13g2_xnor2_1 _3703_ (.Y(_2844_),
    .A(_2402_),
    .B(net973));
 sg13g2_o21ai_1 _3704_ (.B1(_2844_),
    .Y(_2845_),
    .A1(_2827_),
    .A2(_2842_));
 sg13g2_nand2b_1 _3705_ (.Y(_2846_),
    .B(_2826_),
    .A_N(_2845_));
 sg13g2_nand3_1 _3706_ (.B(_2825_),
    .C(_2846_),
    .A(_2823_),
    .Y(_2847_));
 sg13g2_a21oi_2 _3707_ (.B1(_2823_),
    .Y(_2848_),
    .A2(_2846_),
    .A1(_2825_));
 sg13g2_nor2_1 _3708_ (.A(net906),
    .B(_2848_),
    .Y(_2849_));
 sg13g2_a21oi_1 _3709_ (.A1(_2847_),
    .A2(_2849_),
    .Y(_2850_),
    .B1(_2822_));
 sg13g2_a21oi_1 _3710_ (.A1(net889),
    .A2(_2821_),
    .Y(_0291_),
    .B1(_2850_));
 sg13g2_nor2_1 _3711_ (.A(_0029_),
    .B(net937),
    .Y(_0292_));
 sg13g2_nand2b_1 _3712_ (.Y(_0293_),
    .B(net940),
    .A_N(_2780_));
 sg13g2_xnor2_1 _3713_ (.Y(_0294_),
    .A(_0026_),
    .B(net935));
 sg13g2_nand2_1 _3714_ (.Y(_0295_),
    .A(net938),
    .B(_2784_));
 sg13g2_xnor2_1 _3715_ (.Y(_0296_),
    .A(_0018_),
    .B(net938));
 sg13g2_inv_1 _3716_ (.Y(_0297_),
    .A(_0296_));
 sg13g2_nand2b_1 _3717_ (.Y(_0298_),
    .B(_2724_),
    .A_N(_0024_));
 sg13g2_xor2_1 _3718_ (.B(_2724_),
    .A(_0024_),
    .X(_0299_));
 sg13g2_nand2b_1 _3719_ (.Y(_0300_),
    .B(_2705_),
    .A_N(_0025_));
 sg13g2_o21ai_1 _3720_ (.B1(_0298_),
    .Y(_0301_),
    .A1(_0299_),
    .A2(_0300_));
 sg13g2_xnor2_1 _3721_ (.Y(_0302_),
    .A(\i_transform.image_x[2] ),
    .B(_2729_));
 sg13g2_nor2_1 _3722_ (.A(_0023_),
    .B(_2729_),
    .Y(_0303_));
 sg13g2_a21oi_2 _3723_ (.B1(_0303_),
    .Y(_0304_),
    .A2(_0302_),
    .A1(_0301_));
 sg13g2_xnor2_1 _3724_ (.Y(_0305_),
    .A(_0022_),
    .B(_2721_));
 sg13g2_or2_1 _3725_ (.X(_0306_),
    .B(_2721_),
    .A(_2389_));
 sg13g2_o21ai_1 _3726_ (.B1(_0306_),
    .Y(_0307_),
    .A1(_0304_),
    .A2(_0305_));
 sg13g2_xnor2_1 _3727_ (.Y(_0308_),
    .A(\i_transform.image_x[4] ),
    .B(_2735_));
 sg13g2_and2_1 _3728_ (.A(_0307_),
    .B(_0308_),
    .X(_0309_));
 sg13g2_xor2_1 _3729_ (.B(_2717_),
    .A(\i_transform.image_x[5] ),
    .X(_0310_));
 sg13g2_and3_1 _3730_ (.X(_0311_),
    .A(_0307_),
    .B(_0308_),
    .C(_0310_));
 sg13g2_nand3_1 _3731_ (.B(_0308_),
    .C(_0310_),
    .A(_0307_),
    .Y(_0312_));
 sg13g2_nor2_1 _3732_ (.A(_0020_),
    .B(_2735_),
    .Y(_0313_));
 sg13g2_and2_1 _3733_ (.A(_2438_),
    .B(_2717_),
    .X(_0314_));
 sg13g2_a21oi_1 _3734_ (.A1(_0310_),
    .A2(_0313_),
    .Y(_0315_),
    .B1(_0314_));
 sg13g2_a21o_1 _3735_ (.A2(_0313_),
    .A1(_0310_),
    .B1(_0314_),
    .X(_0316_));
 sg13g2_xnor2_1 _3736_ (.Y(_0317_),
    .A(_0021_),
    .B(net938));
 sg13g2_inv_1 _3737_ (.Y(_0318_),
    .A(_0317_));
 sg13g2_a21oi_1 _3738_ (.A1(_0312_),
    .A2(_0315_),
    .Y(_0319_),
    .B1(_0318_));
 sg13g2_nor2_1 _3739_ (.A(_0297_),
    .B(_0318_),
    .Y(_0320_));
 sg13g2_o21ai_1 _3740_ (.B1(_0320_),
    .Y(_0321_),
    .A1(_0311_),
    .A2(_0316_));
 sg13g2_nand2b_1 _3741_ (.Y(_0322_),
    .B(net935),
    .A_N(_0017_));
 sg13g2_nand2_1 _3742_ (.Y(_0323_),
    .A(_0017_),
    .B(net938));
 sg13g2_nand2_1 _3743_ (.Y(_0324_),
    .A(_0322_),
    .B(_0323_));
 sg13g2_inv_1 _3744_ (.Y(_0325_),
    .A(_0324_));
 sg13g2_a21oi_1 _3745_ (.A1(_0295_),
    .A2(_0321_),
    .Y(_0326_),
    .B1(_0325_));
 sg13g2_a221oi_1 _3746_ (.B2(_0323_),
    .C1(_0294_),
    .B1(_0322_),
    .A1(_0295_),
    .Y(_0327_),
    .A2(_0321_));
 sg13g2_nor2_1 _3747_ (.A(_2403_),
    .B(net935),
    .Y(_0328_));
 sg13g2_a21oi_1 _3748_ (.A1(_2403_),
    .A2(_0026_),
    .Y(_0329_),
    .B1(net935));
 sg13g2_xnor2_1 _3749_ (.Y(_0330_),
    .A(_0027_),
    .B(net944));
 sg13g2_o21ai_1 _3750_ (.B1(_0330_),
    .Y(_0331_),
    .A1(_0327_),
    .A2(_0329_));
 sg13g2_xnor2_1 _3751_ (.Y(_0332_),
    .A(_0028_),
    .B(net940));
 sg13g2_inv_1 _3752_ (.Y(_0333_),
    .A(_0332_));
 sg13g2_o21ai_1 _3753_ (.B1(_0293_),
    .Y(_0334_),
    .A1(_0331_),
    .A2(_0333_));
 sg13g2_xnor2_1 _3754_ (.Y(_0335_),
    .A(_0029_),
    .B(net943));
 sg13g2_and2_1 _3755_ (.A(_0334_),
    .B(_0335_),
    .X(_0336_));
 sg13g2_a21oi_1 _3756_ (.A1(_0334_),
    .A2(_0335_),
    .Y(_0337_),
    .B1(_0292_));
 sg13g2_xnor2_1 _3757_ (.Y(_0338_),
    .A(_0030_),
    .B(net942));
 sg13g2_and2_1 _3758_ (.A(_0337_),
    .B(_0338_),
    .X(_0339_));
 sg13g2_o21ai_1 _3759_ (.B1(net876),
    .Y(_0340_),
    .A1(_0337_),
    .A2(_0338_));
 sg13g2_nor2_2 _3760_ (.A(_2645_),
    .B(net902),
    .Y(_0341_));
 sg13g2_nand2b_1 _3761_ (.Y(_0342_),
    .B(net906),
    .A_N(_2645_));
 sg13g2_nand2_2 _3762_ (.Y(_0343_),
    .A(net875),
    .B(_0341_));
 sg13g2_nand2_1 _3763_ (.Y(_0344_),
    .A(net937),
    .B(_2824_));
 sg13g2_nor2_1 _3764_ (.A(_0027_),
    .B(_2717_),
    .Y(_0345_));
 sg13g2_and2_1 _3765_ (.A(net1032),
    .B(_2721_),
    .X(_0346_));
 sg13g2_nand2_1 _3766_ (.Y(_0347_),
    .A(_0019_),
    .B(_2705_));
 sg13g2_xor2_1 _3767_ (.B(_2724_),
    .A(_0021_),
    .X(_0348_));
 sg13g2_a22oi_1 _3768_ (.Y(_0349_),
    .B1(_0347_),
    .B2(_0348_),
    .A2(_2725_),
    .A1(\i_capsule.tf_x[0] ));
 sg13g2_xor2_1 _3769_ (.B(_2729_),
    .A(_0018_),
    .X(_0350_));
 sg13g2_nand2_1 _3770_ (.Y(_0351_),
    .A(\i_bitmap.in[0] ),
    .B(_2729_));
 sg13g2_o21ai_1 _3771_ (.B1(_0351_),
    .Y(_0352_),
    .A1(_0349_),
    .A2(_0350_));
 sg13g2_xnor2_1 _3772_ (.Y(_0353_),
    .A(_2403_),
    .B(_2721_));
 sg13g2_a21oi_1 _3773_ (.A1(_0352_),
    .A2(_0353_),
    .Y(_0354_),
    .B1(_0346_));
 sg13g2_xor2_1 _3774_ (.B(_2735_),
    .A(_0026_),
    .X(_0355_));
 sg13g2_nand2_1 _3775_ (.Y(_0356_),
    .A(\i_bitmap.in[2] ),
    .B(_2735_));
 sg13g2_o21ai_1 _3776_ (.B1(_0356_),
    .Y(_0357_),
    .A1(_0354_),
    .A2(_0355_));
 sg13g2_xnor2_1 _3777_ (.Y(_0358_),
    .A(_0027_),
    .B(_2717_));
 sg13g2_nor2b_1 _3778_ (.A(_0358_),
    .B_N(_0357_),
    .Y(_0359_));
 sg13g2_nand2_1 _3779_ (.Y(_0360_),
    .A(\i_bitmap.in[4] ),
    .B(_2698_));
 sg13g2_xnor2_1 _3780_ (.Y(_0361_),
    .A(\i_bitmap.in[4] ),
    .B(net940));
 sg13g2_o21ai_1 _3781_ (.B1(_0361_),
    .Y(_0362_),
    .A1(_0345_),
    .A2(_0359_));
 sg13g2_xnor2_1 _3782_ (.Y(_0363_),
    .A(\i_bitmap.in[5] ),
    .B(net943));
 sg13g2_nand2b_1 _3783_ (.Y(_0364_),
    .B(_0363_),
    .A_N(_0362_));
 sg13g2_xnor2_1 _3784_ (.Y(_0365_),
    .A(_2401_),
    .B(net942));
 sg13g2_nand3_1 _3785_ (.B(_0364_),
    .C(_0365_),
    .A(_0344_),
    .Y(_0366_));
 sg13g2_a21o_1 _3786_ (.A2(_0364_),
    .A1(_0344_),
    .B1(_0365_),
    .X(_0367_));
 sg13g2_nand3_1 _3787_ (.B(_0366_),
    .C(_0367_),
    .A(_0341_),
    .Y(_0368_));
 sg13g2_nand2_1 _3788_ (.Y(_0369_),
    .A(_0343_),
    .B(_0368_));
 sg13g2_o21ai_1 _3789_ (.B1(_0369_),
    .Y(_0370_),
    .A1(_0339_),
    .A2(_0340_));
 sg13g2_nor2b_1 _3790_ (.A(_0291_),
    .B_N(_0370_),
    .Y(_0371_));
 sg13g2_nand2b_1 _3791_ (.Y(_0372_),
    .B(_2695_),
    .A_N(_0030_));
 sg13g2_nand3b_1 _3792_ (.B(_0370_),
    .C(_0372_),
    .Y(_0373_),
    .A_N(_0291_));
 sg13g2_and2_1 _3793_ (.A(net986),
    .B(net826),
    .X(_0374_));
 sg13g2_nand2_2 _3794_ (.Y(_0375_),
    .A(net986),
    .B(net826));
 sg13g2_and2_1 _3795_ (.A(\i_bitmap.in[3] ),
    .B(net968),
    .X(_0376_));
 sg13g2_o21ai_1 _3796_ (.B1(_2816_),
    .Y(_0377_),
    .A1(_2815_),
    .A2(_0376_));
 sg13g2_or3_1 _3797_ (.A(_2815_),
    .B(_2816_),
    .C(_0376_),
    .X(_0378_));
 sg13g2_nand3_1 _3798_ (.B(_0377_),
    .C(_0378_),
    .A(net887),
    .Y(_0379_));
 sg13g2_or3_1 _3799_ (.A(_2827_),
    .B(_2842_),
    .C(_2844_),
    .X(_0380_));
 sg13g2_nand3_1 _3800_ (.B(_2845_),
    .C(_0380_),
    .A(net902),
    .Y(_0381_));
 sg13g2_nand2b_1 _3801_ (.Y(_0382_),
    .B(_0381_),
    .A_N(_2822_));
 sg13g2_nand2_1 _3802_ (.Y(_0383_),
    .A(\i_bitmap.in[3] ),
    .B(net944));
 sg13g2_a21o_1 _3803_ (.A2(_0383_),
    .A1(_0331_),
    .B1(_0332_),
    .X(_0384_));
 sg13g2_nand3_1 _3804_ (.B(_0332_),
    .C(_0383_),
    .A(_0331_),
    .Y(_0385_));
 sg13g2_nand3_1 _3805_ (.B(_0384_),
    .C(_0385_),
    .A(net876),
    .Y(_0386_));
 sg13g2_or3_1 _3806_ (.A(_0345_),
    .B(_0359_),
    .C(_0361_),
    .X(_0387_));
 sg13g2_nand2_1 _3807_ (.Y(_0388_),
    .A(_0362_),
    .B(_0387_));
 sg13g2_a21oi_1 _3808_ (.A1(net880),
    .A2(_0388_),
    .Y(_0389_),
    .B1(net885));
 sg13g2_a22oi_1 _3809_ (.Y(_0390_),
    .B1(_0386_),
    .B2(_0389_),
    .A2(_0382_),
    .A1(_0379_));
 sg13g2_nor2_1 _3810_ (.A(_0028_),
    .B(net895),
    .Y(_0391_));
 sg13g2_a221oi_1 _3811_ (.B2(_0389_),
    .C1(_0391_),
    .B1(_0386_),
    .A1(_0379_),
    .Y(_0392_),
    .A2(_0382_));
 sg13g2_nand2b_2 _3812_ (.Y(_0393_),
    .B(_0390_),
    .A_N(_0391_));
 sg13g2_nor2_1 _3813_ (.A(net981),
    .B(_0392_),
    .Y(_0394_));
 sg13g2_nand2b_1 _3814_ (.Y(_0395_),
    .B(net988),
    .A_N(_0392_));
 sg13g2_and3_1 _3815_ (.X(_0396_),
    .A(_0295_),
    .B(_0321_),
    .C(_0325_));
 sg13g2_nor3_1 _3816_ (.A(net879),
    .B(_0326_),
    .C(_0396_),
    .Y(_0397_));
 sg13g2_xnor2_1 _3817_ (.Y(_0398_),
    .A(_0352_),
    .B(_0353_));
 sg13g2_o21ai_1 _3818_ (.B1(net905),
    .Y(_0399_),
    .A1(_2648_),
    .A2(_0398_));
 sg13g2_nor2_1 _3819_ (.A(_2695_),
    .B(net893),
    .Y(_0400_));
 sg13g2_nand2_2 _3820_ (.Y(_0401_),
    .A(net894),
    .B(net888));
 sg13g2_xnor2_1 _3821_ (.Y(_0402_),
    .A(_2810_),
    .B(_2811_));
 sg13g2_nand3_1 _3822_ (.B(_2836_),
    .C(_2837_),
    .A(_2835_),
    .Y(_0403_));
 sg13g2_nor2_1 _3823_ (.A(net886),
    .B(_2838_),
    .Y(_0404_));
 sg13g2_a21oi_1 _3824_ (.A1(_0403_),
    .A2(_0404_),
    .Y(_0405_),
    .B1(_0341_));
 sg13g2_o21ai_1 _3825_ (.B1(_0405_),
    .Y(_0406_),
    .A1(_0401_),
    .A2(_0402_));
 sg13g2_o21ai_1 _3826_ (.B1(_0406_),
    .Y(_0407_),
    .A1(_0397_),
    .A2(_0399_));
 sg13g2_nand2b_2 _3827_ (.Y(_0408_),
    .B(net897),
    .A_N(_0017_));
 sg13g2_nand2_2 _3828_ (.Y(_0409_),
    .A(_0407_),
    .B(_0408_));
 sg13g2_a21oi_2 _3829_ (.B1(net981),
    .Y(_0410_),
    .A2(_0408_),
    .A1(_0407_));
 sg13g2_a21o_2 _3830_ (.A2(_0408_),
    .A1(_0407_),
    .B1(net981),
    .X(_0411_));
 sg13g2_and2_1 _3831_ (.A(\i_capsule.tf_x[0] ),
    .B(net938),
    .X(_0412_));
 sg13g2_o21ai_1 _3832_ (.B1(_0297_),
    .Y(_0413_),
    .A1(_0319_),
    .A2(_0412_));
 sg13g2_or3_1 _3833_ (.A(_0297_),
    .B(_0319_),
    .C(_0412_),
    .X(_0414_));
 sg13g2_nand3_1 _3834_ (.B(_0413_),
    .C(_0414_),
    .A(net874),
    .Y(_0415_));
 sg13g2_xnor2_1 _3835_ (.Y(_0416_),
    .A(_0349_),
    .B(_0350_));
 sg13g2_a21oi_1 _3836_ (.A1(net878),
    .A2(_0416_),
    .Y(_0417_),
    .B1(net884));
 sg13g2_a22oi_1 _3837_ (.Y(_0418_),
    .B1(_2805_),
    .B2(_2808_),
    .A2(net966),
    .A1(\i_capsule.tf_x[0] ));
 sg13g2_xnor2_1 _3838_ (.Y(_0419_),
    .A(_2806_),
    .B(_0418_));
 sg13g2_or3_1 _3839_ (.A(_2832_),
    .B(_2833_),
    .C(_2834_),
    .X(_0420_));
 sg13g2_a21oi_1 _3840_ (.A1(_2835_),
    .A2(_0420_),
    .Y(_0421_),
    .B1(net886));
 sg13g2_a21oi_1 _3841_ (.A1(net886),
    .A2(_0419_),
    .Y(_0422_),
    .B1(_0421_));
 sg13g2_a22oi_1 _3842_ (.Y(_0423_),
    .B1(_0422_),
    .B2(net901),
    .A2(_0417_),
    .A1(_0415_));
 sg13g2_nor2_1 _3843_ (.A(_0018_),
    .B(net894),
    .Y(_0424_));
 sg13g2_nand2b_1 _3844_ (.Y(_0425_),
    .B(_2695_),
    .A_N(_0018_));
 sg13g2_a221oi_1 _3845_ (.B2(net901),
    .C1(_0424_),
    .B1(_0422_),
    .A1(_0415_),
    .Y(_0426_),
    .A2(_0417_));
 sg13g2_nand2_2 _3846_ (.Y(_0427_),
    .A(_0423_),
    .B(_0425_));
 sg13g2_nor2_2 _3847_ (.A(net981),
    .B(_0426_),
    .Y(_0428_));
 sg13g2_nand2b_2 _3848_ (.Y(_0429_),
    .B(net985),
    .A_N(_0426_));
 sg13g2_nor2_2 _3849_ (.A(_0410_),
    .B(_0428_),
    .Y(_0430_));
 sg13g2_nand2_2 _3850_ (.Y(_0431_),
    .A(net867),
    .B(_0429_));
 sg13g2_xnor2_1 _3851_ (.Y(_0432_),
    .A(_0354_),
    .B(_0355_));
 sg13g2_nand2_1 _3852_ (.Y(_0433_),
    .A(net879),
    .B(_0432_));
 sg13g2_or3_1 _3853_ (.A(_0294_),
    .B(_0326_),
    .C(_0328_),
    .X(_0434_));
 sg13g2_o21ai_1 _3854_ (.B1(_0294_),
    .Y(_0435_),
    .A1(_0326_),
    .A2(_0328_));
 sg13g2_nand3_1 _3855_ (.B(_0434_),
    .C(_0435_),
    .A(net874),
    .Y(_0436_));
 sg13g2_a21oi_2 _3856_ (.B1(net884),
    .Y(_0437_),
    .A2(_0436_),
    .A1(_0433_));
 sg13g2_a21o_1 _3857_ (.A2(_0436_),
    .A1(_0433_),
    .B1(net884),
    .X(_0438_));
 sg13g2_nor2_1 _3858_ (.A(_2782_),
    .B(_2783_),
    .Y(_0439_));
 sg13g2_or3_1 _3859_ (.A(_2829_),
    .B(_2838_),
    .C(_2839_),
    .X(_0440_));
 sg13g2_nor2_2 _3860_ (.A(net977),
    .B(net901),
    .Y(_0441_));
 sg13g2_a21o_1 _3861_ (.A2(_0440_),
    .A1(_2840_),
    .B1(net887),
    .X(_0442_));
 sg13g2_xor2_1 _3862_ (.B(_0439_),
    .A(_2812_),
    .X(_0443_));
 sg13g2_a21oi_1 _3863_ (.A1(net887),
    .A2(_0443_),
    .Y(_0444_),
    .B1(net976));
 sg13g2_a21o_1 _3864_ (.A2(_0444_),
    .A1(_0442_),
    .B1(_0441_),
    .X(_0445_));
 sg13g2_a21oi_2 _3865_ (.B1(_0441_),
    .Y(_0446_),
    .A2(_0444_),
    .A1(_0442_));
 sg13g2_and2_1 _3866_ (.A(_0026_),
    .B(net896),
    .X(_0447_));
 sg13g2_nand2_1 _3867_ (.Y(_0448_),
    .A(_0026_),
    .B(net896));
 sg13g2_nor3_1 _3868_ (.A(_0437_),
    .B(_0446_),
    .C(_0447_),
    .Y(_0449_));
 sg13g2_nand3_1 _3869_ (.B(_0445_),
    .C(_0448_),
    .A(_0438_),
    .Y(_0450_));
 sg13g2_a221oi_1 _3870_ (.B2(_0425_),
    .C1(net981),
    .B1(_0423_),
    .A1(_0407_),
    .Y(_0451_),
    .A2(_0408_));
 sg13g2_nand2_2 _3871_ (.Y(_0452_),
    .A(_0409_),
    .B(_0428_));
 sg13g2_nand2_2 _3872_ (.Y(_0453_),
    .A(net863),
    .B(_0452_));
 sg13g2_nand2_2 _3873_ (.Y(_0454_),
    .A(_0431_),
    .B(net861));
 sg13g2_a21o_2 _3874_ (.A2(_0429_),
    .A1(net867),
    .B1(_0451_),
    .X(_0455_));
 sg13g2_nand2b_2 _3875_ (.Y(_0456_),
    .B(net861),
    .A_N(_0455_));
 sg13g2_o21ai_1 _3876_ (.B1(_2814_),
    .Y(_0457_),
    .A1(_2782_),
    .A2(_2813_));
 sg13g2_nand3b_1 _3877_ (.B(_0400_),
    .C(_0457_),
    .Y(_0458_),
    .A_N(_2815_));
 sg13g2_nand3_1 _3878_ (.B(_2840_),
    .C(_2841_),
    .A(_2828_),
    .Y(_0459_));
 sg13g2_nor2_1 _3879_ (.A(net887),
    .B(_2842_),
    .Y(_0460_));
 sg13g2_a21oi_1 _3880_ (.A1(_0459_),
    .A2(_0460_),
    .Y(_0461_),
    .B1(_0341_));
 sg13g2_or3_1 _3881_ (.A(_0327_),
    .B(_0329_),
    .C(_0330_),
    .X(_0462_));
 sg13g2_nand3_1 _3882_ (.B(_0331_),
    .C(_0462_),
    .A(net874),
    .Y(_0463_));
 sg13g2_nor2b_1 _3883_ (.A(_0357_),
    .B_N(_0358_),
    .Y(_0464_));
 sg13g2_nor3_1 _3884_ (.A(net874),
    .B(_0359_),
    .C(_0464_),
    .Y(_0465_));
 sg13g2_nor2_1 _3885_ (.A(net902),
    .B(_0465_),
    .Y(_0466_));
 sg13g2_a22oi_1 _3886_ (.Y(_0467_),
    .B1(_0463_),
    .B2(_0466_),
    .A2(_0461_),
    .A1(_0458_));
 sg13g2_nor2b_2 _3887_ (.A(_0027_),
    .B_N(net897),
    .Y(_0468_));
 sg13g2_or2_1 _3888_ (.X(_0469_),
    .B(_0468_),
    .A(_0467_));
 sg13g2_inv_1 _3889_ (.Y(_0470_),
    .A(net859));
 sg13g2_and2_1 _3890_ (.A(net985),
    .B(net859),
    .X(_0471_));
 sg13g2_o21ai_1 _3891_ (.B1(net990),
    .Y(_0472_),
    .A1(_0467_),
    .A2(_0468_));
 sg13g2_nand2b_2 _3892_ (.Y(_0473_),
    .B(_0455_),
    .A_N(net855));
 sg13g2_nand2_1 _3893_ (.Y(_0474_),
    .A(_0456_),
    .B(_0473_));
 sg13g2_a22oi_1 _3894_ (.Y(_0475_),
    .B1(net844),
    .B2(_0474_),
    .A2(net826),
    .A1(net986));
 sg13g2_nor4_2 _3895_ (.A(_0409_),
    .B(_0437_),
    .C(_0446_),
    .Y(_0476_),
    .D(_0447_));
 sg13g2_nand2b_2 _3896_ (.Y(_0477_),
    .B(net865),
    .A_N(_0409_));
 sg13g2_nand2_2 _3897_ (.Y(_0478_),
    .A(_0427_),
    .B(_0476_));
 sg13g2_nor2_2 _3898_ (.A(_0411_),
    .B(_0427_),
    .Y(_0479_));
 sg13g2_nand2_2 _3899_ (.Y(_0480_),
    .A(_0410_),
    .B(_0426_));
 sg13g2_and2_1 _3900_ (.A(net853),
    .B(_0480_),
    .X(_0481_));
 sg13g2_nand2_1 _3901_ (.Y(_0482_),
    .A(_0478_),
    .B(_0481_));
 sg13g2_and4_1 _3902_ (.A(_0438_),
    .B(_0445_),
    .C(_0448_),
    .D(_0451_),
    .X(_0483_));
 sg13g2_nor2_2 _3903_ (.A(net851),
    .B(net848),
    .Y(_0484_));
 sg13g2_nor2_2 _3904_ (.A(_0409_),
    .B(_0429_),
    .Y(_0485_));
 sg13g2_nand2b_1 _3905_ (.Y(_0486_),
    .B(_0428_),
    .A_N(_0409_));
 sg13g2_nand2_2 _3906_ (.Y(_0487_),
    .A(net861),
    .B(_0485_));
 sg13g2_a22oi_1 _3907_ (.Y(_0488_),
    .B1(_0484_),
    .B2(_0487_),
    .A2(_0481_),
    .A1(_0478_));
 sg13g2_or2_1 _3908_ (.X(_0489_),
    .B(_0488_),
    .A(net845));
 sg13g2_or3_1 _3909_ (.A(_2699_),
    .B(_2741_),
    .C(_2743_),
    .X(_0490_));
 sg13g2_o21ai_1 _3910_ (.B1(_2699_),
    .Y(_0491_),
    .A1(_2741_),
    .A2(_2743_));
 sg13g2_a21oi_1 _3911_ (.A1(_0490_),
    .A2(_0491_),
    .Y(_0492_),
    .B1(net891));
 sg13g2_or3_1 _3912_ (.A(_2761_),
    .B(_2764_),
    .C(_2765_),
    .X(_0493_));
 sg13g2_and2_1 _3913_ (.A(_2766_),
    .B(_0493_),
    .X(_0494_));
 sg13g2_o21ai_1 _3914_ (.B1(net901),
    .Y(_0495_),
    .A1(net886),
    .A2(_0494_));
 sg13g2_nor2_1 _3915_ (.A(_0492_),
    .B(_0495_),
    .Y(_0496_));
 sg13g2_a21oi_1 _3916_ (.A1(\i_capsule.tf_y[0] ),
    .A2(net966),
    .Y(_0497_),
    .B1(_2592_));
 sg13g2_nand2b_1 _3917_ (.Y(_0498_),
    .B(_2479_),
    .A_N(_0497_));
 sg13g2_a21oi_1 _3918_ (.A1(_2480_),
    .A2(_0497_),
    .Y(_0499_),
    .B1(net878));
 sg13g2_xor2_1 _3919_ (.B(_2686_),
    .A(_2685_),
    .X(_0500_));
 sg13g2_a221oi_1 _3920_ (.B2(net878),
    .C1(net884),
    .B1(_0500_),
    .A1(_0498_),
    .Y(_0501_),
    .A2(_0499_));
 sg13g2_nor2_1 _3921_ (.A(_0031_),
    .B(net894),
    .Y(_0502_));
 sg13g2_or3_2 _3922_ (.A(_0496_),
    .B(_0501_),
    .C(_0502_),
    .X(_0503_));
 sg13g2_and2_1 _3923_ (.A(net985),
    .B(_0503_),
    .X(_0504_));
 sg13g2_nand2_2 _3924_ (.Y(_0505_),
    .A(net988),
    .B(_0503_));
 sg13g2_and3_2 _3925_ (.X(_0506_),
    .A(net860),
    .B(_0452_),
    .C(net849));
 sg13g2_nand3_1 _3926_ (.B(_0452_),
    .C(net852),
    .A(net863),
    .Y(_0507_));
 sg13g2_nand2_1 _3927_ (.Y(_0508_),
    .A(net847),
    .B(_0506_));
 sg13g2_a221oi_1 _3928_ (.B2(net826),
    .C1(_0505_),
    .B1(_0508_),
    .A1(_0475_),
    .Y(_0509_),
    .A2(_0489_));
 sg13g2_xor2_1 _3929_ (.B(_0335_),
    .A(_0334_),
    .X(_0510_));
 sg13g2_a21oi_1 _3930_ (.A1(_0360_),
    .A2(_0362_),
    .Y(_0511_),
    .B1(_0363_));
 sg13g2_nand3_1 _3931_ (.B(_0362_),
    .C(_0363_),
    .A(_0360_),
    .Y(_0512_));
 sg13g2_nor2_1 _3932_ (.A(net875),
    .B(_0511_),
    .Y(_0513_));
 sg13g2_a21oi_1 _3933_ (.A1(_0512_),
    .A2(_0513_),
    .Y(_0514_),
    .B1(net885));
 sg13g2_o21ai_1 _3934_ (.B1(_0514_),
    .Y(_0515_),
    .A1(net881),
    .A2(_0510_));
 sg13g2_nand3_1 _3935_ (.B(_2781_),
    .C(_2817_),
    .A(_2779_),
    .Y(_0516_));
 sg13g2_a21oi_1 _3936_ (.A1(_2818_),
    .A2(_0516_),
    .Y(_0517_),
    .B1(net893));
 sg13g2_a21oi_1 _3937_ (.A1(_2843_),
    .A2(_2845_),
    .Y(_0518_),
    .B1(_2826_));
 sg13g2_and3_1 _3938_ (.X(_0519_),
    .A(_2826_),
    .B(_2843_),
    .C(_2845_));
 sg13g2_nor3_1 _3939_ (.A(net889),
    .B(_0518_),
    .C(_0519_),
    .Y(_0520_));
 sg13g2_or3_1 _3940_ (.A(net906),
    .B(_0517_),
    .C(_0520_),
    .X(_0521_));
 sg13g2_nand2_1 _3941_ (.Y(_0522_),
    .A(_0515_),
    .B(_0521_));
 sg13g2_nand2_1 _3942_ (.Y(_0523_),
    .A(_2439_),
    .B(_2695_));
 sg13g2_nand3_1 _3943_ (.B(_0521_),
    .C(_0523_),
    .A(_0515_),
    .Y(_0524_));
 sg13g2_and2_1 _3944_ (.A(net987),
    .B(net829),
    .X(_0525_));
 sg13g2_nand2_1 _3945_ (.Y(_0526_),
    .A(net987),
    .B(net829));
 sg13g2_nand2_1 _3946_ (.Y(_0527_),
    .A(_0456_),
    .B(_0471_));
 sg13g2_a21o_1 _3947_ (.A2(_0527_),
    .A1(_0482_),
    .B1(net843),
    .X(_0528_));
 sg13g2_nand2_2 _3948_ (.Y(_0529_),
    .A(net865),
    .B(net859));
 sg13g2_nand2_1 _3949_ (.Y(_0530_),
    .A(net847),
    .B(_0529_));
 sg13g2_nor2_2 _3950_ (.A(net842),
    .B(net833),
    .Y(_0531_));
 sg13g2_a221oi_1 _3951_ (.B2(net817),
    .C1(net833),
    .B1(_0530_),
    .A1(_0475_),
    .Y(_0532_),
    .A2(_0528_));
 sg13g2_nor2_1 _3952_ (.A(_0509_),
    .B(_0532_),
    .Y(_0533_));
 sg13g2_and2_1 _3953_ (.A(_0410_),
    .B(net859),
    .X(_0534_));
 sg13g2_o21ai_1 _3954_ (.B1(_0410_),
    .Y(_0535_),
    .A1(_0467_),
    .A2(_0468_));
 sg13g2_nor2_2 _3955_ (.A(net867),
    .B(net866),
    .Y(_0536_));
 sg13g2_nand2_1 _3956_ (.Y(_0537_),
    .A(_0410_),
    .B(net864));
 sg13g2_o21ai_1 _3957_ (.B1(_0531_),
    .Y(_0538_),
    .A1(net828),
    .A2(_0536_));
 sg13g2_nor2_2 _3958_ (.A(net847),
    .B(net831),
    .Y(_0539_));
 sg13g2_nor2_1 _3959_ (.A(_0410_),
    .B(net850),
    .Y(_0540_));
 sg13g2_nand2_1 _3960_ (.Y(_0541_),
    .A(net867),
    .B(net836));
 sg13g2_and2_1 _3961_ (.A(_0454_),
    .B(net854),
    .X(_0542_));
 sg13g2_nand2_1 _3962_ (.Y(_0543_),
    .A(net861),
    .B(net854));
 sg13g2_nand3_1 _3963_ (.B(net861),
    .C(net853),
    .A(_0431_),
    .Y(_0544_));
 sg13g2_nand2_1 _3964_ (.Y(_0545_),
    .A(_0535_),
    .B(_0544_));
 sg13g2_nand3_1 _3965_ (.B(net853),
    .C(_0477_),
    .A(_0454_),
    .Y(_0546_));
 sg13g2_nor2_1 _3966_ (.A(net839),
    .B(net828),
    .Y(_0547_));
 sg13g2_a22oi_1 _3967_ (.Y(_0548_),
    .B1(_0546_),
    .B2(_0547_),
    .A2(_0545_),
    .A1(_0539_));
 sg13g2_nand2_1 _3968_ (.Y(_0549_),
    .A(_0538_),
    .B(_0548_));
 sg13g2_a21oi_2 _3969_ (.B1(net851),
    .Y(_0550_),
    .A2(_0452_),
    .A1(net860));
 sg13g2_nand2_2 _3970_ (.Y(_0551_),
    .A(net862),
    .B(_0479_));
 sg13g2_a21oi_2 _3971_ (.B1(_0485_),
    .Y(_0552_),
    .A2(_0479_),
    .A1(net862));
 sg13g2_nor2_2 _3972_ (.A(net835),
    .B(_0552_),
    .Y(_0553_));
 sg13g2_or4_1 _3973_ (.A(_0373_),
    .B(net844),
    .C(_0550_),
    .D(_0553_),
    .X(_0554_));
 sg13g2_a21oi_1 _3974_ (.A1(_0373_),
    .A2(_0549_),
    .Y(_0555_),
    .B1(net822));
 sg13g2_a22oi_1 _3975_ (.Y(_0556_),
    .B1(_0554_),
    .B2(_0555_),
    .A2(_0533_),
    .A1(net822));
 sg13g2_nand2_1 _3976_ (.Y(_0557_),
    .A(\i_bitmap.in[8] ),
    .B(net966));
 sg13g2_o21ai_1 _3977_ (.B1(_0557_),
    .Y(_0558_),
    .A1(_2594_),
    .A2(_2596_));
 sg13g2_nor2_1 _3978_ (.A(_0035_),
    .B(net970),
    .Y(_0559_));
 sg13g2_nand2_1 _3979_ (.Y(_0560_),
    .A(_0035_),
    .B(net970));
 sg13g2_nand2b_1 _3980_ (.Y(_0561_),
    .B(_0560_),
    .A_N(_0559_));
 sg13g2_a21oi_1 _3981_ (.A1(_0558_),
    .A2(_0561_),
    .Y(_0562_),
    .B1(net879));
 sg13g2_o21ai_1 _3982_ (.B1(_0562_),
    .Y(_0563_),
    .A1(_0558_),
    .A2(_0561_));
 sg13g2_a21o_1 _3983_ (.A2(net898),
    .A1(\i_bitmap.in[8] ),
    .B1(_2691_),
    .X(_0564_));
 sg13g2_xnor2_1 _3984_ (.Y(_0565_),
    .A(_0035_),
    .B(_2585_));
 sg13g2_xnor2_1 _3985_ (.Y(_0566_),
    .A(_0564_),
    .B(_0565_));
 sg13g2_a21oi_1 _3986_ (.A1(net879),
    .A2(_0566_),
    .Y(_0567_),
    .B1(net885));
 sg13g2_a21oi_1 _3987_ (.A1(_2440_),
    .A2(net935),
    .Y(_0568_),
    .B1(_2759_));
 sg13g2_nand2_1 _3988_ (.Y(_0569_),
    .A(\i_bitmap.in[9] ),
    .B(net936));
 sg13g2_nor2_1 _3989_ (.A(\i_bitmap.in[9] ),
    .B(net936),
    .Y(_0570_));
 sg13g2_xnor2_1 _3990_ (.Y(_0571_),
    .A(\i_bitmap.in[9] ),
    .B(net938));
 sg13g2_or2_1 _3991_ (.X(_0572_),
    .B(_0571_),
    .A(_0568_));
 sg13g2_a21oi_1 _3992_ (.A1(_0568_),
    .A2(_0571_),
    .Y(_0573_),
    .B1(net892));
 sg13g2_o21ai_1 _3993_ (.B1(_2770_),
    .Y(_0574_),
    .A1(_0034_),
    .A2(_2721_));
 sg13g2_xor2_1 _3994_ (.B(_2735_),
    .A(\i_bitmap.in[9] ),
    .X(_0575_));
 sg13g2_inv_1 _3995_ (.Y(_0576_),
    .A(_0575_));
 sg13g2_xnor2_1 _3996_ (.Y(_0577_),
    .A(_0574_),
    .B(_0576_));
 sg13g2_a22oi_1 _3997_ (.Y(_0578_),
    .B1(_0577_),
    .B2(net892),
    .A2(_0573_),
    .A1(_0572_));
 sg13g2_a22oi_1 _3998_ (.Y(_0579_),
    .B1(_0578_),
    .B2(net901),
    .A2(_0567_),
    .A1(_0563_));
 sg13g2_o21ai_1 _3999_ (.B1(_0579_),
    .Y(_0580_),
    .A1(_0035_),
    .A2(net894));
 sg13g2_inv_1 _4000_ (.Y(_0581_),
    .A(_0580_));
 sg13g2_nand2_1 _4001_ (.Y(_0582_),
    .A(net987),
    .B(_0580_));
 sg13g2_inv_1 _4002_ (.Y(_0583_),
    .A(_0582_));
 sg13g2_nor2_2 _4003_ (.A(_0430_),
    .B(net864),
    .Y(_0584_));
 sg13g2_and3_2 _4004_ (.X(_0585_),
    .A(_0431_),
    .B(net866),
    .C(net849));
 sg13g2_nand3_1 _4005_ (.B(net866),
    .C(net851),
    .A(_0431_),
    .Y(_0586_));
 sg13g2_nand2_2 _4006_ (.Y(_0587_),
    .A(net867),
    .B(net860));
 sg13g2_and2_2 _4007_ (.A(net867),
    .B(net856),
    .X(_0588_));
 sg13g2_and3_2 _4008_ (.X(_0589_),
    .A(net867),
    .B(net860),
    .C(net849));
 sg13g2_nand2_2 _4009_ (.Y(_0590_),
    .A(net863),
    .B(_0588_));
 sg13g2_nor4_1 _4010_ (.A(net830),
    .B(_0540_),
    .C(_0585_),
    .D(_0589_),
    .Y(_0591_));
 sg13g2_nor4_1 _4011_ (.A(net832),
    .B(_0506_),
    .C(_0540_),
    .D(_0585_),
    .Y(_0592_));
 sg13g2_o21ai_1 _4012_ (.B1(net837),
    .Y(_0593_),
    .A1(_0591_),
    .A2(_0592_));
 sg13g2_o21ai_1 _4013_ (.B1(net849),
    .Y(_0594_),
    .A1(net866),
    .A2(_0451_));
 sg13g2_a21oi_1 _4014_ (.A1(_0456_),
    .A2(net857),
    .Y(_0595_),
    .B1(net828));
 sg13g2_nand2_1 _4015_ (.Y(_0596_),
    .A(net847),
    .B(_0595_));
 sg13g2_nand3_1 _4016_ (.B(_0593_),
    .C(_0596_),
    .A(net817),
    .Y(_0597_));
 sg13g2_nand3_1 _4017_ (.B(net856),
    .C(_0552_),
    .A(net840),
    .Y(_0598_));
 sg13g2_nand2_1 _4018_ (.Y(_0599_),
    .A(net814),
    .B(_0598_));
 sg13g2_a21oi_1 _4019_ (.A1(net814),
    .A2(_0598_),
    .Y(_0600_),
    .B1(net822));
 sg13g2_nand4_1 _4020_ (.B(_0438_),
    .C(_0445_),
    .A(_0409_),
    .Y(_0601_),
    .D(_0448_));
 sg13g2_nor2_2 _4021_ (.A(net860),
    .B(_0535_),
    .Y(_0602_));
 sg13g2_nand2_1 _4022_ (.Y(_0603_),
    .A(net865),
    .B(_0534_));
 sg13g2_nand2_2 _4023_ (.Y(_0604_),
    .A(net859),
    .B(net848));
 sg13g2_nor2_2 _4024_ (.A(net845),
    .B(_0604_),
    .Y(_0605_));
 sg13g2_nand3b_1 _4025_ (.B(net817),
    .C(_0530_),
    .Y(_0606_),
    .A_N(_0605_));
 sg13g2_nand2_1 _4026_ (.Y(_0607_),
    .A(_0455_),
    .B(net850));
 sg13g2_a21oi_2 _4027_ (.B1(net857),
    .Y(_0608_),
    .A2(net861),
    .A1(_0411_));
 sg13g2_a21o_2 _4028_ (.A2(net860),
    .A1(net867),
    .B1(net849),
    .X(_0609_));
 sg13g2_nor2_2 _4029_ (.A(net848),
    .B(_0609_),
    .Y(_0610_));
 sg13g2_o21ai_1 _4030_ (.B1(_0607_),
    .Y(_0611_),
    .A1(net848),
    .A2(_0609_));
 sg13g2_nor2_1 _4031_ (.A(net853),
    .B(_0476_),
    .Y(_0612_));
 sg13g2_a22oi_1 _4032_ (.Y(_0613_),
    .B1(_0612_),
    .B2(_0454_),
    .A2(_0481_),
    .A1(_0478_));
 sg13g2_mux2_1 _4033_ (.A0(_0611_),
    .A1(_0613_),
    .S(net838),
    .X(_0614_));
 sg13g2_a21oi_1 _4034_ (.A1(net814),
    .A2(_0614_),
    .Y(_0615_),
    .B1(net825));
 sg13g2_a22oi_1 _4035_ (.Y(_0616_),
    .B1(_0606_),
    .B2(_0615_),
    .A2(_0600_),
    .A1(_0597_));
 sg13g2_a21oi_1 _4036_ (.A1(net827),
    .A2(_0616_),
    .Y(_0617_),
    .B1(_0582_));
 sg13g2_o21ai_1 _4037_ (.B1(_0617_),
    .Y(_0618_),
    .A1(_2778_),
    .A2(_0556_));
 sg13g2_o21ai_1 _4038_ (.B1(_0569_),
    .Y(_0619_),
    .A1(_0568_),
    .A2(_0570_));
 sg13g2_xnor2_1 _4039_ (.Y(_0620_),
    .A(\i_bitmap.in[10] ),
    .B(net935));
 sg13g2_inv_1 _4040_ (.Y(_0621_),
    .A(_0620_));
 sg13g2_xnor2_1 _4041_ (.Y(_0622_),
    .A(_0619_),
    .B(_0621_));
 sg13g2_nor2_1 _4042_ (.A(_0035_),
    .B(_2735_),
    .Y(_0623_));
 sg13g2_a21oi_2 _4043_ (.B1(_0623_),
    .Y(_0624_),
    .A2(_0576_),
    .A1(_0574_));
 sg13g2_nand2_1 _4044_ (.Y(_0625_),
    .A(\i_bitmap.in[10] ),
    .B(_2717_));
 sg13g2_or2_1 _4045_ (.X(_0626_),
    .B(_2717_),
    .A(\i_bitmap.in[10] ));
 sg13g2_and2_1 _4046_ (.A(_0625_),
    .B(_0626_),
    .X(_0627_));
 sg13g2_o21ai_1 _4047_ (.B1(net892),
    .Y(_0628_),
    .A1(_0624_),
    .A2(_0627_));
 sg13g2_a21oi_1 _4048_ (.A1(_0624_),
    .A2(_0627_),
    .Y(_0629_),
    .B1(_0628_));
 sg13g2_a21oi_1 _4049_ (.A1(net888),
    .A2(_0622_),
    .Y(_0630_),
    .B1(_0629_));
 sg13g2_a21oi_2 _4050_ (.B1(_0559_),
    .Y(_0631_),
    .A2(_0560_),
    .A1(_0558_));
 sg13g2_xnor2_1 _4051_ (.Y(_0632_),
    .A(_0036_),
    .B(net970));
 sg13g2_xnor2_1 _4052_ (.Y(_0633_),
    .A(_0631_),
    .B(_0632_));
 sg13g2_a22oi_1 _4053_ (.Y(_0634_),
    .B1(_0564_),
    .B2(_0565_),
    .A2(_2585_),
    .A1(\i_bitmap.in[9] ));
 sg13g2_nor2_1 _4054_ (.A(_0036_),
    .B(net899),
    .Y(_0635_));
 sg13g2_xnor2_1 _4055_ (.Y(_0636_),
    .A(_2441_),
    .B(net899));
 sg13g2_xnor2_1 _4056_ (.Y(_0637_),
    .A(_0634_),
    .B(_0636_));
 sg13g2_nor2_1 _4057_ (.A(net874),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_a21oi_1 _4058_ (.A1(net874),
    .A2(_0633_),
    .Y(_0639_),
    .B1(_0638_));
 sg13g2_a22oi_1 _4059_ (.Y(_0640_),
    .B1(_0639_),
    .B2(_0341_),
    .A2(_0630_),
    .A1(net902));
 sg13g2_o21ai_1 _4060_ (.B1(_0640_),
    .Y(_0641_),
    .A1(_0036_),
    .A2(net894));
 sg13g2_and2_1 _4061_ (.A(net985),
    .B(_0641_),
    .X(_0642_));
 sg13g2_nand2_1 _4062_ (.Y(_0643_),
    .A(net985),
    .B(_0641_));
 sg13g2_a22oi_1 _4063_ (.Y(_0644_),
    .B1(_0479_),
    .B2(net861),
    .A2(_0469_),
    .A1(net986));
 sg13g2_a21o_1 _4064_ (.A2(_0487_),
    .A1(net835),
    .B1(_0644_),
    .X(_0645_));
 sg13g2_nor2_2 _4065_ (.A(_0431_),
    .B(net866),
    .Y(_0646_));
 sg13g2_nand2_2 _4066_ (.Y(_0647_),
    .A(net865),
    .B(_0452_));
 sg13g2_a21oi_2 _4067_ (.B1(net848),
    .Y(_0648_),
    .A2(net863),
    .A1(_0430_));
 sg13g2_a21o_2 _4068_ (.A2(net863),
    .A1(_0430_),
    .B1(net848),
    .X(_0649_));
 sg13g2_a21oi_2 _4069_ (.B1(net838),
    .Y(_0650_),
    .A2(_0649_),
    .A1(net851));
 sg13g2_nor2_1 _4070_ (.A(net863),
    .B(_0480_),
    .Y(_0651_));
 sg13g2_nand2_2 _4071_ (.Y(_0652_),
    .A(net865),
    .B(_0479_));
 sg13g2_nand2_1 _4072_ (.Y(_0653_),
    .A(net836),
    .B(_0651_));
 sg13g2_mux4_1 _4073_ (.S0(net854),
    .A0(_0487_),
    .A1(_0551_),
    .A2(_0652_),
    .A3(_0648_),
    .S1(net845),
    .X(_0654_));
 sg13g2_or2_1 _4074_ (.X(_0655_),
    .B(_0654_),
    .A(net831));
 sg13g2_and2_2 _4075_ (.A(net850),
    .B(_0601_),
    .X(_0656_));
 sg13g2_nand2_1 _4076_ (.Y(_0657_),
    .A(_0587_),
    .B(_0656_));
 sg13g2_a221oi_1 _4077_ (.B2(_0587_),
    .C1(net839),
    .B1(_0656_),
    .A1(net835),
    .Y(_0658_),
    .A2(_0652_));
 sg13g2_nand2_1 _4078_ (.Y(_0659_),
    .A(net831),
    .B(_0658_));
 sg13g2_nand2b_1 _4079_ (.Y(_0660_),
    .B(net863),
    .A_N(_0535_));
 sg13g2_a21o_1 _4080_ (.A2(_0647_),
    .A1(net836),
    .B1(_0536_),
    .X(_0661_));
 sg13g2_nand3_1 _4081_ (.B(_0660_),
    .C(_0661_),
    .A(_0531_),
    .Y(_0662_));
 sg13g2_nand4_1 _4082_ (.B(_0655_),
    .C(_0659_),
    .A(net815),
    .Y(_0663_),
    .D(_0662_));
 sg13g2_nand2_1 _4083_ (.Y(_0664_),
    .A(net841),
    .B(_0585_));
 sg13g2_nand2_1 _4084_ (.Y(_0665_),
    .A(_0392_),
    .B(_0602_));
 sg13g2_a22oi_1 _4085_ (.Y(_0666_),
    .B1(_0602_),
    .B2(_0392_),
    .A2(_0585_),
    .A1(net841));
 sg13g2_o21ai_1 _4086_ (.B1(_0664_),
    .Y(_0667_),
    .A1(net832),
    .A2(_0665_));
 sg13g2_a21oi_1 _4087_ (.A1(net816),
    .A2(_0667_),
    .Y(_0668_),
    .B1(net824));
 sg13g2_nand2_1 _4088_ (.Y(_0669_),
    .A(_0535_),
    .B(_0650_));
 sg13g2_and2_1 _4089_ (.A(net850),
    .B(_0476_),
    .X(_0670_));
 sg13g2_nand2_2 _4090_ (.Y(_0671_),
    .A(net852),
    .B(_0476_));
 sg13g2_o21ai_1 _4091_ (.B1(_0671_),
    .Y(_0672_),
    .A1(_0483_),
    .A2(_0609_));
 sg13g2_a21oi_1 _4092_ (.A1(net860),
    .A2(_0451_),
    .Y(_0673_),
    .B1(_0476_));
 sg13g2_o21ai_1 _4093_ (.B1(_0609_),
    .Y(_0674_),
    .A1(net836),
    .A2(_0673_));
 sg13g2_a22oi_1 _4094_ (.Y(_0675_),
    .B1(_0674_),
    .B2(_0539_),
    .A2(_0672_),
    .A1(_0531_));
 sg13g2_a21o_1 _4095_ (.A2(_0675_),
    .A1(_0669_),
    .B1(net814),
    .X(_0676_));
 sg13g2_nand2_1 _4096_ (.Y(_0677_),
    .A(net839),
    .B(_0529_));
 sg13g2_nor3_1 _4097_ (.A(_0373_),
    .B(_0553_),
    .C(_0677_),
    .Y(_0678_));
 sg13g2_nor2_1 _4098_ (.A(net822),
    .B(_0678_),
    .Y(_0679_));
 sg13g2_a221oi_1 _4099_ (.B2(_0679_),
    .C1(net827),
    .B1(_0676_),
    .A1(_0663_),
    .Y(_0680_),
    .A2(_0668_));
 sg13g2_o21ai_1 _4100_ (.B1(net842),
    .Y(_0681_),
    .A1(net836),
    .A2(_0584_));
 sg13g2_nand3_1 _4101_ (.B(_0665_),
    .C(_0681_),
    .A(net818),
    .Y(_0682_));
 sg13g2_and2_2 _4102_ (.A(net841),
    .B(net829),
    .X(_0683_));
 sg13g2_nand2_2 _4103_ (.Y(_0684_),
    .A(net845),
    .B(net829));
 sg13g2_nand2b_1 _4104_ (.Y(_0685_),
    .B(net823),
    .A_N(_0588_));
 sg13g2_nand4_1 _4105_ (.B(_0682_),
    .C(_0684_),
    .A(net816),
    .Y(_0686_),
    .D(_0685_));
 sg13g2_nor2_2 _4106_ (.A(net843),
    .B(net820),
    .Y(_0687_));
 sg13g2_nand4_1 _4107_ (.B(net837),
    .C(net829),
    .A(net985),
    .Y(_0688_),
    .D(_0670_));
 sg13g2_o21ai_1 _4108_ (.B1(_0688_),
    .Y(_0689_),
    .A1(net823),
    .A2(_0666_));
 sg13g2_nand3_1 _4109_ (.B(_0503_),
    .C(_0689_),
    .A(net816),
    .Y(_0690_));
 sg13g2_o21ai_1 _4110_ (.B1(_0690_),
    .Y(_0691_),
    .A1(net832),
    .A2(_0686_));
 sg13g2_a21o_1 _4111_ (.A2(_0691_),
    .A1(net827),
    .B1(_0680_),
    .X(_0692_));
 sg13g2_a21oi_1 _4112_ (.A1(_0581_),
    .A2(_0692_),
    .Y(_0693_),
    .B1(_0643_));
 sg13g2_nand2_2 _4113_ (.Y(_0694_),
    .A(_0453_),
    .B(_0484_));
 sg13g2_nor3_1 _4114_ (.A(net842),
    .B(net818),
    .C(_0694_),
    .Y(_0695_));
 sg13g2_nor2_2 _4115_ (.A(net839),
    .B(net829),
    .Y(_0696_));
 sg13g2_or4_1 _4116_ (.A(net837),
    .B(net850),
    .C(net829),
    .D(_0673_),
    .X(_0697_));
 sg13g2_nor2_1 _4117_ (.A(net849),
    .B(_0646_),
    .Y(_0698_));
 sg13g2_a21oi_1 _4118_ (.A1(_0587_),
    .A2(_0656_),
    .Y(_0699_),
    .B1(_0698_));
 sg13g2_o21ai_1 _4119_ (.B1(_0697_),
    .Y(_0700_),
    .A1(_0684_),
    .A2(_0699_));
 sg13g2_or4_1 _4120_ (.A(net814),
    .B(_0689_),
    .C(_0695_),
    .D(_0700_),
    .X(_0701_));
 sg13g2_or2_1 _4121_ (.X(_0702_),
    .B(_0551_),
    .A(net853));
 sg13g2_mux4_1 _4122_ (.S0(net836),
    .A0(_0456_),
    .A1(_0587_),
    .A2(_0648_),
    .A3(_0551_),
    .S1(net845),
    .X(_0703_));
 sg13g2_nand2_1 _4123_ (.Y(_0704_),
    .A(net863),
    .B(_0486_));
 sg13g2_a22oi_1 _4124_ (.Y(_0705_),
    .B1(_0486_),
    .B2(net864),
    .A2(net859),
    .A1(net985));
 sg13g2_a22oi_1 _4125_ (.Y(_0706_),
    .B1(_0601_),
    .B2(_0705_),
    .A2(net828),
    .A1(net860));
 sg13g2_nand3_1 _4126_ (.B(_0646_),
    .C(_0683_),
    .A(net852),
    .Y(_0707_));
 sg13g2_a221oi_1 _4127_ (.B2(_0687_),
    .C1(net816),
    .B1(_0706_),
    .A1(net819),
    .Y(_0708_),
    .A2(_0703_));
 sg13g2_nor2_1 _4128_ (.A(net844),
    .B(net825),
    .Y(_0709_));
 sg13g2_nand2_2 _4129_ (.Y(_0710_),
    .A(net839),
    .B(net820));
 sg13g2_a21oi_1 _4130_ (.A1(_0707_),
    .A2(_0708_),
    .Y(_0711_),
    .B1(net830));
 sg13g2_nor2_2 _4131_ (.A(net839),
    .B(_0589_),
    .Y(_0712_));
 sg13g2_nor2_1 _4132_ (.A(_0589_),
    .B(_0684_),
    .Y(_0713_));
 sg13g2_a221oi_1 _4133_ (.B2(_0702_),
    .C1(net824),
    .B1(_0650_),
    .A1(net838),
    .Y(_0714_),
    .A2(_0645_));
 sg13g2_nor3_1 _4134_ (.A(net866),
    .B(_0452_),
    .C(net851),
    .Y(_0715_));
 sg13g2_o21ai_1 _4135_ (.B1(_0586_),
    .Y(_0716_),
    .A1(_0705_),
    .A2(_0715_));
 sg13g2_nor3_1 _4136_ (.A(net842),
    .B(net818),
    .C(_0716_),
    .Y(_0717_));
 sg13g2_or4_1 _4137_ (.A(net816),
    .B(_0713_),
    .C(_0714_),
    .D(_0717_),
    .X(_0718_));
 sg13g2_a21o_1 _4138_ (.A2(_0646_),
    .A1(net849),
    .B1(_0585_),
    .X(_0719_));
 sg13g2_a221oi_1 _4139_ (.B2(net849),
    .C1(_0585_),
    .B1(_0646_),
    .A1(_0550_),
    .Y(_0720_),
    .A2(_0601_));
 sg13g2_nand2b_1 _4140_ (.Y(_0721_),
    .B(net842),
    .A_N(_0720_));
 sg13g2_and3_1 _4141_ (.X(_0722_),
    .A(net818),
    .B(_0665_),
    .C(_0721_));
 sg13g2_nor2_1 _4142_ (.A(net819),
    .B(_0650_),
    .Y(_0723_));
 sg13g2_nand2b_1 _4143_ (.Y(_0724_),
    .B(net823),
    .A_N(_0650_));
 sg13g2_and2_1 _4144_ (.A(net838),
    .B(_0674_),
    .X(_0725_));
 sg13g2_o21ai_1 _4145_ (.B1(net816),
    .Y(_0726_),
    .A1(_0724_),
    .A2(_0725_));
 sg13g2_o21ai_1 _4146_ (.B1(_0718_),
    .Y(_0727_),
    .A1(_0722_),
    .A2(_0726_));
 sg13g2_a221oi_1 _4147_ (.B2(net830),
    .C1(_2777_),
    .B1(_0727_),
    .A1(_0701_),
    .Y(_0728_),
    .A2(_0711_));
 sg13g2_a21oi_1 _4148_ (.A1(_2776_),
    .A2(_0686_),
    .Y(_0729_),
    .B1(_0582_));
 sg13g2_nand2b_1 _4149_ (.Y(_0730_),
    .B(_0729_),
    .A_N(_0728_));
 sg13g2_nand3_1 _4150_ (.B(_0544_),
    .C(_0660_),
    .A(net838),
    .Y(_0731_));
 sg13g2_a21oi_1 _4151_ (.A1(_0535_),
    .A2(_0607_),
    .Y(_0732_),
    .B1(net837));
 sg13g2_nor2_1 _4152_ (.A(net818),
    .B(_0732_),
    .Y(_0733_));
 sg13g2_nand2_1 _4153_ (.Y(_0734_),
    .A(net830),
    .B(_0697_));
 sg13g2_a221oi_1 _4154_ (.B2(_0733_),
    .C1(_0734_),
    .B1(_0731_),
    .A1(_0506_),
    .Y(_0735_),
    .A2(_0696_));
 sg13g2_a21oi_1 _4155_ (.A1(_0550_),
    .A2(_0601_),
    .Y(_0736_),
    .B1(_0589_));
 sg13g2_o21ai_1 _4156_ (.B1(net819),
    .Y(_0737_),
    .A1(net837),
    .A2(_0736_));
 sg13g2_nand3_1 _4157_ (.B(_0535_),
    .C(_0607_),
    .A(net847),
    .Y(_0738_));
 sg13g2_nand2_1 _4158_ (.Y(_0739_),
    .A(_0392_),
    .B(_0536_));
 sg13g2_nand3_1 _4159_ (.B(_0738_),
    .C(_0739_),
    .A(net823),
    .Y(_0740_));
 sg13g2_a21oi_1 _4160_ (.A1(_0737_),
    .A2(_0740_),
    .Y(_0741_),
    .B1(net830));
 sg13g2_nor3_1 _4161_ (.A(_2777_),
    .B(_0735_),
    .C(_0741_),
    .Y(_0742_));
 sg13g2_nor3_1 _4162_ (.A(net837),
    .B(net832),
    .C(_0736_),
    .Y(_0743_));
 sg13g2_nor3_1 _4163_ (.A(net837),
    .B(net830),
    .C(_0720_),
    .Y(_0744_));
 sg13g2_nor4_1 _4164_ (.A(net823),
    .B(_0605_),
    .C(_0743_),
    .D(_0744_),
    .Y(_0745_));
 sg13g2_nand4_1 _4165_ (.B(_0539_),
    .C(_0541_),
    .A(_0507_),
    .Y(_0746_),
    .D(_0586_));
 sg13g2_nand4_1 _4166_ (.B(_0541_),
    .C(_0586_),
    .A(_0531_),
    .Y(_0747_),
    .D(_0590_));
 sg13g2_and4_1 _4167_ (.A(net823),
    .B(_0738_),
    .C(_0746_),
    .D(_0747_),
    .X(_0748_));
 sg13g2_nor3_1 _4168_ (.A(net827),
    .B(_0745_),
    .C(_0748_),
    .Y(_0749_));
 sg13g2_or3_1 _4169_ (.A(net814),
    .B(_0742_),
    .C(_0749_),
    .X(_0750_));
 sg13g2_nand2_1 _4170_ (.Y(_0751_),
    .A(net866),
    .B(_0455_));
 sg13g2_and2_1 _4171_ (.A(net855),
    .B(_0751_),
    .X(_0752_));
 sg13g2_and3_1 _4172_ (.X(_0753_),
    .A(net854),
    .B(_0587_),
    .C(_0751_));
 sg13g2_nand2_1 _4173_ (.Y(_0754_),
    .A(_0456_),
    .B(_0477_));
 sg13g2_a21oi_1 _4174_ (.A1(net835),
    .A2(_0754_),
    .Y(_0755_),
    .B1(_0753_));
 sg13g2_a21oi_1 _4175_ (.A1(_0687_),
    .A2(_0755_),
    .Y(_0756_),
    .B1(_0713_));
 sg13g2_o21ai_1 _4176_ (.B1(_0531_),
    .Y(_0757_),
    .A1(_0610_),
    .A2(_0644_));
 sg13g2_nand3_1 _4177_ (.B(_0604_),
    .C(_0645_),
    .A(_0539_),
    .Y(_0758_));
 sg13g2_a21oi_1 _4178_ (.A1(_0757_),
    .A2(_0758_),
    .Y(_0759_),
    .B1(_2777_));
 sg13g2_nand4_1 _4179_ (.B(net865),
    .C(_0455_),
    .A(net986),
    .Y(_0760_),
    .D(net859));
 sg13g2_nand4_1 _4180_ (.B(_0586_),
    .C(_0660_),
    .A(_0507_),
    .Y(_0761_),
    .D(_0760_));
 sg13g2_o21ai_1 _4181_ (.B1(net822),
    .Y(_0762_),
    .A1(net839),
    .A2(_0761_));
 sg13g2_o21ai_1 _4182_ (.B1(_0482_),
    .Y(_0763_),
    .A1(net853),
    .A2(_0704_));
 sg13g2_nor2_1 _4183_ (.A(net827),
    .B(net847),
    .Y(_0764_));
 sg13g2_a21o_1 _4184_ (.A2(_0764_),
    .A1(_0763_),
    .B1(_0762_),
    .X(_0765_));
 sg13g2_o21ai_1 _4185_ (.B1(_0756_),
    .Y(_0766_),
    .A1(_0759_),
    .A2(_0765_));
 sg13g2_a21oi_1 _4186_ (.A1(net814),
    .A2(_0766_),
    .Y(_0767_),
    .B1(_0583_));
 sg13g2_a21oi_1 _4187_ (.A1(_0750_),
    .A2(_0767_),
    .Y(_0768_),
    .B1(_0642_));
 sg13g2_a22oi_1 _4188_ (.Y(_0769_),
    .B1(_0619_),
    .B2(_0621_),
    .A2(net935),
    .A1(_2441_));
 sg13g2_xnor2_1 _4189_ (.Y(_0770_),
    .A(\i_bitmap.in[11] ),
    .B(net938));
 sg13g2_o21ai_1 _4190_ (.B1(net887),
    .Y(_0771_),
    .A1(_0769_),
    .A2(_0770_));
 sg13g2_a21oi_1 _4191_ (.A1(_0769_),
    .A2(_0770_),
    .Y(_0772_),
    .B1(_0771_));
 sg13g2_nor2_1 _4192_ (.A(_0037_),
    .B(net935),
    .Y(_0773_));
 sg13g2_xnor2_1 _4193_ (.Y(_0774_),
    .A(_0037_),
    .B(net938));
 sg13g2_nand2_1 _4194_ (.Y(_0775_),
    .A(_0624_),
    .B(_0625_));
 sg13g2_a21oi_1 _4195_ (.A1(_0626_),
    .A2(_0775_),
    .Y(_0776_),
    .B1(_0774_));
 sg13g2_and3_1 _4196_ (.X(_0777_),
    .A(_0626_),
    .B(_0774_),
    .C(_0775_));
 sg13g2_nor2_1 _4197_ (.A(_0776_),
    .B(_0777_),
    .Y(_0778_));
 sg13g2_o21ai_1 _4198_ (.B1(net902),
    .Y(_0779_),
    .A1(net887),
    .A2(_0778_));
 sg13g2_xnor2_1 _4199_ (.Y(_0780_),
    .A(_2418_),
    .B(net972));
 sg13g2_a21oi_1 _4200_ (.A1(_0036_),
    .A2(net899),
    .Y(_0781_),
    .B1(_0634_));
 sg13g2_nor2_1 _4201_ (.A(_0635_),
    .B(_0781_),
    .Y(_0782_));
 sg13g2_nand2b_1 _4202_ (.Y(_0783_),
    .B(_0782_),
    .A_N(_0780_));
 sg13g2_nor2b_1 _4203_ (.A(_0782_),
    .B_N(_0780_),
    .Y(_0784_));
 sg13g2_nand3b_1 _4204_ (.B(net879),
    .C(_0783_),
    .Y(_0785_),
    .A_N(_0784_));
 sg13g2_nand2_1 _4205_ (.Y(_0786_),
    .A(\i_bitmap.in[10] ),
    .B(net966));
 sg13g2_o21ai_1 _4206_ (.B1(_0786_),
    .Y(_0787_),
    .A1(_0631_),
    .A2(_0632_));
 sg13g2_xnor2_1 _4207_ (.Y(_0788_),
    .A(_2442_),
    .B(net970));
 sg13g2_a21oi_1 _4208_ (.A1(_0787_),
    .A2(_0788_),
    .Y(_0789_),
    .B1(net879));
 sg13g2_o21ai_1 _4209_ (.B1(_0789_),
    .Y(_0790_),
    .A1(_0787_),
    .A2(_0788_));
 sg13g2_a21o_1 _4210_ (.A2(_0790_),
    .A1(_0785_),
    .B1(net884),
    .X(_0791_));
 sg13g2_o21ai_1 _4211_ (.B1(_0791_),
    .Y(_0792_),
    .A1(_0772_),
    .A2(_0779_));
 sg13g2_a21oi_2 _4212_ (.B1(_0792_),
    .Y(_0793_),
    .A2(_2695_),
    .A1(_2442_));
 sg13g2_nor2_1 _4213_ (.A(net981),
    .B(_0793_),
    .Y(_0794_));
 sg13g2_nand2b_1 _4214_ (.Y(_0795_),
    .B(net985),
    .A_N(_0793_));
 sg13g2_a221oi_1 _4215_ (.B2(_0768_),
    .C1(_0794_),
    .B1(_0730_),
    .A1(_0618_),
    .Y(_0796_),
    .A2(_0693_));
 sg13g2_nor2_1 _4216_ (.A(net841),
    .B(net828),
    .Y(_0797_));
 sg13g2_nor3_1 _4217_ (.A(net841),
    .B(_0506_),
    .C(net828),
    .Y(_0798_));
 sg13g2_o21ai_1 _4218_ (.B1(net818),
    .Y(_0799_),
    .A1(_0484_),
    .A2(_0719_));
 sg13g2_nor2_1 _4219_ (.A(_0503_),
    .B(_0798_),
    .Y(_0800_));
 sg13g2_nand3_1 _4220_ (.B(_0537_),
    .C(_0647_),
    .A(net851),
    .Y(_0801_));
 sg13g2_inv_1 _4221_ (.Y(_0802_),
    .A(_0801_));
 sg13g2_o21ai_1 _4222_ (.B1(_0801_),
    .Y(_0803_),
    .A1(net852),
    .A2(_0584_));
 sg13g2_a221oi_1 _4223_ (.B2(net818),
    .C1(net830),
    .B1(_0803_),
    .A1(_0590_),
    .Y(_0804_),
    .A2(_0797_));
 sg13g2_a21oi_1 _4224_ (.A1(_0799_),
    .A2(_0800_),
    .Y(_0805_),
    .B1(_0804_));
 sg13g2_nand2_1 _4225_ (.Y(_0806_),
    .A(net816),
    .B(_0805_));
 sg13g2_a21oi_1 _4226_ (.A1(net815),
    .A2(_0763_),
    .Y(_0807_),
    .B1(_0710_));
 sg13g2_a21oi_1 _4227_ (.A1(net842),
    .A2(_0611_),
    .Y(_0808_),
    .B1(net824));
 sg13g2_nor2_1 _4228_ (.A(_0599_),
    .B(_0808_),
    .Y(_0809_));
 sg13g2_o21ai_1 _4229_ (.B1(net827),
    .Y(_0810_),
    .A1(_0595_),
    .A2(_0684_));
 sg13g2_nor3_1 _4230_ (.A(_0807_),
    .B(_0809_),
    .C(_0810_),
    .Y(_0811_));
 sg13g2_nand3_1 _4231_ (.B(net851),
    .C(_0476_),
    .A(_0428_),
    .Y(_0812_));
 sg13g2_a21oi_2 _4232_ (.B1(_0671_),
    .Y(_0813_),
    .A2(net830),
    .A1(_0429_));
 sg13g2_nor3_1 _4233_ (.A(net843),
    .B(_0542_),
    .C(_0550_),
    .Y(_0814_));
 sg13g2_nor3_1 _4234_ (.A(net822),
    .B(_0677_),
    .C(_0813_),
    .Y(_0815_));
 sg13g2_nor2_1 _4235_ (.A(net817),
    .B(_0815_),
    .Y(_0816_));
 sg13g2_o21ai_1 _4236_ (.B1(net834),
    .Y(_0817_),
    .A1(_0658_),
    .A2(_0814_));
 sg13g2_o21ai_1 _4237_ (.B1(_0817_),
    .Y(_0818_),
    .A1(net834),
    .A2(_0654_));
 sg13g2_o21ai_1 _4238_ (.B1(_0816_),
    .Y(_0819_),
    .A1(net825),
    .A2(_0818_));
 sg13g2_nor3_1 _4239_ (.A(net837),
    .B(_0602_),
    .C(_0656_),
    .Y(_0820_));
 sg13g2_or2_1 _4240_ (.X(_0821_),
    .B(_0820_),
    .A(net823));
 sg13g2_nand2b_1 _4241_ (.Y(_0822_),
    .B(_0687_),
    .A_N(_0610_));
 sg13g2_nand3_1 _4242_ (.B(_0649_),
    .C(_0683_),
    .A(_0529_),
    .Y(_0823_));
 sg13g2_nand4_1 _4243_ (.B(_0821_),
    .C(_0822_),
    .A(net833),
    .Y(_0824_),
    .D(_0823_));
 sg13g2_nand2_2 _4244_ (.Y(_0825_),
    .A(net845),
    .B(_0543_));
 sg13g2_a221oi_1 _4245_ (.B2(net819),
    .C1(net833),
    .B1(_0825_),
    .A1(_0609_),
    .Y(_0826_),
    .A2(_0723_));
 sg13g2_nor2_1 _4246_ (.A(net814),
    .B(_0826_),
    .Y(_0827_));
 sg13g2_a21oi_1 _4247_ (.A1(_0824_),
    .A2(_0827_),
    .Y(_0828_),
    .B1(net827));
 sg13g2_a22oi_1 _4248_ (.Y(_0829_),
    .B1(_0819_),
    .B2(_0828_),
    .A2(_0811_),
    .A1(_0806_));
 sg13g2_nor4_1 _4249_ (.A(_0580_),
    .B(_0641_),
    .C(_0795_),
    .D(_0829_),
    .Y(_0830_));
 sg13g2_nand3_1 _4250_ (.B(_0621_),
    .C(_0770_),
    .A(_0619_),
    .Y(_0831_));
 sg13g2_a21oi_1 _4251_ (.A1(_2418_),
    .A2(_2441_),
    .Y(_0832_),
    .B1(_2442_));
 sg13g2_o21ai_1 _4252_ (.B1(_0831_),
    .Y(_0833_),
    .A1(net941),
    .A2(_0832_));
 sg13g2_and2_1 _4253_ (.A(\i_bitmap.in[12] ),
    .B(net937),
    .X(_0834_));
 sg13g2_nand2_1 _4254_ (.Y(_0835_),
    .A(\i_bitmap.in[12] ),
    .B(net941));
 sg13g2_xnor2_1 _4255_ (.Y(_0836_),
    .A(\i_bitmap.in[12] ),
    .B(net941));
 sg13g2_xor2_1 _4256_ (.B(_0836_),
    .A(_0833_),
    .X(_0837_));
 sg13g2_nor2_2 _4257_ (.A(net977),
    .B(net906),
    .Y(_0838_));
 sg13g2_nand2_2 _4258_ (.Y(_0839_),
    .A(net984),
    .B(net901));
 sg13g2_xnor2_1 _4259_ (.Y(_0840_),
    .A(_0038_),
    .B(net941));
 sg13g2_or3_1 _4260_ (.A(_0773_),
    .B(_0777_),
    .C(_0840_),
    .X(_0841_));
 sg13g2_o21ai_1 _4261_ (.B1(_0840_),
    .Y(_0842_),
    .A1(_0773_),
    .A2(_0777_));
 sg13g2_a21oi_1 _4262_ (.A1(_0841_),
    .A2(_0842_),
    .Y(_0843_),
    .B1(net888));
 sg13g2_nor2_1 _4263_ (.A(_0839_),
    .B(_0843_),
    .Y(_0844_));
 sg13g2_o21ai_1 _4264_ (.B1(_0844_),
    .Y(_0845_),
    .A1(net893),
    .A2(_0837_));
 sg13g2_a21oi_1 _4265_ (.A1(\i_bitmap.in[11] ),
    .A2(net972),
    .Y(_0846_),
    .B1(_0784_));
 sg13g2_xnor2_1 _4266_ (.Y(_0847_),
    .A(\i_bitmap.in[12] ),
    .B(net972));
 sg13g2_inv_1 _4267_ (.Y(_0848_),
    .A(_0847_));
 sg13g2_xnor2_1 _4268_ (.Y(_0849_),
    .A(_0846_),
    .B(_0848_));
 sg13g2_a22oi_1 _4269_ (.Y(_0850_),
    .B1(_0787_),
    .B2(_0788_),
    .A2(net968),
    .A1(\i_bitmap.in[11] ));
 sg13g2_xnor2_1 _4270_ (.Y(_0851_),
    .A(_0038_),
    .B(net972));
 sg13g2_nand2_1 _4271_ (.Y(_0852_),
    .A(_0850_),
    .B(_0851_));
 sg13g2_nor2_1 _4272_ (.A(_0850_),
    .B(_0851_),
    .Y(_0853_));
 sg13g2_nor2_1 _4273_ (.A(net880),
    .B(_0853_),
    .Y(_0854_));
 sg13g2_a22oi_1 _4274_ (.Y(_0855_),
    .B1(_0852_),
    .B2(_0854_),
    .A2(_0849_),
    .A1(net880));
 sg13g2_nor2_1 _4275_ (.A(net982),
    .B(net885),
    .Y(_0856_));
 sg13g2_nand2_1 _4276_ (.Y(_0857_),
    .A(net990),
    .B(_0341_));
 sg13g2_o21ai_1 _4277_ (.B1(_0845_),
    .Y(_0858_),
    .A1(_0855_),
    .A2(net883));
 sg13g2_nor2_2 _4278_ (.A(net976),
    .B(net894),
    .Y(_0859_));
 sg13g2_a21oi_2 _4279_ (.B1(_0858_),
    .Y(_0860_),
    .A2(net882),
    .A1(_2443_));
 sg13g2_o21ai_1 _4280_ (.B1(_0860_),
    .Y(_0861_),
    .A1(_0796_),
    .A2(_0830_));
 sg13g2_o21ai_1 _4281_ (.B1(_0684_),
    .Y(_0862_),
    .A1(net822),
    .A2(_0608_));
 sg13g2_o21ai_1 _4282_ (.B1(net834),
    .Y(_0863_),
    .A1(net829),
    .A2(_0653_));
 sg13g2_a221oi_1 _4283_ (.B2(_0669_),
    .C1(_0863_),
    .B1(_0862_),
    .A1(net819),
    .Y(_0864_),
    .A2(_0825_));
 sg13g2_nand3_1 _4284_ (.B(net824),
    .C(_0694_),
    .A(net838),
    .Y(_0865_));
 sg13g2_nand3_1 _4285_ (.B(_0657_),
    .C(_0683_),
    .A(_0541_),
    .Y(_0866_));
 sg13g2_nand4_1 _4286_ (.B(_0821_),
    .C(_0865_),
    .A(net831),
    .Y(_0867_),
    .D(_0866_));
 sg13g2_nand2b_1 _4287_ (.Y(_0868_),
    .B(_0867_),
    .A_N(_0864_));
 sg13g2_a21oi_1 _4288_ (.A1(_0431_),
    .A2(_0587_),
    .Y(_0869_),
    .B1(net835));
 sg13g2_and2_1 _4289_ (.A(_0477_),
    .B(_0550_),
    .X(_0870_));
 sg13g2_o21ai_1 _4290_ (.B1(_0539_),
    .Y(_0871_),
    .A1(_0869_),
    .A2(_0870_));
 sg13g2_o21ai_1 _4291_ (.B1(_0531_),
    .Y(_0872_),
    .A1(net828),
    .A2(_0588_));
 sg13g2_nand2_1 _4292_ (.Y(_0873_),
    .A(_0871_),
    .B(_0872_));
 sg13g2_o21ai_1 _4293_ (.B1(net825),
    .Y(_0874_),
    .A1(_0712_),
    .A2(_0873_));
 sg13g2_a221oi_1 _4294_ (.B2(net986),
    .C1(_0479_),
    .B1(_0469_),
    .A1(_0427_),
    .Y(_0875_),
    .A2(net865));
 sg13g2_nor3_1 _4295_ (.A(_0608_),
    .B(_0710_),
    .C(_0875_),
    .Y(_0876_));
 sg13g2_a21oi_1 _4296_ (.A1(_0696_),
    .A2(_0761_),
    .Y(_0877_),
    .B1(net817));
 sg13g2_nor2b_1 _4297_ (.A(_0876_),
    .B_N(_0877_),
    .Y(_0878_));
 sg13g2_a22oi_1 _4298_ (.Y(_0879_),
    .B1(_0874_),
    .B2(_0878_),
    .A2(_0868_),
    .A1(net817));
 sg13g2_or2_1 _4299_ (.X(_0880_),
    .B(_0879_),
    .A(_2776_));
 sg13g2_nor4_1 _4300_ (.A(net841),
    .B(net832),
    .C(net828),
    .D(_0589_),
    .Y(_0881_));
 sg13g2_a21oi_1 _4301_ (.A1(net832),
    .A2(_0798_),
    .Y(_0882_),
    .B1(_0881_));
 sg13g2_nor2_1 _4302_ (.A(net832),
    .B(_0801_),
    .Y(_0883_));
 sg13g2_a21oi_1 _4303_ (.A1(net832),
    .A2(_0719_),
    .Y(_0884_),
    .B1(_0883_));
 sg13g2_a21oi_1 _4304_ (.A1(_0480_),
    .A2(_0587_),
    .Y(_0885_),
    .B1(net851));
 sg13g2_nor2_1 _4305_ (.A(net823),
    .B(_0885_),
    .Y(_0886_));
 sg13g2_a22oi_1 _4306_ (.Y(_0887_),
    .B1(_0884_),
    .B2(_0886_),
    .A2(_0882_),
    .A1(_0733_));
 sg13g2_a21oi_1 _4307_ (.A1(net862),
    .A2(_0534_),
    .Y(_0888_),
    .B1(_0875_));
 sg13g2_nand2_1 _4308_ (.Y(_0889_),
    .A(_0756_),
    .B(_0877_));
 sg13g2_o21ai_1 _4309_ (.B1(_0889_),
    .Y(_0890_),
    .A1(net815),
    .A2(_0887_));
 sg13g2_o21ai_1 _4310_ (.B1(_0709_),
    .Y(_0891_),
    .A1(_0888_),
    .A2(_0889_));
 sg13g2_nand3_1 _4311_ (.B(_0890_),
    .C(_0891_),
    .A(_2777_),
    .Y(_0892_));
 sg13g2_nand3_1 _4312_ (.B(_0880_),
    .C(_0892_),
    .A(_0794_),
    .Y(_0893_));
 sg13g2_a21oi_1 _4313_ (.A1(_0580_),
    .A2(_0893_),
    .Y(_0894_),
    .B1(_0643_));
 sg13g2_o21ai_1 _4314_ (.B1(_0712_),
    .Y(_0895_),
    .A1(net855),
    .A2(_0648_));
 sg13g2_nor2_1 _4315_ (.A(net836),
    .B(_0652_),
    .Y(_0896_));
 sg13g2_a22oi_1 _4316_ (.Y(_0897_),
    .B1(_0651_),
    .B2(net853),
    .A2(_0536_),
    .A1(_0470_));
 sg13g2_o21ai_1 _4317_ (.B1(_0897_),
    .Y(_0898_),
    .A1(net855),
    .A2(_0478_));
 sg13g2_o21ai_1 _4318_ (.B1(_0604_),
    .Y(_0899_),
    .A1(_0456_),
    .A2(net854));
 sg13g2_nor3_1 _4319_ (.A(_0684_),
    .B(_0752_),
    .C(_0899_),
    .Y(_0900_));
 sg13g2_a221oi_1 _4320_ (.B2(_0687_),
    .C1(_0900_),
    .B1(_0898_),
    .A1(net821),
    .Y(_0901_),
    .A2(_0895_));
 sg13g2_o21ai_1 _4321_ (.B1(_0897_),
    .Y(_0902_),
    .A1(net854),
    .A2(_0647_));
 sg13g2_nand4_1 _4322_ (.B(_0411_),
    .C(net861),
    .A(net986),
    .Y(_0903_),
    .D(net859));
 sg13g2_nand4_1 _4323_ (.B(_0603_),
    .C(_0801_),
    .A(net843),
    .Y(_0904_),
    .D(_0903_));
 sg13g2_nand2_1 _4324_ (.Y(_0905_),
    .A(_0453_),
    .B(_0455_));
 sg13g2_a21oi_1 _4325_ (.A1(_0527_),
    .A2(_0905_),
    .Y(_0906_),
    .B1(_0684_));
 sg13g2_a22oi_1 _4326_ (.Y(_0907_),
    .B1(_0904_),
    .B2(net820),
    .A2(_0902_),
    .A1(_0687_));
 sg13g2_nor2_1 _4327_ (.A(_0505_),
    .B(_0906_),
    .Y(_0908_));
 sg13g2_a221oi_1 _4328_ (.B2(_0908_),
    .C1(net815),
    .B1(_0907_),
    .A1(net831),
    .Y(_0909_),
    .A2(_0901_));
 sg13g2_nor2b_1 _4329_ (.A(_0584_),
    .B_N(_0550_),
    .Y(_0910_));
 sg13g2_o21ai_1 _4330_ (.B1(net839),
    .Y(_0911_),
    .A1(net835),
    .A2(_0647_));
 sg13g2_nand3_1 _4331_ (.B(_0478_),
    .C(_0480_),
    .A(net835),
    .Y(_0912_));
 sg13g2_inv_1 _4332_ (.Y(_0913_),
    .A(_0912_));
 sg13g2_nand3_1 _4333_ (.B(_0590_),
    .C(_0912_),
    .A(_0586_),
    .Y(_0914_));
 sg13g2_o21ai_1 _4334_ (.B1(net834),
    .Y(_0915_),
    .A1(_0910_),
    .A2(_0911_));
 sg13g2_a21oi_1 _4335_ (.A1(net845),
    .A2(_0914_),
    .Y(_0916_),
    .B1(_0915_));
 sg13g2_o21ai_1 _4336_ (.B1(net853),
    .Y(_0917_),
    .A1(net865),
    .A2(_0452_));
 sg13g2_nand3_1 _4337_ (.B(_0912_),
    .C(_0917_),
    .A(net845),
    .Y(_0918_));
 sg13g2_o21ai_1 _4338_ (.B1(_0812_),
    .Y(_0919_),
    .A1(_0431_),
    .A2(_0529_));
 sg13g2_a21oi_1 _4339_ (.A1(_0531_),
    .A2(_0919_),
    .Y(_0920_),
    .B1(_0525_));
 sg13g2_o21ai_1 _4340_ (.B1(_0920_),
    .Y(_0921_),
    .A1(_0503_),
    .A2(_0918_));
 sg13g2_or4_2 _4341_ (.A(net841),
    .B(net818),
    .C(_0602_),
    .D(_0705_),
    .X(_0922_));
 sg13g2_o21ai_1 _4342_ (.B1(_0922_),
    .Y(_0923_),
    .A1(_0916_),
    .A2(_0921_));
 sg13g2_o21ai_1 _4343_ (.B1(net827),
    .Y(_0924_),
    .A1(net816),
    .A2(_0923_));
 sg13g2_o21ai_1 _4344_ (.B1(_0583_),
    .Y(_0925_),
    .A1(_0909_),
    .A2(_0924_));
 sg13g2_a221oi_1 _4345_ (.B2(net856),
    .C1(net840),
    .B1(_0754_),
    .A1(_0455_),
    .Y(_0926_),
    .A2(_0550_));
 sg13g2_nor3_1 _4346_ (.A(_0393_),
    .B(_0608_),
    .C(_0705_),
    .Y(_0927_));
 sg13g2_nor2_1 _4347_ (.A(net821),
    .B(_0927_),
    .Y(_0928_));
 sg13g2_nand2_1 _4348_ (.Y(_0929_),
    .A(net843),
    .B(_0473_));
 sg13g2_o21ai_1 _4349_ (.B1(net821),
    .Y(_0930_),
    .A1(_0588_),
    .A2(_0929_));
 sg13g2_nor2_1 _4350_ (.A(net854),
    .B(_0552_),
    .Y(_0931_));
 sg13g2_nor2b_1 _4351_ (.A(_0931_),
    .B_N(_0897_),
    .Y(_0932_));
 sg13g2_or2_1 _4352_ (.X(_0933_),
    .B(_0932_),
    .A(net844));
 sg13g2_and2_1 _4353_ (.A(_0760_),
    .B(_0903_),
    .X(_0934_));
 sg13g2_nand2_1 _4354_ (.Y(_0935_),
    .A(_0760_),
    .B(_0903_));
 sg13g2_o21ai_1 _4355_ (.B1(_0709_),
    .Y(_0936_),
    .A1(_0553_),
    .A2(_0935_));
 sg13g2_o21ai_1 _4356_ (.B1(net833),
    .Y(_0937_),
    .A1(_0753_),
    .A2(_0899_));
 sg13g2_nand3b_1 _4357_ (.B(_0694_),
    .C(_0505_),
    .Y(_0938_),
    .A_N(_0869_));
 sg13g2_nand3_1 _4358_ (.B(_0937_),
    .C(_0938_),
    .A(_0683_),
    .Y(_0939_));
 sg13g2_o21ai_1 _4359_ (.B1(_0375_),
    .Y(_0940_),
    .A1(_0926_),
    .A2(_0928_));
 sg13g2_a21o_1 _4360_ (.A2(_0933_),
    .A1(_0930_),
    .B1(net815),
    .X(_0941_));
 sg13g2_nand4_1 _4361_ (.B(_0939_),
    .C(_0940_),
    .A(_0936_),
    .Y(_0942_),
    .D(_0941_));
 sg13g2_a21oi_1 _4362_ (.A1(_2777_),
    .A2(_0942_),
    .Y(_0943_),
    .B1(_0793_));
 sg13g2_a21oi_1 _4363_ (.A1(_0925_),
    .A2(_0943_),
    .Y(_0944_),
    .B1(_0642_));
 sg13g2_nand2_1 _4364_ (.Y(_0945_),
    .A(_0543_),
    .B(_0551_));
 sg13g2_a21o_1 _4365_ (.A2(_0945_),
    .A1(_0696_),
    .B1(net826),
    .X(_0946_));
 sg13g2_a21oi_1 _4366_ (.A1(_0812_),
    .A2(_0934_),
    .Y(_0947_),
    .B1(_0710_));
 sg13g2_a21oi_1 _4367_ (.A1(_0647_),
    .A2(_0705_),
    .Y(_0948_),
    .B1(net843));
 sg13g2_a21oi_1 _4368_ (.A1(_0603_),
    .A2(_0948_),
    .Y(_0949_),
    .B1(net820));
 sg13g2_nor3_1 _4369_ (.A(_0946_),
    .B(_0947_),
    .C(_0949_),
    .Y(_0950_));
 sg13g2_nor2_1 _4370_ (.A(net843),
    .B(_0896_),
    .Y(_0951_));
 sg13g2_o21ai_1 _4371_ (.B1(_0951_),
    .Y(_0952_),
    .A1(net855),
    .A2(_0552_));
 sg13g2_a21o_1 _4372_ (.A2(_0647_),
    .A1(net854),
    .B1(_0649_),
    .X(_0953_));
 sg13g2_a21oi_1 _4373_ (.A1(net847),
    .A2(_0953_),
    .Y(_0954_),
    .B1(net820));
 sg13g2_a221oi_1 _4374_ (.B2(_0954_),
    .C1(net815),
    .B1(_0952_),
    .A1(net820),
    .Y(_0955_),
    .A2(_0895_));
 sg13g2_nor3_1 _4375_ (.A(net831),
    .B(_0950_),
    .C(_0955_),
    .Y(_0956_));
 sg13g2_nand3_1 _4376_ (.B(_0454_),
    .C(_0543_),
    .A(net843),
    .Y(_0957_));
 sg13g2_nand3_1 _4377_ (.B(_0671_),
    .C(_0934_),
    .A(net840),
    .Y(_0958_));
 sg13g2_a21o_1 _4378_ (.A2(_0958_),
    .A1(_0957_),
    .B1(net825),
    .X(_0959_));
 sg13g2_nand3_1 _4379_ (.B(_0687_),
    .C(_0801_),
    .A(_0603_),
    .Y(_0960_));
 sg13g2_a21oi_1 _4380_ (.A1(_0959_),
    .A2(_0960_),
    .Y(_0961_),
    .B1(net826));
 sg13g2_nor2_1 _4381_ (.A(net848),
    .B(_0594_),
    .Y(_0962_));
 sg13g2_o21ai_1 _4382_ (.B1(net841),
    .Y(_0963_),
    .A1(_0698_),
    .A2(_0962_));
 sg13g2_nand4_1 _4383_ (.B(_0473_),
    .C(_0544_),
    .A(net840),
    .Y(_0964_),
    .D(_0751_));
 sg13g2_a21oi_1 _4384_ (.A1(_0963_),
    .A2(_0964_),
    .Y(_0965_),
    .B1(net820));
 sg13g2_a221oi_1 _4385_ (.B2(_0904_),
    .C1(_0965_),
    .B1(net821),
    .A1(_0371_),
    .Y(_0966_),
    .A2(_0372_));
 sg13g2_nor3_1 _4386_ (.A(net833),
    .B(_0961_),
    .C(_0966_),
    .Y(_0967_));
 sg13g2_or3_1 _4387_ (.A(_2776_),
    .B(_0956_),
    .C(_0967_),
    .X(_0968_));
 sg13g2_nor2_1 _4388_ (.A(net844),
    .B(_0553_),
    .Y(_0969_));
 sg13g2_a221oi_1 _4389_ (.B2(_0760_),
    .C1(net825),
    .B1(_0969_),
    .A1(net847),
    .Y(_0970_),
    .A2(_0913_));
 sg13g2_nor3_1 _4390_ (.A(net826),
    .B(_0928_),
    .C(_0970_),
    .Y(_0971_));
 sg13g2_a221oi_1 _4391_ (.B2(_0712_),
    .C1(net820),
    .B1(_0953_),
    .A1(net840),
    .Y(_0972_),
    .A2(_0932_));
 sg13g2_nand2_1 _4392_ (.Y(_0973_),
    .A(net817),
    .B(_0930_));
 sg13g2_nor2_1 _4393_ (.A(_0972_),
    .B(_0973_),
    .Y(_0974_));
 sg13g2_o21ai_1 _4394_ (.B1(_2776_),
    .Y(_0975_),
    .A1(_0971_),
    .A2(_0974_));
 sg13g2_and3_1 _4395_ (.X(_0976_),
    .A(_0793_),
    .B(_0968_),
    .C(_0975_));
 sg13g2_and3_1 _4396_ (.X(_0977_),
    .A(_0375_),
    .B(_0473_),
    .C(_0917_));
 sg13g2_o21ai_1 _4397_ (.B1(_0524_),
    .Y(_0978_),
    .A1(_0610_),
    .A2(_0656_));
 sg13g2_nor2_1 _4398_ (.A(net831),
    .B(_0977_),
    .Y(_0979_));
 sg13g2_nand2b_1 _4399_ (.Y(_0980_),
    .B(_0375_),
    .A_N(_0914_));
 sg13g2_a221oi_1 _4400_ (.B2(net835),
    .C1(net822),
    .B1(_0649_),
    .A1(_0470_),
    .Y(_0981_),
    .A2(net848));
 sg13g2_nor2_1 _4401_ (.A(net833),
    .B(_0981_),
    .Y(_0982_));
 sg13g2_a221oi_1 _4402_ (.B2(_0982_),
    .C1(net840),
    .B1(_0980_),
    .A1(_0978_),
    .Y(_0983_),
    .A2(_0979_));
 sg13g2_o21ai_1 _4403_ (.B1(net821),
    .Y(_0984_),
    .A1(_0802_),
    .A2(_0929_));
 sg13g2_a21oi_1 _4404_ (.A1(_0933_),
    .A2(_0984_),
    .Y(_0985_),
    .B1(net815));
 sg13g2_nor3_1 _4405_ (.A(_0393_),
    .B(_0584_),
    .C(_0705_),
    .Y(_0986_));
 sg13g2_nor3_1 _4406_ (.A(net826),
    .B(net821),
    .C(_0986_),
    .Y(_0987_));
 sg13g2_a221oi_1 _4407_ (.B2(_0431_),
    .C1(_0710_),
    .B1(_0608_),
    .A1(_0477_),
    .Y(_0988_),
    .A2(_0542_));
 sg13g2_nor4_2 _4408_ (.A(_0983_),
    .B(_0985_),
    .C(_0987_),
    .Y(_0989_),
    .D(_0988_));
 sg13g2_nor3_1 _4409_ (.A(_2776_),
    .B(_0580_),
    .C(_0989_),
    .Y(_0990_));
 sg13g2_or4_1 _4410_ (.A(_0860_),
    .B(_0944_),
    .C(_0976_),
    .D(_0990_),
    .X(_0991_));
 sg13g2_o21ai_1 _4411_ (.B1(_0861_),
    .Y(_0000_),
    .A1(_0894_),
    .A2(_0991_));
 sg13g2_and2_1 _4412_ (.A(\i_orchestrator.vga_x[1] ),
    .B(net326),
    .X(_0992_));
 sg13g2_and2_1 _4413_ (.A(net346),
    .B(_0992_),
    .X(_0993_));
 sg13g2_and2_1 _4414_ (.A(net463),
    .B(_0993_),
    .X(_0994_));
 sg13g2_and2_1 _4415_ (.A(net538),
    .B(_0994_),
    .X(_0995_));
 sg13g2_nand2_1 _4416_ (.Y(_0996_),
    .A(net1060),
    .B(\i_orchestrator.vga_x[8] ));
 sg13g2_nor4_1 _4417_ (.A(\i_orchestrator.vga_x[5] ),
    .B(net1061),
    .C(\i_orchestrator.vga_x[6] ),
    .D(_0996_),
    .Y(_0997_));
 sg13g2_and2_1 _4418_ (.A(_0995_),
    .B(_0997_),
    .X(_0998_));
 sg13g2_nor2_2 _4419_ (.A(net1068),
    .B(_0998_),
    .Y(_0999_));
 sg13g2_nand2b_1 _4420_ (.Y(_1000_),
    .B(net1074),
    .A_N(_0998_));
 sg13g2_and2_1 _4421_ (.A(net244),
    .B(_0999_),
    .X(_0075_));
 sg13g2_nor2_1 _4422_ (.A(\i_orchestrator.vga_x[1] ),
    .B(net326),
    .Y(_1001_));
 sg13g2_nor3_1 _4423_ (.A(_0992_),
    .B(net908),
    .C(net327),
    .Y(_0076_));
 sg13g2_nor2_1 _4424_ (.A(net346),
    .B(_0992_),
    .Y(_1002_));
 sg13g2_nor3_1 _4425_ (.A(net1068),
    .B(_0993_),
    .C(net347),
    .Y(_0077_));
 sg13g2_o21ai_1 _4426_ (.B1(net1078),
    .Y(_1003_),
    .A1(net463),
    .A2(_0993_));
 sg13g2_nor2_1 _4427_ (.A(_0994_),
    .B(_1003_),
    .Y(_0078_));
 sg13g2_o21ai_1 _4428_ (.B1(net1078),
    .Y(_1004_),
    .A1(net495),
    .A2(_0994_));
 sg13g2_nor2_1 _4429_ (.A(_0995_),
    .B(_1004_),
    .Y(_0079_));
 sg13g2_o21ai_1 _4430_ (.B1(_0999_),
    .Y(_1005_),
    .A1(net1062),
    .A2(_0995_));
 sg13g2_a21oi_1 _4431_ (.A1(net1062),
    .A2(_0995_),
    .Y(_0080_),
    .B1(_1005_));
 sg13g2_a21oi_1 _4432_ (.A1(net1062),
    .A2(_0995_),
    .Y(_1006_),
    .B1(net307));
 sg13g2_and2_1 _4433_ (.A(_2472_),
    .B(_0994_),
    .X(_1007_));
 sg13g2_nor3_1 _4434_ (.A(net908),
    .B(net308),
    .C(_1007_),
    .Y(_0081_));
 sg13g2_xnor2_1 _4435_ (.Y(_1008_),
    .A(net1061),
    .B(_1007_));
 sg13g2_nor2_1 _4436_ (.A(net908),
    .B(_1008_),
    .Y(_0082_));
 sg13g2_a21oi_1 _4437_ (.A1(net1061),
    .A2(_1007_),
    .Y(_1009_),
    .B1(net417));
 sg13g2_and3_1 _4438_ (.X(_1010_),
    .A(net1061),
    .B(\i_orchestrator.vga_x[8] ),
    .C(_1007_));
 sg13g2_nor3_1 _4439_ (.A(net908),
    .B(net418),
    .C(_1010_),
    .Y(_0083_));
 sg13g2_a21oi_1 _4440_ (.A1(net1060),
    .A2(_1010_),
    .Y(_1011_),
    .B1(net907));
 sg13g2_o21ai_1 _4441_ (.B1(_1011_),
    .Y(_1012_),
    .A1(net1060),
    .A2(_1010_));
 sg13g2_inv_1 _4442_ (.Y(_0084_),
    .A(_1012_));
 sg13g2_nor2_2 _4443_ (.A(_2399_),
    .B(\i_bitmap.in[5] ),
    .Y(_1013_));
 sg13g2_inv_1 _4444_ (.Y(_1014_),
    .A(_1013_));
 sg13g2_nor2_1 _4445_ (.A(\i_bitmap.in[4] ),
    .B(_1013_),
    .Y(_1015_));
 sg13g2_nor2b_1 _4446_ (.A(net1031),
    .B_N(\i_bitmap.in[5] ),
    .Y(_1016_));
 sg13g2_nand2_2 _4447_ (.Y(_1017_),
    .A(_2399_),
    .B(\i_bitmap.in[5] ));
 sg13g2_nand2_1 _4448_ (.Y(_1018_),
    .A(\i_bitmap.in[4] ),
    .B(_1017_));
 sg13g2_nor2b_1 _4449_ (.A(_1015_),
    .B_N(_1018_),
    .Y(_1019_));
 sg13g2_nand2b_2 _4450_ (.Y(_1020_),
    .B(_1018_),
    .A_N(_1015_));
 sg13g2_nor2_1 _4451_ (.A(\i_bitmap.in[3] ),
    .B(_1013_),
    .Y(_1021_));
 sg13g2_nand2_1 _4452_ (.Y(_1022_),
    .A(\i_bitmap.in[3] ),
    .B(_1017_));
 sg13g2_nor2b_2 _4453_ (.A(_1021_),
    .B_N(_1022_),
    .Y(_1023_));
 sg13g2_nand2b_2 _4454_ (.Y(_1024_),
    .B(_1022_),
    .A_N(_1021_));
 sg13g2_xor2_1 _4455_ (.B(\i_bitmap.in[2] ),
    .A(net1031),
    .X(_1025_));
 sg13g2_xnor2_1 _4456_ (.Y(_1026_),
    .A(net1031),
    .B(\i_bitmap.in[2] ));
 sg13g2_a21oi_1 _4457_ (.A1(_1014_),
    .A2(_1017_),
    .Y(_1027_),
    .B1(_1026_));
 sg13g2_o21ai_1 _4458_ (.B1(_1025_),
    .Y(_1028_),
    .A1(_1013_),
    .A2(_1016_));
 sg13g2_xor2_1 _4459_ (.B(\i_bitmap.in[0] ),
    .A(net1031),
    .X(_1029_));
 sg13g2_o21ai_1 _4460_ (.B1(_1029_),
    .Y(_1030_),
    .A1(_1013_),
    .A2(_1016_));
 sg13g2_nand2_1 _4461_ (.Y(_1031_),
    .A(\i_bitmap.in[1] ),
    .B(_1017_));
 sg13g2_o21ai_1 _4462_ (.B1(_1031_),
    .Y(_1032_),
    .A1(net1032),
    .A2(_1013_));
 sg13g2_and2_1 _4463_ (.A(_1030_),
    .B(_1032_),
    .X(_1033_));
 sg13g2_nand2_2 _4464_ (.Y(_1034_),
    .A(_1030_),
    .B(net915));
 sg13g2_a21oi_1 _4465_ (.A1(net916),
    .A2(_1034_),
    .Y(_1035_),
    .B1(_1023_));
 sg13g2_nor2_1 _4466_ (.A(_1020_),
    .B(_1035_),
    .Y(_1036_));
 sg13g2_nor2b_1 _4467_ (.A(net915),
    .B_N(_1029_),
    .Y(_1037_));
 sg13g2_nand2b_1 _4468_ (.Y(_1038_),
    .B(_1029_),
    .A_N(net915));
 sg13g2_nand3_1 _4469_ (.B(net916),
    .C(_1038_),
    .A(_1023_),
    .Y(_1039_));
 sg13g2_nand2_1 _4470_ (.Y(_1040_),
    .A(_1036_),
    .B(_1039_));
 sg13g2_xnor2_1 _4471_ (.Y(_1041_),
    .A(net1051),
    .B(\i_bitmap.in[10] ));
 sg13g2_a21oi_1 _4472_ (.A1(net916),
    .A2(_1029_),
    .Y(_1042_),
    .B1(_1024_));
 sg13g2_nand2_1 _4473_ (.Y(_1043_),
    .A(_1034_),
    .B(_1042_));
 sg13g2_xor2_1 _4474_ (.B(\i_capsule.tf_x[0] ),
    .A(net1031),
    .X(_1044_));
 sg13g2_o21ai_1 _4475_ (.B1(_1044_),
    .Y(_1045_),
    .A1(_1013_),
    .A2(_1016_));
 sg13g2_nor2_1 _4476_ (.A(_1038_),
    .B(_1045_),
    .Y(_1046_));
 sg13g2_nand3_1 _4477_ (.B(_1025_),
    .C(_1046_),
    .A(_1023_),
    .Y(_1047_));
 sg13g2_a22oi_1 _4478_ (.Y(_1048_),
    .B1(_1047_),
    .B2(_1020_),
    .A2(_1043_),
    .A1(_1036_));
 sg13g2_xor2_1 _4479_ (.B(\i_bitmap.in[9] ),
    .A(net1051),
    .X(_1049_));
 sg13g2_a21oi_1 _4480_ (.A1(net916),
    .A2(_1038_),
    .Y(_1050_),
    .B1(_1023_));
 sg13g2_nand2_1 _4481_ (.Y(_1051_),
    .A(_1030_),
    .B(_1045_));
 sg13g2_nand2b_2 _4482_ (.Y(_1052_),
    .B(_1051_),
    .A_N(net915));
 sg13g2_nand2_1 _4483_ (.Y(_1053_),
    .A(_1034_),
    .B(_1052_));
 sg13g2_nand3_1 _4484_ (.B(_1034_),
    .C(_1052_),
    .A(_1028_),
    .Y(_1054_));
 sg13g2_inv_1 _4485_ (.Y(_1055_),
    .A(_1054_));
 sg13g2_nor2_1 _4486_ (.A(_1024_),
    .B(_1055_),
    .Y(_1056_));
 sg13g2_nor2_1 _4487_ (.A(_1028_),
    .B(_1046_),
    .Y(_1057_));
 sg13g2_nand2_1 _4488_ (.Y(_1058_),
    .A(_1053_),
    .B(_1057_));
 sg13g2_a21oi_1 _4489_ (.A1(_1056_),
    .A2(_1058_),
    .Y(_1059_),
    .B1(_1050_));
 sg13g2_nor2_1 _4490_ (.A(net915),
    .B(_1044_),
    .Y(_1060_));
 sg13g2_nor3_1 _4491_ (.A(_1033_),
    .B(_1037_),
    .C(_1060_),
    .Y(_1061_));
 sg13g2_nor2_1 _4492_ (.A(net916),
    .B(_1061_),
    .Y(_1062_));
 sg13g2_nor2_1 _4493_ (.A(_1023_),
    .B(_1028_),
    .Y(_1063_));
 sg13g2_a21oi_1 _4494_ (.A1(_1027_),
    .A2(_1060_),
    .Y(_1064_),
    .B1(_1024_));
 sg13g2_nor2_1 _4495_ (.A(_1029_),
    .B(net915),
    .Y(_1065_));
 sg13g2_nor2_1 _4496_ (.A(_1045_),
    .B(_1065_),
    .Y(_1066_));
 sg13g2_o21ai_1 _4497_ (.B1(_1066_),
    .Y(_1067_),
    .A1(_1063_),
    .A2(_1064_));
 sg13g2_o21ai_1 _4498_ (.B1(_1028_),
    .Y(_1068_),
    .A1(net915),
    .A2(_1051_));
 sg13g2_a221oi_1 _4499_ (.B2(_1068_),
    .C1(_1020_),
    .B1(_1064_),
    .A1(_1024_),
    .Y(_1069_),
    .A2(_1062_));
 sg13g2_xor2_1 _4500_ (.B(\i_capsule.tf_y[0] ),
    .A(\i_capsule.tf_y[9] ),
    .X(_1070_));
 sg13g2_o21ai_1 _4501_ (.B1(_1070_),
    .Y(_1071_),
    .A1(_1019_),
    .A2(_1059_));
 sg13g2_a21oi_1 _4502_ (.A1(_1067_),
    .A2(_1069_),
    .Y(_1072_),
    .B1(_1071_));
 sg13g2_a21oi_1 _4503_ (.A1(net915),
    .A2(_1045_),
    .Y(_1073_),
    .B1(_1028_));
 sg13g2_and2_1 _4504_ (.A(_1052_),
    .B(_1073_),
    .X(_1074_));
 sg13g2_o21ai_1 _4505_ (.B1(_1023_),
    .Y(_1075_),
    .A1(_1062_),
    .A2(_1074_));
 sg13g2_a221oi_1 _4506_ (.B2(_1030_),
    .C1(_1020_),
    .B1(_1063_),
    .A1(_1024_),
    .Y(_1076_),
    .A2(_1055_));
 sg13g2_a21oi_1 _4507_ (.A1(net916),
    .A2(_1033_),
    .Y(_1077_),
    .B1(_1024_));
 sg13g2_o21ai_1 _4508_ (.B1(_1077_),
    .Y(_1078_),
    .A1(_1052_),
    .A2(_1057_));
 sg13g2_a21oi_1 _4509_ (.A1(_1037_),
    .A2(_1063_),
    .Y(_1079_),
    .B1(_1019_));
 sg13g2_a22oi_1 _4510_ (.Y(_1080_),
    .B1(_1078_),
    .B2(_1079_),
    .A2(_1076_),
    .A1(_1075_));
 sg13g2_xor2_1 _4511_ (.B(\i_bitmap.in[7] ),
    .A(\i_capsule.tf_y[9] ),
    .X(_1081_));
 sg13g2_a21oi_1 _4512_ (.A1(_1080_),
    .A2(_1081_),
    .Y(_1082_),
    .B1(_1072_));
 sg13g2_xor2_1 _4513_ (.B(\i_bitmap.in[8] ),
    .A(\i_capsule.tf_y[9] ),
    .X(_1083_));
 sg13g2_o21ai_1 _4514_ (.B1(net916),
    .Y(_1084_),
    .A1(_1033_),
    .A2(_1060_));
 sg13g2_a22oi_1 _4515_ (.Y(_1085_),
    .B1(_1084_),
    .B2(_1056_),
    .A2(_1063_),
    .A1(_1033_));
 sg13g2_a21oi_1 _4516_ (.A1(net916),
    .A2(_1046_),
    .Y(_1086_),
    .B1(_1019_));
 sg13g2_a22oi_1 _4517_ (.Y(_1087_),
    .B1(_1028_),
    .B2(_1052_),
    .A2(_1024_),
    .A1(_1020_));
 sg13g2_o21ai_1 _4518_ (.B1(_1087_),
    .Y(_1088_),
    .A1(_1050_),
    .A2(_1086_));
 sg13g2_o21ai_1 _4519_ (.B1(_1088_),
    .Y(_1089_),
    .A1(_1020_),
    .A2(_1085_));
 sg13g2_or2_1 _4520_ (.X(_1090_),
    .B(_1081_),
    .A(_1080_));
 sg13g2_o21ai_1 _4521_ (.B1(_1090_),
    .Y(_1091_),
    .A1(_1083_),
    .A2(_1089_));
 sg13g2_a22oi_1 _4522_ (.Y(_1092_),
    .B1(_1083_),
    .B2(_1089_),
    .A2(_1049_),
    .A1(_1048_));
 sg13g2_o21ai_1 _4523_ (.B1(_1092_),
    .Y(_1093_),
    .A1(_1082_),
    .A2(_1091_));
 sg13g2_o21ai_1 _4524_ (.B1(_1093_),
    .Y(_1094_),
    .A1(_1048_),
    .A2(_1049_));
 sg13g2_o21ai_1 _4525_ (.B1(_1094_),
    .Y(_1095_),
    .A1(_1040_),
    .A2(_1041_));
 sg13g2_nor3_1 _4526_ (.A(_1020_),
    .B(_1024_),
    .C(_1026_),
    .Y(_1096_));
 sg13g2_xor2_1 _4527_ (.B(\i_bitmap.in[11] ),
    .A(net1051),
    .X(_1097_));
 sg13g2_nor2_1 _4528_ (.A(_1096_),
    .B(_1097_),
    .Y(_1098_));
 sg13g2_a21oi_1 _4529_ (.A1(_1040_),
    .A2(_1041_),
    .Y(_1099_),
    .B1(_1098_));
 sg13g2_a21oi_1 _4530_ (.A1(\i_capsule.tf_x[8] ),
    .A2(\i_bitmap.in[6] ),
    .Y(_1100_),
    .B1(_2399_));
 sg13g2_a21oi_1 _4531_ (.A1(_2400_),
    .A2(_2401_),
    .Y(_1101_),
    .B1(net1031));
 sg13g2_nor2_1 _4532_ (.A(net1051),
    .B(\i_bitmap.in[12] ),
    .Y(_1102_));
 sg13g2_a21oi_2 _4533_ (.B1(_1102_),
    .Y(_1103_),
    .A2(\i_capsule.tf_y[7] ),
    .A1(\i_capsule.tf_y[8] ));
 sg13g2_a22oi_1 _4534_ (.Y(_1104_),
    .B1(\i_bitmap.in[12] ),
    .B2(net1051),
    .A2(_2417_),
    .A1(_2416_));
 sg13g2_or4_1 _4535_ (.A(_1100_),
    .B(_1101_),
    .C(_1103_),
    .D(_1104_),
    .X(_1105_));
 sg13g2_a221oi_1 _4536_ (.B2(_1095_),
    .C1(_1105_),
    .B1(_1099_),
    .A1(_1096_),
    .Y(_1106_),
    .A2(_1097_));
 sg13g2_nand2_1 _4537_ (.Y(_1107_),
    .A(net920),
    .B(_1106_));
 sg13g2_nor2b_1 _4538_ (.A(net6),
    .B_N(net415),
    .Y(_1108_));
 sg13g2_nand2b_2 _4539_ (.Y(_1109_),
    .B(net415),
    .A_N(net6));
 sg13g2_o21ai_1 _4540_ (.B1(_1108_),
    .Y(_1110_),
    .A1(_2386_),
    .A2(_2387_));
 sg13g2_o21ai_1 _4541_ (.B1(net413),
    .Y(_1111_),
    .A1(net329),
    .A2(_1109_));
 sg13g2_a21oi_1 _4542_ (.A1(_1110_),
    .A2(_1111_),
    .Y(_0085_),
    .B1(_1107_));
 sg13g2_nor2b_2 _4543_ (.A(net8),
    .B_N(handle_impact),
    .Y(_1112_));
 sg13g2_xnor2_1 _4544_ (.Y(_1113_),
    .A(net369),
    .B(net1020));
 sg13g2_o21ai_1 _4545_ (.B1(net1071),
    .Y(_1114_),
    .A1(net391),
    .A2(_1112_));
 sg13g2_a21oi_1 _4546_ (.A1(_1112_),
    .A2(_1113_),
    .Y(_0086_),
    .B1(_1114_));
 sg13g2_xnor2_1 _4547_ (.Y(_1115_),
    .A(net1062),
    .B(\i_orchestrator.vga_y[5] ));
 sg13g2_nor2_1 _4548_ (.A(net5),
    .B(_1115_),
    .Y(_1116_));
 sg13g2_nand3_1 _4549_ (.B(\capsule_color[3] ),
    .C(net1019),
    .A(\i_colors.capsule_color[4] ),
    .Y(_1117_));
 sg13g2_and2_1 _4550_ (.A(net358),
    .B(_1108_),
    .X(_1118_));
 sg13g2_a22oi_1 _4551_ (.Y(_1119_),
    .B1(_1117_),
    .B2(_1118_),
    .A2(_1109_),
    .A1(net393));
 sg13g2_o21ai_1 _4552_ (.B1(net920),
    .Y(_1120_),
    .A1(net868),
    .A2(_1116_));
 sg13g2_a21oi_1 _4553_ (.A1(net868),
    .A2(_1119_),
    .Y(_0087_),
    .B1(_1120_));
 sg13g2_nor4_2 _4554_ (.A(\i_orchestrator.vga_y[7] ),
    .B(\i_orchestrator.vga_y[6] ),
    .C(net1053),
    .Y(_1121_),
    .D(net1052));
 sg13g2_nor2_1 _4555_ (.A(\i_orchestrator.vga_y[8] ),
    .B(_2469_),
    .Y(_1122_));
 sg13g2_nand4_1 _4556_ (.B(_2468_),
    .C(_1121_),
    .A(\i_orchestrator.vga_y[9] ),
    .Y(_1123_),
    .D(_1122_));
 sg13g2_nand2_1 _4557_ (.Y(_1124_),
    .A(net1074),
    .B(_1123_));
 sg13g2_and3_1 _4558_ (.X(_1125_),
    .A(net1074),
    .B(_0998_),
    .C(_1123_));
 sg13g2_a22oi_1 _4559_ (.Y(_1126_),
    .B1(_1125_),
    .B2(net249),
    .A2(_0999_),
    .A1(\i_orchestrator.vga_y[0] ));
 sg13g2_inv_1 _4560_ (.Y(_0088_),
    .A(net250));
 sg13g2_nor2b_1 _4561_ (.A(net1058),
    .B_N(net1059),
    .Y(_1127_));
 sg13g2_xor2_1 _4562_ (.B(net1057),
    .A(net481),
    .X(_1128_));
 sg13g2_a22oi_1 _4563_ (.Y(_1129_),
    .B1(_1125_),
    .B2(_1128_),
    .A2(_0999_),
    .A1(net1057));
 sg13g2_inv_1 _4564_ (.Y(_0089_),
    .A(_1129_));
 sg13g2_nand3_1 _4565_ (.B(net1058),
    .C(net907),
    .A(net1059),
    .Y(_1130_));
 sg13g2_nand4_1 _4566_ (.B(net1057),
    .C(net1056),
    .A(net1059),
    .Y(_1131_),
    .D(net907));
 sg13g2_and2_2 _4567_ (.A(net907),
    .B(_1124_),
    .X(_1132_));
 sg13g2_xor2_1 _4568_ (.B(_1130_),
    .A(net1056),
    .X(_1133_));
 sg13g2_nor2_1 _4569_ (.A(_1132_),
    .B(_1133_),
    .Y(_0090_));
 sg13g2_and4_2 _4570_ (.A(net1059),
    .B(net1057),
    .C(net1056),
    .D(net1055),
    .X(_1134_));
 sg13g2_nor2_1 _4571_ (.A(_1124_),
    .B(_1134_),
    .Y(_1135_));
 sg13g2_a221oi_1 _4572_ (.B2(net907),
    .C1(_1132_),
    .B1(_1134_),
    .A1(_2423_),
    .Y(_0091_),
    .A2(_1131_));
 sg13g2_o21ai_1 _4573_ (.B1(net1054),
    .Y(_1136_),
    .A1(_0999_),
    .A2(_1135_));
 sg13g2_nand2_1 _4574_ (.Y(_1137_),
    .A(_1125_),
    .B(_1134_));
 sg13g2_o21ai_1 _4575_ (.B1(_1136_),
    .Y(_0092_),
    .A1(net1054),
    .A2(_1137_));
 sg13g2_and2_1 _4576_ (.A(net1053),
    .B(_1134_),
    .X(_1138_));
 sg13g2_a21oi_1 _4577_ (.A1(net907),
    .A2(_1138_),
    .Y(_1139_),
    .B1(net1052));
 sg13g2_and3_1 _4578_ (.X(_1140_),
    .A(net1052),
    .B(net907),
    .C(_1138_));
 sg13g2_nand3_1 _4579_ (.B(net907),
    .C(_1138_),
    .A(net1052),
    .Y(_1141_));
 sg13g2_nor3_1 _4580_ (.A(_1132_),
    .B(_1139_),
    .C(_1140_),
    .Y(_0093_));
 sg13g2_nand3b_1 _4581_ (.B(_1141_),
    .C(net428),
    .Y(_1142_),
    .A_N(_1132_));
 sg13g2_nand2b_1 _4582_ (.Y(_1143_),
    .B(net1052),
    .A_N(net428));
 sg13g2_nand3_1 _4583_ (.B(_1125_),
    .C(_1134_),
    .A(net1053),
    .Y(_1144_));
 sg13g2_o21ai_1 _4584_ (.B1(_1142_),
    .Y(_0094_),
    .A1(_1143_),
    .A2(_1144_));
 sg13g2_a21oi_1 _4585_ (.A1(\i_orchestrator.vga_y[6] ),
    .A2(_1140_),
    .Y(_1145_),
    .B1(net399));
 sg13g2_nor2_1 _4586_ (.A(_2458_),
    .B(_1141_),
    .Y(_1146_));
 sg13g2_nor3_1 _4587_ (.A(_1132_),
    .B(net400),
    .C(_1146_),
    .Y(_0095_));
 sg13g2_a21oi_1 _4588_ (.A1(net470),
    .A2(_1146_),
    .Y(_1147_),
    .B1(_1132_));
 sg13g2_o21ai_1 _4589_ (.B1(_1147_),
    .Y(_1148_),
    .A1(net470),
    .A2(_1146_));
 sg13g2_inv_1 _4590_ (.Y(_0096_),
    .A(_1148_));
 sg13g2_nand2_1 _4591_ (.Y(_1149_),
    .A(net382),
    .B(_1147_));
 sg13g2_o21ai_1 _4592_ (.B1(net383),
    .Y(_0097_),
    .A1(_2461_),
    .A2(_1144_));
 sg13g2_nor2_2 _4593_ (.A(net978),
    .B(_2822_),
    .Y(_1150_));
 sg13g2_or2_1 _4594_ (.X(_1151_),
    .B(net978),
    .A(_0057_));
 sg13g2_o21ai_1 _4595_ (.B1(_1151_),
    .Y(_1152_),
    .A1(\center_y[0] ),
    .A2(_2475_));
 sg13g2_nand2_1 _4596_ (.Y(_1153_),
    .A(net309),
    .B(_1150_));
 sg13g2_o21ai_1 _4597_ (.B1(_1153_),
    .Y(_0098_),
    .A1(_1150_),
    .A2(_1152_));
 sg13g2_nand2_1 _4598_ (.Y(_1154_),
    .A(net309),
    .B(\i_transform.track_y[1] ));
 sg13g2_nor2_1 _4599_ (.A(net978),
    .B(_2752_),
    .Y(_1155_));
 sg13g2_a22oi_1 _4600_ (.Y(_1156_),
    .B1(_1154_),
    .B2(_1155_),
    .A2(net977),
    .A1(net437));
 sg13g2_nand2_1 _4601_ (.Y(_1157_),
    .A(net445),
    .B(_1150_));
 sg13g2_o21ai_1 _4602_ (.B1(_1157_),
    .Y(_0099_),
    .A1(_1150_),
    .A2(_1156_));
 sg13g2_nor2_1 _4603_ (.A(net317),
    .B(net984),
    .Y(_1158_));
 sg13g2_nand3_1 _4604_ (.B(\i_transform.track_y[1] ),
    .C(_2822_),
    .A(\i_transform.track_y[0] ),
    .Y(_1159_));
 sg13g2_xor2_1 _4605_ (.B(_1159_),
    .A(\i_transform.track_y[2] ),
    .X(_1160_));
 sg13g2_a21oi_1 _4606_ (.A1(net984),
    .A2(_1160_),
    .Y(_0100_),
    .B1(_1158_));
 sg13g2_nand2_1 _4607_ (.Y(_1161_),
    .A(net297),
    .B(_1150_));
 sg13g2_nand3_1 _4608_ (.B(\i_transform.track_y[1] ),
    .C(\i_transform.track_y[2] ),
    .A(\i_transform.track_y[0] ),
    .Y(_1162_));
 sg13g2_nand2b_1 _4609_ (.Y(_1163_),
    .B(_1162_),
    .A_N(\i_transform.track_y[3] ));
 sg13g2_nand4_1 _4610_ (.B(\i_transform.track_y[1] ),
    .C(\i_transform.track_y[3] ),
    .A(\i_transform.track_y[0] ),
    .Y(_1164_),
    .D(\i_transform.track_y[2] ));
 sg13g2_a21o_1 _4611_ (.A2(_1164_),
    .A1(_1163_),
    .B1(net978),
    .X(_1165_));
 sg13g2_o21ai_1 _4612_ (.B1(_1165_),
    .Y(_1166_),
    .A1(\center_y[3] ),
    .A2(net984));
 sg13g2_o21ai_1 _4613_ (.B1(_1161_),
    .Y(_0101_),
    .A1(_1150_),
    .A2(_1166_));
 sg13g2_xnor2_1 _4614_ (.Y(_1167_),
    .A(net314),
    .B(_1164_));
 sg13g2_nand3_1 _4615_ (.B(_0838_),
    .C(_1167_),
    .A(net887),
    .Y(_1168_));
 sg13g2_a22oi_1 _4616_ (.Y(_1169_),
    .B1(_1150_),
    .B2(net314),
    .A2(net977),
    .A1(\center_y[4] ));
 sg13g2_nand2_1 _4617_ (.Y(_0102_),
    .A(_1168_),
    .B(net315));
 sg13g2_nand3_1 _4618_ (.B(_2587_),
    .C(_2588_),
    .A(_2568_),
    .Y(_1170_));
 sg13g2_a21oi_1 _4619_ (.A1(_2589_),
    .A2(_1170_),
    .Y(_1171_),
    .B1(net877));
 sg13g2_xor2_1 _4620_ (.B(net909),
    .A(_0033_),
    .X(_1172_));
 sg13g2_a21oi_1 _4621_ (.A1(net877),
    .A2(_1172_),
    .Y(_1173_),
    .B1(net884));
 sg13g2_nand2b_1 _4622_ (.Y(_1174_),
    .B(_1173_),
    .A_N(_1171_));
 sg13g2_or3_1 _4623_ (.A(_2720_),
    .B(_2737_),
    .C(_2738_),
    .X(_1175_));
 sg13g2_a21o_1 _4624_ (.A2(_1175_),
    .A1(_2739_),
    .B1(net891),
    .X(_1176_));
 sg13g2_xnor2_1 _4625_ (.Y(_1177_),
    .A(_0033_),
    .B(_2704_));
 sg13g2_a21oi_1 _4626_ (.A1(net891),
    .A2(_1177_),
    .Y(_1178_),
    .B1(net904));
 sg13g2_a22oi_1 _4627_ (.Y(_1179_),
    .B1(_1176_),
    .B2(_1178_),
    .A2(_2695_),
    .A1(net412));
 sg13g2_a21oi_1 _4628_ (.A1(_1174_),
    .A2(_1179_),
    .Y(_0103_),
    .B1(net976));
 sg13g2_nand3_1 _4629_ (.B(_2739_),
    .C(_2740_),
    .A(_2718_),
    .Y(_1180_));
 sg13g2_xor2_1 _4630_ (.B(_2763_),
    .A(_2762_),
    .X(_1181_));
 sg13g2_nor2b_1 _4631_ (.A(_2741_),
    .B_N(_1180_),
    .Y(_1182_));
 sg13g2_a21oi_1 _4632_ (.A1(net891),
    .A2(_1181_),
    .Y(_1183_),
    .B1(net903));
 sg13g2_o21ai_1 _4633_ (.B1(_1183_),
    .Y(_1184_),
    .A1(net891),
    .A2(_1182_));
 sg13g2_xor2_1 _4634_ (.B(_2683_),
    .A(_2682_),
    .X(_1185_));
 sg13g2_and3_1 _4635_ (.X(_1186_),
    .A(_2567_),
    .B(_2589_),
    .C(_2591_));
 sg13g2_o21ai_1 _4636_ (.B1(net874),
    .Y(_1187_),
    .A1(_2592_),
    .A2(_1186_));
 sg13g2_a21oi_1 _4637_ (.A1(net878),
    .A2(_1185_),
    .Y(_1188_),
    .B1(net884));
 sg13g2_a22oi_1 _4638_ (.Y(_1189_),
    .B1(_1187_),
    .B2(_1188_),
    .A2(net896),
    .A1(\i_capsule.tf_y[0] ));
 sg13g2_a21oi_1 _4639_ (.A1(_1184_),
    .A2(_1189_),
    .Y(_0104_),
    .B1(net976));
 sg13g2_o21ai_1 _4640_ (.B1(net984),
    .Y(_1190_),
    .A1(_0496_),
    .A2(_0501_));
 sg13g2_nand2_1 _4641_ (.Y(_1191_),
    .A(net548),
    .B(net882));
 sg13g2_nand2_1 _4642_ (.Y(_0105_),
    .A(_1190_),
    .B(_1191_));
 sg13g2_nand2_1 _4643_ (.Y(_1192_),
    .A(net527),
    .B(net896));
 sg13g2_a21oi_1 _4644_ (.A1(_2775_),
    .A2(_1192_),
    .Y(_0106_),
    .B1(net976));
 sg13g2_nand2_1 _4645_ (.Y(_1193_),
    .A(net529),
    .B(net896));
 sg13g2_a21oi_1 _4646_ (.A1(_0579_),
    .A2(_1193_),
    .Y(_0107_),
    .B1(net979));
 sg13g2_nand2_1 _4647_ (.Y(_1194_),
    .A(net482),
    .B(net896));
 sg13g2_a21oi_1 _4648_ (.A1(_0640_),
    .A2(_1194_),
    .Y(_0108_),
    .B1(net976));
 sg13g2_a22oi_1 _4649_ (.Y(_1195_),
    .B1(net882),
    .B2(net431),
    .A2(_0792_),
    .A1(net990));
 sg13g2_inv_1 _4650_ (.Y(_0109_),
    .A(_1195_));
 sg13g2_a21o_1 _4651_ (.A2(net882),
    .A1(net503),
    .B1(_0858_),
    .X(_0110_));
 sg13g2_xnor2_1 _4652_ (.Y(_1196_),
    .A(\i_capsule.tf_y[7] ),
    .B(net941));
 sg13g2_inv_1 _4653_ (.Y(_1197_),
    .A(_1196_));
 sg13g2_a21oi_1 _4654_ (.A1(_0833_),
    .A2(_0836_),
    .Y(_1198_),
    .B1(_0834_));
 sg13g2_nor2_1 _4655_ (.A(_1197_),
    .B(_1198_),
    .Y(_1199_));
 sg13g2_xnor2_1 _4656_ (.Y(_1200_),
    .A(_1197_),
    .B(_1198_));
 sg13g2_nor2_1 _4657_ (.A(_0040_),
    .B(net937),
    .Y(_1201_));
 sg13g2_nor2_1 _4658_ (.A(_0040_),
    .B(net940),
    .Y(_1202_));
 sg13g2_xnor2_1 _4659_ (.Y(_1203_),
    .A(_0040_),
    .B(net937));
 sg13g2_a21o_1 _4660_ (.A2(_0842_),
    .A1(_0835_),
    .B1(_1203_),
    .X(_1204_));
 sg13g2_nand3_1 _4661_ (.B(_0842_),
    .C(_1203_),
    .A(_0835_),
    .Y(_1205_));
 sg13g2_nand3_1 _4662_ (.B(_1204_),
    .C(_1205_),
    .A(net893),
    .Y(_1206_));
 sg13g2_o21ai_1 _4663_ (.B1(_1206_),
    .Y(_1207_),
    .A1(net893),
    .A2(_1200_));
 sg13g2_a22oi_1 _4664_ (.Y(_1208_),
    .B1(_1207_),
    .B2(_0838_),
    .A2(_0859_),
    .A1(net501));
 sg13g2_a21oi_1 _4665_ (.A1(_2443_),
    .A2(net968),
    .Y(_1209_),
    .B1(_0853_));
 sg13g2_xnor2_1 _4666_ (.Y(_1210_),
    .A(_0040_),
    .B(net972));
 sg13g2_or2_1 _4667_ (.X(_1211_),
    .B(_1210_),
    .A(_1209_));
 sg13g2_a21oi_1 _4668_ (.A1(_1209_),
    .A2(_1210_),
    .Y(_1212_),
    .B1(net880));
 sg13g2_o21ai_1 _4669_ (.B1(_0038_),
    .Y(_1213_),
    .A1(\i_bitmap.in[12] ),
    .A2(_2418_));
 sg13g2_a22oi_1 _4670_ (.Y(_1214_),
    .B1(_1213_),
    .B2(net972),
    .A2(_0848_),
    .A1(_0784_));
 sg13g2_nand2_1 _4671_ (.Y(_1215_),
    .A(\i_capsule.tf_y[7] ),
    .B(net968));
 sg13g2_xnor2_1 _4672_ (.Y(_1216_),
    .A(\i_capsule.tf_y[7] ),
    .B(net973));
 sg13g2_or2_1 _4673_ (.X(_1217_),
    .B(_1216_),
    .A(_1214_));
 sg13g2_a21oi_1 _4674_ (.A1(_1214_),
    .A2(_1216_),
    .Y(_1218_),
    .B1(net876));
 sg13g2_a22oi_1 _4675_ (.Y(_1219_),
    .B1(_1217_),
    .B2(_1218_),
    .A2(_1212_),
    .A1(_1211_));
 sg13g2_o21ai_1 _4676_ (.B1(_1208_),
    .Y(_0111_),
    .A1(_0857_),
    .A2(_1219_));
 sg13g2_nor2_1 _4677_ (.A(_0041_),
    .B(net968),
    .Y(_1220_));
 sg13g2_xnor2_1 _4678_ (.Y(_1221_),
    .A(_0041_),
    .B(net973));
 sg13g2_a21oi_1 _4679_ (.A1(_1211_),
    .A2(_1215_),
    .Y(_1222_),
    .B1(_1221_));
 sg13g2_nand3_1 _4680_ (.B(_1215_),
    .C(_1221_),
    .A(_1211_),
    .Y(_1223_));
 sg13g2_nor2b_1 _4681_ (.A(_1222_),
    .B_N(_1223_),
    .Y(_1224_));
 sg13g2_xnor2_1 _4682_ (.Y(_1225_),
    .A(_2416_),
    .B(net973));
 sg13g2_o21ai_1 _4683_ (.B1(_1217_),
    .Y(_1226_),
    .A1(_2417_),
    .A2(net968));
 sg13g2_o21ai_1 _4684_ (.B1(net880),
    .Y(_1227_),
    .A1(_1225_),
    .A2(_1226_));
 sg13g2_a21oi_1 _4685_ (.A1(_1225_),
    .A2(_1226_),
    .Y(_1228_),
    .B1(_1227_));
 sg13g2_a21oi_1 _4686_ (.A1(net876),
    .A2(_1224_),
    .Y(_1229_),
    .B1(_1228_));
 sg13g2_xnor2_1 _4687_ (.Y(_1230_),
    .A(_0041_),
    .B(net940));
 sg13g2_nand2b_1 _4688_ (.Y(_1231_),
    .B(_1204_),
    .A_N(_1201_));
 sg13g2_a21oi_1 _4689_ (.A1(_1230_),
    .A2(_1231_),
    .Y(_1232_),
    .B1(net889));
 sg13g2_o21ai_1 _4690_ (.B1(_1232_),
    .Y(_1233_),
    .A1(_1230_),
    .A2(_1231_));
 sg13g2_xnor2_1 _4691_ (.Y(_1234_),
    .A(\i_capsule.tf_y[8] ),
    .B(net940));
 sg13g2_nor3_1 _4692_ (.A(_1199_),
    .B(_1202_),
    .C(_1234_),
    .Y(_1235_));
 sg13g2_o21ai_1 _4693_ (.B1(_1234_),
    .Y(_1236_),
    .A1(_1199_),
    .A2(_1202_));
 sg13g2_nand2_1 _4694_ (.Y(_1237_),
    .A(net889),
    .B(_1236_));
 sg13g2_o21ai_1 _4695_ (.B1(_1233_),
    .Y(_1238_),
    .A1(_1235_),
    .A2(_1237_));
 sg13g2_a22oi_1 _4696_ (.Y(_1239_),
    .B1(_1238_),
    .B2(_0838_),
    .A2(_0859_),
    .A1(net498));
 sg13g2_o21ai_1 _4697_ (.B1(_1239_),
    .Y(_0112_),
    .A1(net883),
    .A2(_1229_));
 sg13g2_a21oi_1 _4698_ (.A1(\i_capsule.tf_y[8] ),
    .A2(net968),
    .Y(_1240_),
    .B1(_1222_));
 sg13g2_xnor2_1 _4699_ (.Y(_1241_),
    .A(_0042_),
    .B(net969));
 sg13g2_xnor2_1 _4700_ (.Y(_1242_),
    .A(_1240_),
    .B(_1241_));
 sg13g2_nor2b_1 _4701_ (.A(_1217_),
    .B_N(_1225_),
    .Y(_1243_));
 sg13g2_nor3_1 _4702_ (.A(\i_capsule.tf_y[8] ),
    .B(_2417_),
    .C(net968),
    .Y(_1244_));
 sg13g2_nor3_1 _4703_ (.A(_1220_),
    .B(_1243_),
    .C(_1244_),
    .Y(_1245_));
 sg13g2_xnor2_1 _4704_ (.Y(_1246_),
    .A(net1051),
    .B(net973));
 sg13g2_or2_1 _4705_ (.X(_1247_),
    .B(_1246_),
    .A(_1245_));
 sg13g2_a21oi_1 _4706_ (.A1(_1245_),
    .A2(_1246_),
    .Y(_1248_),
    .B1(net876));
 sg13g2_a221oi_1 _4707_ (.B2(_1248_),
    .C1(net885),
    .B1(_1247_),
    .A1(net876),
    .Y(_1249_),
    .A2(_1242_));
 sg13g2_o21ai_1 _4708_ (.B1(_1236_),
    .Y(_1250_),
    .A1(_0041_),
    .A2(net940));
 sg13g2_xnor2_1 _4709_ (.Y(_1251_),
    .A(net1051),
    .B(net937));
 sg13g2_xnor2_1 _4710_ (.Y(_1252_),
    .A(_1250_),
    .B(_1251_));
 sg13g2_nor2b_1 _4711_ (.A(_1204_),
    .B_N(_1230_),
    .Y(_1253_));
 sg13g2_a221oi_1 _4712_ (.B2(_0041_),
    .C1(_1253_),
    .B1(_1201_),
    .A1(\i_capsule.tf_y[8] ),
    .Y(_1254_),
    .A2(net940));
 sg13g2_xnor2_1 _4713_ (.Y(_1255_),
    .A(_0042_),
    .B(net937));
 sg13g2_or2_1 _4714_ (.X(_1256_),
    .B(_1255_),
    .A(_1254_));
 sg13g2_a21oi_1 _4715_ (.A1(_1254_),
    .A2(_1255_),
    .Y(_1257_),
    .B1(net889));
 sg13g2_a221oi_1 _4716_ (.B2(_1257_),
    .C1(net906),
    .B1(_1256_),
    .A1(net889),
    .Y(_1258_),
    .A2(_1252_));
 sg13g2_o21ai_1 _4717_ (.B1(net990),
    .Y(_1259_),
    .A1(net1051),
    .A2(net895));
 sg13g2_nor3_1 _4718_ (.A(_1249_),
    .B(_1258_),
    .C(_1259_),
    .Y(_0113_));
 sg13g2_nor4_1 _4719_ (.A(\i_orchestrator.vga_x[3] ),
    .B(net1061),
    .C(net1060),
    .D(\i_orchestrator.vga_x[8] ),
    .Y(_1260_));
 sg13g2_nand4_1 _4720_ (.B(_2473_),
    .C(_1001_),
    .A(_2421_),
    .Y(_1261_),
    .D(_1260_));
 sg13g2_nor3_2 _4721_ (.A(net1053),
    .B(_2461_),
    .C(_1261_),
    .Y(_1262_));
 sg13g2_nand4_1 _4722_ (.B(_2423_),
    .C(_1127_),
    .A(net1056),
    .Y(_1263_),
    .D(_1262_));
 sg13g2_nor2_1 _4723_ (.A(net381),
    .B(net338),
    .Y(_1264_));
 sg13g2_nor2_1 _4724_ (.A(\i_orchestrator.hit_left ),
    .B(\i_orchestrator.hit_bottom ),
    .Y(_1265_));
 sg13g2_nand3_1 _4725_ (.B(_0055_),
    .C(_1265_),
    .A(_2405_),
    .Y(_1266_));
 sg13g2_nor2_1 _4726_ (.A(_1263_),
    .B(_1266_),
    .Y(_1267_));
 sg13g2_nor2_2 _4727_ (.A(\collision_impact[1] ),
    .B(\collision_impact[0] ),
    .Y(_1268_));
 sg13g2_nor2_1 _4728_ (.A(_1263_),
    .B(_1268_),
    .Y(_1269_));
 sg13g2_nor2_1 _4729_ (.A(net426),
    .B(_1269_),
    .Y(_1270_));
 sg13g2_nor3_1 _4730_ (.A(net1069),
    .B(_1267_),
    .C(_1270_),
    .Y(_0114_));
 sg13g2_nor4_2 _4731_ (.A(net1059),
    .B(net1058),
    .C(net1056),
    .Y(_1271_),
    .D(net1055));
 sg13g2_and2_1 _4732_ (.A(_1262_),
    .B(_1271_),
    .X(_1272_));
 sg13g2_nand2_1 _4733_ (.Y(_1273_),
    .A(_1262_),
    .B(_1271_));
 sg13g2_o21ai_1 _4734_ (.B1(net1074),
    .Y(_1274_),
    .A1(\i_orchestrator.hit_priority[0] ),
    .A2(net914));
 sg13g2_a21oi_1 _4735_ (.A1(_2415_),
    .A2(net914),
    .Y(_0115_),
    .B1(_1274_));
 sg13g2_a21oi_1 _4736_ (.A1(\i_orchestrator.hit_priority[0] ),
    .A2(net914),
    .Y(_1275_),
    .B1(net348));
 sg13g2_and3_1 _4737_ (.X(_1276_),
    .A(net348),
    .B(\i_orchestrator.hit_priority[0] ),
    .C(net914));
 sg13g2_nor3_1 _4738_ (.A(net1069),
    .B(net349),
    .C(_1276_),
    .Y(_0116_));
 sg13g2_xor2_1 _4739_ (.B(\i_orchestrator.lfsr[6] ),
    .A(\color_entropy[1] ),
    .X(_1277_));
 sg13g2_a21oi_1 _4740_ (.A1(net914),
    .A2(_1277_),
    .Y(_1278_),
    .B1(net1068));
 sg13g2_o21ai_1 _4741_ (.B1(_1278_),
    .Y(_0117_),
    .A1(_2414_),
    .A2(net914));
 sg13g2_a21oi_1 _4742_ (.A1(net271),
    .A2(_1273_),
    .Y(_1279_),
    .B1(net1069));
 sg13g2_o21ai_1 _4743_ (.B1(_1279_),
    .Y(_0118_),
    .A1(_2414_),
    .A2(_1273_));
 sg13g2_a21oi_1 _4744_ (.A1(net271),
    .A2(net914),
    .Y(_1280_),
    .B1(net1067));
 sg13g2_o21ai_1 _4745_ (.B1(_1280_),
    .Y(_0119_),
    .A1(_2413_),
    .A2(net914));
 sg13g2_a21oi_1 _4746_ (.A1(net270),
    .A2(net912),
    .Y(_1281_),
    .B1(net1067));
 sg13g2_o21ai_1 _4747_ (.B1(_1281_),
    .Y(_0120_),
    .A1(_2412_),
    .A2(net912));
 sg13g2_a21oi_1 _4748_ (.A1(net266),
    .A2(net913),
    .Y(_1282_),
    .B1(net1067));
 sg13g2_o21ai_1 _4749_ (.B1(_1282_),
    .Y(_0121_),
    .A1(_2411_),
    .A2(net912));
 sg13g2_a21oi_1 _4750_ (.A1(\i_orchestrator.lfsr[4] ),
    .A2(net912),
    .Y(_1283_),
    .B1(net1066));
 sg13g2_o21ai_1 _4751_ (.B1(_1283_),
    .Y(_0122_),
    .A1(_2410_),
    .A2(net912));
 sg13g2_a21oi_1 _4752_ (.A1(net268),
    .A2(net912),
    .Y(_1284_),
    .B1(net1067));
 sg13g2_o21ai_1 _4753_ (.B1(_1284_),
    .Y(_0123_),
    .A1(_2409_),
    .A2(net912));
 sg13g2_a21oi_1 _4754_ (.A1(\i_orchestrator.lfsr[6] ),
    .A2(net912),
    .Y(_1285_),
    .B1(net1066));
 sg13g2_o21ai_1 _4755_ (.B1(_1285_),
    .Y(_0124_),
    .A1(_2408_),
    .A2(net913));
 sg13g2_a21oi_1 _4756_ (.A1(net279),
    .A2(net913),
    .Y(_1286_),
    .B1(net1066));
 sg13g2_o21ai_1 _4757_ (.B1(_1286_),
    .Y(_0125_),
    .A1(_2407_),
    .A2(net913));
 sg13g2_nand2_2 _4758_ (.Y(_1287_),
    .A(net1077),
    .B(net913));
 sg13g2_a22oi_1 _4759_ (.Y(_1288_),
    .B1(_1287_),
    .B2(_2449_),
    .A2(net913),
    .A1(net295));
 sg13g2_inv_1 _4760_ (.Y(_0126_),
    .A(_1288_));
 sg13g2_and2_1 _4761_ (.A(_1134_),
    .B(_1262_),
    .X(_1289_));
 sg13g2_nand2b_1 _4762_ (.Y(_1290_),
    .B(net1074),
    .A_N(_1289_));
 sg13g2_nand3_1 _4763_ (.B(net919),
    .C(_1007_),
    .A(\i_orchestrator.vga_x[9] ),
    .Y(_1291_));
 sg13g2_nand2b_1 _4764_ (.Y(_1292_),
    .B(_1291_),
    .A_N(_1289_));
 sg13g2_or2_1 _4765_ (.X(_1293_),
    .B(_1292_),
    .A(net868));
 sg13g2_nand2b_1 _4766_ (.Y(_1294_),
    .B(net928),
    .A_N(_1261_));
 sg13g2_nand2b_1 _4767_ (.Y(_1295_),
    .B(_1294_),
    .A_N(_1292_));
 sg13g2_nor3_1 _4768_ (.A(_2422_),
    .B(net1052),
    .C(_2458_),
    .Y(_1296_));
 sg13g2_nand4_1 _4769_ (.B(_2599_),
    .C(_1134_),
    .A(_2460_),
    .Y(_1297_),
    .D(_1296_));
 sg13g2_nand2b_1 _4770_ (.Y(_1298_),
    .B(_1297_),
    .A_N(_1295_));
 sg13g2_nand4_1 _4771_ (.B(_1293_),
    .C(_1294_),
    .A(_1291_),
    .Y(_1299_),
    .D(_1298_));
 sg13g2_a21oi_1 _4772_ (.A1(_2406_),
    .A2(_1299_),
    .Y(_0127_),
    .B1(_1290_));
 sg13g2_nand4_1 _4773_ (.B(_2599_),
    .C(_1121_),
    .A(_2464_),
    .Y(_1300_),
    .D(_1271_));
 sg13g2_or3_1 _4774_ (.A(net868),
    .B(_1298_),
    .C(_1300_),
    .X(_1301_));
 sg13g2_nand2b_1 _4775_ (.Y(_1302_),
    .B(_1300_),
    .A_N(_1292_));
 sg13g2_or2_1 _4776_ (.X(_1303_),
    .B(_1261_),
    .A(_2463_));
 sg13g2_and4_1 _4777_ (.A(_1263_),
    .B(_1273_),
    .C(_1291_),
    .D(_1303_),
    .X(_1304_));
 sg13g2_nand4_1 _4778_ (.B(_1301_),
    .C(_1302_),
    .A(_1294_),
    .Y(_1305_),
    .D(_1304_));
 sg13g2_a21oi_1 _4779_ (.A1(_2405_),
    .A2(_1305_),
    .Y(_0128_),
    .B1(_1290_));
 sg13g2_a21oi_1 _4780_ (.A1(net868),
    .A2(_1292_),
    .Y(_1306_),
    .B1(net322));
 sg13g2_nor2_1 _4781_ (.A(_1290_),
    .B(_1306_),
    .Y(_0129_));
 sg13g2_nand3_1 _4782_ (.B(_1295_),
    .C(_1304_),
    .A(_1293_),
    .Y(_1307_));
 sg13g2_a21oi_1 _4783_ (.A1(_2404_),
    .A2(_1307_),
    .Y(_0130_),
    .B1(_1290_));
 sg13g2_nand4_1 _4784_ (.B(net283),
    .C(_1266_),
    .A(net1074),
    .Y(_1308_),
    .D(_1269_));
 sg13g2_inv_1 _4785_ (.Y(_0131_),
    .A(net284));
 sg13g2_nor4_1 _4786_ (.A(\i_orchestrator.sample_counter[2] ),
    .B(\i_orchestrator.sample_counter[5] ),
    .C(\i_orchestrator.sample_counter[4] ),
    .D(\i_orchestrator.sample_counter[7] ),
    .Y(_1309_));
 sg13g2_nor2_1 _4787_ (.A(net373),
    .B(\i_orchestrator.sample_counter[1] ),
    .Y(_1310_));
 sg13g2_nand4_1 _4788_ (.B(_2435_),
    .C(_1309_),
    .A(net1076),
    .Y(_1311_),
    .D(_1310_));
 sg13g2_nor4_2 _4789_ (.A(\i_orchestrator.sample_counter[6] ),
    .B(net242),
    .C(\i_orchestrator.sample_counter[8] ),
    .Y(_0132_),
    .D(_1311_));
 sg13g2_and2_1 _4790_ (.A(net1074),
    .B(_1289_),
    .X(_0133_));
 sg13g2_nor3_1 _4791_ (.A(net1069),
    .B(net1),
    .C(_1303_),
    .Y(_0134_));
 sg13g2_o21ai_1 _4792_ (.B1(net245),
    .Y(_1312_),
    .A1(_2404_),
    .A2(\i_orchestrator.hit_right ));
 sg13g2_a21o_1 _4793_ (.A2(_1312_),
    .A1(net247),
    .B1(net348),
    .X(_1313_));
 sg13g2_nand2_1 _4794_ (.Y(_1314_),
    .A(\i_orchestrator.hit_left ),
    .B(_2406_));
 sg13g2_nor2b_1 _4795_ (.A(\i_orchestrator.hit_top ),
    .B_N(\i_orchestrator.hit_priority[1] ),
    .Y(_1315_));
 sg13g2_a21oi_1 _4796_ (.A1(_1314_),
    .A2(_1315_),
    .Y(_1316_),
    .B1(\i_orchestrator.hit_priority[0] ));
 sg13g2_a21o_1 _4797_ (.A2(\i_orchestrator.hit_priority[1] ),
    .A1(\i_orchestrator.hit_right ),
    .B1(_2405_),
    .X(_1317_));
 sg13g2_nand2_1 _4798_ (.Y(_1318_),
    .A(\i_orchestrator.hit_bottom ),
    .B(net353));
 sg13g2_a21oi_1 _4799_ (.A1(_0055_),
    .A2(_1318_),
    .Y(_1319_),
    .B1(net348));
 sg13g2_a21oi_1 _4800_ (.A1(net353),
    .A2(_1317_),
    .Y(_1320_),
    .B1(_1319_));
 sg13g2_a22oi_1 _4801_ (.Y(_1321_),
    .B1(net354),
    .B2(\i_orchestrator.hit_priority[0] ),
    .A2(_1316_),
    .A1(_1313_));
 sg13g2_nor2_1 _4802_ (.A(_1287_),
    .B(net355),
    .Y(_0135_));
 sg13g2_nor2_1 _4803_ (.A(net365),
    .B(net322),
    .Y(_1322_));
 sg13g2_nor2_1 _4804_ (.A(net476),
    .B(_1264_),
    .Y(_1323_));
 sg13g2_nor3_1 _4805_ (.A(_1287_),
    .B(_1322_),
    .C(_1323_),
    .Y(_0136_));
 sg13g2_nor3_1 _4806_ (.A(\i_orchestrator.hit_left ),
    .B(\i_orchestrator.hit_right ),
    .C(\i_orchestrator.hit_bottom ),
    .Y(_1324_));
 sg13g2_a21oi_1 _4807_ (.A1(net245),
    .A2(_1324_),
    .Y(_0137_),
    .B1(_1287_));
 sg13g2_or2_1 _4808_ (.X(_1325_),
    .B(net434),
    .A(net356));
 sg13g2_nand2_1 _4809_ (.Y(_1326_),
    .A(net356),
    .B(net434));
 sg13g2_and3_1 _4810_ (.X(_0138_),
    .A(net1073),
    .B(_1325_),
    .C(_1326_));
 sg13g2_xnor2_1 _4811_ (.Y(_1327_),
    .A(net552),
    .B(net475));
 sg13g2_and2_1 _4812_ (.A(_1326_),
    .B(_1327_),
    .X(_1328_));
 sg13g2_nor2_1 _4813_ (.A(_1326_),
    .B(_1327_),
    .Y(_1329_));
 sg13g2_nor3_1 _4814_ (.A(net1070),
    .B(_1328_),
    .C(_1329_),
    .Y(_0139_));
 sg13g2_xnor2_1 _4815_ (.Y(_1330_),
    .A(net438),
    .B(net530));
 sg13g2_a21oi_1 _4816_ (.A1(net490),
    .A2(net475),
    .Y(_1331_),
    .B1(_1329_));
 sg13g2_and2_1 _4817_ (.A(_1330_),
    .B(_1331_),
    .X(_1332_));
 sg13g2_nor2_1 _4818_ (.A(_1330_),
    .B(_1331_),
    .Y(_1333_));
 sg13g2_nor3_1 _4819_ (.A(net1070),
    .B(_1332_),
    .C(_1333_),
    .Y(_0140_));
 sg13g2_nand2_1 _4820_ (.Y(_1334_),
    .A(\i_delta_sigma.sample[3] ),
    .B(\i_delta_sigma.acc[3] ));
 sg13g2_xnor2_1 _4821_ (.Y(_1335_),
    .A(\i_delta_sigma.sample[3] ),
    .B(net409));
 sg13g2_a21oi_1 _4822_ (.A1(\i_delta_sigma.sample[2] ),
    .A2(\i_delta_sigma.acc[2] ),
    .Y(_1336_),
    .B1(_1333_));
 sg13g2_or2_1 _4823_ (.X(_1337_),
    .B(_1336_),
    .A(_1335_));
 sg13g2_nand2_1 _4824_ (.Y(_1338_),
    .A(net1071),
    .B(_1337_));
 sg13g2_a21oi_1 _4825_ (.A1(net410),
    .A2(_1336_),
    .Y(_0141_),
    .B1(_1338_));
 sg13g2_nand2_1 _4826_ (.Y(_1339_),
    .A(\i_delta_sigma.sample[4] ),
    .B(net366));
 sg13g2_xnor2_1 _4827_ (.Y(_1340_),
    .A(\i_delta_sigma.sample[4] ),
    .B(net366));
 sg13g2_and2_1 _4828_ (.A(_1334_),
    .B(_1337_),
    .X(_1341_));
 sg13g2_or2_1 _4829_ (.X(_1342_),
    .B(_1341_),
    .A(_1340_));
 sg13g2_nand2_1 _4830_ (.Y(_1343_),
    .A(net1072),
    .B(_1342_));
 sg13g2_a21oi_1 _4831_ (.A1(net367),
    .A2(_1341_),
    .Y(_0142_),
    .B1(_1343_));
 sg13g2_and2_1 _4832_ (.A(_1339_),
    .B(_1342_),
    .X(_1344_));
 sg13g2_nor2_1 _4833_ (.A(\i_delta_sigma.sample[5] ),
    .B(net496),
    .Y(_1345_));
 sg13g2_nand2_1 _4834_ (.Y(_1346_),
    .A(\i_delta_sigma.sample[5] ),
    .B(net496));
 sg13g2_nand2b_1 _4835_ (.Y(_1347_),
    .B(_1346_),
    .A_N(_1345_));
 sg13g2_o21ai_1 _4836_ (.B1(net1072),
    .Y(_1348_),
    .A1(_1344_),
    .A2(_1347_));
 sg13g2_a21oi_1 _4837_ (.A1(_1344_),
    .A2(_1347_),
    .Y(_0143_),
    .B1(_1348_));
 sg13g2_xor2_1 _4838_ (.B(net520),
    .A(\i_delta_sigma.sample[6] ),
    .X(_1349_));
 sg13g2_o21ai_1 _4839_ (.B1(_1346_),
    .Y(_1350_),
    .A1(_1344_),
    .A2(_1345_));
 sg13g2_and2_1 _4840_ (.A(_1349_),
    .B(_1350_),
    .X(_1351_));
 sg13g2_o21ai_1 _4841_ (.B1(net1072),
    .Y(_1352_),
    .A1(_1349_),
    .A2(_1350_));
 sg13g2_nor2_1 _4842_ (.A(_1351_),
    .B(_1352_),
    .Y(_0144_));
 sg13g2_a21oi_1 _4843_ (.A1(\i_delta_sigma.sample[6] ),
    .A2(\i_delta_sigma.acc[6] ),
    .Y(_1353_),
    .B1(_1351_));
 sg13g2_xnor2_1 _4844_ (.Y(_1354_),
    .A(\i_delta_sigma.sample[7] ),
    .B(net505));
 sg13g2_nor2_1 _4845_ (.A(_1353_),
    .B(_1354_),
    .Y(_1355_));
 sg13g2_a21oi_1 _4846_ (.A1(_1353_),
    .A2(_1354_),
    .Y(_1356_),
    .B1(net1070));
 sg13g2_nor2b_1 _4847_ (.A(net506),
    .B_N(_1356_),
    .Y(_0145_));
 sg13g2_a21oi_1 _4848_ (.A1(\i_delta_sigma.sample[7] ),
    .A2(\i_delta_sigma.acc[7] ),
    .Y(_1357_),
    .B1(_1355_));
 sg13g2_xnor2_1 _4849_ (.Y(_1358_),
    .A(\i_delta_sigma.sample[8] ),
    .B(net378));
 sg13g2_or2_1 _4850_ (.X(_1359_),
    .B(_1358_),
    .A(_1357_));
 sg13g2_nand2_1 _4851_ (.Y(_1360_),
    .A(net1072),
    .B(_1359_));
 sg13g2_a21oi_1 _4852_ (.A1(_1357_),
    .A2(net379),
    .Y(_0146_),
    .B1(_1360_));
 sg13g2_o21ai_1 _4853_ (.B1(_1359_),
    .Y(_1361_),
    .A1(_2381_),
    .A2(_2420_));
 sg13g2_nor2_1 _4854_ (.A(net1014),
    .B(net473),
    .Y(_1362_));
 sg13g2_xor2_1 _4855_ (.B(net473),
    .A(\i_delta_sigma.sample[9] ),
    .X(_1363_));
 sg13g2_o21ai_1 _4856_ (.B1(net1073),
    .Y(_1364_),
    .A1(_1361_),
    .A2(net474));
 sg13g2_a21oi_1 _4857_ (.A1(_1361_),
    .A2(net474),
    .Y(_0147_),
    .B1(_1364_));
 sg13g2_xor2_1 _4858_ (.B(net531),
    .A(net1013),
    .X(_1365_));
 sg13g2_a21oi_1 _4859_ (.A1(net1014),
    .A2(net473),
    .Y(_1366_),
    .B1(_1361_));
 sg13g2_nor2_1 _4860_ (.A(_1362_),
    .B(_1366_),
    .Y(_1367_));
 sg13g2_nand2_1 _4861_ (.Y(_1368_),
    .A(_1365_),
    .B(_1367_));
 sg13g2_o21ai_1 _4862_ (.B1(net1073),
    .Y(_1369_),
    .A1(_1365_),
    .A2(_1367_));
 sg13g2_nor2b_1 _4863_ (.A(_1369_),
    .B_N(_1368_),
    .Y(_0148_));
 sg13g2_xor2_1 _4864_ (.B(\i_delta_sigma.acc[11] ),
    .A(net1018),
    .X(_1370_));
 sg13g2_o21ai_1 _4865_ (.B1(_1368_),
    .Y(_1371_),
    .A1(_2380_),
    .A2(_2419_));
 sg13g2_xnor2_1 _4866_ (.Y(_1372_),
    .A(_1370_),
    .B(_1371_));
 sg13g2_and2_1 _4867_ (.A(net1077),
    .B(_1372_),
    .X(_0149_));
 sg13g2_xnor2_1 _4868_ (.Y(_1373_),
    .A(net1018),
    .B(\i_delta_sigma.acc[12] ));
 sg13g2_a21o_1 _4869_ (.A2(\i_delta_sigma.acc[11] ),
    .A1(net1018),
    .B1(_1371_),
    .X(_1374_));
 sg13g2_o21ai_1 _4870_ (.B1(_1374_),
    .Y(_1375_),
    .A1(net1018),
    .A2(\i_delta_sigma.acc[11] ));
 sg13g2_xor2_1 _4871_ (.B(_1375_),
    .A(_1373_),
    .X(_1376_));
 sg13g2_inv_1 _4872_ (.Y(_1377_),
    .A(_1376_));
 sg13g2_xnor2_1 _4873_ (.Y(_1378_),
    .A(net364),
    .B(_1376_));
 sg13g2_or2_1 _4874_ (.X(_1379_),
    .B(_1378_),
    .A(_1372_));
 sg13g2_nand2_1 _4875_ (.Y(_1380_),
    .A(net1077),
    .B(_1379_));
 sg13g2_a21oi_1 _4876_ (.A1(_1372_),
    .A2(_1378_),
    .Y(_0150_),
    .B1(_1380_));
 sg13g2_o21ai_1 _4877_ (.B1(_1379_),
    .Y(_1381_),
    .A1(net524),
    .A2(_1377_));
 sg13g2_xor2_1 _4878_ (.B(_0054_),
    .A(\i_delta_sigma.acc[13] ),
    .X(_1382_));
 sg13g2_nand2_1 _4879_ (.Y(_1383_),
    .A(net1018),
    .B(\i_delta_sigma.acc[12] ));
 sg13g2_o21ai_1 _4880_ (.B1(_1383_),
    .Y(_1384_),
    .A1(_1373_),
    .A2(_1375_));
 sg13g2_xnor2_1 _4881_ (.Y(_1385_),
    .A(net1018),
    .B(_1382_));
 sg13g2_xnor2_1 _4882_ (.Y(_1386_),
    .A(_1384_),
    .B(_1385_));
 sg13g2_o21ai_1 _4883_ (.B1(net1077),
    .Y(_1387_),
    .A1(_1381_),
    .A2(_1386_));
 sg13g2_a21oi_1 _4884_ (.A1(_1381_),
    .A2(_1386_),
    .Y(_0151_),
    .B1(_1387_));
 sg13g2_a21oi_1 _4885_ (.A1(_2800_),
    .A2(_2801_),
    .Y(_1388_),
    .B1(_2803_));
 sg13g2_a21oi_1 _4886_ (.A1(_2786_),
    .A2(_1388_),
    .Y(_1389_),
    .B1(net891));
 sg13g2_o21ai_1 _4887_ (.B1(_1389_),
    .Y(_1390_),
    .A1(_2786_),
    .A2(_1388_));
 sg13g2_xnor2_1 _4888_ (.Y(_1391_),
    .A(_0019_),
    .B(net909));
 sg13g2_o21ai_1 _4889_ (.B1(_1390_),
    .Y(_1392_),
    .A1(net886),
    .A2(_1391_));
 sg13g2_nor2_1 _4890_ (.A(_0309_),
    .B(_0313_),
    .Y(_1393_));
 sg13g2_a21oi_1 _4891_ (.A1(_0310_),
    .A2(_1393_),
    .Y(_1394_),
    .B1(net877));
 sg13g2_o21ai_1 _4892_ (.B1(_1394_),
    .Y(_1395_),
    .A1(_0310_),
    .A2(_1393_));
 sg13g2_xnor2_1 _4893_ (.Y(_1396_),
    .A(_0019_),
    .B(_2704_));
 sg13g2_a21oi_1 _4894_ (.A1(net877),
    .A2(_1396_),
    .Y(_1397_),
    .B1(net883));
 sg13g2_a22oi_1 _4895_ (.Y(_1398_),
    .B1(_1395_),
    .B2(_1397_),
    .A2(net882),
    .A1(net344));
 sg13g2_o21ai_1 _4896_ (.B1(_1398_),
    .Y(_0152_),
    .A1(_0839_),
    .A2(_1392_));
 sg13g2_xor2_1 _4897_ (.B(_2831_),
    .A(_2830_),
    .X(_1399_));
 sg13g2_xnor2_1 _4898_ (.Y(_1400_),
    .A(_2805_),
    .B(_2808_));
 sg13g2_nand2_1 _4899_ (.Y(_1401_),
    .A(net886),
    .B(_1400_));
 sg13g2_a21oi_1 _4900_ (.A1(net891),
    .A2(_1399_),
    .Y(_1402_),
    .B1(net905));
 sg13g2_xnor2_1 _4901_ (.Y(_1403_),
    .A(_0347_),
    .B(_0348_));
 sg13g2_nor3_1 _4902_ (.A(_0311_),
    .B(_0316_),
    .C(_0317_),
    .Y(_1404_));
 sg13g2_nor2_1 _4903_ (.A(_0319_),
    .B(_1404_),
    .Y(_1405_));
 sg13g2_a22oi_1 _4904_ (.Y(_1406_),
    .B1(_1401_),
    .B2(_1402_),
    .A2(net896),
    .A1(net551));
 sg13g2_a21oi_1 _4905_ (.A1(net877),
    .A2(_1403_),
    .Y(_1407_),
    .B1(net884));
 sg13g2_o21ai_1 _4906_ (.B1(_1407_),
    .Y(_1408_),
    .A1(net878),
    .A2(_1405_));
 sg13g2_a21oi_1 _4907_ (.A1(_1406_),
    .A2(_1408_),
    .Y(_0153_),
    .B1(net976));
 sg13g2_nand2_1 _4908_ (.Y(_1409_),
    .A(net504),
    .B(net896));
 sg13g2_a21oi_1 _4909_ (.A1(_0423_),
    .A2(_1409_),
    .Y(_0154_),
    .B1(net979));
 sg13g2_nand2_1 _4910_ (.Y(_1410_),
    .A(net1032),
    .B(net897));
 sg13g2_a21oi_1 _4911_ (.A1(_0407_),
    .A2(_1410_),
    .Y(_0155_),
    .B1(net979));
 sg13g2_nor2_1 _4912_ (.A(net502),
    .B(net895),
    .Y(_1411_));
 sg13g2_nor3_1 _4913_ (.A(_0437_),
    .B(_0446_),
    .C(_1411_),
    .Y(_0156_));
 sg13g2_a22oi_1 _4914_ (.Y(_1412_),
    .B1(net882),
    .B2(net407),
    .A2(_0467_),
    .A1(net990));
 sg13g2_inv_1 _4915_ (.Y(_0157_),
    .A(net408));
 sg13g2_nand2_1 _4916_ (.Y(_1413_),
    .A(net493),
    .B(net897));
 sg13g2_a21oi_1 _4917_ (.A1(_0390_),
    .A2(_1413_),
    .Y(_0158_),
    .B1(net981));
 sg13g2_a22oi_1 _4918_ (.Y(_1414_),
    .B1(net882),
    .B2(net460),
    .A2(_0522_),
    .A1(net986));
 sg13g2_inv_1 _4919_ (.Y(_0159_),
    .A(_1414_));
 sg13g2_nand2_1 _4920_ (.Y(_1415_),
    .A(net440),
    .B(net897));
 sg13g2_a21oi_1 _4921_ (.A1(_0371_),
    .A2(_1415_),
    .Y(_0160_),
    .B1(net981));
 sg13g2_a21oi_1 _4922_ (.A1(_2439_),
    .A2(_0030_),
    .Y(_1416_),
    .B1(\i_bitmap.in[6] ));
 sg13g2_inv_1 _4923_ (.Y(_1417_),
    .A(_1416_));
 sg13g2_nand2_1 _4924_ (.Y(_1418_),
    .A(net969),
    .B(_1417_));
 sg13g2_o21ai_1 _4925_ (.B1(_1418_),
    .Y(_1419_),
    .A1(_2818_),
    .A2(_2820_));
 sg13g2_nor2_1 _4926_ (.A(_0039_),
    .B(net969),
    .Y(_1420_));
 sg13g2_xnor2_1 _4927_ (.Y(_1421_),
    .A(_0039_),
    .B(net969));
 sg13g2_nand2_1 _4928_ (.Y(_1422_),
    .A(_1419_),
    .B(_1421_));
 sg13g2_nor2_1 _4929_ (.A(\i_capsule.tf_x[8] ),
    .B(net969),
    .Y(_1423_));
 sg13g2_xnor2_1 _4930_ (.Y(_1424_),
    .A(_2400_),
    .B(net974));
 sg13g2_a21o_1 _4931_ (.A2(net974),
    .A1(\i_bitmap.in[6] ),
    .B1(_2848_),
    .X(_1425_));
 sg13g2_o21ai_1 _4932_ (.B1(net890),
    .Y(_1426_),
    .A1(_1419_),
    .A2(_1421_));
 sg13g2_nand2b_1 _4933_ (.Y(_1427_),
    .B(_1422_),
    .A_N(_1426_));
 sg13g2_a21oi_1 _4934_ (.A1(_1424_),
    .A2(_1425_),
    .Y(_1428_),
    .B1(net890));
 sg13g2_o21ai_1 _4935_ (.B1(_1428_),
    .Y(_1429_),
    .A1(_1424_),
    .A2(_1425_));
 sg13g2_a21oi_1 _4936_ (.A1(_1427_),
    .A2(_1429_),
    .Y(_1430_),
    .B1(_0839_));
 sg13g2_a22oi_1 _4937_ (.Y(_1431_),
    .B1(_1417_),
    .B2(net943),
    .A2(_0338_),
    .A1(_0336_));
 sg13g2_inv_1 _4938_ (.Y(_1432_),
    .A(_1431_));
 sg13g2_nor2_1 _4939_ (.A(_0039_),
    .B(net942),
    .Y(_1433_));
 sg13g2_xnor2_1 _4940_ (.Y(_1434_),
    .A(_0039_),
    .B(net942));
 sg13g2_xor2_1 _4941_ (.B(_1434_),
    .A(_1431_),
    .X(_1435_));
 sg13g2_nand2_1 _4942_ (.Y(_1436_),
    .A(net875),
    .B(_1435_));
 sg13g2_xnor2_1 _4943_ (.Y(_1437_),
    .A(\i_capsule.tf_x[8] ),
    .B(net942));
 sg13g2_o21ai_1 _4944_ (.B1(_0367_),
    .Y(_1438_),
    .A1(_2401_),
    .A2(net942));
 sg13g2_xnor2_1 _4945_ (.Y(_1439_),
    .A(_1437_),
    .B(_1438_));
 sg13g2_a21oi_1 _4946_ (.A1(net880),
    .A2(_1439_),
    .Y(_1440_),
    .B1(net883));
 sg13g2_a221oi_1 _4947_ (.B2(_1440_),
    .C1(_1430_),
    .B1(_1436_),
    .A1(net532),
    .Y(_1441_),
    .A2(net882));
 sg13g2_inv_1 _4948_ (.Y(_0161_),
    .A(_1441_));
 sg13g2_nor2b_1 _4949_ (.A(_0367_),
    .B_N(_1437_),
    .Y(_1442_));
 sg13g2_nor3_1 _4950_ (.A(\i_capsule.tf_x[8] ),
    .B(_2401_),
    .C(net942),
    .Y(_1443_));
 sg13g2_nor3_1 _4951_ (.A(_1433_),
    .B(_1442_),
    .C(_1443_),
    .Y(_1444_));
 sg13g2_xnor2_1 _4952_ (.Y(_1445_),
    .A(_2399_),
    .B(net943));
 sg13g2_a21oi_1 _4953_ (.A1(_1444_),
    .A2(_1445_),
    .Y(_1446_),
    .B1(net875));
 sg13g2_o21ai_1 _4954_ (.B1(_1446_),
    .Y(_1447_),
    .A1(_1444_),
    .A2(_1445_));
 sg13g2_a22oi_1 _4955_ (.Y(_1448_),
    .B1(_1432_),
    .B2(_1434_),
    .A2(net942),
    .A1(\i_capsule.tf_x[8] ));
 sg13g2_xnor2_1 _4956_ (.Y(_1449_),
    .A(_0056_),
    .B(net937));
 sg13g2_xnor2_1 _4957_ (.Y(_1450_),
    .A(_1448_),
    .B(_1449_));
 sg13g2_o21ai_1 _4958_ (.B1(_1447_),
    .Y(_1451_),
    .A1(net880),
    .A2(_1450_));
 sg13g2_a221oi_1 _4959_ (.B2(_2848_),
    .C1(_1420_),
    .B1(_1424_),
    .A1(\i_bitmap.in[6] ),
    .Y(_1452_),
    .A2(_1423_));
 sg13g2_xnor2_1 _4960_ (.Y(_1453_),
    .A(net1031),
    .B(net974));
 sg13g2_a21oi_1 _4961_ (.A1(_1452_),
    .A2(_1453_),
    .Y(_1454_),
    .B1(net889));
 sg13g2_o21ai_1 _4962_ (.B1(_1454_),
    .Y(_1455_),
    .A1(_1452_),
    .A2(_1453_));
 sg13g2_o21ai_1 _4963_ (.B1(_1422_),
    .Y(_1456_),
    .A1(_2400_),
    .A2(net974));
 sg13g2_xnor2_1 _4964_ (.Y(_1457_),
    .A(_0056_),
    .B(net974));
 sg13g2_xnor2_1 _4965_ (.Y(_1458_),
    .A(_1456_),
    .B(_1457_));
 sg13g2_nand2_1 _4966_ (.Y(_1459_),
    .A(net889),
    .B(_1458_));
 sg13g2_a21oi_1 _4967_ (.A1(_1455_),
    .A2(_1459_),
    .Y(_1460_),
    .B1(_0839_));
 sg13g2_a221oi_1 _4968_ (.B2(_0856_),
    .C1(_1460_),
    .B1(_1451_),
    .A1(net1031),
    .Y(_1461_),
    .A2(_0859_));
 sg13g2_inv_1 _4969_ (.Y(_0162_),
    .A(_1461_));
 sg13g2_nand2b_1 _4970_ (.Y(_1462_),
    .B(_2751_),
    .A_N(_0060_));
 sg13g2_nor2_1 _4971_ (.A(_0061_),
    .B(_1164_),
    .Y(_1463_));
 sg13g2_xnor2_1 _4972_ (.Y(_1464_),
    .A(_2425_),
    .B(_1463_));
 sg13g2_o21ai_1 _4973_ (.B1(_1462_),
    .Y(_1465_),
    .A1(net892),
    .A2(_1464_));
 sg13g2_nor2_1 _4974_ (.A(\center_y[5] ),
    .B(net984),
    .Y(_1466_));
 sg13g2_a221oi_1 _4975_ (.B2(_1465_),
    .C1(_1466_),
    .B1(_0838_),
    .A1(_2425_),
    .Y(_0163_),
    .A2(_0441_));
 sg13g2_nor4_1 _4976_ (.A(_2425_),
    .B(_2426_),
    .C(net891),
    .D(_1164_),
    .Y(_1467_));
 sg13g2_a21oi_1 _4977_ (.A1(_2425_),
    .A2(net892),
    .Y(_1468_),
    .B1(_1467_));
 sg13g2_and2_1 _4978_ (.A(_2424_),
    .B(_1468_),
    .X(_1469_));
 sg13g2_o21ai_1 _4979_ (.B1(_0838_),
    .Y(_1470_),
    .A1(_2424_),
    .A2(_1468_));
 sg13g2_a22oi_1 _4980_ (.Y(_1471_),
    .B1(_0441_),
    .B2(net484),
    .A2(net977),
    .A1(net451));
 sg13g2_o21ai_1 _4981_ (.B1(_1471_),
    .Y(_0164_),
    .A1(_1469_),
    .A2(_1470_));
 sg13g2_nor3_1 _4982_ (.A(\i_transform.track_y[6] ),
    .B(\i_transform.track_y[5] ),
    .C(net887),
    .Y(_1472_));
 sg13g2_and2_1 _4983_ (.A(\i_transform.track_y[6] ),
    .B(_1467_),
    .X(_1473_));
 sg13g2_nor2_1 _4984_ (.A(_1472_),
    .B(_1473_),
    .Y(_1474_));
 sg13g2_xor2_1 _4985_ (.B(_1474_),
    .A(net489),
    .X(_1475_));
 sg13g2_a22oi_1 _4986_ (.Y(_1476_),
    .B1(_0441_),
    .B2(net489),
    .A2(net977),
    .A1(net447));
 sg13g2_o21ai_1 _4987_ (.B1(_1476_),
    .Y(_0165_),
    .A1(_0839_),
    .A2(_1475_));
 sg13g2_nand2b_1 _4988_ (.Y(_1477_),
    .B(_1472_),
    .A_N(\i_transform.track_y[7] ));
 sg13g2_nand2_1 _4989_ (.Y(_1478_),
    .A(\i_transform.track_y[7] ),
    .B(_1473_));
 sg13g2_nand2_1 _4990_ (.Y(_1479_),
    .A(_1477_),
    .B(_1478_));
 sg13g2_a21oi_1 _4991_ (.A1(\i_transform.track_y[8] ),
    .A2(_1479_),
    .Y(_1480_),
    .B1(_0839_));
 sg13g2_o21ai_1 _4992_ (.B1(_1480_),
    .Y(_1481_),
    .A1(net396),
    .A2(_1479_));
 sg13g2_a22oi_1 _4993_ (.Y(_1482_),
    .B1(_0441_),
    .B2(net396),
    .A2(net977),
    .A1(net390));
 sg13g2_nand2_1 _4994_ (.Y(_0166_),
    .A(_1481_),
    .B(_1482_));
 sg13g2_nand3_1 _4995_ (.B(\i_transform.track_y[8] ),
    .C(_1473_),
    .A(\i_transform.track_y[7] ),
    .Y(_1483_));
 sg13g2_o21ai_1 _4996_ (.B1(_1483_),
    .Y(_1484_),
    .A1(\i_transform.track_y[8] ),
    .A2(_1477_));
 sg13g2_xnor2_1 _4997_ (.Y(_1485_),
    .A(net293),
    .B(_1484_));
 sg13g2_a22oi_1 _4998_ (.Y(_1486_),
    .B1(_0441_),
    .B2(net293),
    .A2(net977),
    .A1(\center_y[9] ));
 sg13g2_o21ai_1 _4999_ (.B1(net294),
    .Y(_0167_),
    .A1(_0839_),
    .A2(_1485_));
 sg13g2_nor2_1 _5000_ (.A(net3),
    .B(_1308_),
    .Y(_1487_));
 sg13g2_and2_1 _5001_ (.A(net256),
    .B(_1487_),
    .X(_0168_));
 sg13g2_and2_1 _5002_ (.A(net262),
    .B(_1487_),
    .X(_0169_));
 sg13g2_nor2b_1 _5003_ (.A(net1034),
    .B_N(net256),
    .Y(_1488_));
 sg13g2_nor2_1 _5004_ (.A(\i_collision.vy[1] ),
    .B(net1035),
    .Y(_1489_));
 sg13g2_nand2b_1 _5005_ (.Y(_1490_),
    .B(net1036),
    .A_N(\i_collision.vx[1] ));
 sg13g2_nor2b_2 _5006_ (.A(_1489_),
    .B_N(_1490_),
    .Y(_1491_));
 sg13g2_nand2b_2 _5007_ (.Y(_1492_),
    .B(_1490_),
    .A_N(_1489_));
 sg13g2_nor2_1 _5008_ (.A(net999),
    .B(net1023),
    .Y(_1493_));
 sg13g2_xor2_1 _5009_ (.B(net1035),
    .A(net1020),
    .X(_1494_));
 sg13g2_xnor2_1 _5010_ (.Y(_1495_),
    .A(net1020),
    .B(net1035));
 sg13g2_nor2_1 _5011_ (.A(net1035),
    .B(_0008_),
    .Y(_1496_));
 sg13g2_nand2_1 _5012_ (.Y(_1497_),
    .A(net1036),
    .B(_2434_));
 sg13g2_nor2b_1 _5013_ (.A(_1496_),
    .B_N(_1497_),
    .Y(_1498_));
 sg13g2_nand2b_1 _5014_ (.Y(_1499_),
    .B(_1497_),
    .A_N(_1496_));
 sg13g2_and2_1 _5015_ (.A(net999),
    .B(net1023),
    .X(_1500_));
 sg13g2_nand2_1 _5016_ (.Y(_1501_),
    .A(net999),
    .B(net1023));
 sg13g2_o21ai_1 _5017_ (.B1(net925),
    .Y(_1502_),
    .A1(_1493_),
    .A2(net951));
 sg13g2_a21oi_1 _5018_ (.A1(net951),
    .A2(_1501_),
    .Y(_1503_),
    .B1(_1502_));
 sg13g2_nand2_1 _5019_ (.Y(_1504_),
    .A(net1023),
    .B(net951));
 sg13g2_nor2_2 _5020_ (.A(_2374_),
    .B(net951),
    .Y(_1505_));
 sg13g2_nand2_1 _5021_ (.Y(_1506_),
    .A(net1002),
    .B(net953));
 sg13g2_nand3b_1 _5022_ (.B(_1504_),
    .C(_1506_),
    .Y(_1507_),
    .A_N(_1493_));
 sg13g2_nor2_1 _5023_ (.A(net925),
    .B(_1507_),
    .Y(_1508_));
 sg13g2_o21ai_1 _5024_ (.B1(_1491_),
    .Y(_1509_),
    .A1(_1503_),
    .A2(_1508_));
 sg13g2_nor2_1 _5025_ (.A(net995),
    .B(net1005),
    .Y(_1510_));
 sg13g2_nor2_1 _5026_ (.A(_1491_),
    .B(net924),
    .Y(_1511_));
 sg13g2_nand3_1 _5027_ (.B(_1510_),
    .C(_1511_),
    .A(_1507_),
    .Y(_1512_));
 sg13g2_nand2_2 _5028_ (.Y(_1513_),
    .A(_1492_),
    .B(net924));
 sg13g2_nor2_1 _5029_ (.A(_2444_),
    .B(net951),
    .Y(_1514_));
 sg13g2_nand2_1 _5030_ (.Y(_1515_),
    .A(_2373_),
    .B(net1024));
 sg13g2_o21ai_1 _5031_ (.B1(net949),
    .Y(_1516_),
    .A1(net1023),
    .A2(net951));
 sg13g2_o21ai_1 _5032_ (.B1(_1516_),
    .Y(_1517_),
    .A1(_0050_),
    .A2(net953));
 sg13g2_a21oi_1 _5033_ (.A1(net1002),
    .A2(_1517_),
    .Y(_1518_),
    .B1(_1513_));
 sg13g2_o21ai_1 _5034_ (.B1(_1504_),
    .Y(_1519_),
    .A1(net949),
    .A2(_1514_));
 sg13g2_o21ai_1 _5035_ (.B1(_1518_),
    .Y(_1520_),
    .A1(net1002),
    .A2(_1519_));
 sg13g2_nand3_1 _5036_ (.B(_1512_),
    .C(_1520_),
    .A(_1509_),
    .Y(_1521_));
 sg13g2_nor2_1 _5037_ (.A(net1030),
    .B(net1036),
    .Y(_1522_));
 sg13g2_a21oi_2 _5038_ (.B1(_1522_),
    .Y(_1523_),
    .A2(net1036),
    .A1(_2396_));
 sg13g2_xor2_1 _5039_ (.B(_1523_),
    .A(\i_collision.mirror ),
    .X(_1524_));
 sg13g2_xnor2_1 _5040_ (.Y(_1525_),
    .A(\i_collision.mirror ),
    .B(_1523_));
 sg13g2_nor2_2 _5041_ (.A(net1002),
    .B(net953),
    .Y(_1526_));
 sg13g2_o21ai_1 _5042_ (.B1(_1504_),
    .Y(_1527_),
    .A1(_1500_),
    .A2(_1526_));
 sg13g2_nor3_1 _5043_ (.A(net949),
    .B(_1525_),
    .C(_1527_),
    .Y(_1528_));
 sg13g2_mux2_1 _5044_ (.A0(net921),
    .A1(_1528_),
    .S(_1521_),
    .X(_1529_));
 sg13g2_a21oi_1 _5045_ (.A1(net1033),
    .A2(_1529_),
    .Y(_1530_),
    .B1(_1488_));
 sg13g2_nor2_1 _5046_ (.A(net1070),
    .B(_1530_),
    .Y(_0170_));
 sg13g2_nand2b_1 _5047_ (.Y(_1531_),
    .B(net262),
    .A_N(net1033));
 sg13g2_or2_1 _5048_ (.X(_1532_),
    .B(net1024),
    .A(net995));
 sg13g2_nand2_1 _5049_ (.Y(_1533_),
    .A(net952),
    .B(_1532_));
 sg13g2_nand2_1 _5050_ (.Y(_1534_),
    .A(net1005),
    .B(net952));
 sg13g2_a21oi_1 _5051_ (.A1(\i_collision.i_coll_table.in[1] ),
    .A2(net949),
    .Y(_1535_),
    .B1(_2374_));
 sg13g2_nand2_1 _5052_ (.Y(_1536_),
    .A(_1533_),
    .B(_1534_));
 sg13g2_o21ai_1 _5053_ (.B1(_1506_),
    .Y(_1537_),
    .A1(_1535_),
    .A2(_1536_));
 sg13g2_nor3_1 _5054_ (.A(_1491_),
    .B(net924),
    .C(_1537_),
    .Y(_1538_));
 sg13g2_o21ai_1 _5055_ (.B1(_1505_),
    .Y(_1539_),
    .A1(net997),
    .A2(_0050_));
 sg13g2_o21ai_1 _5056_ (.B1(_1526_),
    .Y(_1540_),
    .A1(net997),
    .A2(_2444_));
 sg13g2_nand3_1 _5057_ (.B(_1539_),
    .C(_1540_),
    .A(net925),
    .Y(_1541_));
 sg13g2_o21ai_1 _5058_ (.B1(net1004),
    .Y(_1542_),
    .A1(_1505_),
    .A2(_1526_));
 sg13g2_nand3b_1 _5059_ (.B(_1542_),
    .C(_1492_),
    .Y(_1543_),
    .A_N(_1541_));
 sg13g2_nor2_1 _5060_ (.A(_1492_),
    .B(net923),
    .Y(_1544_));
 sg13g2_nand2b_1 _5061_ (.Y(_1545_),
    .B(_1544_),
    .A_N(_1507_));
 sg13g2_nand4_1 _5062_ (.B(net921),
    .C(_1543_),
    .A(net1033),
    .Y(_1546_),
    .D(_1545_));
 sg13g2_o21ai_1 _5063_ (.B1(_1531_),
    .Y(_1547_),
    .A1(_1538_),
    .A2(_1546_));
 sg13g2_and2_1 _5064_ (.A(net1071),
    .B(_1547_),
    .X(_0171_));
 sg13g2_nor2b_2 _5065_ (.A(net1035),
    .B_N(net1034),
    .Y(_1548_));
 sg13g2_nor2_1 _5066_ (.A(net922),
    .B(_1527_),
    .Y(_1549_));
 sg13g2_nand2b_2 _5067_ (.Y(_1550_),
    .B(net997),
    .A_N(net1003));
 sg13g2_inv_1 _5068_ (.Y(_1551_),
    .A(_1550_));
 sg13g2_nand3_1 _5069_ (.B(net1050),
    .C(_1492_),
    .A(net1004),
    .Y(_1552_));
 sg13g2_o21ai_1 _5070_ (.B1(_1552_),
    .Y(_1553_),
    .A1(net1050),
    .A2(_1550_));
 sg13g2_nand2_1 _5071_ (.Y(_1554_),
    .A(_1549_),
    .B(_1553_));
 sg13g2_o21ai_1 _5072_ (.B1(net924),
    .Y(_1555_),
    .A1(_2373_),
    .A2(net1050));
 sg13g2_a221oi_1 _5073_ (.B2(_1491_),
    .C1(net921),
    .B1(_1555_),
    .A1(_0053_),
    .Y(_1556_),
    .A2(net923));
 sg13g2_nor2_2 _5074_ (.A(net1024),
    .B(_2414_),
    .Y(_1557_));
 sg13g2_nor2_1 _5075_ (.A(net953),
    .B(_1557_),
    .Y(_1558_));
 sg13g2_o21ai_1 _5076_ (.B1(net950),
    .Y(_1559_),
    .A1(net1024),
    .A2(_2414_));
 sg13g2_a21oi_2 _5077_ (.B1(net950),
    .Y(_1560_),
    .A2(_2414_),
    .A1(net1024));
 sg13g2_nand3b_1 _5078_ (.B(net996),
    .C(_1559_),
    .Y(_1561_),
    .A_N(_1560_));
 sg13g2_nor2_1 _5079_ (.A(net1004),
    .B(_1558_),
    .Y(_1562_));
 sg13g2_a21oi_1 _5080_ (.A1(_2373_),
    .A2(_1558_),
    .Y(_1563_),
    .B1(net1003));
 sg13g2_a221oi_1 _5081_ (.B2(_1563_),
    .C1(net1000),
    .B1(_1561_),
    .A1(net1003),
    .Y(_1564_),
    .A2(_1560_));
 sg13g2_nor2_1 _5082_ (.A(net1024),
    .B(net1049),
    .Y(_1565_));
 sg13g2_or2_1 _5083_ (.X(_1566_),
    .B(_1565_),
    .A(net953));
 sg13g2_nand2_2 _5084_ (.Y(_1567_),
    .A(net1024),
    .B(net1049));
 sg13g2_and2_1 _5085_ (.A(net953),
    .B(_1567_),
    .X(_1568_));
 sg13g2_nand2_1 _5086_ (.Y(_1569_),
    .A(net952),
    .B(_1567_));
 sg13g2_nand3_1 _5087_ (.B(_1566_),
    .C(_1569_),
    .A(net996),
    .Y(_1570_));
 sg13g2_a21oi_1 _5088_ (.A1(_2373_),
    .A2(_1568_),
    .Y(_1571_),
    .B1(net1003));
 sg13g2_nand2_2 _5089_ (.Y(_1572_),
    .A(net1003),
    .B(net950));
 sg13g2_o21ai_1 _5090_ (.B1(net1000),
    .Y(_1573_),
    .A1(_1565_),
    .A2(_1572_));
 sg13g2_a21oi_1 _5091_ (.A1(_1570_),
    .A2(_1571_),
    .Y(_1574_),
    .B1(_1573_));
 sg13g2_o21ai_1 _5092_ (.B1(_1511_),
    .Y(_1575_),
    .A1(_1564_),
    .A2(_1574_));
 sg13g2_o21ai_1 _5093_ (.B1(_2374_),
    .Y(_1576_),
    .A1(net1049),
    .A2(_1532_));
 sg13g2_nand2_1 _5094_ (.Y(_1577_),
    .A(net995),
    .B(net950));
 sg13g2_nor2_1 _5095_ (.A(_1557_),
    .B(_1577_),
    .Y(_1578_));
 sg13g2_o21ai_1 _5096_ (.B1(net1000),
    .Y(_1579_),
    .A1(net1049),
    .A2(_1515_));
 sg13g2_nand3_1 _5097_ (.B(net952),
    .C(_1567_),
    .A(net996),
    .Y(_1580_));
 sg13g2_nand2b_1 _5098_ (.Y(_1581_),
    .B(_1580_),
    .A_N(_1579_));
 sg13g2_o21ai_1 _5099_ (.B1(_1581_),
    .Y(_1582_),
    .A1(_1576_),
    .A2(_1578_));
 sg13g2_o21ai_1 _5100_ (.B1(_1560_),
    .Y(_1583_),
    .A1(net1000),
    .A2(_2414_));
 sg13g2_a21o_1 _5101_ (.A2(net1049),
    .A1(net1000),
    .B1(_1566_),
    .X(_1584_));
 sg13g2_nand3_1 _5102_ (.B(_1583_),
    .C(_1584_),
    .A(net922),
    .Y(_1585_));
 sg13g2_nand2_1 _5103_ (.Y(_1586_),
    .A(_1491_),
    .B(_1585_));
 sg13g2_a21oi_1 _5104_ (.A1(net924),
    .A2(_1582_),
    .Y(_1587_),
    .B1(_1586_));
 sg13g2_xnor2_1 _5105_ (.Y(_1588_),
    .A(_2373_),
    .B(_1567_));
 sg13g2_nor2_1 _5106_ (.A(_1572_),
    .B(_1588_),
    .Y(_1589_));
 sg13g2_nor3_1 _5107_ (.A(net1003),
    .B(_0051_),
    .C(net952),
    .Y(_1590_));
 sg13g2_nor3_1 _5108_ (.A(net1001),
    .B(_1589_),
    .C(_1590_),
    .Y(_1591_));
 sg13g2_nor2_1 _5109_ (.A(_2414_),
    .B(_1532_),
    .Y(_1592_));
 sg13g2_xnor2_1 _5110_ (.Y(_1593_),
    .A(net995),
    .B(_1557_));
 sg13g2_nor2_1 _5111_ (.A(net950),
    .B(_1550_),
    .Y(_1594_));
 sg13g2_o21ai_1 _5112_ (.B1(net1000),
    .Y(_1595_),
    .A1(_1534_),
    .A2(_1593_));
 sg13g2_nor2_1 _5113_ (.A(_1594_),
    .B(_1595_),
    .Y(_1596_));
 sg13g2_nor3_1 _5114_ (.A(_1513_),
    .B(_1591_),
    .C(_1596_),
    .Y(_1597_));
 sg13g2_nor3_1 _5115_ (.A(_1524_),
    .B(_1587_),
    .C(_1597_),
    .Y(_1598_));
 sg13g2_a22oi_1 _5116_ (.Y(_1599_),
    .B1(_1575_),
    .B2(_1598_),
    .A2(_1556_),
    .A1(_1554_));
 sg13g2_a21oi_1 _5117_ (.A1(_1548_),
    .A2(_1599_),
    .Y(_1600_),
    .B1(net1070));
 sg13g2_o21ai_1 _5118_ (.B1(_1600_),
    .Y(_0172_),
    .A1(_2398_),
    .A2(_1548_));
 sg13g2_nand2_1 _5119_ (.Y(_1601_),
    .A(_1492_),
    .B(_1524_));
 sg13g2_nor2_1 _5120_ (.A(_0052_),
    .B(net922),
    .Y(_1602_));
 sg13g2_nor2_1 _5121_ (.A(net1049),
    .B(_1527_),
    .Y(_1603_));
 sg13g2_a21oi_1 _5122_ (.A1(_1602_),
    .A2(_1603_),
    .Y(_1604_),
    .B1(_1601_));
 sg13g2_nand2_1 _5123_ (.Y(_1605_),
    .A(_1559_),
    .B(_1569_));
 sg13g2_o21ai_1 _5124_ (.B1(_1605_),
    .Y(_1606_),
    .A1(_1505_),
    .A2(_1526_));
 sg13g2_a21oi_1 _5125_ (.A1(net923),
    .A2(_1606_),
    .Y(_1607_),
    .B1(_1492_));
 sg13g2_nand2_1 _5126_ (.Y(_1608_),
    .A(_1541_),
    .B(_1607_));
 sg13g2_o21ai_1 _5127_ (.B1(_1542_),
    .Y(_1609_),
    .A1(_0051_),
    .A2(_1606_));
 sg13g2_o21ai_1 _5128_ (.B1(_1526_),
    .Y(_1610_),
    .A1(net997),
    .A2(_1567_));
 sg13g2_o21ai_1 _5129_ (.B1(_1610_),
    .Y(_1611_),
    .A1(_1506_),
    .A2(_1592_));
 sg13g2_nor2_1 _5130_ (.A(_0052_),
    .B(_1513_),
    .Y(_1612_));
 sg13g2_a221oi_1 _5131_ (.B2(_1612_),
    .C1(_1524_),
    .B1(_1611_),
    .A1(_1511_),
    .Y(_1613_),
    .A2(_1609_));
 sg13g2_a21oi_2 _5132_ (.B1(_1604_),
    .Y(_1614_),
    .A2(_1613_),
    .A1(_1608_));
 sg13g2_nor2b_1 _5133_ (.A(_1614_),
    .B_N(_1548_),
    .Y(_1615_));
 sg13g2_o21ai_1 _5134_ (.B1(net1071),
    .Y(_1616_),
    .A1(net516),
    .A2(_1548_));
 sg13g2_nor2_1 _5135_ (.A(_1615_),
    .B(_1616_),
    .Y(_0173_));
 sg13g2_a22oi_1 _5136_ (.Y(_1617_),
    .B1(_1537_),
    .B2(_1492_),
    .A2(_1513_),
    .A1(_1507_));
 sg13g2_nor2_1 _5137_ (.A(\i_collision.mirror ),
    .B(_1617_),
    .Y(_1618_));
 sg13g2_a21oi_1 _5138_ (.A1(_1523_),
    .A2(_1617_),
    .Y(_1619_),
    .B1(_1618_));
 sg13g2_o21ai_1 _5139_ (.B1(net1071),
    .Y(_1620_),
    .A1(net1030),
    .A2(_1548_));
 sg13g2_a21oi_1 _5140_ (.A1(_1548_),
    .A2(_1619_),
    .Y(_0174_),
    .B1(_1620_));
 sg13g2_nand2_1 _5141_ (.Y(_1621_),
    .A(net1034),
    .B(net1035));
 sg13g2_o21ai_1 _5142_ (.B1(net1071),
    .Y(_1622_),
    .A1(_1599_),
    .A2(_1621_));
 sg13g2_a21oi_1 _5143_ (.A1(_2397_),
    .A2(_1621_),
    .Y(_0175_),
    .B1(_1622_));
 sg13g2_nand3_1 _5144_ (.B(net1035),
    .C(_1614_),
    .A(net1034),
    .Y(_1623_));
 sg13g2_a21oi_1 _5145_ (.A1(net499),
    .A2(_1621_),
    .Y(_1624_),
    .B1(net1070));
 sg13g2_nand2_1 _5146_ (.Y(_0176_),
    .A(_1623_),
    .B(_1624_));
 sg13g2_nand3_1 _5147_ (.B(net1035),
    .C(_1619_),
    .A(net1034),
    .Y(_1625_));
 sg13g2_nand2_1 _5148_ (.Y(_1626_),
    .A(net1071),
    .B(_1625_));
 sg13g2_a21oi_1 _5149_ (.A1(_2396_),
    .A2(_1621_),
    .Y(_0177_),
    .B1(_1626_));
 sg13g2_and3_1 _5150_ (.X(_1627_),
    .A(net1040),
    .B(\i_collision.vy[1] ),
    .C(\i_collision.vy[0] ));
 sg13g2_nor2_2 _5151_ (.A(net1069),
    .B(net2),
    .Y(_1628_));
 sg13g2_nand2b_2 _5152_ (.Y(_1629_),
    .B(net1074),
    .A_N(net2));
 sg13g2_o21ai_1 _5153_ (.B1(net947),
    .Y(_1630_),
    .A1(net252),
    .A2(_1627_));
 sg13g2_a21oi_1 _5154_ (.A1(net252),
    .A2(_1627_),
    .Y(_0178_),
    .B1(_1630_));
 sg13g2_nand3_1 _5155_ (.B(\i_collision.vy[1] ),
    .C(\i_collision.vy[0] ),
    .A(net252),
    .Y(_1631_));
 sg13g2_nor2_1 _5156_ (.A(\i_collision.vy[1] ),
    .B(\i_collision.vy[0] ),
    .Y(_1632_));
 sg13g2_nor2b_1 _5157_ (.A(net1030),
    .B_N(\i_collision.vy[1] ),
    .Y(_1633_));
 sg13g2_nor2b_1 _5158_ (.A(\i_collision.vy[0] ),
    .B_N(\i_collision.vy[1] ),
    .Y(_1634_));
 sg13g2_a21oi_1 _5159_ (.A1(\i_collision.vy[0] ),
    .A2(_1633_),
    .Y(_1635_),
    .B1(_1632_));
 sg13g2_nand2_1 _5160_ (.Y(_1636_),
    .A(\i_kinematics.center_y_lo[1] ),
    .B(_1635_));
 sg13g2_xnor2_1 _5161_ (.Y(_1637_),
    .A(net362),
    .B(_1635_));
 sg13g2_or2_1 _5162_ (.X(_1638_),
    .B(_1637_),
    .A(_1631_));
 sg13g2_xnor2_1 _5163_ (.Y(_1639_),
    .A(_1631_),
    .B(_1637_));
 sg13g2_o21ai_1 _5164_ (.B1(net947),
    .Y(_1640_),
    .A1(net1040),
    .A2(net362));
 sg13g2_a21oi_1 _5165_ (.A1(net1040),
    .A2(_1639_),
    .Y(_0179_),
    .B1(_1640_));
 sg13g2_and3_1 _5166_ (.X(_1641_),
    .A(net1045),
    .B(\i_collision.vx[1] ),
    .C(\i_collision.vx[0] ));
 sg13g2_o21ai_1 _5167_ (.B1(net948),
    .Y(_1642_),
    .A1(net254),
    .A2(_1641_));
 sg13g2_a21oi_1 _5168_ (.A1(net254),
    .A2(_1641_),
    .Y(_0180_),
    .B1(_1642_));
 sg13g2_nand3_1 _5169_ (.B(\i_collision.vx[1] ),
    .C(\i_collision.vx[0] ),
    .A(net254),
    .Y(_1643_));
 sg13g2_nor2_1 _5170_ (.A(\i_collision.vx[1] ),
    .B(\i_collision.vx[0] ),
    .Y(_1644_));
 sg13g2_nor2b_1 _5171_ (.A(net1027),
    .B_N(\i_collision.vx[1] ),
    .Y(_1645_));
 sg13g2_a21oi_1 _5172_ (.A1(\i_collision.vx[0] ),
    .A2(_1645_),
    .Y(_1646_),
    .B1(_1644_));
 sg13g2_nand2_1 _5173_ (.Y(_1647_),
    .A(\i_kinematics.center_x_lo[1] ),
    .B(_1646_));
 sg13g2_xnor2_1 _5174_ (.Y(_1648_),
    .A(net360),
    .B(_1646_));
 sg13g2_or2_1 _5175_ (.X(_1649_),
    .B(_1648_),
    .A(_1643_));
 sg13g2_xnor2_1 _5176_ (.Y(_1650_),
    .A(_1643_),
    .B(_1648_));
 sg13g2_o21ai_1 _5177_ (.B1(net948),
    .Y(_1651_),
    .A1(net1045),
    .A2(net360));
 sg13g2_a21oi_1 _5178_ (.A1(net1045),
    .A2(_1650_),
    .Y(_0181_),
    .B1(_1651_));
 sg13g2_nor2_1 _5179_ (.A(net1030),
    .B(_0008_),
    .Y(_1652_));
 sg13g2_a21oi_1 _5180_ (.A1(net1030),
    .A2(_1634_),
    .Y(_1653_),
    .B1(_1652_));
 sg13g2_nor2b_1 _5181_ (.A(_1653_),
    .B_N(\center_y[0] ),
    .Y(_1654_));
 sg13g2_xnor2_1 _5182_ (.Y(_1655_),
    .A(\center_y[0] ),
    .B(_1653_));
 sg13g2_inv_1 _5183_ (.Y(_1656_),
    .A(_1655_));
 sg13g2_and3_1 _5184_ (.X(_1657_),
    .A(_1636_),
    .B(_1638_),
    .C(_1656_));
 sg13g2_a21oi_1 _5185_ (.A1(_1636_),
    .A2(_1638_),
    .Y(_1658_),
    .B1(_1656_));
 sg13g2_or2_1 _5186_ (.X(_1659_),
    .B(_1658_),
    .A(_1657_));
 sg13g2_o21ai_1 _5187_ (.B1(net947),
    .Y(_1660_),
    .A1(net1041),
    .A2(net459));
 sg13g2_a21oi_1 _5188_ (.A1(net1041),
    .A2(_1659_),
    .Y(_0182_),
    .B1(_1660_));
 sg13g2_xor2_1 _5189_ (.B(\i_collision.vy[1] ),
    .A(net1030),
    .X(_1661_));
 sg13g2_nand2b_1 _5190_ (.Y(_1662_),
    .B(_1661_),
    .A_N(_1632_));
 sg13g2_nand2_1 _5191_ (.Y(_1663_),
    .A(\center_y[1] ),
    .B(_1662_));
 sg13g2_xor2_1 _5192_ (.B(_1662_),
    .A(\center_y[1] ),
    .X(_1664_));
 sg13g2_or3_1 _5193_ (.A(_1654_),
    .B(_1658_),
    .C(_1664_),
    .X(_1665_));
 sg13g2_o21ai_1 _5194_ (.B1(_1664_),
    .Y(_1666_),
    .A1(_1654_),
    .A2(_1658_));
 sg13g2_a21oi_1 _5195_ (.A1(_1665_),
    .A2(_1666_),
    .Y(_1667_),
    .B1(net992));
 sg13g2_o21ai_1 _5196_ (.B1(net947),
    .Y(_1668_),
    .A1(net1045),
    .A2(net437));
 sg13g2_nor2_1 _5197_ (.A(_1667_),
    .B(_1668_),
    .Y(_0183_));
 sg13g2_xnor2_1 _5198_ (.Y(_1669_),
    .A(\center_y[2] ),
    .B(_1661_));
 sg13g2_and3_1 _5199_ (.X(_1670_),
    .A(_1663_),
    .B(_1666_),
    .C(_1669_));
 sg13g2_a21oi_1 _5200_ (.A1(_1663_),
    .A2(_1666_),
    .Y(_1671_),
    .B1(_1669_));
 sg13g2_o21ai_1 _5201_ (.B1(net1041),
    .Y(_1672_),
    .A1(_1670_),
    .A2(_1671_));
 sg13g2_o21ai_1 _5202_ (.B1(_1672_),
    .Y(_1673_),
    .A1(net1041),
    .A2(net317));
 sg13g2_nor2_1 _5203_ (.A(net1065),
    .B(_1673_),
    .Y(_0184_));
 sg13g2_a21oi_1 _5204_ (.A1(net387),
    .A2(_1661_),
    .Y(_1674_),
    .B1(_1671_));
 sg13g2_or2_1 _5205_ (.X(_1675_),
    .B(net1029),
    .A(\center_y[3] ));
 sg13g2_nand2_1 _5206_ (.Y(_1676_),
    .A(\center_y[3] ),
    .B(net1029));
 sg13g2_nand2_1 _5207_ (.Y(_1677_),
    .A(_1675_),
    .B(_1676_));
 sg13g2_xnor2_1 _5208_ (.Y(_1678_),
    .A(_1674_),
    .B(_1677_));
 sg13g2_o21ai_1 _5209_ (.B1(net947),
    .Y(_1679_),
    .A1(net1040),
    .A2(net406));
 sg13g2_a21oi_1 _5210_ (.A1(net1040),
    .A2(_1678_),
    .Y(_0185_),
    .B1(_1679_));
 sg13g2_nand2_1 _5211_ (.Y(_1680_),
    .A(\center_y[4] ),
    .B(net1029));
 sg13g2_xor2_1 _5212_ (.B(net1029),
    .A(net461),
    .X(_1681_));
 sg13g2_nand2_1 _5213_ (.Y(_1682_),
    .A(_1674_),
    .B(_1676_));
 sg13g2_a21oi_1 _5214_ (.A1(_1675_),
    .A2(_1682_),
    .Y(_1683_),
    .B1(_1681_));
 sg13g2_nand3_1 _5215_ (.B(_1681_),
    .C(_1682_),
    .A(_1675_),
    .Y(_1684_));
 sg13g2_nand2_1 _5216_ (.Y(_1685_),
    .A(net1040),
    .B(_1684_));
 sg13g2_a21oi_1 _5217_ (.A1(net991),
    .A2(net461),
    .Y(_1686_),
    .B1(net1065));
 sg13g2_o21ai_1 _5218_ (.B1(_1686_),
    .Y(_0186_),
    .A1(_1683_),
    .A2(_1685_));
 sg13g2_and2_1 _5219_ (.A(_1680_),
    .B(_1684_),
    .X(_1687_));
 sg13g2_nor2_1 _5220_ (.A(\center_y[5] ),
    .B(net1028),
    .Y(_1688_));
 sg13g2_nand2_1 _5221_ (.Y(_1689_),
    .A(\center_y[5] ),
    .B(net1028));
 sg13g2_nand2b_1 _5222_ (.Y(_1690_),
    .B(_1689_),
    .A_N(_1688_));
 sg13g2_xnor2_1 _5223_ (.Y(_1691_),
    .A(_1687_),
    .B(_1690_));
 sg13g2_a21oi_1 _5224_ (.A1(net991),
    .A2(net465),
    .Y(_1692_),
    .B1(net1065));
 sg13g2_o21ai_1 _5225_ (.B1(_1692_),
    .Y(_0187_),
    .A1(net991),
    .A2(_1691_));
 sg13g2_and2_1 _5226_ (.A(\center_y[6] ),
    .B(net1028),
    .X(_1693_));
 sg13g2_xor2_1 _5227_ (.B(net1028),
    .A(\center_y[6] ),
    .X(_1694_));
 sg13g2_o21ai_1 _5228_ (.B1(_1689_),
    .Y(_1695_),
    .A1(_1687_),
    .A2(_1688_));
 sg13g2_xnor2_1 _5229_ (.Y(_1696_),
    .A(_1694_),
    .B(_1695_));
 sg13g2_a21oi_1 _5230_ (.A1(net991),
    .A2(net451),
    .Y(_1697_),
    .B1(net1065));
 sg13g2_o21ai_1 _5231_ (.B1(_1697_),
    .Y(_0188_),
    .A1(net991),
    .A2(_1696_));
 sg13g2_a21o_1 _5232_ (.A2(_1695_),
    .A1(_1694_),
    .B1(_1693_),
    .X(_1698_));
 sg13g2_xor2_1 _5233_ (.B(net1028),
    .A(\center_y[7] ),
    .X(_1699_));
 sg13g2_xnor2_1 _5234_ (.Y(_1700_),
    .A(_1698_),
    .B(_1699_));
 sg13g2_a21oi_1 _5235_ (.A1(net991),
    .A2(net447),
    .Y(_1701_),
    .B1(net1065));
 sg13g2_o21ai_1 _5236_ (.B1(_1701_),
    .Y(_0189_),
    .A1(net991),
    .A2(_1700_));
 sg13g2_nand2b_1 _5237_ (.Y(_1702_),
    .B(net1029),
    .A_N(\center_y[8] ));
 sg13g2_xnor2_1 _5238_ (.Y(_1703_),
    .A(\center_y[8] ),
    .B(net1028));
 sg13g2_a21o_1 _5239_ (.A2(net1028),
    .A1(\center_y[7] ),
    .B1(_1698_),
    .X(_1704_));
 sg13g2_o21ai_1 _5240_ (.B1(_1704_),
    .Y(_1705_),
    .A1(\center_y[7] ),
    .A2(net1028));
 sg13g2_nor2_1 _5241_ (.A(_1703_),
    .B(_1705_),
    .Y(_1706_));
 sg13g2_xnor2_1 _5242_ (.Y(_1707_),
    .A(_1703_),
    .B(_1705_));
 sg13g2_o21ai_1 _5243_ (.B1(net947),
    .Y(_1708_),
    .A1(net1040),
    .A2(net390));
 sg13g2_a21oi_1 _5244_ (.A1(net1040),
    .A2(_1707_),
    .Y(_0190_),
    .B1(_1708_));
 sg13g2_mux2_1 _5245_ (.A0(_1702_),
    .A1(net1029),
    .S(_1706_),
    .X(_1709_));
 sg13g2_nor2_1 _5246_ (.A(net991),
    .B(_1709_),
    .Y(_1710_));
 sg13g2_xnor2_1 _5247_ (.Y(_1711_),
    .A(net296),
    .B(_1710_));
 sg13g2_nor2_1 _5248_ (.A(net1065),
    .B(_1711_),
    .Y(_0191_));
 sg13g2_and2_1 _5249_ (.A(net1027),
    .B(\i_collision.vx[1] ),
    .X(_1712_));
 sg13g2_a22oi_1 _5250_ (.Y(_1713_),
    .B1(_1712_),
    .B2(_2397_),
    .A2(_2434_),
    .A1(_2396_));
 sg13g2_nor2b_1 _5251_ (.A(_1713_),
    .B_N(\center_x[0] ),
    .Y(_1714_));
 sg13g2_xnor2_1 _5252_ (.Y(_1715_),
    .A(\center_x[0] ),
    .B(_1713_));
 sg13g2_inv_1 _5253_ (.Y(_1716_),
    .A(_1715_));
 sg13g2_and3_1 _5254_ (.X(_1717_),
    .A(_1647_),
    .B(_1649_),
    .C(_1716_));
 sg13g2_a21oi_1 _5255_ (.A1(_1647_),
    .A2(_1649_),
    .Y(_1718_),
    .B1(_1716_));
 sg13g2_or2_1 _5256_ (.X(_1719_),
    .B(_1718_),
    .A(_1717_));
 sg13g2_o21ai_1 _5257_ (.B1(net948),
    .Y(_1720_),
    .A1(net1045),
    .A2(net497));
 sg13g2_a21oi_1 _5258_ (.A1(net1045),
    .A2(_1719_),
    .Y(_0192_),
    .B1(_1720_));
 sg13g2_xor2_1 _5259_ (.B(\i_collision.vx[1] ),
    .A(net1027),
    .X(_1721_));
 sg13g2_nand2b_1 _5260_ (.Y(_1722_),
    .B(_1721_),
    .A_N(_1644_));
 sg13g2_nand2_1 _5261_ (.Y(_1723_),
    .A(\center_x[1] ),
    .B(_1722_));
 sg13g2_xor2_1 _5262_ (.B(_1722_),
    .A(\center_x[1] ),
    .X(_1724_));
 sg13g2_or3_1 _5263_ (.A(_1714_),
    .B(_1718_),
    .C(_1724_),
    .X(_1725_));
 sg13g2_o21ai_1 _5264_ (.B1(_1724_),
    .Y(_1726_),
    .A1(_1714_),
    .A2(_1718_));
 sg13g2_a21oi_1 _5265_ (.A1(_1725_),
    .A2(_1726_),
    .Y(_1727_),
    .B1(net993));
 sg13g2_o21ai_1 _5266_ (.B1(net948),
    .Y(_1728_),
    .A1(net1045),
    .A2(net521));
 sg13g2_nor2_1 _5267_ (.A(_1727_),
    .B(_1728_),
    .Y(_0193_));
 sg13g2_xnor2_1 _5268_ (.Y(_1729_),
    .A(\center_x[2] ),
    .B(_1721_));
 sg13g2_and3_1 _5269_ (.X(_1730_),
    .A(_1723_),
    .B(_1726_),
    .C(_1729_));
 sg13g2_a21oi_1 _5270_ (.A1(_1723_),
    .A2(_1726_),
    .Y(_1731_),
    .B1(_1729_));
 sg13g2_o21ai_1 _5271_ (.B1(net1044),
    .Y(_1732_),
    .A1(_1730_),
    .A2(_1731_));
 sg13g2_o21ai_1 _5272_ (.B1(_1732_),
    .Y(_1733_),
    .A1(net1044),
    .A2(net435));
 sg13g2_nor2_1 _5273_ (.A(_1629_),
    .B(_1733_),
    .Y(_0194_));
 sg13g2_a21oi_2 _5274_ (.B1(_1731_),
    .Y(_1734_),
    .A2(_1721_),
    .A1(\center_x[2] ));
 sg13g2_xnor2_1 _5275_ (.Y(_1735_),
    .A(\center_x[3] ),
    .B(net1027));
 sg13g2_xnor2_1 _5276_ (.Y(_1736_),
    .A(_1734_),
    .B(_1735_));
 sg13g2_o21ai_1 _5277_ (.B1(net948),
    .Y(_1737_),
    .A1(net1044),
    .A2(net508));
 sg13g2_a21oi_1 _5278_ (.A1(net1044),
    .A2(_1736_),
    .Y(_0195_),
    .B1(_1737_));
 sg13g2_xnor2_1 _5279_ (.Y(_1738_),
    .A(\center_x[4] ),
    .B(net1025));
 sg13g2_o21ai_1 _5280_ (.B1(_1734_),
    .Y(_1739_),
    .A1(_2395_),
    .A2(_2396_));
 sg13g2_o21ai_1 _5281_ (.B1(_1739_),
    .Y(_1740_),
    .A1(\center_x[3] ),
    .A2(net1026));
 sg13g2_nor2_1 _5282_ (.A(_1738_),
    .B(_1740_),
    .Y(_1741_));
 sg13g2_xnor2_1 _5283_ (.Y(_1742_),
    .A(_1738_),
    .B(_1740_));
 sg13g2_o21ai_1 _5284_ (.B1(_1628_),
    .Y(_1743_),
    .A1(net1043),
    .A2(net441));
 sg13g2_a21oi_1 _5285_ (.A1(net1043),
    .A2(_1742_),
    .Y(_0196_),
    .B1(_1743_));
 sg13g2_nor2_1 _5286_ (.A(\center_x[5] ),
    .B(net1026),
    .Y(_1744_));
 sg13g2_a21oi_1 _5287_ (.A1(\center_x[4] ),
    .A2(net1025),
    .Y(_1745_),
    .B1(_1741_));
 sg13g2_nand2_1 _5288_ (.Y(_1746_),
    .A(\center_x[5] ),
    .B(net1026));
 sg13g2_and2_1 _5289_ (.A(_1745_),
    .B(_1746_),
    .X(_1747_));
 sg13g2_nand2b_1 _5290_ (.Y(_1748_),
    .B(_1746_),
    .A_N(_1744_));
 sg13g2_xnor2_1 _5291_ (.Y(_1749_),
    .A(_1745_),
    .B(_1748_));
 sg13g2_o21ai_1 _5292_ (.B1(net948),
    .Y(_1750_),
    .A1(net1043),
    .A2(net443));
 sg13g2_a21oi_1 _5293_ (.A1(net1043),
    .A2(_1749_),
    .Y(_0197_),
    .B1(_1750_));
 sg13g2_xnor2_1 _5294_ (.Y(_1751_),
    .A(\center_x[6] ),
    .B(net1025));
 sg13g2_o21ai_1 _5295_ (.B1(_1751_),
    .Y(_1752_),
    .A1(_1744_),
    .A2(_1747_));
 sg13g2_nor3_1 _5296_ (.A(_1744_),
    .B(_1747_),
    .C(_1751_),
    .Y(_1753_));
 sg13g2_nand2_1 _5297_ (.Y(_1754_),
    .A(net1043),
    .B(_1752_));
 sg13g2_a21oi_1 _5298_ (.A1(net993),
    .A2(net477),
    .Y(_1755_),
    .B1(_1629_));
 sg13g2_o21ai_1 _5299_ (.B1(_1755_),
    .Y(_0198_),
    .A1(_1753_),
    .A2(_1754_));
 sg13g2_a21o_1 _5300_ (.A2(net1025),
    .A1(\center_x[6] ),
    .B1(_1753_),
    .X(_1756_));
 sg13g2_a21o_1 _5301_ (.A2(net1025),
    .A1(\center_x[7] ),
    .B1(_1756_),
    .X(_1757_));
 sg13g2_xor2_1 _5302_ (.B(net1025),
    .A(\center_x[7] ),
    .X(_1758_));
 sg13g2_xnor2_1 _5303_ (.Y(_1759_),
    .A(_1756_),
    .B(_1758_));
 sg13g2_o21ai_1 _5304_ (.B1(net948),
    .Y(_1760_),
    .A1(net1043),
    .A2(net479));
 sg13g2_a21oi_1 _5305_ (.A1(net1043),
    .A2(_1759_),
    .Y(_0199_),
    .B1(_1760_));
 sg13g2_nand2b_1 _5306_ (.Y(_1761_),
    .B(net1025),
    .A_N(\center_x[8] ));
 sg13g2_nand2_1 _5307_ (.Y(_1762_),
    .A(\center_x[8] ),
    .B(_2396_));
 sg13g2_nand2_1 _5308_ (.Y(_1763_),
    .A(_1761_),
    .B(_1762_));
 sg13g2_o21ai_1 _5309_ (.B1(_1757_),
    .Y(_1764_),
    .A1(\center_x[7] ),
    .A2(net1025));
 sg13g2_xor2_1 _5310_ (.B(_1764_),
    .A(_1763_),
    .X(_1765_));
 sg13g2_a21oi_1 _5311_ (.A1(net993),
    .A2(net469),
    .Y(_1766_),
    .B1(_1629_));
 sg13g2_o21ai_1 _5312_ (.B1(_1766_),
    .Y(_0200_),
    .A1(net993),
    .A2(_1765_));
 sg13g2_or2_1 _5313_ (.X(_1767_),
    .B(_1764_),
    .A(_1762_));
 sg13g2_o21ai_1 _5314_ (.B1(_1767_),
    .Y(_1768_),
    .A1(_1757_),
    .A2(_1761_));
 sg13g2_and2_1 _5315_ (.A(net1043),
    .B(_1768_),
    .X(_1769_));
 sg13g2_o21ai_1 _5316_ (.B1(net948),
    .Y(_1770_),
    .A1(net304),
    .A2(_1769_));
 sg13g2_a21oi_1 _5317_ (.A1(net304),
    .A2(_1769_),
    .Y(_0201_),
    .B1(_1770_));
 sg13g2_and2_1 _5318_ (.A(net995),
    .B(net1005),
    .X(_1771_));
 sg13g2_and2_1 _5319_ (.A(net1042),
    .B(_1771_),
    .X(_1772_));
 sg13g2_o21ai_1 _5320_ (.B1(net947),
    .Y(_1773_),
    .A1(net251),
    .A2(_1772_));
 sg13g2_a21oi_1 _5321_ (.A1(net251),
    .A2(_1772_),
    .Y(_0202_),
    .B1(_1773_));
 sg13g2_nand2_1 _5322_ (.Y(_1774_),
    .A(net251),
    .B(_1771_));
 sg13g2_a21o_1 _5323_ (.A2(_1771_),
    .A1(_2374_),
    .B1(net949),
    .X(_1775_));
 sg13g2_or2_1 _5324_ (.X(_1776_),
    .B(_1775_),
    .A(_2394_));
 sg13g2_xnor2_1 _5325_ (.Y(_1777_),
    .A(_2394_),
    .B(_1775_));
 sg13g2_or2_1 _5326_ (.X(_1778_),
    .B(_1777_),
    .A(_1774_));
 sg13g2_xnor2_1 _5327_ (.Y(_1779_),
    .A(_1774_),
    .B(_1777_));
 sg13g2_o21ai_1 _5328_ (.B1(net946),
    .Y(_1780_),
    .A1(net1038),
    .A2(net305));
 sg13g2_a21oi_1 _5329_ (.A1(net1038),
    .A2(_1779_),
    .Y(_0203_),
    .B1(_1780_));
 sg13g2_and2_1 _5330_ (.A(net1001),
    .B(net1005),
    .X(_1781_));
 sg13g2_nand2_1 _5331_ (.Y(_1782_),
    .A(_2373_),
    .B(_1781_));
 sg13g2_o21ai_1 _5332_ (.B1(_1782_),
    .Y(_1783_),
    .A1(net1001),
    .A2(_0051_));
 sg13g2_and2_1 _5333_ (.A(\i_kinematics.phi[2] ),
    .B(_1783_),
    .X(_1784_));
 sg13g2_xor2_1 _5334_ (.B(_1783_),
    .A(\i_kinematics.phi[2] ),
    .X(_1785_));
 sg13g2_inv_1 _5335_ (.Y(_1786_),
    .A(_1785_));
 sg13g2_and3_1 _5336_ (.X(_1787_),
    .A(_1776_),
    .B(_1778_),
    .C(_1786_));
 sg13g2_a21oi_1 _5337_ (.A1(_1776_),
    .A2(_1778_),
    .Y(_1788_),
    .B1(_1786_));
 sg13g2_or2_1 _5338_ (.X(_1789_),
    .B(_1788_),
    .A(_1787_));
 sg13g2_o21ai_1 _5339_ (.B1(net946),
    .Y(_1790_),
    .A1(net1038),
    .A2(net333));
 sg13g2_a21oi_1 _5340_ (.A1(net1038),
    .A2(_1789_),
    .Y(_0204_),
    .B1(_1790_));
 sg13g2_xnor2_1 _5341_ (.Y(_1791_),
    .A(net998),
    .B(net1005));
 sg13g2_inv_1 _5342_ (.Y(_1792_),
    .A(_1791_));
 sg13g2_nor3_1 _5343_ (.A(\i_kinematics.phi[3] ),
    .B(net949),
    .C(_1791_),
    .Y(_1793_));
 sg13g2_o21ai_1 _5344_ (.B1(\i_kinematics.phi[3] ),
    .Y(_1794_),
    .A1(net949),
    .A2(_1791_));
 sg13g2_nor2b_1 _5345_ (.A(_1793_),
    .B_N(_1794_),
    .Y(_1795_));
 sg13g2_or3_1 _5346_ (.A(_1784_),
    .B(_1788_),
    .C(_1795_),
    .X(_1796_));
 sg13g2_o21ai_1 _5347_ (.B1(_1795_),
    .Y(_1797_),
    .A1(_1784_),
    .A2(_1788_));
 sg13g2_a21oi_1 _5348_ (.A1(_1796_),
    .A2(_1797_),
    .Y(_1798_),
    .B1(net992));
 sg13g2_o21ai_1 _5349_ (.B1(net946),
    .Y(_1799_),
    .A1(net1037),
    .A2(net518));
 sg13g2_nor2_1 _5350_ (.A(_1798_),
    .B(_1799_),
    .Y(_0205_));
 sg13g2_xor2_1 _5351_ (.B(_1791_),
    .A(\i_kinematics.phi[4] ),
    .X(_1800_));
 sg13g2_and3_1 _5352_ (.X(_1801_),
    .A(_1794_),
    .B(_1797_),
    .C(_1800_));
 sg13g2_a21oi_1 _5353_ (.A1(_1794_),
    .A2(_1797_),
    .Y(_1802_),
    .B1(_1800_));
 sg13g2_o21ai_1 _5354_ (.B1(net1037),
    .Y(_1803_),
    .A1(_1801_),
    .A2(_1802_));
 sg13g2_o21ai_1 _5355_ (.B1(_1803_),
    .Y(_1804_),
    .A1(net1038),
    .A2(net514));
 sg13g2_nor2_1 _5356_ (.A(net1065),
    .B(_1804_),
    .Y(_0206_));
 sg13g2_a21oi_1 _5357_ (.A1(\i_kinematics.phi[4] ),
    .A2(_1792_),
    .Y(_1805_),
    .B1(_1802_));
 sg13g2_xnor2_1 _5358_ (.Y(_1806_),
    .A(net998),
    .B(\i_kinematics.phi[5] ));
 sg13g2_xnor2_1 _5359_ (.Y(_1807_),
    .A(_1805_),
    .B(_1806_));
 sg13g2_o21ai_1 _5360_ (.B1(net946),
    .Y(_1808_),
    .A1(net1037),
    .A2(net494));
 sg13g2_a21oi_1 _5361_ (.A1(net1037),
    .A2(_1807_),
    .Y(_0207_),
    .B1(_1808_));
 sg13g2_nand2_1 _5362_ (.Y(_1809_),
    .A(net998),
    .B(\i_kinematics.phi[6] ));
 sg13g2_xnor2_1 _5363_ (.Y(_1810_),
    .A(net998),
    .B(\i_kinematics.phi[6] ));
 sg13g2_o21ai_1 _5364_ (.B1(_1805_),
    .Y(_1811_),
    .A1(_2374_),
    .A2(_2393_));
 sg13g2_o21ai_1 _5365_ (.B1(_1811_),
    .Y(_1812_),
    .A1(net998),
    .A2(\i_kinematics.phi[5] ));
 sg13g2_xnor2_1 _5366_ (.Y(_1813_),
    .A(_1810_),
    .B(_1812_));
 sg13g2_o21ai_1 _5367_ (.B1(net946),
    .Y(_1814_),
    .A1(net1037),
    .A2(net458));
 sg13g2_a21oi_1 _5368_ (.A1(net1037),
    .A2(_1813_),
    .Y(_0208_),
    .B1(_1814_));
 sg13g2_xor2_1 _5369_ (.B(\i_kinematics.phi[7] ),
    .A(net998),
    .X(_1815_));
 sg13g2_o21ai_1 _5370_ (.B1(_1809_),
    .Y(_1816_),
    .A1(_1810_),
    .A2(_1812_));
 sg13g2_xnor2_1 _5371_ (.Y(_1817_),
    .A(_1815_),
    .B(_1816_));
 sg13g2_o21ai_1 _5372_ (.B1(net946),
    .Y(_1818_),
    .A1(net1037),
    .A2(net492));
 sg13g2_a21oi_1 _5373_ (.A1(net1037),
    .A2(_1817_),
    .Y(_0209_),
    .B1(_1818_));
 sg13g2_nor2_1 _5374_ (.A(_1493_),
    .B(_1500_),
    .Y(_1819_));
 sg13g2_o21ai_1 _5375_ (.B1(_1816_),
    .Y(_1820_),
    .A1(net998),
    .A2(\i_kinematics.phi[7] ));
 sg13g2_inv_1 _5376_ (.Y(_1821_),
    .A(_1820_));
 sg13g2_a21oi_1 _5377_ (.A1(net999),
    .A2(\i_kinematics.phi[7] ),
    .Y(_1822_),
    .B1(_1821_));
 sg13g2_nand2b_1 _5378_ (.Y(_1823_),
    .B(_1819_),
    .A_N(_1822_));
 sg13g2_xor2_1 _5379_ (.B(_1822_),
    .A(_1819_),
    .X(_1824_));
 sg13g2_a21oi_1 _5380_ (.A1(net992),
    .A2(net1023),
    .Y(_1825_),
    .B1(net1065));
 sg13g2_o21ai_1 _5381_ (.B1(_1825_),
    .Y(_0210_),
    .A1(net992),
    .A2(_1824_));
 sg13g2_nand2_1 _5382_ (.Y(_1826_),
    .A(_1501_),
    .B(_1823_));
 sg13g2_xor2_1 _5383_ (.B(net543),
    .A(net999),
    .X(_1827_));
 sg13g2_nand2_1 _5384_ (.Y(_1828_),
    .A(net1039),
    .B(_1827_));
 sg13g2_o21ai_1 _5385_ (.B1(net946),
    .Y(_1829_),
    .A1(net1039),
    .A2(net1020));
 sg13g2_nor3_1 _5386_ (.A(net992),
    .B(_1826_),
    .C(_1827_),
    .Y(_1830_));
 sg13g2_a21oi_1 _5387_ (.A1(_1501_),
    .A2(_1823_),
    .Y(_1831_),
    .B1(_1828_));
 sg13g2_nor3_1 _5388_ (.A(_1829_),
    .B(_1830_),
    .C(_1831_),
    .Y(_0211_));
 sg13g2_a221oi_1 _5389_ (.B2(_2392_),
    .C1(_1828_),
    .B1(_1826_),
    .A1(_2374_),
    .Y(_1832_),
    .A2(_1823_));
 sg13g2_o21ai_1 _5390_ (.B1(net946),
    .Y(_1833_),
    .A1(net369),
    .A2(_1832_));
 sg13g2_a21oi_1 _5391_ (.A1(net369),
    .A2(_1832_),
    .Y(_0212_),
    .B1(_1833_));
 sg13g2_a21oi_1 _5392_ (.A1(net877),
    .A2(net903),
    .Y(_1834_),
    .B1(_0401_));
 sg13g2_nand2_1 _5393_ (.Y(_1835_),
    .A(net909),
    .B(net904));
 sg13g2_o21ai_1 _5394_ (.B1(_1835_),
    .Y(_1836_),
    .A1(net904),
    .A2(_2704_));
 sg13g2_xor2_1 _5395_ (.B(_1836_),
    .A(_0012_),
    .X(_1837_));
 sg13g2_o21ai_1 _5396_ (.B1(net983),
    .Y(_1838_),
    .A1(net311),
    .A2(net869));
 sg13g2_a21oi_1 _5397_ (.A1(net869),
    .A2(_1837_),
    .Y(_0213_),
    .B1(_1838_));
 sg13g2_nand3_1 _5398_ (.B(_2705_),
    .C(_2727_),
    .A(_0012_),
    .Y(_1839_));
 sg13g2_nand3_1 _5399_ (.B(_2728_),
    .C(_1839_),
    .A(net900),
    .Y(_1840_));
 sg13g2_xnor2_1 _5400_ (.Y(_1841_),
    .A(_2572_),
    .B(_2575_));
 sg13g2_nor2_1 _5401_ (.A(net900),
    .B(_1841_),
    .Y(_1842_));
 sg13g2_nand2_1 _5402_ (.Y(_1843_),
    .A(net869),
    .B(_1840_));
 sg13g2_nor2_1 _5403_ (.A(_1842_),
    .B(_1843_),
    .Y(_1844_));
 sg13g2_o21ai_1 _5404_ (.B1(net983),
    .Y(_1845_),
    .A1(net336),
    .A2(net869));
 sg13g2_nor2_1 _5405_ (.A(_1844_),
    .B(_1845_),
    .Y(_0214_));
 sg13g2_nor2_1 _5406_ (.A(_2577_),
    .B(_2580_),
    .Y(_1846_));
 sg13g2_nand3_1 _5407_ (.B(_2728_),
    .C(_2730_),
    .A(_2726_),
    .Y(_1847_));
 sg13g2_and2_1 _5408_ (.A(net900),
    .B(_2731_),
    .X(_1848_));
 sg13g2_nor2_1 _5409_ (.A(net900),
    .B(_1846_),
    .Y(_1849_));
 sg13g2_a22oi_1 _5410_ (.Y(_1850_),
    .B1(_1849_),
    .B2(_2581_),
    .A2(_1848_),
    .A1(_1847_));
 sg13g2_o21ai_1 _5411_ (.B1(net983),
    .Y(_1851_),
    .A1(net377),
    .A2(net870));
 sg13g2_a21oi_1 _5412_ (.A1(net870),
    .A2(_1850_),
    .Y(_0215_),
    .B1(_1851_));
 sg13g2_a21oi_1 _5413_ (.A1(_2571_),
    .A2(_2583_),
    .Y(_1852_),
    .B1(net900));
 sg13g2_nand2b_1 _5414_ (.Y(_1853_),
    .B(_1852_),
    .A_N(_2584_));
 sg13g2_nand3_1 _5415_ (.B(_2732_),
    .C(_2733_),
    .A(_2731_),
    .Y(_1854_));
 sg13g2_nand3_1 _5416_ (.B(_2734_),
    .C(_1854_),
    .A(net900),
    .Y(_1855_));
 sg13g2_nand3_1 _5417_ (.B(_1853_),
    .C(_1855_),
    .A(net871),
    .Y(_1856_));
 sg13g2_o21ai_1 _5418_ (.B1(_1856_),
    .Y(_1857_),
    .A1(net320),
    .A2(net871));
 sg13g2_nor2_1 _5419_ (.A(net976),
    .B(_1857_),
    .Y(_0216_));
 sg13g2_and3_1 _5420_ (.X(_1858_),
    .A(_2722_),
    .B(_2734_),
    .C(_2736_));
 sg13g2_nor3_1 _5421_ (.A(net903),
    .B(_2737_),
    .C(_1858_),
    .Y(_1859_));
 sg13g2_nor3_1 _5422_ (.A(_2570_),
    .B(_2584_),
    .C(_2586_),
    .Y(_1860_));
 sg13g2_nand2_1 _5423_ (.Y(_1861_),
    .A(_2587_),
    .B(net903));
 sg13g2_o21ai_1 _5424_ (.B1(net871),
    .Y(_1862_),
    .A1(_1860_),
    .A2(_1861_));
 sg13g2_nor2_1 _5425_ (.A(net313),
    .B(net871),
    .Y(_1863_));
 sg13g2_o21ai_1 _5426_ (.B1(net983),
    .Y(_1864_),
    .A1(_1859_),
    .A2(_1862_));
 sg13g2_nor2_1 _5427_ (.A(_1863_),
    .B(_1864_),
    .Y(_0217_));
 sg13g2_nand2_1 _5428_ (.Y(_1865_),
    .A(net909),
    .B(net900));
 sg13g2_o21ai_1 _5429_ (.B1(_1865_),
    .Y(_1866_),
    .A1(net900),
    .A2(_2704_));
 sg13g2_xor2_1 _5430_ (.B(_1866_),
    .A(_0025_),
    .X(_1867_));
 sg13g2_o21ai_1 _5431_ (.B1(net983),
    .Y(_1868_),
    .A1(net285),
    .A2(net869));
 sg13g2_a21oi_1 _5432_ (.A1(net869),
    .A2(_1867_),
    .Y(_0218_),
    .B1(_1868_));
 sg13g2_a21oi_1 _5433_ (.A1(_2788_),
    .A2(_2790_),
    .Y(_1869_),
    .B1(net904));
 sg13g2_o21ai_1 _5434_ (.B1(_1869_),
    .Y(_1870_),
    .A1(_2788_),
    .A2(_2790_));
 sg13g2_o21ai_1 _5435_ (.B1(net904),
    .Y(_1871_),
    .A1(_0299_),
    .A2(_0300_));
 sg13g2_a21o_1 _5436_ (.A2(_0300_),
    .A1(_0299_),
    .B1(_1871_),
    .X(_1872_));
 sg13g2_and3_1 _5437_ (.X(_1873_),
    .A(net869),
    .B(_1870_),
    .C(_1872_));
 sg13g2_o21ai_1 _5438_ (.B1(net983),
    .Y(_1874_),
    .A1(net321),
    .A2(net869));
 sg13g2_nor2_1 _5439_ (.A(_1873_),
    .B(_1874_),
    .Y(_0219_));
 sg13g2_a21o_1 _5440_ (.A2(_2792_),
    .A1(_2791_),
    .B1(net904),
    .X(_1875_));
 sg13g2_o21ai_1 _5441_ (.B1(net870),
    .Y(_1876_),
    .A1(_2793_),
    .A2(_1875_));
 sg13g2_xor2_1 _5442_ (.B(_0302_),
    .A(_0301_),
    .X(_1877_));
 sg13g2_a21oi_1 _5443_ (.A1(net904),
    .A2(_1877_),
    .Y(_1878_),
    .B1(_1876_));
 sg13g2_o21ai_1 _5444_ (.B1(net983),
    .Y(_1879_),
    .A1(net436),
    .A2(net870));
 sg13g2_nor2_1 _5445_ (.A(_1878_),
    .B(_1879_),
    .Y(_0220_));
 sg13g2_nor2_1 _5446_ (.A(_2795_),
    .B(_2796_),
    .Y(_1880_));
 sg13g2_nor2_1 _5447_ (.A(net903),
    .B(_1880_),
    .Y(_1881_));
 sg13g2_a221oi_1 _5448_ (.B2(_1881_),
    .C1(_0401_),
    .B1(_2797_),
    .A1(net877),
    .Y(_1882_),
    .A2(net903));
 sg13g2_o21ai_1 _5449_ (.B1(net903),
    .Y(_1883_),
    .A1(_0304_),
    .A2(_0305_));
 sg13g2_a21o_1 _5450_ (.A2(_0305_),
    .A1(_0304_),
    .B1(_1883_),
    .X(_1884_));
 sg13g2_o21ai_1 _5451_ (.B1(net984),
    .Y(_1885_),
    .A1(net342),
    .A2(net871));
 sg13g2_a21oi_1 _5452_ (.A1(_1882_),
    .A2(_1884_),
    .Y(_0221_),
    .B1(net343));
 sg13g2_nor2_1 _5453_ (.A(_0307_),
    .B(_0308_),
    .Y(_1886_));
 sg13g2_nor3_1 _5454_ (.A(net901),
    .B(_0309_),
    .C(_1886_),
    .Y(_1887_));
 sg13g2_xor2_1 _5455_ (.B(_2801_),
    .A(_2799_),
    .X(_1888_));
 sg13g2_o21ai_1 _5456_ (.B1(net871),
    .Y(_1889_),
    .A1(net903),
    .A2(_1888_));
 sg13g2_nor2_1 _5457_ (.A(_1887_),
    .B(_1889_),
    .Y(_1890_));
 sg13g2_o21ai_1 _5458_ (.B1(net983),
    .Y(_1891_),
    .A1(net389),
    .A2(net871));
 sg13g2_nor2_1 _5459_ (.A(_1890_),
    .B(_1891_),
    .Y(_0222_));
 sg13g2_nand2_2 _5460_ (.Y(_1892_),
    .A(net989),
    .B(_0343_));
 sg13g2_or2_1 _5461_ (.X(_1893_),
    .B(net980),
    .A(_0063_));
 sg13g2_o21ai_1 _5462_ (.B1(_1893_),
    .Y(_1894_),
    .A1(\center_x[0] ),
    .A2(net989));
 sg13g2_nor2_1 _5463_ (.A(net351),
    .B(_1892_),
    .Y(_1895_));
 sg13g2_a21oi_1 _5464_ (.A1(_1892_),
    .A2(_1894_),
    .Y(_0223_),
    .B1(_1895_));
 sg13g2_o21ai_1 _5465_ (.B1(net989),
    .Y(_1896_),
    .A1(\i_transform.track_x[0] ),
    .A2(\i_transform.track_x[1] ));
 sg13g2_a21oi_1 _5466_ (.A1(net351),
    .A2(net471),
    .Y(_1897_),
    .B1(_1896_));
 sg13g2_a21oi_1 _5467_ (.A1(\center_x[1] ),
    .A2(net980),
    .Y(_1898_),
    .B1(_1897_));
 sg13g2_nor2_1 _5468_ (.A(net471),
    .B(_1892_),
    .Y(_1899_));
 sg13g2_a21oi_1 _5469_ (.A1(_1892_),
    .A2(_1898_),
    .Y(_0224_),
    .B1(_1899_));
 sg13g2_and4_1 _5470_ (.A(\i_transform.track_x[0] ),
    .B(\i_transform.track_x[1] ),
    .C(net875),
    .D(_0341_),
    .X(_1900_));
 sg13g2_nand3_1 _5471_ (.B(\i_transform.track_x[1] ),
    .C(\i_transform.track_x[2] ),
    .A(\i_transform.track_x[0] ),
    .Y(_1901_));
 sg13g2_nor2_2 _5472_ (.A(net435),
    .B(net990),
    .Y(_1902_));
 sg13g2_xnor2_1 _5473_ (.Y(_1903_),
    .A(net453),
    .B(_1900_));
 sg13g2_a21oi_1 _5474_ (.A1(net989),
    .A2(net454),
    .Y(_0225_),
    .B1(_1902_));
 sg13g2_or2_2 _5475_ (.X(_1904_),
    .B(_1901_),
    .A(_2429_));
 sg13g2_a21oi_1 _5476_ (.A1(_2429_),
    .A2(_1901_),
    .Y(_1905_),
    .B1(net980));
 sg13g2_a22oi_1 _5477_ (.Y(_1906_),
    .B1(_1904_),
    .B2(_1905_),
    .A2(net980),
    .A1(\center_x[3] ));
 sg13g2_nor2_1 _5478_ (.A(net264),
    .B(_1892_),
    .Y(_1907_));
 sg13g2_a21oi_1 _5479_ (.A1(_1892_),
    .A2(_1906_),
    .Y(_0226_),
    .B1(_1907_));
 sg13g2_nor2_1 _5480_ (.A(\center_x[4] ),
    .B(net989),
    .Y(_1908_));
 sg13g2_nor2_1 _5481_ (.A(_0343_),
    .B(_1904_),
    .Y(_1909_));
 sg13g2_xnor2_1 _5482_ (.Y(_1910_),
    .A(net401),
    .B(_1909_));
 sg13g2_a21oi_1 _5483_ (.A1(net989),
    .A2(_1910_),
    .Y(_0227_),
    .B1(_1908_));
 sg13g2_and2_1 _5484_ (.A(net1076),
    .B(net239),
    .X(_0228_));
 sg13g2_and2_1 _5485_ (.A(net373),
    .B(\i_orchestrator.sample_counter[1] ),
    .X(_1911_));
 sg13g2_nor3_1 _5486_ (.A(net1066),
    .B(net374),
    .C(_1911_),
    .Y(_0229_));
 sg13g2_nor2_1 _5487_ (.A(net301),
    .B(_1911_),
    .Y(_1912_));
 sg13g2_nand2_1 _5488_ (.Y(_1913_),
    .A(net301),
    .B(_1911_));
 sg13g2_nand2_1 _5489_ (.Y(_1914_),
    .A(net1076),
    .B(_1913_));
 sg13g2_nor2_1 _5490_ (.A(net302),
    .B(_1914_),
    .Y(_0230_));
 sg13g2_or2_1 _5491_ (.X(_1915_),
    .B(_1913_),
    .A(_2435_));
 sg13g2_nand2_1 _5492_ (.Y(_1916_),
    .A(net1076),
    .B(_1915_));
 sg13g2_a21oi_1 _5493_ (.A1(_2435_),
    .A2(_1913_),
    .Y(_0231_),
    .B1(_1916_));
 sg13g2_and2_1 _5494_ (.A(_2436_),
    .B(_1915_),
    .X(_1917_));
 sg13g2_nor2_1 _5495_ (.A(_2436_),
    .B(_1915_),
    .Y(_1918_));
 sg13g2_nor3_1 _5496_ (.A(net1066),
    .B(_1917_),
    .C(_1918_),
    .Y(_0232_));
 sg13g2_and2_1 _5497_ (.A(net334),
    .B(_1918_),
    .X(_1919_));
 sg13g2_o21ai_1 _5498_ (.B1(net1076),
    .Y(_1920_),
    .A1(net334),
    .A2(_1918_));
 sg13g2_nor2_1 _5499_ (.A(_1919_),
    .B(net335),
    .Y(_0233_));
 sg13g2_xnor2_1 _5500_ (.Y(_1921_),
    .A(net319),
    .B(_1919_));
 sg13g2_nor2_1 _5501_ (.A(net1066),
    .B(_1921_),
    .Y(_0234_));
 sg13g2_a21oi_1 _5502_ (.A1(\i_orchestrator.sample_counter[6] ),
    .A2(_1919_),
    .Y(_1922_),
    .B1(net274));
 sg13g2_nand3_1 _5503_ (.B(\i_orchestrator.sample_counter[6] ),
    .C(_1919_),
    .A(net274),
    .Y(_1923_));
 sg13g2_nand2_1 _5504_ (.Y(_1924_),
    .A(net1076),
    .B(_1923_));
 sg13g2_nor2_1 _5505_ (.A(net275),
    .B(_1924_),
    .Y(_0235_));
 sg13g2_or2_1 _5506_ (.X(_1925_),
    .B(_1923_),
    .A(_2437_));
 sg13g2_nand2_1 _5507_ (.Y(_1926_),
    .A(net1077),
    .B(_1925_));
 sg13g2_a21oi_1 _5508_ (.A1(_2437_),
    .A2(_1923_),
    .Y(_0236_),
    .B1(_1926_));
 sg13g2_xor2_1 _5509_ (.B(_1925_),
    .A(net242),
    .X(_1927_));
 sg13g2_nor2_1 _5510_ (.A(net1066),
    .B(_1927_),
    .Y(_0237_));
 sg13g2_and2_1 _5511_ (.A(_1264_),
    .B(_1322_),
    .X(_1928_));
 sg13g2_nor4_2 _5512_ (.A(\i_orchestrator.trigger_debounce ),
    .B(_1267_),
    .C(_1270_),
    .Y(_1929_),
    .D(_1928_));
 sg13g2_o21ai_1 _5513_ (.B1(net1078),
    .Y(_1930_),
    .A1(\i_orchestrator.tension[1] ),
    .A2(_1929_));
 sg13g2_a21oi_1 _5514_ (.A1(_2388_),
    .A2(_1929_),
    .Y(_0238_),
    .B1(_1930_));
 sg13g2_nand2_1 _5515_ (.Y(_1931_),
    .A(_1265_),
    .B(_1929_));
 sg13g2_nand3_1 _5516_ (.B(_1265_),
    .C(_1929_),
    .A(net322),
    .Y(_1932_));
 sg13g2_o21ai_1 _5517_ (.B1(net1078),
    .Y(_1933_),
    .A1(net258),
    .A2(_1929_));
 sg13g2_nor2b_1 _5518_ (.A(_1933_),
    .B_N(net323),
    .Y(_0239_));
 sg13g2_nand2b_1 _5519_ (.Y(_1934_),
    .B(net260),
    .A_N(_1929_));
 sg13g2_a21oi_1 _5520_ (.A1(_1931_),
    .A2(_1934_),
    .Y(_0240_),
    .B1(net1069));
 sg13g2_nor3_1 _5521_ (.A(\i_colors.channel[1] ),
    .B(\i_colors.channel[2] ),
    .C(_2446_),
    .Y(_1935_));
 sg13g2_inv_1 _5522_ (.Y(_1936_),
    .A(_1935_));
 sg13g2_nand2_1 _5523_ (.Y(_1937_),
    .A(\i_colors.channel[0] ),
    .B(_1935_));
 sg13g2_a21oi_1 _5524_ (.A1(net329),
    .A2(_1937_),
    .Y(_1938_),
    .B1(net1068));
 sg13g2_o21ai_1 _5525_ (.B1(_1938_),
    .Y(_0241_),
    .A1(net329),
    .A2(_1936_));
 sg13g2_o21ai_1 _5526_ (.B1(net329),
    .Y(_1939_),
    .A1(\capsule_color[1] ),
    .A2(_0044_));
 sg13g2_o21ai_1 _5527_ (.B1(\color_entropy[0] ),
    .Y(_1940_),
    .A1(\capsule_color[3] ),
    .A2(\capsule_color[2] ));
 sg13g2_nand2_1 _5528_ (.Y(_1941_),
    .A(\i_colors.capsule_color[5] ),
    .B(\color_entropy[0] ));
 sg13g2_nand3_1 _5529_ (.B(_1940_),
    .C(_1941_),
    .A(net413),
    .Y(_1942_));
 sg13g2_a21oi_1 _5530_ (.A1(_1939_),
    .A2(_1942_),
    .Y(_1943_),
    .B1(_1937_));
 sg13g2_a21oi_1 _5531_ (.A1(net413),
    .A2(_1936_),
    .Y(_1944_),
    .B1(_1943_));
 sg13g2_nor2_1 _5532_ (.A(net1068),
    .B(net414),
    .Y(_0242_));
 sg13g2_nor3_1 _5533_ (.A(net423),
    .B(net432),
    .C(_2446_),
    .Y(_1945_));
 sg13g2_inv_1 _5534_ (.Y(_1946_),
    .A(_1945_));
 sg13g2_nand2_1 _5535_ (.Y(_1947_),
    .A(net449),
    .B(_1945_));
 sg13g2_a21oi_1 _5536_ (.A1(net1019),
    .A2(_1947_),
    .Y(_1948_),
    .B1(net1068));
 sg13g2_o21ai_1 _5537_ (.B1(_1948_),
    .Y(_0243_),
    .A1(net1019),
    .A2(_1946_));
 sg13g2_a21o_1 _5538_ (.A2(\capsule_color[1] ),
    .A1(_2387_),
    .B1(net358),
    .X(_1949_));
 sg13g2_a21oi_1 _5539_ (.A1(\capsule_color[3] ),
    .A2(net1019),
    .Y(_1950_),
    .B1(_2407_));
 sg13g2_a221oi_1 _5540_ (.B2(_1950_),
    .C1(_1947_),
    .B1(_1949_),
    .A1(_2386_),
    .Y(_1951_),
    .A2(_2387_));
 sg13g2_a21oi_1 _5541_ (.A1(net425),
    .A2(_1946_),
    .Y(_1952_),
    .B1(_1951_));
 sg13g2_nor2_1 _5542_ (.A(net1068),
    .B(_1952_),
    .Y(_0244_));
 sg13g2_or3_1 _5543_ (.A(\i_colors.channel[2] ),
    .B(\i_colors.channel[0] ),
    .C(_2446_),
    .X(_1953_));
 sg13g2_o21ai_1 _5544_ (.B1(\i_colors.capsule_color[4] ),
    .Y(_1954_),
    .A1(net339),
    .A2(_1953_));
 sg13g2_or2_1 _5545_ (.X(_1955_),
    .B(_1953_),
    .A(\i_colors.capsule_color[4] ));
 sg13g2_nand3_1 _5546_ (.B(net340),
    .C(_1955_),
    .A(net1075),
    .Y(_0245_));
 sg13g2_nor2_1 _5547_ (.A(\capsule_color[3] ),
    .B(\capsule_color[1] ),
    .Y(_1956_));
 sg13g2_or2_1 _5548_ (.X(_1957_),
    .B(_1956_),
    .A(_1940_));
 sg13g2_o21ai_1 _5549_ (.B1(net358),
    .Y(_1958_),
    .A1(_1955_),
    .A2(_1957_));
 sg13g2_a21oi_1 _5550_ (.A1(\i_colors.capsule_color[4] ),
    .A2(_0044_),
    .Y(_1959_),
    .B1(net339));
 sg13g2_o21ai_1 _5551_ (.B1(net1076),
    .Y(_1960_),
    .A1(_1953_),
    .A2(_1959_));
 sg13g2_nand2b_1 _5552_ (.Y(_0246_),
    .B(_1958_),
    .A_N(_1960_));
 sg13g2_nor2_2 _5553_ (.A(net980),
    .B(_0341_),
    .Y(_1961_));
 sg13g2_nand2b_1 _5554_ (.Y(_1962_),
    .B(_1961_),
    .A_N(\i_transform.track_x[5] ));
 sg13g2_o21ai_1 _5555_ (.B1(_1962_),
    .Y(_1963_),
    .A1(\center_x[5] ),
    .A2(net989));
 sg13g2_nand2_1 _5556_ (.Y(_1964_),
    .A(net287),
    .B(net881));
 sg13g2_nor2_1 _5557_ (.A(_0067_),
    .B(_1904_),
    .Y(_1965_));
 sg13g2_xor2_1 _5558_ (.B(_1965_),
    .A(\i_transform.track_x[5] ),
    .X(_1966_));
 sg13g2_a21oi_1 _5559_ (.A1(net875),
    .A2(_1966_),
    .Y(_1967_),
    .B1(net883));
 sg13g2_a21oi_1 _5560_ (.A1(_1964_),
    .A2(_1967_),
    .Y(_0247_),
    .B1(_1963_));
 sg13g2_a22oi_1 _5561_ (.Y(_1968_),
    .B1(_1961_),
    .B2(net525),
    .A2(net982),
    .A1(net477));
 sg13g2_nand2_1 _5562_ (.Y(_1969_),
    .A(\i_transform.track_x[5] ),
    .B(\i_transform.track_x[4] ));
 sg13g2_nor3_2 _5563_ (.A(net880),
    .B(_1904_),
    .C(_1969_),
    .Y(_1970_));
 sg13g2_nor2_1 _5564_ (.A(\i_transform.track_x[5] ),
    .B(net875),
    .Y(_1971_));
 sg13g2_nor3_1 _5565_ (.A(\i_transform.track_x[6] ),
    .B(_1970_),
    .C(_1971_),
    .Y(_1972_));
 sg13g2_o21ai_1 _5566_ (.B1(net525),
    .Y(_1973_),
    .A1(_1970_),
    .A2(_1971_));
 sg13g2_nand2_1 _5567_ (.Y(_1974_),
    .A(_0856_),
    .B(_1973_));
 sg13g2_o21ai_1 _5568_ (.B1(_1968_),
    .Y(_0248_),
    .A1(_1972_),
    .A2(_1974_));
 sg13g2_a22oi_1 _5569_ (.Y(_1975_),
    .B1(_1961_),
    .B2(net455),
    .A2(net980),
    .A1(\center_x[7] ));
 sg13g2_and2_1 _5570_ (.A(\i_transform.track_x[6] ),
    .B(_1970_),
    .X(_1976_));
 sg13g2_nor3_1 _5571_ (.A(\i_transform.track_x[6] ),
    .B(\i_transform.track_x[5] ),
    .C(net875),
    .Y(_1977_));
 sg13g2_nor2_1 _5572_ (.A(_1976_),
    .B(_1977_),
    .Y(_1978_));
 sg13g2_xor2_1 _5573_ (.B(_1978_),
    .A(net455),
    .X(_1979_));
 sg13g2_o21ai_1 _5574_ (.B1(net456),
    .Y(_0249_),
    .A1(net883),
    .A2(_1979_));
 sg13g2_a22oi_1 _5575_ (.Y(_1980_),
    .B1(_1961_),
    .B2(net467),
    .A2(net980),
    .A1(\center_x[8] ));
 sg13g2_nand2_1 _5576_ (.Y(_1981_),
    .A(\i_transform.track_x[7] ),
    .B(_1976_));
 sg13g2_nor2b_1 _5577_ (.A(\i_transform.track_x[7] ),
    .B_N(_1977_),
    .Y(_1982_));
 sg13g2_nor2_1 _5578_ (.A(\i_transform.track_x[8] ),
    .B(_1982_),
    .Y(_1983_));
 sg13g2_a21oi_1 _5579_ (.A1(\i_transform.track_x[7] ),
    .A2(_1976_),
    .Y(_1984_),
    .B1(_1982_));
 sg13g2_xor2_1 _5580_ (.B(_1984_),
    .A(net467),
    .X(_1985_));
 sg13g2_o21ai_1 _5581_ (.B1(net468),
    .Y(_0250_),
    .A1(net883),
    .A2(_1985_));
 sg13g2_a22oi_1 _5582_ (.Y(_1986_),
    .B1(_1961_),
    .B2(net299),
    .A2(net980),
    .A1(\center_x[9] ));
 sg13g2_a21oi_1 _5583_ (.A1(\i_transform.track_x[8] ),
    .A2(_1981_),
    .Y(_1987_),
    .B1(_1983_));
 sg13g2_a21oi_1 _5584_ (.A1(net299),
    .A2(_1987_),
    .Y(_1988_),
    .B1(net883));
 sg13g2_o21ai_1 _5585_ (.B1(_1988_),
    .Y(_1989_),
    .A1(net299),
    .A2(_1987_));
 sg13g2_nand2_1 _5586_ (.Y(_0251_),
    .A(net300),
    .B(_1989_));
 sg13g2_o21ai_1 _5587_ (.B1(net358),
    .Y(_1990_),
    .A1(net393),
    .A2(_1109_));
 sg13g2_a21oi_1 _5588_ (.A1(_1110_),
    .A2(net394),
    .Y(_0252_),
    .B1(_1107_));
 sg13g2_nor3_2 _5589_ (.A(\i_resonator.counter[3] ),
    .B(\i_resonator.counter[2] ),
    .C(\i_resonator.counter[1] ),
    .Y(_1991_));
 sg13g2_or3_1 _5590_ (.A(\i_resonator.counter[3] ),
    .B(\i_resonator.counter[2] ),
    .C(\i_resonator.counter[1] ),
    .X(_1992_));
 sg13g2_nand3_1 _5591_ (.B(_2433_),
    .C(_1991_),
    .A(\i_resonator.counter[0] ),
    .Y(_1993_));
 sg13g2_nor2_1 _5592_ (.A(net1008),
    .B(net1015),
    .Y(_1994_));
 sg13g2_or2_1 _5593_ (.X(_1995_),
    .B(net1014),
    .A(net1007));
 sg13g2_xnor2_1 _5594_ (.Y(_1996_),
    .A(net1006),
    .B(\i_delta_sigma.sample[7] ));
 sg13g2_xnor2_1 _5595_ (.Y(_1997_),
    .A(net1006),
    .B(\i_delta_sigma.sample[6] ));
 sg13g2_nand2_1 _5596_ (.Y(_1998_),
    .A(net1006),
    .B(\i_delta_sigma.sample[5] ));
 sg13g2_xnor2_1 _5597_ (.Y(_1999_),
    .A(net1006),
    .B(\i_delta_sigma.sample[5] ));
 sg13g2_xnor2_1 _5598_ (.Y(_2000_),
    .A(\i_resonator.v[14] ),
    .B(\i_delta_sigma.sample[4] ));
 sg13g2_nand2_1 _5599_ (.Y(_2001_),
    .A(net1011),
    .B(\i_delta_sigma.sample[3] ));
 sg13g2_xnor2_1 _5600_ (.Y(_2002_),
    .A(net1011),
    .B(\i_delta_sigma.sample[3] ));
 sg13g2_and2_1 _5601_ (.A(\i_resonator.v[12] ),
    .B(\i_delta_sigma.sample[2] ),
    .X(_2003_));
 sg13g2_xor2_1 _5602_ (.B(\i_delta_sigma.sample[2] ),
    .A(\i_resonator.v[12] ),
    .X(_2004_));
 sg13g2_nand2_1 _5603_ (.Y(_2005_),
    .A(\i_resonator.v[11] ),
    .B(\i_delta_sigma.sample[1] ));
 sg13g2_nand2_1 _5604_ (.Y(_2006_),
    .A(net1012),
    .B(\i_delta_sigma.sample[0] ));
 sg13g2_xnor2_1 _5605_ (.Y(_2007_),
    .A(\i_resonator.v[11] ),
    .B(\i_delta_sigma.sample[1] ));
 sg13g2_o21ai_1 _5606_ (.B1(_2005_),
    .Y(_2008_),
    .A1(_2006_),
    .A2(_2007_));
 sg13g2_a21oi_1 _5607_ (.A1(_2004_),
    .A2(_2008_),
    .Y(_2009_),
    .B1(_2003_));
 sg13g2_or2_1 _5608_ (.X(_2010_),
    .B(_2009_),
    .A(_2002_));
 sg13g2_a21oi_1 _5609_ (.A1(_2001_),
    .A2(_2010_),
    .Y(_2011_),
    .B1(_2000_));
 sg13g2_a21oi_1 _5610_ (.A1(\i_resonator.v[14] ),
    .A2(\i_delta_sigma.sample[4] ),
    .Y(_2012_),
    .B1(_2011_));
 sg13g2_or2_1 _5611_ (.X(_2013_),
    .B(_2012_),
    .A(_1999_));
 sg13g2_a21oi_1 _5612_ (.A1(_1998_),
    .A2(_2013_),
    .Y(_2014_),
    .B1(_1997_));
 sg13g2_nand2b_1 _5613_ (.Y(_2015_),
    .B(_2014_),
    .A_N(_1996_));
 sg13g2_o21ai_1 _5614_ (.B1(net1006),
    .Y(_2016_),
    .A1(\i_delta_sigma.sample[7] ),
    .A2(\i_delta_sigma.sample[6] ));
 sg13g2_xnor2_1 _5615_ (.Y(_2017_),
    .A(net1006),
    .B(\i_delta_sigma.sample[8] ));
 sg13g2_a21oi_1 _5616_ (.A1(_2015_),
    .A2(_2016_),
    .Y(_2018_),
    .B1(_2017_));
 sg13g2_a21o_1 _5617_ (.A2(net1014),
    .A1(net1007),
    .B1(_2018_),
    .X(_2019_));
 sg13g2_xnor2_1 _5618_ (.Y(_2020_),
    .A(net1007),
    .B(net1014));
 sg13g2_a22oi_1 _5619_ (.Y(_2021_),
    .B1(_1995_),
    .B2(_2019_),
    .A2(\i_delta_sigma.sample[8] ),
    .A1(net1007));
 sg13g2_xor2_1 _5620_ (.B(net1013),
    .A(net1008),
    .X(_2022_));
 sg13g2_nor2b_2 _5621_ (.A(_2021_),
    .B_N(_2022_),
    .Y(_2023_));
 sg13g2_a21oi_1 _5622_ (.A1(net1008),
    .A2(net1013),
    .Y(_2024_),
    .B1(_2023_));
 sg13g2_xnor2_1 _5623_ (.Y(_2025_),
    .A(net1009),
    .B(net1015));
 sg13g2_nor2_1 _5624_ (.A(_2024_),
    .B(_2025_),
    .Y(_2026_));
 sg13g2_nor2_2 _5625_ (.A(_1994_),
    .B(_2026_),
    .Y(_2027_));
 sg13g2_nand2b_2 _5626_ (.Y(_2028_),
    .B(net1075),
    .A_N(net4));
 sg13g2_or3_2 _5627_ (.A(\i_orchestrator.trigger_resonator[1] ),
    .B(\i_orchestrator.trigger_resonator[0] ),
    .C(net1064),
    .X(_2029_));
 sg13g2_inv_1 _5628_ (.Y(_2030_),
    .A(_2029_));
 sg13g2_mux2_1 _5629_ (.A0(_2027_),
    .A1(net1018),
    .S(_1993_),
    .X(_2031_));
 sg13g2_and2_1 _5630_ (.A(net934),
    .B(_2031_),
    .X(_0253_));
 sg13g2_xnor2_1 _5631_ (.Y(_2032_),
    .A(net1012),
    .B(\i_delta_sigma.sample[0] ));
 sg13g2_nor4_2 _5632_ (.A(net994),
    .B(net1013),
    .C(_2385_),
    .Y(_2033_),
    .D(_2023_));
 sg13g2_nor2_1 _5633_ (.A(_2032_),
    .B(_2033_),
    .Y(_2034_));
 sg13g2_and2_1 _5634_ (.A(_1994_),
    .B(_2023_),
    .X(_2035_));
 sg13g2_o21ai_1 _5635_ (.B1(_2432_),
    .Y(_2036_),
    .A1(_2034_),
    .A2(net872));
 sg13g2_nand2b_1 _5636_ (.Y(_2037_),
    .B(net289),
    .A_N(\i_resonator.counter[0] ));
 sg13g2_nor3_1 _5637_ (.A(\i_resonator.counter[2] ),
    .B(\i_resonator.counter[1] ),
    .C(\i_resonator.counter[0] ),
    .Y(_2038_));
 sg13g2_a21oi_1 _5638_ (.A1(\i_resonator.counter[3] ),
    .A2(_2038_),
    .Y(_2039_),
    .B1(_2037_));
 sg13g2_nor3_2 _5639_ (.A(net1048),
    .B(_1992_),
    .C(_2039_),
    .Y(_2040_));
 sg13g2_nor3_1 _5640_ (.A(\i_orchestrator.trigger_resonator[1] ),
    .B(\i_orchestrator.trigger_resonator[0] ),
    .C(_2040_),
    .Y(_2041_));
 sg13g2_nor2_2 _5641_ (.A(net519),
    .B(net910),
    .Y(_2042_));
 sg13g2_a221oi_1 _5642_ (.B2(_2036_),
    .C1(net1064),
    .B1(_2042_),
    .A1(_2384_),
    .Y(_0254_),
    .A2(net911));
 sg13g2_xnor2_1 _5643_ (.Y(_2043_),
    .A(_2006_),
    .B(_2007_));
 sg13g2_nor2_1 _5644_ (.A(_2033_),
    .B(_2043_),
    .Y(_2044_));
 sg13g2_o21ai_1 _5645_ (.B1(_2042_),
    .Y(_2045_),
    .A1(_2035_),
    .A2(_2044_));
 sg13g2_a21oi_1 _5646_ (.A1(net490),
    .A2(net911),
    .Y(_2046_),
    .B1(net486));
 sg13g2_a21oi_1 _5647_ (.A1(_2045_),
    .A2(_2046_),
    .Y(_0255_),
    .B1(net1064));
 sg13g2_xnor2_1 _5648_ (.Y(_2047_),
    .A(_2004_),
    .B(_2008_));
 sg13g2_nor2_1 _5649_ (.A(_2033_),
    .B(_2047_),
    .Y(_2048_));
 sg13g2_and2_2 _5650_ (.A(_2432_),
    .B(_2040_),
    .X(_2049_));
 sg13g2_o21ai_1 _5651_ (.B1(_2049_),
    .Y(_2050_),
    .A1(_2035_),
    .A2(_2048_));
 sg13g2_a21oi_1 _5652_ (.A1(net438),
    .A2(net911),
    .Y(_2051_),
    .B1(\i_orchestrator.trigger_resonator[1] ));
 sg13g2_a21oi_1 _5653_ (.A1(_2050_),
    .A2(net439),
    .Y(_0256_),
    .B1(net1064));
 sg13g2_xnor2_1 _5654_ (.Y(_2052_),
    .A(_2002_),
    .B(_2009_));
 sg13g2_nor2_1 _5655_ (.A(net873),
    .B(_2052_),
    .Y(_2053_));
 sg13g2_o21ai_1 _5656_ (.B1(_2042_),
    .Y(_2054_),
    .A1(net872),
    .A2(_2053_));
 sg13g2_a21oi_1 _5657_ (.A1(net488),
    .A2(net910),
    .Y(_2055_),
    .B1(net486));
 sg13g2_a21oi_1 _5658_ (.A1(_2054_),
    .A2(_2055_),
    .Y(_0257_),
    .B1(net1063));
 sg13g2_and3_1 _5659_ (.X(_2056_),
    .A(_2000_),
    .B(_2001_),
    .C(_2010_));
 sg13g2_nor3_1 _5660_ (.A(_2011_),
    .B(net873),
    .C(_2056_),
    .Y(_2057_));
 sg13g2_o21ai_1 _5661_ (.B1(_2049_),
    .Y(_2058_),
    .A1(net872),
    .A2(_2057_));
 sg13g2_a21oi_1 _5662_ (.A1(\i_delta_sigma.sample[4] ),
    .A2(net910),
    .Y(_2059_),
    .B1(net510));
 sg13g2_a21oi_1 _5663_ (.A1(_2058_),
    .A2(net511),
    .Y(_0258_),
    .B1(net1063));
 sg13g2_xnor2_1 _5664_ (.Y(_2060_),
    .A(_1999_),
    .B(_2012_));
 sg13g2_nor2_1 _5665_ (.A(net873),
    .B(_2060_),
    .Y(_2061_));
 sg13g2_o21ai_1 _5666_ (.B1(_2042_),
    .Y(_2062_),
    .A1(net872),
    .A2(_2061_));
 sg13g2_a21oi_1 _5667_ (.A1(\i_delta_sigma.sample[5] ),
    .A2(net910),
    .Y(_2063_),
    .B1(net486));
 sg13g2_a21oi_1 _5668_ (.A1(_2062_),
    .A2(net487),
    .Y(_0259_),
    .B1(net1063));
 sg13g2_and3_1 _5669_ (.X(_2064_),
    .A(_1997_),
    .B(_1998_),
    .C(_2013_));
 sg13g2_nor3_1 _5670_ (.A(_2014_),
    .B(net873),
    .C(_2064_),
    .Y(_2065_));
 sg13g2_o21ai_1 _5671_ (.B1(_2049_),
    .Y(_2066_),
    .A1(net872),
    .A2(_2065_));
 sg13g2_a21oi_1 _5672_ (.A1(net534),
    .A2(net910),
    .Y(_2067_),
    .B1(net510));
 sg13g2_a21oi_1 _5673_ (.A1(_2066_),
    .A2(_2067_),
    .Y(_0260_),
    .B1(net1063));
 sg13g2_a21oi_1 _5674_ (.A1(net1006),
    .A2(\i_delta_sigma.sample[6] ),
    .Y(_2068_),
    .B1(_2014_));
 sg13g2_xnor2_1 _5675_ (.Y(_2069_),
    .A(_1996_),
    .B(_2068_));
 sg13g2_nor2_1 _5676_ (.A(net873),
    .B(_2069_),
    .Y(_2070_));
 sg13g2_o21ai_1 _5677_ (.B1(_2042_),
    .Y(_2071_),
    .A1(net872),
    .A2(_2070_));
 sg13g2_a21oi_1 _5678_ (.A1(net515),
    .A2(net910),
    .Y(_2072_),
    .B1(net486));
 sg13g2_a21oi_1 _5679_ (.A1(_2071_),
    .A2(_2072_),
    .Y(_0261_),
    .B1(net1063));
 sg13g2_and3_1 _5680_ (.X(_2073_),
    .A(_2015_),
    .B(_2016_),
    .C(_2017_));
 sg13g2_nor3_1 _5681_ (.A(_2018_),
    .B(net873),
    .C(_2073_),
    .Y(_2074_));
 sg13g2_o21ai_1 _5682_ (.B1(_2049_),
    .Y(_2075_),
    .A1(net872),
    .A2(_2074_));
 sg13g2_a21oi_1 _5683_ (.A1(net528),
    .A2(net910),
    .Y(_2076_),
    .B1(net510));
 sg13g2_a21oi_1 _5684_ (.A1(_2075_),
    .A2(_2076_),
    .Y(_0262_),
    .B1(net1063));
 sg13g2_a21oi_1 _5685_ (.A1(net1006),
    .A2(\i_delta_sigma.sample[8] ),
    .Y(_2077_),
    .B1(_2018_));
 sg13g2_xnor2_1 _5686_ (.Y(_2078_),
    .A(_2020_),
    .B(_2077_));
 sg13g2_nor2_1 _5687_ (.A(net873),
    .B(_2078_),
    .Y(_2079_));
 sg13g2_o21ai_1 _5688_ (.B1(_2042_),
    .Y(_2080_),
    .A1(net872),
    .A2(_2079_));
 sg13g2_a21oi_1 _5689_ (.A1(net1014),
    .A2(net911),
    .Y(_2081_),
    .B1(net486));
 sg13g2_a21oi_1 _5690_ (.A1(_2080_),
    .A2(_2081_),
    .Y(_0263_),
    .B1(net1063));
 sg13g2_nor2b_1 _5691_ (.A(_2022_),
    .B_N(_2021_),
    .Y(_2082_));
 sg13g2_nor3_1 _5692_ (.A(_2023_),
    .B(net873),
    .C(_2082_),
    .Y(_2083_));
 sg13g2_o21ai_1 _5693_ (.B1(_2049_),
    .Y(_2084_),
    .A1(_2035_),
    .A2(_2083_));
 sg13g2_a21oi_1 _5694_ (.A1(net1013),
    .A2(net910),
    .Y(_2085_),
    .B1(net510));
 sg13g2_a21oi_1 _5695_ (.A1(_2084_),
    .A2(_2085_),
    .Y(_0264_),
    .B1(net1063));
 sg13g2_a21oi_1 _5696_ (.A1(\i_orchestrator.vga_x[4] ),
    .A2(net1054),
    .Y(_2086_),
    .B1(net5));
 sg13g2_o21ai_1 _5697_ (.B1(_2086_),
    .Y(_2087_),
    .A1(\i_orchestrator.vga_x[4] ),
    .A2(net1054));
 sg13g2_nor3_1 _5698_ (.A(_2386_),
    .B(net1019),
    .C(_1109_),
    .Y(_2088_));
 sg13g2_a21oi_1 _5699_ (.A1(net1019),
    .A2(_1109_),
    .Y(_2089_),
    .B1(_2088_));
 sg13g2_mux2_1 _5700_ (.A0(_2087_),
    .A1(_2089_),
    .S(net868),
    .X(_2090_));
 sg13g2_nor2_1 _5701_ (.A(_2601_),
    .B(_2090_),
    .Y(_0265_));
 sg13g2_and2_1 _5702_ (.A(_0069_),
    .B(_1991_),
    .X(_2091_));
 sg13g2_nand2_1 _5703_ (.Y(_2092_),
    .A(net289),
    .B(_1991_));
 sg13g2_nand2_1 _5704_ (.Y(_2093_),
    .A(\i_resonator.v[7] ),
    .B(_2385_));
 sg13g2_xor2_1 _5705_ (.B(net1017),
    .A(\i_resonator.v[7] ),
    .X(_2094_));
 sg13g2_nand2_1 _5706_ (.Y(_2095_),
    .A(\i_resonator.v[6] ),
    .B(_2380_));
 sg13g2_xnor2_1 _5707_ (.Y(_2096_),
    .A(\i_resonator.v[6] ),
    .B(\i_delta_sigma.sample[10] ));
 sg13g2_nor2b_1 _5708_ (.A(\i_delta_sigma.sample[9] ),
    .B_N(\i_resonator.v[5] ),
    .Y(_2097_));
 sg13g2_xnor2_1 _5709_ (.Y(_2098_),
    .A(\i_resonator.v[5] ),
    .B(\i_delta_sigma.sample[9] ));
 sg13g2_xor2_1 _5710_ (.B(\i_delta_sigma.sample[8] ),
    .A(\i_resonator.v[4] ),
    .X(_2099_));
 sg13g2_xor2_1 _5711_ (.B(\i_delta_sigma.sample[7] ),
    .A(\i_resonator.v[3] ),
    .X(_2100_));
 sg13g2_xor2_1 _5712_ (.B(\i_delta_sigma.sample[6] ),
    .A(\i_resonator.v[2] ),
    .X(_2101_));
 sg13g2_nor2b_1 _5713_ (.A(\i_delta_sigma.sample[5] ),
    .B_N(\i_resonator.v[1] ),
    .Y(_2102_));
 sg13g2_nand2b_1 _5714_ (.Y(_2103_),
    .B(\i_delta_sigma.sample[4] ),
    .A_N(\i_resonator.v[0] ));
 sg13g2_xnor2_1 _5715_ (.Y(_2104_),
    .A(\i_resonator.v[1] ),
    .B(\i_delta_sigma.sample[5] ));
 sg13g2_a21oi_1 _5716_ (.A1(_2103_),
    .A2(_2104_),
    .Y(_2105_),
    .B1(_2102_));
 sg13g2_nor2_1 _5717_ (.A(_2101_),
    .B(_2105_),
    .Y(_2106_));
 sg13g2_a21oi_1 _5718_ (.A1(\i_resonator.v[2] ),
    .A2(_2383_),
    .Y(_2107_),
    .B1(_2106_));
 sg13g2_nor2_1 _5719_ (.A(_2100_),
    .B(_2107_),
    .Y(_2108_));
 sg13g2_a21oi_1 _5720_ (.A1(\i_resonator.v[3] ),
    .A2(_2382_),
    .Y(_2109_),
    .B1(_2108_));
 sg13g2_nor2_1 _5721_ (.A(_2099_),
    .B(_2109_),
    .Y(_2110_));
 sg13g2_a21oi_2 _5722_ (.B1(_2110_),
    .Y(_2111_),
    .A2(_2381_),
    .A1(\i_resonator.v[4] ));
 sg13g2_nor2b_1 _5723_ (.A(_2111_),
    .B_N(_2098_),
    .Y(_2112_));
 sg13g2_o21ai_1 _5724_ (.B1(_2096_),
    .Y(_2113_),
    .A1(_2097_),
    .A2(_2112_));
 sg13g2_and2_1 _5725_ (.A(_2095_),
    .B(_2113_),
    .X(_2114_));
 sg13g2_o21ai_1 _5726_ (.B1(_2093_),
    .Y(_2115_),
    .A1(_2094_),
    .A2(_2114_));
 sg13g2_xnor2_1 _5727_ (.Y(_2116_),
    .A(\i_resonator.v[8] ),
    .B(net1017));
 sg13g2_and2_1 _5728_ (.A(_2115_),
    .B(_2116_),
    .X(_2117_));
 sg13g2_xor2_1 _5729_ (.B(net1017),
    .A(\i_resonator.v[9] ),
    .X(_2118_));
 sg13g2_inv_1 _5730_ (.Y(_2119_),
    .A(_2118_));
 sg13g2_nand2_1 _5731_ (.Y(_2120_),
    .A(_2117_),
    .B(_2119_));
 sg13g2_nand2_1 _5732_ (.Y(_2121_),
    .A(net1012),
    .B(_2385_));
 sg13g2_xor2_1 _5733_ (.B(net1017),
    .A(\i_resonator.v[10] ),
    .X(_2122_));
 sg13g2_xor2_1 _5734_ (.B(net1017),
    .A(\i_resonator.v[11] ),
    .X(_2123_));
 sg13g2_nor3_2 _5735_ (.A(_2120_),
    .B(_2122_),
    .C(_2123_),
    .Y(_2124_));
 sg13g2_nor3_1 _5736_ (.A(net1009),
    .B(\i_resonator.v[14] ),
    .C(\i_resonator.v[13] ),
    .Y(_2125_));
 sg13g2_nand3_1 _5737_ (.B(\i_resonator.v[14] ),
    .C(\i_resonator.v[13] ),
    .A(net1009),
    .Y(_2126_));
 sg13g2_nand2b_1 _5738_ (.Y(_2127_),
    .B(_2126_),
    .A_N(_2125_));
 sg13g2_xnor2_1 _5739_ (.Y(_2128_),
    .A(\i_resonator.v[12] ),
    .B(net1016));
 sg13g2_nand2b_1 _5740_ (.Y(_2129_),
    .B(net1015),
    .A_N(net1011));
 sg13g2_nor2b_1 _5741_ (.A(net1015),
    .B_N(net1011),
    .Y(_2130_));
 sg13g2_xnor2_1 _5742_ (.Y(_2131_),
    .A(net1011),
    .B(net1016));
 sg13g2_nand4_1 _5743_ (.B(_2127_),
    .C(_2128_),
    .A(_2124_),
    .Y(_2132_),
    .D(_2131_));
 sg13g2_a21oi_1 _5744_ (.A1(_2378_),
    .A2(_2379_),
    .Y(_2133_),
    .B1(net1017));
 sg13g2_a21oi_1 _5745_ (.A1(\i_resonator.v[11] ),
    .A2(_2385_),
    .Y(_2134_),
    .B1(_2133_));
 sg13g2_nand2_2 _5746_ (.Y(_2135_),
    .A(_2121_),
    .B(_2134_));
 sg13g2_a21oi_1 _5747_ (.A1(_2377_),
    .A2(_2125_),
    .Y(_2136_),
    .B1(net1016));
 sg13g2_nor2_1 _5748_ (.A(_2135_),
    .B(_2136_),
    .Y(_2137_));
 sg13g2_xor2_1 _5749_ (.B(net1015),
    .A(\i_resonator.v[14] ),
    .X(_2138_));
 sg13g2_o21ai_1 _5750_ (.B1(_2128_),
    .Y(_2139_),
    .A1(_2124_),
    .A2(_2135_));
 sg13g2_o21ai_1 _5751_ (.B1(_2139_),
    .Y(_2140_),
    .A1(_2377_),
    .A2(net1015));
 sg13g2_o21ai_1 _5752_ (.B1(_2129_),
    .Y(_2141_),
    .A1(_2130_),
    .A2(_2140_));
 sg13g2_nor2_1 _5753_ (.A(_2138_),
    .B(_2141_),
    .Y(_2142_));
 sg13g2_a21oi_1 _5754_ (.A1(\i_resonator.v[14] ),
    .A2(_2385_),
    .Y(_2143_),
    .B1(_2142_));
 sg13g2_a21oi_1 _5755_ (.A1(_2132_),
    .A2(_2137_),
    .Y(_2144_),
    .B1(_2025_));
 sg13g2_a21oi_2 _5756_ (.B1(_2144_),
    .Y(_2145_),
    .A2(_2143_),
    .A1(_2025_));
 sg13g2_xnor2_1 _5757_ (.Y(_2146_),
    .A(_2025_),
    .B(_2143_));
 sg13g2_nand2_2 _5758_ (.Y(_2147_),
    .A(_2145_),
    .B(_2146_));
 sg13g2_inv_1 _5759_ (.Y(_2148_),
    .A(_2147_));
 sg13g2_nor2_2 _5760_ (.A(net1048),
    .B(_2148_),
    .Y(_2149_));
 sg13g2_nor2_2 _5761_ (.A(_2145_),
    .B(_2146_),
    .Y(_2150_));
 sg13g2_xnor2_1 _5762_ (.Y(_2151_),
    .A(net331),
    .B(\i_delta_sigma.sample[4] ));
 sg13g2_o21ai_1 _5763_ (.B1(_2149_),
    .Y(_2152_),
    .A1(_2150_),
    .A2(_2151_));
 sg13g2_and3_1 _5764_ (.X(_2153_),
    .A(net1013),
    .B(net1014),
    .C(net1015));
 sg13g2_nor3_1 _5765_ (.A(net1013),
    .B(net1014),
    .C(net1015),
    .Y(_2154_));
 sg13g2_o21ai_1 _5766_ (.B1(_2127_),
    .Y(_2155_),
    .A1(_2153_),
    .A2(_2154_));
 sg13g2_mux2_1 _5767_ (.A0(_0047_),
    .A1(_0046_),
    .S(_2155_),
    .X(_2156_));
 sg13g2_inv_1 _5768_ (.Y(_2157_),
    .A(_2156_));
 sg13g2_nand2_2 _5769_ (.Y(_2158_),
    .A(_0045_),
    .B(_2157_));
 sg13g2_o21ai_1 _5770_ (.B1(net1046),
    .Y(_2159_),
    .A1(_0045_),
    .A2(_2157_));
 sg13g2_nand2b_1 _5771_ (.Y(_2160_),
    .B(_2158_),
    .A_N(_2159_));
 sg13g2_a21oi_1 _5772_ (.A1(_2152_),
    .A2(_2160_),
    .Y(_2161_),
    .B1(net930));
 sg13g2_o21ai_1 _5773_ (.B1(net934),
    .Y(_2162_),
    .A1(net331),
    .A2(net929));
 sg13g2_nor2_1 _5774_ (.A(_2161_),
    .B(_2162_),
    .Y(_0266_));
 sg13g2_xnor2_1 _5775_ (.Y(_2163_),
    .A(_2103_),
    .B(_2104_));
 sg13g2_o21ai_1 _5776_ (.B1(_2149_),
    .Y(_2164_),
    .A1(_2150_),
    .A2(_2163_));
 sg13g2_nor2_1 _5777_ (.A(net1012),
    .B(_2155_),
    .Y(_2165_));
 sg13g2_a21oi_2 _5778_ (.B1(_2165_),
    .Y(_2166_),
    .A2(_2155_),
    .A1(_2377_));
 sg13g2_nor2b_1 _5779_ (.A(_2166_),
    .B_N(\i_resonator.v[1] ),
    .Y(_2167_));
 sg13g2_xnor2_1 _5780_ (.Y(_2168_),
    .A(\i_resonator.v[1] ),
    .B(_2166_));
 sg13g2_xnor2_1 _5781_ (.Y(_2169_),
    .A(_2158_),
    .B(_2168_));
 sg13g2_a21oi_1 _5782_ (.A1(net1046),
    .A2(_2169_),
    .Y(_2170_),
    .B1(net930));
 sg13g2_a22oi_1 _5783_ (.Y(_2171_),
    .B1(_2164_),
    .B2(_2170_),
    .A2(net930),
    .A1(net403));
 sg13g2_nor2_1 _5784_ (.A(net945),
    .B(net404),
    .Y(_0267_));
 sg13g2_xnor2_1 _5785_ (.Y(_2172_),
    .A(_2101_),
    .B(_2105_));
 sg13g2_o21ai_1 _5786_ (.B1(_2149_),
    .Y(_2173_),
    .A1(_2150_),
    .A2(_2172_));
 sg13g2_mux2_1 _5787_ (.A0(_0046_),
    .A1(_0048_),
    .S(_2155_),
    .X(_2174_));
 sg13g2_xor2_1 _5788_ (.B(_2174_),
    .A(\i_resonator.v[2] ),
    .X(_2175_));
 sg13g2_a21oi_1 _5789_ (.A1(_2158_),
    .A2(_2168_),
    .Y(_2176_),
    .B1(_2167_));
 sg13g2_nor2b_1 _5790_ (.A(_2176_),
    .B_N(_2175_),
    .Y(_2177_));
 sg13g2_xor2_1 _5791_ (.B(_2176_),
    .A(_2175_),
    .X(_2178_));
 sg13g2_a21oi_1 _5792_ (.A1(net1046),
    .A2(_2178_),
    .Y(_2179_),
    .B1(net930));
 sg13g2_a22oi_1 _5793_ (.Y(_2180_),
    .B1(_2173_),
    .B2(_2179_),
    .A2(net930),
    .A1(net422));
 sg13g2_nor2_1 _5794_ (.A(net945),
    .B(_2180_),
    .Y(_0268_));
 sg13g2_xnor2_1 _5795_ (.Y(_2181_),
    .A(_2100_),
    .B(_2107_));
 sg13g2_o21ai_1 _5796_ (.B1(_2149_),
    .Y(_2182_),
    .A1(_2150_),
    .A2(_2181_));
 sg13g2_nor2_1 _5797_ (.A(\i_resonator.v[12] ),
    .B(_2155_),
    .Y(_2183_));
 sg13g2_a21oi_2 _5798_ (.B1(_2183_),
    .Y(_2184_),
    .A2(_2155_),
    .A1(_2376_));
 sg13g2_nor2b_1 _5799_ (.A(_2184_),
    .B_N(\i_resonator.v[3] ),
    .Y(_2185_));
 sg13g2_xnor2_1 _5800_ (.Y(_2186_),
    .A(\i_resonator.v[3] ),
    .B(_2184_));
 sg13g2_a21o_1 _5801_ (.A2(_2174_),
    .A1(\i_resonator.v[2] ),
    .B1(_2177_),
    .X(_2187_));
 sg13g2_xnor2_1 _5802_ (.Y(_2188_),
    .A(_2186_),
    .B(_2187_));
 sg13g2_a21oi_1 _5803_ (.A1(net1046),
    .A2(_2188_),
    .Y(_2189_),
    .B1(net930));
 sg13g2_a22oi_1 _5804_ (.Y(_2190_),
    .B1(_2182_),
    .B2(_2189_),
    .A2(net930),
    .A1(net421));
 sg13g2_nor2_1 _5805_ (.A(net945),
    .B(_2190_),
    .Y(_0269_));
 sg13g2_xnor2_1 _5806_ (.Y(_2191_),
    .A(_2099_),
    .B(_2109_));
 sg13g2_o21ai_1 _5807_ (.B1(_2149_),
    .Y(_2192_),
    .A1(_2150_),
    .A2(_2191_));
 sg13g2_mux2_1 _5808_ (.A0(_0048_),
    .A1(_0049_),
    .S(_2155_),
    .X(_2193_));
 sg13g2_xor2_1 _5809_ (.B(_2193_),
    .A(\i_resonator.v[4] ),
    .X(_2194_));
 sg13g2_a21oi_1 _5810_ (.A1(_2186_),
    .A2(_2187_),
    .Y(_2195_),
    .B1(_2185_));
 sg13g2_nor2b_1 _5811_ (.A(_2195_),
    .B_N(_2194_),
    .Y(_2196_));
 sg13g2_xor2_1 _5812_ (.B(_2195_),
    .A(_2194_),
    .X(_2197_));
 sg13g2_a21oi_1 _5813_ (.A1(net1046),
    .A2(_2197_),
    .Y(_2198_),
    .B1(net931));
 sg13g2_a22oi_1 _5814_ (.Y(_2199_),
    .B1(_2192_),
    .B2(_2198_),
    .A2(net930),
    .A1(net398));
 sg13g2_nor2_1 _5815_ (.A(net945),
    .B(_2199_),
    .Y(_0270_));
 sg13g2_xnor2_1 _5816_ (.Y(_2200_),
    .A(_2098_),
    .B(_2111_));
 sg13g2_nor2_1 _5817_ (.A(net1046),
    .B(_2150_),
    .Y(_2201_));
 sg13g2_nand2b_1 _5818_ (.Y(_2202_),
    .B(net1009),
    .A_N(\i_resonator.v[5] ));
 sg13g2_nand2_1 _5819_ (.Y(_2203_),
    .A(net994),
    .B(\i_resonator.v[5] ));
 sg13g2_inv_1 _5820_ (.Y(_2204_),
    .A(_2203_));
 sg13g2_a21o_2 _5821_ (.A2(_2193_),
    .A1(\i_resonator.v[4] ),
    .B1(_2196_),
    .X(_2205_));
 sg13g2_nand3_1 _5822_ (.B(_2203_),
    .C(_2205_),
    .A(_2202_),
    .Y(_2206_));
 sg13g2_a21oi_1 _5823_ (.A1(_2202_),
    .A2(_2203_),
    .Y(_2207_),
    .B1(_2205_));
 sg13g2_nand2_1 _5824_ (.Y(_2208_),
    .A(net1048),
    .B(_2206_));
 sg13g2_o21ai_1 _5825_ (.B1(net929),
    .Y(_2209_),
    .A1(_2207_),
    .A2(_2208_));
 sg13g2_a221oi_1 _5826_ (.B2(net813),
    .C1(_2209_),
    .B1(_2200_),
    .A1(_2433_),
    .Y(_2210_),
    .A2(_2148_));
 sg13g2_o21ai_1 _5827_ (.B1(net934),
    .Y(_2211_),
    .A1(net430),
    .A2(net929));
 sg13g2_nor2_1 _5828_ (.A(_2210_),
    .B(_2211_),
    .Y(_0271_));
 sg13g2_or3_1 _5829_ (.A(_2096_),
    .B(_2097_),
    .C(_2112_),
    .X(_2212_));
 sg13g2_nand2_1 _5830_ (.Y(_2213_),
    .A(_2113_),
    .B(_2212_));
 sg13g2_o21ai_1 _5831_ (.B1(_2149_),
    .Y(_2214_),
    .A1(_2150_),
    .A2(_2213_));
 sg13g2_nand2_1 _5832_ (.Y(_2215_),
    .A(net994),
    .B(\i_resonator.v[6] ));
 sg13g2_xor2_1 _5833_ (.B(\i_resonator.v[6] ),
    .A(net1010),
    .X(_2216_));
 sg13g2_a21oi_1 _5834_ (.A1(_2202_),
    .A2(_2205_),
    .Y(_2217_),
    .B1(_2204_));
 sg13g2_xnor2_1 _5835_ (.Y(_2218_),
    .A(_2216_),
    .B(_2217_));
 sg13g2_a21oi_1 _5836_ (.A1(net1047),
    .A2(_2218_),
    .Y(_2219_),
    .B1(net933));
 sg13g2_a22oi_1 _5837_ (.Y(_2220_),
    .B1(_2214_),
    .B2(_2219_),
    .A2(net932),
    .A1(net405));
 sg13g2_nor2_1 _5838_ (.A(net945),
    .B(_2220_),
    .Y(_0272_));
 sg13g2_xnor2_1 _5839_ (.Y(_2221_),
    .A(_2094_),
    .B(_2114_));
 sg13g2_nand2_1 _5840_ (.Y(_2222_),
    .A(_2147_),
    .B(_2221_));
 sg13g2_nand2b_1 _5841_ (.Y(_2223_),
    .B(net1010),
    .A_N(\i_resonator.v[7] ));
 sg13g2_nand2_1 _5842_ (.Y(_2224_),
    .A(_2375_),
    .B(\i_resonator.v[7] ));
 sg13g2_o21ai_1 _5843_ (.B1(_2215_),
    .Y(_2225_),
    .A1(_2216_),
    .A2(_2217_));
 sg13g2_a21oi_1 _5844_ (.A1(_2223_),
    .A2(_2224_),
    .Y(_2226_),
    .B1(_2225_));
 sg13g2_nand3_1 _5845_ (.B(_2224_),
    .C(_2225_),
    .A(_2223_),
    .Y(_2227_));
 sg13g2_nor2_1 _5846_ (.A(_2433_),
    .B(_2226_),
    .Y(_2228_));
 sg13g2_a221oi_1 _5847_ (.B2(_2228_),
    .C1(net933),
    .B1(_2227_),
    .A1(net813),
    .Y(_2229_),
    .A2(_2222_));
 sg13g2_o21ai_1 _5848_ (.B1(net934),
    .Y(_2230_),
    .A1(net457),
    .A2(_2092_));
 sg13g2_nor2_1 _5849_ (.A(_2229_),
    .B(_2230_),
    .Y(_0273_));
 sg13g2_nor2_1 _5850_ (.A(_2115_),
    .B(_2116_),
    .Y(_2231_));
 sg13g2_o21ai_1 _5851_ (.B1(_2147_),
    .Y(_2232_),
    .A1(_2117_),
    .A2(_2231_));
 sg13g2_xor2_1 _5852_ (.B(\i_resonator.v[8] ),
    .A(net1010),
    .X(_2233_));
 sg13g2_nand2_1 _5853_ (.Y(_2234_),
    .A(_2223_),
    .B(_2225_));
 sg13g2_and2_1 _5854_ (.A(_2224_),
    .B(_2234_),
    .X(_2235_));
 sg13g2_nor2_1 _5855_ (.A(_2233_),
    .B(_2235_),
    .Y(_2236_));
 sg13g2_or2_1 _5856_ (.X(_2237_),
    .B(_2235_),
    .A(_2233_));
 sg13g2_a21oi_1 _5857_ (.A1(_2233_),
    .A2(_2235_),
    .Y(_2238_),
    .B1(_2433_));
 sg13g2_a221oi_1 _5858_ (.B2(_2238_),
    .C1(net933),
    .B1(_2237_),
    .A1(net813),
    .Y(_2239_),
    .A2(_2232_));
 sg13g2_o21ai_1 _5859_ (.B1(_2030_),
    .Y(_2240_),
    .A1(net517),
    .A2(net929));
 sg13g2_nor2_1 _5860_ (.A(_2239_),
    .B(_2240_),
    .Y(_0274_));
 sg13g2_a21oi_1 _5861_ (.A1(\i_resonator.v[8] ),
    .A2(_2385_),
    .Y(_2241_),
    .B1(_2117_));
 sg13g2_xnor2_1 _5862_ (.Y(_2242_),
    .A(_2118_),
    .B(_2241_));
 sg13g2_nand2_1 _5863_ (.Y(_2243_),
    .A(_2147_),
    .B(_2242_));
 sg13g2_xor2_1 _5864_ (.B(\i_resonator.v[9] ),
    .A(net1010),
    .X(_2244_));
 sg13g2_a21oi_1 _5865_ (.A1(_2375_),
    .A2(\i_resonator.v[8] ),
    .Y(_2245_),
    .B1(_2236_));
 sg13g2_or2_1 _5866_ (.X(_2246_),
    .B(_2245_),
    .A(_2244_));
 sg13g2_a21oi_1 _5867_ (.A1(_2244_),
    .A2(_2245_),
    .Y(_2247_),
    .B1(_2433_));
 sg13g2_a221oi_1 _5868_ (.B2(_2247_),
    .C1(net932),
    .B1(_2246_),
    .A1(_2201_),
    .Y(_2248_),
    .A2(_2243_));
 sg13g2_o21ai_1 _5869_ (.B1(_2030_),
    .Y(_2249_),
    .A1(net466),
    .A2(net929));
 sg13g2_nor2_1 _5870_ (.A(_2248_),
    .B(_2249_),
    .Y(_0275_));
 sg13g2_a21oi_1 _5871_ (.A1(_2117_),
    .A2(_2119_),
    .Y(_2250_),
    .B1(_2133_));
 sg13g2_xnor2_1 _5872_ (.Y(_2251_),
    .A(_2122_),
    .B(_2250_));
 sg13g2_nand2_1 _5873_ (.Y(_2252_),
    .A(_2147_),
    .B(_2251_));
 sg13g2_nand2_1 _5874_ (.Y(_2253_),
    .A(_2375_),
    .B(net1012));
 sg13g2_xnor2_1 _5875_ (.Y(_2254_),
    .A(net1010),
    .B(net1012));
 sg13g2_inv_1 _5876_ (.Y(_2255_),
    .A(_2254_));
 sg13g2_o21ai_1 _5877_ (.B1(net994),
    .Y(_2256_),
    .A1(\i_resonator.v[9] ),
    .A2(\i_resonator.v[8] ));
 sg13g2_o21ai_1 _5878_ (.B1(_2256_),
    .Y(_2257_),
    .A1(_2237_),
    .A2(_2244_));
 sg13g2_nand2_1 _5879_ (.Y(_2258_),
    .A(_2254_),
    .B(_2257_));
 sg13g2_o21ai_1 _5880_ (.B1(net1047),
    .Y(_2259_),
    .A1(_2254_),
    .A2(_2257_));
 sg13g2_inv_1 _5881_ (.Y(_2260_),
    .A(_2259_));
 sg13g2_a221oi_1 _5882_ (.B2(_2260_),
    .C1(net932),
    .B1(_2258_),
    .A1(net813),
    .Y(_2261_),
    .A2(_2252_));
 sg13g2_o21ai_1 _5883_ (.B1(net934),
    .Y(_2262_),
    .A1(net1012),
    .A2(net929));
 sg13g2_nor2_1 _5884_ (.A(_2261_),
    .B(_2262_),
    .Y(_0276_));
 sg13g2_o21ai_1 _5885_ (.B1(_2121_),
    .Y(_2263_),
    .A1(_2122_),
    .A2(_2250_));
 sg13g2_xor2_1 _5886_ (.B(_2263_),
    .A(_2123_),
    .X(_2264_));
 sg13g2_nand2_1 _5887_ (.Y(_2265_),
    .A(_2147_),
    .B(_2264_));
 sg13g2_xor2_1 _5888_ (.B(\i_resonator.v[11] ),
    .A(net1010),
    .X(_2266_));
 sg13g2_nand3_1 _5889_ (.B(_2258_),
    .C(_2266_),
    .A(_2253_),
    .Y(_2267_));
 sg13g2_a21oi_1 _5890_ (.A1(_2253_),
    .A2(_2258_),
    .Y(_2268_),
    .B1(_2266_));
 sg13g2_nor2_1 _5891_ (.A(_2433_),
    .B(_2268_),
    .Y(_2269_));
 sg13g2_a221oi_1 _5892_ (.B2(_2269_),
    .C1(net932),
    .B1(_2267_),
    .A1(net813),
    .Y(_2270_),
    .A2(_2265_));
 sg13g2_o21ai_1 _5893_ (.B1(net934),
    .Y(_2271_),
    .A1(net537),
    .A2(net929));
 sg13g2_nor2_1 _5894_ (.A(_2270_),
    .B(_2271_),
    .Y(_0277_));
 sg13g2_or3_1 _5895_ (.A(_2124_),
    .B(_2128_),
    .C(_2135_),
    .X(_2272_));
 sg13g2_and2_1 _5896_ (.A(_2139_),
    .B(_2272_),
    .X(_2273_));
 sg13g2_o21ai_1 _5897_ (.B1(net813),
    .Y(_2274_),
    .A1(_2148_),
    .A2(_2273_));
 sg13g2_nand2_1 _5898_ (.Y(_2275_),
    .A(net994),
    .B(\i_resonator.v[12] ));
 sg13g2_xnor2_1 _5899_ (.Y(_2276_),
    .A(net1009),
    .B(\i_resonator.v[12] ));
 sg13g2_or4_1 _5900_ (.A(_2237_),
    .B(_2244_),
    .C(_2255_),
    .D(_2266_),
    .X(_2277_));
 sg13g2_o21ai_1 _5901_ (.B1(net994),
    .Y(_2278_),
    .A1(\i_resonator.v[11] ),
    .A2(net1012));
 sg13g2_nand3_1 _5902_ (.B(_2277_),
    .C(_2278_),
    .A(_2256_),
    .Y(_2279_));
 sg13g2_nand2_2 _5903_ (.Y(_2280_),
    .A(_2276_),
    .B(_2279_));
 sg13g2_o21ai_1 _5904_ (.B1(net1046),
    .Y(_2281_),
    .A1(_2276_),
    .A2(_2279_));
 sg13g2_inv_1 _5905_ (.Y(_2282_),
    .A(_2281_));
 sg13g2_a21oi_1 _5906_ (.A1(_2280_),
    .A2(_2282_),
    .Y(_2283_),
    .B1(net932));
 sg13g2_a221oi_1 _5907_ (.B2(_2283_),
    .C1(net945),
    .B1(_2274_),
    .A1(_2377_),
    .Y(_0278_),
    .A2(net932));
 sg13g2_xnor2_1 _5908_ (.Y(_2284_),
    .A(net1009),
    .B(net1011));
 sg13g2_inv_1 _5909_ (.Y(_2285_),
    .A(_2284_));
 sg13g2_a21oi_1 _5910_ (.A1(_2275_),
    .A2(_2280_),
    .Y(_2286_),
    .B1(_2285_));
 sg13g2_nand3_1 _5911_ (.B(_2280_),
    .C(_2285_),
    .A(_2275_),
    .Y(_2287_));
 sg13g2_nor2_1 _5912_ (.A(_2433_),
    .B(_2286_),
    .Y(_2288_));
 sg13g2_xnor2_1 _5913_ (.Y(_2289_),
    .A(_2131_),
    .B(_2140_));
 sg13g2_nand2_1 _5914_ (.Y(_2290_),
    .A(_2147_),
    .B(_2289_));
 sg13g2_a221oi_1 _5915_ (.B2(net813),
    .C1(net932),
    .B1(_2290_),
    .A1(_2287_),
    .Y(_2291_),
    .A2(_2288_));
 sg13g2_o21ai_1 _5916_ (.B1(net934),
    .Y(_2292_),
    .A1(net1011),
    .A2(net929));
 sg13g2_nor2_1 _5917_ (.A(_2291_),
    .B(_2292_),
    .Y(_0279_));
 sg13g2_xnor2_1 _5918_ (.Y(_2293_),
    .A(net1009),
    .B(\i_resonator.v[14] ));
 sg13g2_o21ai_1 _5919_ (.B1(net994),
    .Y(_2294_),
    .A1(net1011),
    .A2(\i_resonator.v[12] ));
 sg13g2_o21ai_1 _5920_ (.B1(_2294_),
    .Y(_2295_),
    .A1(_2280_),
    .A2(_2285_));
 sg13g2_a21oi_1 _5921_ (.A1(_2293_),
    .A2(_2295_),
    .Y(_2296_),
    .B1(_2433_));
 sg13g2_o21ai_1 _5922_ (.B1(_2296_),
    .Y(_2297_),
    .A1(_2293_),
    .A2(_2295_));
 sg13g2_xnor2_1 _5923_ (.Y(_2298_),
    .A(_2138_),
    .B(_2141_));
 sg13g2_nand2_1 _5924_ (.Y(_2299_),
    .A(_2147_),
    .B(_2298_));
 sg13g2_a21oi_1 _5925_ (.A1(net813),
    .A2(_2299_),
    .Y(_2300_),
    .B1(net932));
 sg13g2_a221oi_1 _5926_ (.B2(_2300_),
    .C1(net945),
    .B1(_2297_),
    .A1(_2376_),
    .Y(_0280_),
    .A2(net931));
 sg13g2_o21ai_1 _5927_ (.B1(_2296_),
    .Y(_2301_),
    .A1(net1009),
    .A2(_2376_));
 sg13g2_nor2_1 _5928_ (.A(net1046),
    .B(_2145_),
    .Y(_2302_));
 sg13g2_nor2_1 _5929_ (.A(net931),
    .B(_2302_),
    .Y(_2303_));
 sg13g2_a221oi_1 _5930_ (.B2(_2303_),
    .C1(net945),
    .B1(_2301_),
    .A1(net994),
    .Y(_0281_),
    .A2(net931));
 sg13g2_nor3_1 _5931_ (.A(_1991_),
    .B(_2029_),
    .C(net290),
    .Y(_0282_));
 sg13g2_xnor2_1 _5932_ (.Y(_2304_),
    .A(\i_resonator.counter[1] ),
    .B(\i_resonator.counter[0] ));
 sg13g2_nor2_1 _5933_ (.A(net1047),
    .B(_1991_),
    .Y(_2305_));
 sg13g2_a22oi_1 _5934_ (.Y(_2306_),
    .B1(_2304_),
    .B2(_2305_),
    .A2(net1047),
    .A1(net277));
 sg13g2_o21ai_1 _5935_ (.B1(net934),
    .Y(_2307_),
    .A1(_1992_),
    .A2(_2037_));
 sg13g2_nor2_1 _5936_ (.A(net278),
    .B(_2307_),
    .Y(_0283_));
 sg13g2_o21ai_1 _5937_ (.B1(\i_resonator.counter[2] ),
    .Y(_2308_),
    .A1(\i_resonator.counter[1] ),
    .A2(\i_resonator.counter[0] ));
 sg13g2_nand2b_1 _5938_ (.Y(_2309_),
    .B(_2308_),
    .A_N(_2038_));
 sg13g2_a22oi_1 _5939_ (.Y(_2310_),
    .B1(_2305_),
    .B2(_2309_),
    .A2(net1047),
    .A1(net258));
 sg13g2_nor2_1 _5940_ (.A(_2307_),
    .B(net259),
    .Y(_0284_));
 sg13g2_nor2b_1 _5941_ (.A(_2038_),
    .B_N(net388),
    .Y(_2311_));
 sg13g2_nand2b_1 _5942_ (.Y(_2312_),
    .B(net1047),
    .A_N(net260));
 sg13g2_o21ai_1 _5943_ (.B1(_2312_),
    .Y(_2313_),
    .A1(net1047),
    .A2(_2311_));
 sg13g2_nor2_1 _5944_ (.A(_2307_),
    .B(_2313_),
    .Y(_0285_));
 sg13g2_nor2_1 _5945_ (.A(_0051_),
    .B(net924),
    .Y(_2314_));
 sg13g2_a221oi_1 _5946_ (.B2(_2314_),
    .C1(net1000),
    .B1(_1560_),
    .A1(net1003),
    .Y(_2315_),
    .A2(net952));
 sg13g2_o21ai_1 _5947_ (.B1(_1572_),
    .Y(_2316_),
    .A1(_0051_),
    .A2(_1566_));
 sg13g2_a22oi_1 _5948_ (.Y(_2317_),
    .B1(_2316_),
    .B2(net923),
    .A2(_1602_),
    .A1(net950));
 sg13g2_a21oi_1 _5949_ (.A1(net1002),
    .A2(_2317_),
    .Y(_2318_),
    .B1(_2315_));
 sg13g2_a21oi_1 _5950_ (.A1(net952),
    .A2(_1515_),
    .Y(_2319_),
    .B1(_1579_));
 sg13g2_a21oi_1 _5951_ (.A1(net950),
    .A2(_1532_),
    .Y(_2320_),
    .B1(_1576_));
 sg13g2_o21ai_1 _5952_ (.B1(net924),
    .Y(_2321_),
    .A1(_2319_),
    .A2(_2320_));
 sg13g2_a21oi_1 _5953_ (.A1(_1607_),
    .A2(_2321_),
    .Y(_2322_),
    .B1(_1524_));
 sg13g2_o21ai_1 _5954_ (.B1(_2322_),
    .Y(_2323_),
    .A1(_1491_),
    .A2(_2318_));
 sg13g2_nor2_1 _5955_ (.A(_2373_),
    .B(_2414_),
    .Y(_2324_));
 sg13g2_nor2_1 _5956_ (.A(_0052_),
    .B(_1549_),
    .Y(_2325_));
 sg13g2_a21oi_1 _5957_ (.A1(_0052_),
    .A2(net924),
    .Y(_2326_),
    .B1(_1601_));
 sg13g2_o21ai_1 _5958_ (.B1(_2326_),
    .Y(_2327_),
    .A1(_2324_),
    .A2(_2325_));
 sg13g2_nand3_1 _5959_ (.B(_2323_),
    .C(_2327_),
    .A(net1033),
    .Y(_2328_));
 sg13g2_o21ai_1 _5960_ (.B1(_2328_),
    .Y(_2329_),
    .A1(net1004),
    .A2(net1033));
 sg13g2_nor2_1 _5961_ (.A(net1070),
    .B(_2329_),
    .Y(_0286_));
 sg13g2_a21oi_1 _5962_ (.A1(_2386_),
    .A2(_1109_),
    .Y(_0287_),
    .B1(_1107_));
 sg13g2_xnor2_1 _5963_ (.Y(_2330_),
    .A(net554),
    .B(net1055));
 sg13g2_nor2_1 _5964_ (.A(net5),
    .B(_2330_),
    .Y(_2331_));
 sg13g2_nand3_1 _5965_ (.B(net1019),
    .C(net329),
    .A(\capsule_color[3] ),
    .Y(_2332_));
 sg13g2_and2_1 _5966_ (.A(net413),
    .B(_1108_),
    .X(_2333_));
 sg13g2_a22oi_1 _5967_ (.Y(_2334_),
    .B1(_2332_),
    .B2(_2333_),
    .A2(_1109_),
    .A1(net329));
 sg13g2_o21ai_1 _5968_ (.B1(net920),
    .Y(_2335_),
    .A1(net868),
    .A2(_2331_));
 sg13g2_a21oi_1 _5969_ (.A1(net868),
    .A2(_2334_),
    .Y(_0288_),
    .B1(_2335_));
 sg13g2_nand2_1 _5970_ (.Y(_2336_),
    .A(net997),
    .B(net925));
 sg13g2_a22oi_1 _5971_ (.Y(_2337_),
    .B1(_2336_),
    .B2(_1491_),
    .A2(net949),
    .A1(net923));
 sg13g2_nor2b_1 _5972_ (.A(net1023),
    .B_N(_2337_),
    .Y(_2338_));
 sg13g2_nand3_1 _5973_ (.B(net953),
    .C(net921),
    .A(net1033),
    .Y(_2339_));
 sg13g2_o21ai_1 _5974_ (.B1(net1002),
    .Y(_2340_),
    .A1(_2338_),
    .A2(_2339_));
 sg13g2_nand2_1 _5975_ (.Y(_2341_),
    .A(net1023),
    .B(_2337_));
 sg13g2_nand4_1 _5976_ (.B(net951),
    .C(net921),
    .A(net1033),
    .Y(_2342_),
    .D(_2341_));
 sg13g2_a21oi_1 _5977_ (.A1(_2340_),
    .A2(_2342_),
    .Y(_0289_),
    .B1(net1070));
 sg13g2_a21oi_1 _5978_ (.A1(_0070_),
    .A2(net951),
    .Y(_2343_),
    .B1(_1505_));
 sg13g2_nand3_1 _5979_ (.B(_1612_),
    .C(_2343_),
    .A(net921),
    .Y(_2344_));
 sg13g2_and2_1 _5980_ (.A(net1033),
    .B(_2344_),
    .X(_2345_));
 sg13g2_o21ai_1 _5981_ (.B1(_1551_),
    .Y(_2346_),
    .A1(net1050),
    .A2(_1527_));
 sg13g2_o21ai_1 _5982_ (.B1(_1577_),
    .Y(_2347_),
    .A1(net950),
    .A2(_1588_));
 sg13g2_nand3_1 _5983_ (.B(net1005),
    .C(net952),
    .A(net995),
    .Y(_2348_));
 sg13g2_o21ai_1 _5984_ (.B1(_2348_),
    .Y(_2349_),
    .A1(_1572_),
    .A2(_1593_));
 sg13g2_a221oi_1 _5985_ (.B2(_2374_),
    .C1(net922),
    .B1(_2349_),
    .A1(_1781_),
    .Y(_2350_),
    .A2(_2347_));
 sg13g2_o21ai_1 _5986_ (.B1(net922),
    .Y(_2351_),
    .A1(net1049),
    .A2(_1550_));
 sg13g2_a21oi_1 _5987_ (.A1(net1050),
    .A2(_1550_),
    .Y(_2352_),
    .B1(_2351_));
 sg13g2_a21oi_1 _5988_ (.A1(_2346_),
    .A2(_2350_),
    .Y(_2353_),
    .B1(_2352_));
 sg13g2_a221oi_1 _5989_ (.B2(_1492_),
    .C1(net921),
    .B1(_2353_),
    .A1(_1544_),
    .Y(_2354_),
    .A2(_2324_));
 sg13g2_a21oi_1 _5990_ (.A1(net995),
    .A2(_1559_),
    .Y(_2355_),
    .B1(_1576_));
 sg13g2_a21oi_1 _5991_ (.A1(net995),
    .A2(_1569_),
    .Y(_2356_),
    .B1(_1579_));
 sg13g2_nor3_1 _5992_ (.A(net922),
    .B(_2355_),
    .C(_2356_),
    .Y(_2357_));
 sg13g2_nor2_1 _5993_ (.A(_2373_),
    .B(_1566_),
    .Y(_2358_));
 sg13g2_nor3_1 _5994_ (.A(net1004),
    .B(_1568_),
    .C(_2358_),
    .Y(_2359_));
 sg13g2_nand2_1 _5995_ (.Y(_2360_),
    .A(net996),
    .B(_1560_));
 sg13g2_a221oi_1 _5996_ (.B2(_2360_),
    .C1(net1000),
    .B1(_1562_),
    .A1(net1003),
    .Y(_2361_),
    .A2(_1560_));
 sg13g2_o21ai_1 _5997_ (.B1(net922),
    .Y(_2362_),
    .A1(_1573_),
    .A2(_2359_));
 sg13g2_nor2_1 _5998_ (.A(net1001),
    .B(_1594_),
    .Y(_2363_));
 sg13g2_o21ai_1 _5999_ (.B1(_2363_),
    .Y(_2364_),
    .A1(_1567_),
    .A2(_1572_));
 sg13g2_nand2b_1 _6000_ (.Y(_2365_),
    .B(_1557_),
    .A_N(_1534_));
 sg13g2_nor2_1 _6001_ (.A(_2374_),
    .B(_1590_),
    .Y(_2366_));
 sg13g2_a21oi_1 _6002_ (.A1(_2365_),
    .A2(_2366_),
    .Y(_2367_),
    .B1(net922));
 sg13g2_a21oi_1 _6003_ (.A1(_2364_),
    .A2(_2367_),
    .Y(_2368_),
    .B1(_1491_));
 sg13g2_o21ai_1 _6004_ (.B1(_2368_),
    .Y(_2369_),
    .A1(_2361_),
    .A2(_2362_));
 sg13g2_o21ai_1 _6005_ (.B1(_2369_),
    .Y(_2370_),
    .A1(_1586_),
    .A2(_2357_));
 sg13g2_o21ai_1 _6006_ (.B1(net1071),
    .Y(_2371_),
    .A1(net997),
    .A2(_2345_));
 sg13g2_a21o_1 _6007_ (.A2(_2370_),
    .A1(net921),
    .B1(_2354_),
    .X(_2372_));
 sg13g2_a21oi_1 _6008_ (.A1(_2345_),
    .A2(_2372_),
    .Y(_0290_),
    .B1(_2371_));
 sg13g2_dfrbp_1 _6009_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net24),
    .D(_0075_),
    .Q_N(_0074_),
    .Q(\i_orchestrator.vga_x[0] ));
 sg13g2_dfrbp_1 _6010_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net136),
    .D(net328),
    .Q_N(_3000_),
    .Q(\i_orchestrator.vga_x[1] ));
 sg13g2_dfrbp_1 _6011_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net135),
    .D(_0077_),
    .Q_N(_2999_),
    .Q(\i_orchestrator.vga_x[2] ));
 sg13g2_dfrbp_1 _6012_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net134),
    .D(_0078_),
    .Q_N(_2998_),
    .Q(\i_orchestrator.vga_x[3] ));
 sg13g2_dfrbp_1 _6013_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net133),
    .D(_0079_),
    .Q_N(_2997_),
    .Q(\i_orchestrator.vga_x[4] ));
 sg13g2_dfrbp_1 _6014_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net132),
    .D(_0080_),
    .Q_N(_2996_),
    .Q(\i_orchestrator.vga_x[5] ));
 sg13g2_dfrbp_1 _6015_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net131),
    .D(_0081_),
    .Q_N(_2995_),
    .Q(\i_orchestrator.vga_x[6] ));
 sg13g2_dfrbp_1 _6016_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net130),
    .D(_0082_),
    .Q_N(_2994_),
    .Q(\i_orchestrator.vga_x[7] ));
 sg13g2_dfrbp_1 _6017_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net129),
    .D(net419),
    .Q_N(_2993_),
    .Q(\i_orchestrator.vga_x[8] ));
 sg13g2_dfrbp_1 _6018_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net128),
    .D(_0084_),
    .Q_N(_2992_),
    .Q(\i_orchestrator.vga_x[9] ));
 sg13g2_dfrbp_1 _6019_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net127),
    .D(_0085_),
    .Q_N(_2991_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _6020_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net126),
    .D(net392),
    .Q_N(_2990_),
    .Q(orient));
 sg13g2_dfrbp_1 _6021_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net124),
    .D(_0087_),
    .Q_N(_2989_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _6022_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net123),
    .D(_0088_),
    .Q_N(_0073_),
    .Q(\i_orchestrator.vga_y[0] ));
 sg13g2_dfrbp_1 _6023_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net121),
    .D(_0089_),
    .Q_N(_2988_),
    .Q(\i_orchestrator.vga_y[1] ));
 sg13g2_dfrbp_1 _6024_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net119),
    .D(_0090_),
    .Q_N(_2987_),
    .Q(\i_orchestrator.vga_y[2] ));
 sg13g2_dfrbp_1 _6025_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net117),
    .D(_0091_),
    .Q_N(_2986_),
    .Q(\i_orchestrator.vga_y[3] ));
 sg13g2_dfrbp_1 _6026_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net115),
    .D(_0092_),
    .Q_N(_2985_),
    .Q(\i_orchestrator.vga_y[4] ));
 sg13g2_dfrbp_1 _6027_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net113),
    .D(_0093_),
    .Q_N(_2984_),
    .Q(\i_orchestrator.vga_y[5] ));
 sg13g2_dfrbp_1 _6028_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net111),
    .D(net429),
    .Q_N(_2983_),
    .Q(\i_orchestrator.vga_y[6] ));
 sg13g2_dfrbp_1 _6029_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net109),
    .D(_0095_),
    .Q_N(_2982_),
    .Q(\i_orchestrator.vga_y[7] ));
 sg13g2_dfrbp_1 _6030_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net107),
    .D(_0096_),
    .Q_N(_2981_),
    .Q(\i_orchestrator.vga_y[8] ));
 sg13g2_dfrbp_1 _6031_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net105),
    .D(net384),
    .Q_N(_2980_),
    .Q(\i_orchestrator.vga_y[9] ));
 sg13g2_dfrbp_1 _6032_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net103),
    .D(net310),
    .Q_N(_0057_),
    .Q(\i_transform.track_y[0] ));
 sg13g2_dfrbp_1 _6033_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net102),
    .D(_0099_),
    .Q_N(_2979_),
    .Q(\i_transform.track_y[1] ));
 sg13g2_dfrbp_1 _6034_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net101),
    .D(net318),
    .Q_N(_2978_),
    .Q(\i_transform.track_y[2] ));
 sg13g2_dfrbp_1 _6035_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net100),
    .D(net298),
    .Q_N(_0058_),
    .Q(\i_transform.track_y[3] ));
 sg13g2_dfrbp_1 _6036_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net25),
    .D(net316),
    .Q_N(_0061_),
    .Q(\i_transform.track_y[4] ));
 sg13g2_dfrbp_1 _6037_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net75),
    .D(_0007_),
    .Q_N(_3001_),
    .Q(\i_vga_beam.vsync ));
 sg13g2_dfrbp_1 _6038_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net99),
    .D(_0006_),
    .Q_N(_2977_),
    .Q(hsync));
 sg13g2_dfrbp_1 _6039_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net98),
    .D(_0103_),
    .Q_N(_0033_),
    .Q(\i_transform.image_y[5] ));
 sg13g2_dfrbp_1 _6040_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net93),
    .D(_0104_),
    .Q_N(_0032_),
    .Q(\i_capsule.tf_y[0] ));
 sg13g2_dfrbp_1 _6041_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net91),
    .D(_0105_),
    .Q_N(_0031_),
    .Q(\i_bitmap.in[7] ));
 sg13g2_dfrbp_1 _6042_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net89),
    .D(_0106_),
    .Q_N(_0034_),
    .Q(\i_bitmap.in[8] ));
 sg13g2_dfrbp_1 _6043_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net87),
    .D(_0107_),
    .Q_N(_0035_),
    .Q(\i_bitmap.in[9] ));
 sg13g2_dfrbp_1 _6044_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net85),
    .D(_0108_),
    .Q_N(_0036_),
    .Q(\i_bitmap.in[10] ));
 sg13g2_dfrbp_1 _6045_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net83),
    .D(_0109_),
    .Q_N(_0037_),
    .Q(\i_bitmap.in[11] ));
 sg13g2_dfrbp_1 _6046_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net81),
    .D(_0110_),
    .Q_N(_0038_),
    .Q(\i_bitmap.in[12] ));
 sg13g2_dfrbp_1 _6047_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net79),
    .D(_0111_),
    .Q_N(_0040_),
    .Q(\i_capsule.tf_y[7] ));
 sg13g2_dfrbp_1 _6048_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net77),
    .D(_0112_),
    .Q_N(_0041_),
    .Q(\i_capsule.tf_y[8] ));
 sg13g2_dfrbp_1 _6049_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net74),
    .D(_0113_),
    .Q_N(_0042_),
    .Q(\i_capsule.tf_y[9] ));
 sg13g2_dfrbp_1 _6050_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net72),
    .D(net427),
    .Q_N(_0004_),
    .Q(\i_orchestrator.trigger_debounce ));
 sg13g2_dfrbp_1 _6051_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net70),
    .D(net241),
    .Q_N(_0072_),
    .Q(\i_orchestrator.hit_priority[0] ));
 sg13g2_dfrbp_1 _6052_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net68),
    .D(net350),
    .Q_N(_2976_),
    .Q(\i_orchestrator.hit_priority[1] ));
 sg13g2_dfrbp_1 _6053_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net66),
    .D(_0117_),
    .Q_N(_0053_),
    .Q(\i_collision.i_coll_table.in[0] ));
 sg13g2_dfrbp_1 _6054_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net64),
    .D(_0118_),
    .Q_N(_2975_),
    .Q(\i_orchestrator.lfsr[1] ));
 sg13g2_dfrbp_1 _6055_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net62),
    .D(_0119_),
    .Q_N(_2974_),
    .Q(\i_orchestrator.lfsr[2] ));
 sg13g2_dfrbp_1 _6056_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net60),
    .D(_0120_),
    .Q_N(_2973_),
    .Q(\i_orchestrator.lfsr[3] ));
 sg13g2_dfrbp_1 _6057_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net58),
    .D(net267),
    .Q_N(_2972_),
    .Q(\i_orchestrator.lfsr[4] ));
 sg13g2_dfrbp_1 _6058_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net56),
    .D(net269),
    .Q_N(_2971_),
    .Q(\i_orchestrator.lfsr[5] ));
 sg13g2_dfrbp_1 _6059_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net54),
    .D(_0123_),
    .Q_N(_2970_),
    .Q(\i_orchestrator.lfsr[6] ));
 sg13g2_dfrbp_1 _6060_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net52),
    .D(net280),
    .Q_N(_2969_),
    .Q(\i_orchestrator.lfsr[7] ));
 sg13g2_dfrbp_1 _6061_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net50),
    .D(_0125_),
    .Q_N(_0044_),
    .Q(\color_entropy[0] ));
 sg13g2_dfrbp_1 _6062_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net48),
    .D(_0126_),
    .Q_N(_2968_),
    .Q(\color_entropy[1] ));
 sg13g2_dfrbp_1 _6063_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net46),
    .D(_0127_),
    .Q_N(_0005_),
    .Q(\i_orchestrator.hit_bottom ));
 sg13g2_dfrbp_1 _6064_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net44),
    .D(_0128_),
    .Q_N(_0010_),
    .Q(\i_orchestrator.hit_top ));
 sg13g2_dfrbp_1 _6065_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net42),
    .D(_0129_),
    .Q_N(_0055_),
    .Q(\i_orchestrator.hit_right ));
 sg13g2_dfrbp_1 _6066_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net40),
    .D(_0130_),
    .Q_N(_0011_),
    .Q(\i_orchestrator.hit_left ));
 sg13g2_dfrbp_1 _6067_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net38),
    .D(_0131_),
    .Q_N(_2967_),
    .Q(handle_impact));
 sg13g2_dfrbp_1 _6068_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net37),
    .D(net243),
    .Q_N(_0069_),
    .Q(\i_orchestrator.update_resonator ));
 sg13g2_dfrbp_1 _6069_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net36),
    .D(_0133_),
    .Q_N(_2966_),
    .Q(\i_orchestrator.update_transform ));
 sg13g2_dfrbp_1 _6070_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net35),
    .D(_0134_),
    .Q_N(_2965_),
    .Q(\i_kinematics.update ));
 sg13g2_dfrbp_1 _6071_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net34),
    .D(_0135_),
    .Q_N(_2964_),
    .Q(\i_collision.mirror ));
 sg13g2_dfrbp_1 _6072_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net33),
    .D(_0136_),
    .Q_N(_2963_),
    .Q(\i_collision.rotate ));
 sg13g2_dfrbp_1 _6073_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net32),
    .D(net246),
    .Q_N(_2962_),
    .Q(\i_collision.update ));
 sg13g2_dfrbp_1 _6074_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net31),
    .D(_0138_),
    .Q_N(_2961_),
    .Q(\i_delta_sigma.acc[0] ));
 sg13g2_dfrbp_1 _6075_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net30),
    .D(_0139_),
    .Q_N(_2960_),
    .Q(\i_delta_sigma.acc[1] ));
 sg13g2_dfrbp_1 _6076_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net29),
    .D(_0140_),
    .Q_N(_2959_),
    .Q(\i_delta_sigma.acc[2] ));
 sg13g2_dfrbp_1 _6077_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net28),
    .D(net411),
    .Q_N(_2958_),
    .Q(\i_delta_sigma.acc[3] ));
 sg13g2_dfrbp_1 _6078_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net27),
    .D(net368),
    .Q_N(_2957_),
    .Q(\i_delta_sigma.acc[4] ));
 sg13g2_dfrbp_1 _6079_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net26),
    .D(_0143_),
    .Q_N(_2956_),
    .Q(\i_delta_sigma.acc[5] ));
 sg13g2_dfrbp_1 _6080_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net23),
    .D(_0144_),
    .Q_N(_2955_),
    .Q(\i_delta_sigma.acc[6] ));
 sg13g2_dfrbp_1 _6081_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net22),
    .D(net507),
    .Q_N(_2954_),
    .Q(\i_delta_sigma.acc[7] ));
 sg13g2_dfrbp_1 _6082_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net21),
    .D(net380),
    .Q_N(_2953_),
    .Q(\i_delta_sigma.acc[8] ));
 sg13g2_dfrbp_1 _6083_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net20),
    .D(_0147_),
    .Q_N(_2952_),
    .Q(\i_delta_sigma.acc[9] ));
 sg13g2_dfrbp_1 _6084_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net19),
    .D(_0148_),
    .Q_N(_2951_),
    .Q(\i_delta_sigma.acc[10] ));
 sg13g2_dfrbp_1 _6085_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net18),
    .D(_0149_),
    .Q_N(_2950_),
    .Q(\i_delta_sigma.acc[11] ));
 sg13g2_dfrbp_1 _6086_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net17),
    .D(_0150_),
    .Q_N(_2949_),
    .Q(\i_delta_sigma.acc[12] ));
 sg13g2_dfrbp_1 _6087_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net94),
    .D(_0151_),
    .Q_N(_0054_),
    .Q(\i_delta_sigma.acc[13] ));
 sg13g2_dfrbp_1 _6088_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net16),
    .D(_0000_),
    .Q_N(_2948_),
    .Q(bitmap_pixel));
 sg13g2_dfrbp_1 _6089_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net15),
    .D(net345),
    .Q_N(_0019_),
    .Q(\i_transform.image_x[5] ));
 sg13g2_dfrbp_1 _6090_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net13),
    .D(_0153_),
    .Q_N(_0021_),
    .Q(\i_capsule.tf_x[0] ));
 sg13g2_dfrbp_1 _6091_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net11),
    .D(_0154_),
    .Q_N(_0018_),
    .Q(\i_bitmap.in[0] ));
 sg13g2_dfrbp_1 _6092_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net9),
    .D(_0155_),
    .Q_N(_0017_),
    .Q(\i_bitmap.in[1] ));
 sg13g2_dfrbp_1 _6093_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net229),
    .D(_0156_),
    .Q_N(_0026_),
    .Q(\i_bitmap.in[2] ));
 sg13g2_dfrbp_1 _6094_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net227),
    .D(_0157_),
    .Q_N(_0027_),
    .Q(\i_bitmap.in[3] ));
 sg13g2_dfrbp_1 _6095_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net225),
    .D(_0158_),
    .Q_N(_0028_),
    .Q(\i_bitmap.in[4] ));
 sg13g2_dfrbp_1 _6096_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net223),
    .D(_0159_),
    .Q_N(_0029_),
    .Q(\i_bitmap.in[5] ));
 sg13g2_dfrbp_1 _6097_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net221),
    .D(_0160_),
    .Q_N(_0030_),
    .Q(\i_bitmap.in[6] ));
 sg13g2_dfrbp_1 _6098_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net219),
    .D(_0161_),
    .Q_N(_0039_),
    .Q(\i_capsule.tf_x[8] ));
 sg13g2_dfrbp_1 _6099_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net217),
    .D(_0162_),
    .Q_N(_0056_),
    .Q(\i_capsule.tf_x[9] ));
 sg13g2_dfrbp_1 _6100_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net215),
    .D(net371),
    .Q_N(_0060_),
    .Q(\i_transform.track_y[5] ));
 sg13g2_dfrbp_1 _6101_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net214),
    .D(net485),
    .Q_N(_2947_),
    .Q(\i_transform.track_y[6] ));
 sg13g2_dfrbp_1 _6102_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net213),
    .D(_0165_),
    .Q_N(_0059_),
    .Q(\i_transform.track_y[7] ));
 sg13g2_dfrbp_1 _6103_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net212),
    .D(net397),
    .Q_N(_2946_),
    .Q(\i_transform.track_y[8] ));
 sg13g2_dfrbp_1 _6104_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net211),
    .D(_0167_),
    .Q_N(_0062_),
    .Q(\i_transform.track_y[9] ));
 sg13g2_dfrbp_1 _6105_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net210),
    .D(net257),
    .Q_N(_2945_),
    .Q(\i_orchestrator.trigger_resonator[0] ));
 sg13g2_dfrbp_1 _6106_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net95),
    .D(net263),
    .Q_N(_3002_),
    .Q(\i_orchestrator.trigger_resonator[1] ));
 sg13g2_dfrbp_1 _6107_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net96),
    .D(_0001_),
    .Q_N(_3003_),
    .Q(\i_colors.channel[0] ));
 sg13g2_dfrbp_1 _6108_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net53),
    .D(net424),
    .Q_N(_0043_),
    .Q(\i_colors.channel[1] ));
 sg13g2_dfrbp_1 _6109_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net209),
    .D(net433),
    .Q_N(_2944_),
    .Q(\i_colors.channel[2] ));
 sg13g2_dfrbp_1 _6110_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net208),
    .D(_0170_),
    .Q_N(_2943_),
    .Q(\collision_impact[0] ));
 sg13g2_dfrbp_1 _6111_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net206),
    .D(_0171_),
    .Q_N(_2942_),
    .Q(\collision_impact[1] ));
 sg13g2_dfrbp_1 _6112_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net204),
    .D(_0172_),
    .Q_N(_0008_),
    .Q(\i_collision.vy[0] ));
 sg13g2_dfrbp_1 _6113_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net202),
    .D(_0173_),
    .Q_N(_2941_),
    .Q(\i_collision.vy[1] ));
 sg13g2_dfrbp_1 _6114_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net200),
    .D(net523),
    .Q_N(_2940_),
    .Q(\i_collision.vy[2] ));
 sg13g2_dfrbp_1 _6115_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net198),
    .D(net386),
    .Q_N(_0009_),
    .Q(\i_collision.vx[0] ));
 sg13g2_dfrbp_1 _6116_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net196),
    .D(net500),
    .Q_N(_2939_),
    .Q(\i_collision.vx[1] ));
 sg13g2_dfrbp_1 _6117_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net194),
    .D(net545),
    .Q_N(_2938_),
    .Q(\i_collision.vx[2] ));
 sg13g2_dfrbp_1 _6118_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net192),
    .D(net253),
    .Q_N(_2937_),
    .Q(\i_kinematics.center_y_lo[0] ));
 sg13g2_dfrbp_1 _6119_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net190),
    .D(net363),
    .Q_N(_2936_),
    .Q(\i_kinematics.center_y_lo[1] ));
 sg13g2_dfrbp_1 _6120_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net188),
    .D(net255),
    .Q_N(_2935_),
    .Q(\i_kinematics.center_x_lo[0] ));
 sg13g2_dfrbp_1 _6121_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net186),
    .D(net361),
    .Q_N(_2934_),
    .Q(\i_kinematics.center_x_lo[1] ));
 sg13g2_dfrbp_1 _6122_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net184),
    .D(_0182_),
    .Q_N(_2933_),
    .Q(\center_y[0] ));
 sg13g2_dfrbp_1 _6123_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net182),
    .D(_0183_),
    .Q_N(_2932_),
    .Q(\center_y[1] ));
 sg13g2_dfrbp_1 _6124_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net180),
    .D(_0184_),
    .Q_N(_2931_),
    .Q(\center_y[2] ));
 sg13g2_dfrbp_1 _6125_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net178),
    .D(_0185_),
    .Q_N(_2930_),
    .Q(\center_y[3] ));
 sg13g2_dfrbp_1 _6126_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net176),
    .D(net462),
    .Q_N(_2929_),
    .Q(\center_y[4] ));
 sg13g2_dfrbp_1 _6127_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net174),
    .D(_0187_),
    .Q_N(_2928_),
    .Q(\center_y[5] ));
 sg13g2_dfrbp_1 _6128_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net172),
    .D(net452),
    .Q_N(_2927_),
    .Q(\center_y[6] ));
 sg13g2_dfrbp_1 _6129_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net170),
    .D(net448),
    .Q_N(_2926_),
    .Q(\center_y[7] ));
 sg13g2_dfrbp_1 _6130_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net168),
    .D(_0190_),
    .Q_N(_2925_),
    .Q(\center_y[8] ));
 sg13g2_dfrbp_1 _6131_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net166),
    .D(_0191_),
    .Q_N(_2924_),
    .Q(\center_y[9] ));
 sg13g2_dfrbp_1 _6132_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net164),
    .D(_0192_),
    .Q_N(_2923_),
    .Q(\center_x[0] ));
 sg13g2_dfrbp_1 _6133_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net162),
    .D(_0193_),
    .Q_N(_2922_),
    .Q(\center_x[1] ));
 sg13g2_dfrbp_1 _6134_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net160),
    .D(_0194_),
    .Q_N(_2921_),
    .Q(\center_x[2] ));
 sg13g2_dfrbp_1 _6135_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net158),
    .D(net509),
    .Q_N(_2920_),
    .Q(\center_x[3] ));
 sg13g2_dfrbp_1 _6136_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net156),
    .D(net442),
    .Q_N(_2919_),
    .Q(\center_x[4] ));
 sg13g2_dfrbp_1 _6137_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net154),
    .D(net444),
    .Q_N(_2918_),
    .Q(\center_x[5] ));
 sg13g2_dfrbp_1 _6138_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net152),
    .D(net478),
    .Q_N(_2917_),
    .Q(\center_x[6] ));
 sg13g2_dfrbp_1 _6139_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net150),
    .D(net480),
    .Q_N(_2916_),
    .Q(\center_x[7] ));
 sg13g2_dfrbp_1 _6140_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net148),
    .D(_0200_),
    .Q_N(_2915_),
    .Q(\center_x[8] ));
 sg13g2_dfrbp_1 _6141_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net146),
    .D(_0201_),
    .Q_N(_2914_),
    .Q(\center_x[9] ));
 sg13g2_dfrbp_1 _6142_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net144),
    .D(_0202_),
    .Q_N(_2913_),
    .Q(\i_kinematics.phi[0] ));
 sg13g2_dfrbp_1 _6143_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net142),
    .D(_0203_),
    .Q_N(_2912_),
    .Q(\i_kinematics.phi[1] ));
 sg13g2_dfrbp_1 _6144_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net140),
    .D(_0204_),
    .Q_N(_2911_),
    .Q(\i_kinematics.phi[2] ));
 sg13g2_dfrbp_1 _6145_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net138),
    .D(_0205_),
    .Q_N(_2910_),
    .Q(\i_kinematics.phi[3] ));
 sg13g2_dfrbp_1 _6146_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net125),
    .D(_0206_),
    .Q_N(_2909_),
    .Q(\i_kinematics.phi[4] ));
 sg13g2_dfrbp_1 _6147_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net120),
    .D(_0207_),
    .Q_N(_2908_),
    .Q(\i_kinematics.phi[5] ));
 sg13g2_dfrbp_1 _6148_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net116),
    .D(_0208_),
    .Q_N(_2907_),
    .Q(\i_kinematics.phi[6] ));
 sg13g2_dfrbp_1 _6149_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net112),
    .D(_0209_),
    .Q_N(_2906_),
    .Q(\i_kinematics.phi[7] ));
 sg13g2_dfrbp_1 _6150_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net108),
    .D(_0210_),
    .Q_N(_0050_),
    .Q(\i_collision.i_coll_table.in[1] ));
 sg13g2_dfrbp_1 _6151_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net104),
    .D(_0211_),
    .Q_N(_2905_),
    .Q(\i_collision.phi[1] ));
 sg13g2_dfrbp_1 _6152_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net92),
    .D(_0212_),
    .Q_N(_2904_),
    .Q(\i_kinematics.phi[10] ));
 sg13g2_dfrbp_1 _6153_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net88),
    .D(net312),
    .Q_N(_0012_),
    .Q(\i_transform.image_y[0] ));
 sg13g2_dfrbp_1 _6154_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net84),
    .D(_0214_),
    .Q_N(_0013_),
    .Q(\i_transform.image_y[1] ));
 sg13g2_dfrbp_1 _6155_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net80),
    .D(_0215_),
    .Q_N(_0014_),
    .Q(\i_transform.image_y[2] ));
 sg13g2_dfrbp_1 _6156_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net76),
    .D(_0216_),
    .Q_N(_0015_),
    .Q(\i_transform.image_y[3] ));
 sg13g2_dfrbp_1 _6157_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net71),
    .D(_0217_),
    .Q_N(_0016_),
    .Q(\i_transform.image_y[4] ));
 sg13g2_dfrbp_1 _6158_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net67),
    .D(net286),
    .Q_N(_0025_),
    .Q(\i_transform.image_x[0] ));
 sg13g2_dfrbp_1 _6159_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net63),
    .D(_0219_),
    .Q_N(_0024_),
    .Q(\i_transform.image_x[1] ));
 sg13g2_dfrbp_1 _6160_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net59),
    .D(_0220_),
    .Q_N(_0023_),
    .Q(\i_transform.image_x[2] ));
 sg13g2_dfrbp_1 _6161_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net55),
    .D(_0221_),
    .Q_N(_0022_),
    .Q(\i_transform.image_x[3] ));
 sg13g2_dfrbp_1 _6162_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net51),
    .D(_0222_),
    .Q_N(_0020_),
    .Q(\i_transform.image_x[4] ));
 sg13g2_dfrbp_1 _6163_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net47),
    .D(net352),
    .Q_N(_0063_),
    .Q(\i_transform.track_x[0] ));
 sg13g2_dfrbp_1 _6164_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net45),
    .D(net472),
    .Q_N(_2903_),
    .Q(\i_transform.track_x[1] ));
 sg13g2_dfrbp_1 _6165_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net43),
    .D(_0225_),
    .Q_N(_2902_),
    .Q(\i_transform.track_x[2] ));
 sg13g2_dfrbp_1 _6166_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net41),
    .D(net265),
    .Q_N(_0064_),
    .Q(\i_transform.track_x[3] ));
 sg13g2_dfrbp_1 _6167_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net39),
    .D(net402),
    .Q_N(_0067_),
    .Q(\i_transform.track_x[4] ));
 sg13g2_dfrbp_1 _6168_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net14),
    .D(_0228_),
    .Q_N(_0071_),
    .Q(\i_orchestrator.sample_counter[0] ));
 sg13g2_dfrbp_1 _6169_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net12),
    .D(net375),
    .Q_N(_2901_),
    .Q(\i_orchestrator.sample_counter[1] ));
 sg13g2_dfrbp_1 _6170_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net10),
    .D(_0230_),
    .Q_N(_2900_),
    .Q(\i_orchestrator.sample_counter[2] ));
 sg13g2_dfrbp_1 _6171_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net230),
    .D(net273),
    .Q_N(_2899_),
    .Q(\i_orchestrator.sample_counter[3] ));
 sg13g2_dfrbp_1 _6172_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net228),
    .D(_0232_),
    .Q_N(_2898_),
    .Q(\i_orchestrator.sample_counter[4] ));
 sg13g2_dfrbp_1 _6173_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net226),
    .D(_0233_),
    .Q_N(_2897_),
    .Q(\i_orchestrator.sample_counter[5] ));
 sg13g2_dfrbp_1 _6174_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net224),
    .D(_0234_),
    .Q_N(_2896_),
    .Q(\i_orchestrator.sample_counter[6] ));
 sg13g2_dfrbp_1 _6175_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net222),
    .D(net276),
    .Q_N(_2895_),
    .Q(\i_orchestrator.sample_counter[7] ));
 sg13g2_dfrbp_1 _6176_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net220),
    .D(net282),
    .Q_N(_2894_),
    .Q(\i_orchestrator.sample_counter[8] ));
 sg13g2_dfrbp_1 _6177_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net218),
    .D(_0237_),
    .Q_N(_2893_),
    .Q(\i_orchestrator.sample_counter[9] ));
 sg13g2_dfrbp_1 _6178_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net216),
    .D(net248),
    .Q_N(_2892_),
    .Q(\i_orchestrator.tension[1] ));
 sg13g2_dfrbp_1 _6179_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net205),
    .D(net324),
    .Q_N(_2891_),
    .Q(\i_orchestrator.tension[2] ));
 sg13g2_dfrbp_1 _6180_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net201),
    .D(net261),
    .Q_N(_2890_),
    .Q(\i_orchestrator.tension[3] ));
 sg13g2_dfrbp_1 _6181_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net197),
    .D(net330),
    .Q_N(_2889_),
    .Q(\capsule_color[0] ));
 sg13g2_dfrbp_1 _6182_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net193),
    .D(_0242_),
    .Q_N(_2888_),
    .Q(\capsule_color[1] ));
 sg13g2_dfrbp_1 _6183_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net189),
    .D(_0243_),
    .Q_N(_2887_),
    .Q(\capsule_color[2] ));
 sg13g2_dfrbp_1 _6184_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net185),
    .D(_0244_),
    .Q_N(_2886_),
    .Q(\capsule_color[3] ));
 sg13g2_dfrbp_1 _6185_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net181),
    .D(net341),
    .Q_N(_2885_),
    .Q(\i_colors.capsule_color[4] ));
 sg13g2_dfrbp_1 _6186_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net177),
    .D(net359),
    .Q_N(_2884_),
    .Q(\i_colors.capsule_color[5] ));
 sg13g2_dfrbp_1 _6187_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net173),
    .D(net288),
    .Q_N(_0066_),
    .Q(\i_transform.track_x[5] ));
 sg13g2_dfrbp_1 _6188_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net171),
    .D(net526),
    .Q_N(_2883_),
    .Q(\i_transform.track_x[6] ));
 sg13g2_dfrbp_1 _6189_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net169),
    .D(_0249_),
    .Q_N(_0065_),
    .Q(\i_transform.track_x[7] ));
 sg13g2_dfrbp_1 _6190_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net167),
    .D(_0250_),
    .Q_N(_2882_),
    .Q(\i_transform.track_x[8] ));
 sg13g2_dfrbp_1 _6191_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net165),
    .D(_0251_),
    .Q_N(_0068_),
    .Q(\i_transform.track_x[9] ));
 sg13g2_dfrbp_1 _6192_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net163),
    .D(net395),
    .Q_N(_2881_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _6193_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net161),
    .D(_0253_),
    .Q_N(_2880_),
    .Q(\i_delta_sigma.sample[11] ));
 sg13g2_dfrbp_1 _6194_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net157),
    .D(net357),
    .Q_N(_2879_),
    .Q(\i_delta_sigma.sample[0] ));
 sg13g2_dfrbp_1 _6195_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net153),
    .D(_0255_),
    .Q_N(_2878_),
    .Q(\i_delta_sigma.sample[1] ));
 sg13g2_dfrbp_1 _6196_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net149),
    .D(_0256_),
    .Q_N(_2877_),
    .Q(\i_delta_sigma.sample[2] ));
 sg13g2_dfrbp_1 _6197_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net145),
    .D(_0257_),
    .Q_N(_2876_),
    .Q(\i_delta_sigma.sample[3] ));
 sg13g2_dfrbp_1 _6198_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net141),
    .D(_0258_),
    .Q_N(_2875_),
    .Q(\i_delta_sigma.sample[4] ));
 sg13g2_dfrbp_1 _6199_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net137),
    .D(_0259_),
    .Q_N(_2874_),
    .Q(\i_delta_sigma.sample[5] ));
 sg13g2_dfrbp_1 _6200_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net118),
    .D(_0260_),
    .Q_N(_2873_),
    .Q(\i_delta_sigma.sample[6] ));
 sg13g2_dfrbp_1 _6201_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net110),
    .D(_0261_),
    .Q_N(_2872_),
    .Q(\i_delta_sigma.sample[7] ));
 sg13g2_dfrbp_1 _6202_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net97),
    .D(_0262_),
    .Q_N(_2871_),
    .Q(\i_delta_sigma.sample[8] ));
 sg13g2_dfrbp_1 _6203_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net86),
    .D(_0263_),
    .Q_N(_2870_),
    .Q(\i_delta_sigma.sample[9] ));
 sg13g2_dfrbp_1 _6204_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net78),
    .D(_0264_),
    .Q_N(_2869_),
    .Q(\i_delta_sigma.sample[10] ));
 sg13g2_dfrbp_1 _6205_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net69),
    .D(_0265_),
    .Q_N(_2868_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _6206_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net65),
    .D(net332),
    .Q_N(_0045_),
    .Q(\i_resonator.v[0] ));
 sg13g2_dfrbp_1 _6207_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net57),
    .D(_0267_),
    .Q_N(_2867_),
    .Q(\i_resonator.v[1] ));
 sg13g2_dfrbp_1 _6208_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net49),
    .D(_0268_),
    .Q_N(_2866_),
    .Q(\i_resonator.v[2] ));
 sg13g2_dfrbp_1 _6209_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net203),
    .D(_0269_),
    .Q_N(_2865_),
    .Q(\i_resonator.v[3] ));
 sg13g2_dfrbp_1 _6210_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net195),
    .D(_0270_),
    .Q_N(_2864_),
    .Q(\i_resonator.v[4] ));
 sg13g2_dfrbp_1 _6211_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net187),
    .D(_0271_),
    .Q_N(_2863_),
    .Q(\i_resonator.v[5] ));
 sg13g2_dfrbp_1 _6212_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net179),
    .D(_0272_),
    .Q_N(_2862_),
    .Q(\i_resonator.v[6] ));
 sg13g2_dfrbp_1 _6213_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net159),
    .D(_0273_),
    .Q_N(_2861_),
    .Q(\i_resonator.v[7] ));
 sg13g2_dfrbp_1 _6214_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net151),
    .D(_0274_),
    .Q_N(_2860_),
    .Q(\i_resonator.v[8] ));
 sg13g2_dfrbp_1 _6215_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net143),
    .D(_0275_),
    .Q_N(_0047_),
    .Q(\i_resonator.v[9] ));
 sg13g2_dfrbp_1 _6216_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net122),
    .D(_0276_),
    .Q_N(_2859_),
    .Q(\i_resonator.v[10] ));
 sg13g2_dfrbp_1 _6217_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net106),
    .D(_0277_),
    .Q_N(_0046_),
    .Q(\i_resonator.v[11] ));
 sg13g2_dfrbp_1 _6218_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net82),
    .D(_0278_),
    .Q_N(_2858_),
    .Q(\i_resonator.v[12] ));
 sg13g2_dfrbp_1 _6219_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net61),
    .D(_0279_),
    .Q_N(_0048_),
    .Q(\i_resonator.v[13] ));
 sg13g2_dfrbp_1 _6220_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net207),
    .D(_0280_),
    .Q_N(_2857_),
    .Q(\i_resonator.v[14] ));
 sg13g2_dfrbp_1 _6221_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net191),
    .D(_0281_),
    .Q_N(_0049_),
    .Q(\i_resonator.v[15] ));
 sg13g2_dfrbp_1 _6222_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net175),
    .D(net291),
    .Q_N(_2856_),
    .Q(\i_resonator.counter[0] ));
 sg13g2_dfrbp_1 _6223_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net147),
    .D(_0283_),
    .Q_N(_2855_),
    .Q(\i_resonator.counter[1] ));
 sg13g2_dfrbp_1 _6224_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net114),
    .D(_0284_),
    .Q_N(_2854_),
    .Q(\i_resonator.counter[2] ));
 sg13g2_dfrbp_1 _6225_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net73),
    .D(_0285_),
    .Q_N(_2853_),
    .Q(\i_resonator.counter[3] ));
 sg13g2_dfrbp_1 _6226_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net199),
    .D(_0286_),
    .Q_N(_0052_),
    .Q(\i_collision.i_coll_table.in[4] ));
 sg13g2_dfrbp_1 _6227_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net155),
    .D(net416),
    .Q_N(_2852_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _6228_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net139),
    .D(_0288_),
    .Q_N(_2851_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _6229_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net90),
    .D(_0289_),
    .Q_N(_0070_),
    .Q(\i_collision.i_coll_table.in[5] ));
 sg13g2_dfrbp_1 _6230_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net183),
    .D(net513),
    .Q_N(_0051_),
    .Q(\i_collision.i_coll_table.in[3] ));
 sg13g2_tiehi _6170__10 (.L_HI(net10));
 sg13g2_tiehi _6091__11 (.L_HI(net11));
 sg13g2_tiehi _6169__12 (.L_HI(net12));
 sg13g2_tiehi _6090__13 (.L_HI(net13));
 sg13g2_tiehi _6168__14 (.L_HI(net14));
 sg13g2_tiehi _6089__15 (.L_HI(net15));
 sg13g2_tiehi _6088__16 (.L_HI(net16));
 sg13g2_tiehi _6086__17 (.L_HI(net17));
 sg13g2_tiehi _6085__18 (.L_HI(net18));
 sg13g2_tiehi _6084__19 (.L_HI(net19));
 sg13g2_tiehi _6083__20 (.L_HI(net20));
 sg13g2_tiehi _6082__21 (.L_HI(net21));
 sg13g2_tiehi _6081__22 (.L_HI(net22));
 sg13g2_tiehi _6080__23 (.L_HI(net23));
 sg13g2_tiehi _6009__24 (.L_HI(net24));
 sg13g2_tiehi _6036__25 (.L_HI(net25));
 sg13g2_tiehi _6079__26 (.L_HI(net26));
 sg13g2_tiehi _6078__27 (.L_HI(net27));
 sg13g2_tiehi _6077__28 (.L_HI(net28));
 sg13g2_tiehi _6076__29 (.L_HI(net29));
 sg13g2_tiehi _6075__30 (.L_HI(net30));
 sg13g2_tiehi _6074__31 (.L_HI(net31));
 sg13g2_tiehi _6073__32 (.L_HI(net32));
 sg13g2_tiehi _6072__33 (.L_HI(net33));
 sg13g2_tiehi _6071__34 (.L_HI(net34));
 sg13g2_tiehi _6070__35 (.L_HI(net35));
 sg13g2_tiehi _6069__36 (.L_HI(net36));
 sg13g2_tiehi _6068__37 (.L_HI(net37));
 sg13g2_tiehi _6067__38 (.L_HI(net38));
 sg13g2_tiehi _6167__39 (.L_HI(net39));
 sg13g2_tiehi _6066__40 (.L_HI(net40));
 sg13g2_tiehi _6166__41 (.L_HI(net41));
 sg13g2_tiehi _6065__42 (.L_HI(net42));
 sg13g2_tiehi _6165__43 (.L_HI(net43));
 sg13g2_tiehi _6064__44 (.L_HI(net44));
 sg13g2_tiehi _6164__45 (.L_HI(net45));
 sg13g2_tiehi _6063__46 (.L_HI(net46));
 sg13g2_tiehi _6163__47 (.L_HI(net47));
 sg13g2_tiehi _6062__48 (.L_HI(net48));
 sg13g2_tiehi _6208__49 (.L_HI(net49));
 sg13g2_tiehi _6061__50 (.L_HI(net50));
 sg13g2_tiehi _6162__51 (.L_HI(net51));
 sg13g2_tiehi _6060__52 (.L_HI(net52));
 sg13g2_tiehi _6108__53 (.L_HI(net53));
 sg13g2_tiehi _6059__54 (.L_HI(net54));
 sg13g2_tiehi _6161__55 (.L_HI(net55));
 sg13g2_tiehi _6058__56 (.L_HI(net56));
 sg13g2_tiehi _6207__57 (.L_HI(net57));
 sg13g2_tiehi _6057__58 (.L_HI(net58));
 sg13g2_tiehi _6160__59 (.L_HI(net59));
 sg13g2_tiehi _6056__60 (.L_HI(net60));
 sg13g2_tiehi _6219__61 (.L_HI(net61));
 sg13g2_tiehi _6055__62 (.L_HI(net62));
 sg13g2_tiehi _6159__63 (.L_HI(net63));
 sg13g2_tiehi _6054__64 (.L_HI(net64));
 sg13g2_tiehi _6206__65 (.L_HI(net65));
 sg13g2_tiehi _6053__66 (.L_HI(net66));
 sg13g2_tiehi _6158__67 (.L_HI(net67));
 sg13g2_tiehi _6052__68 (.L_HI(net68));
 sg13g2_tiehi _6205__69 (.L_HI(net69));
 sg13g2_tiehi _6051__70 (.L_HI(net70));
 sg13g2_tiehi _6157__71 (.L_HI(net71));
 sg13g2_tiehi _6050__72 (.L_HI(net72));
 sg13g2_tiehi _6225__73 (.L_HI(net73));
 sg13g2_tiehi _6049__74 (.L_HI(net74));
 sg13g2_tiehi _6037__75 (.L_HI(net75));
 sg13g2_tiehi _6156__76 (.L_HI(net76));
 sg13g2_tiehi _6048__77 (.L_HI(net77));
 sg13g2_tiehi _6204__78 (.L_HI(net78));
 sg13g2_tiehi _6047__79 (.L_HI(net79));
 sg13g2_tiehi _6155__80 (.L_HI(net80));
 sg13g2_tiehi _6046__81 (.L_HI(net81));
 sg13g2_tiehi _6218__82 (.L_HI(net82));
 sg13g2_tiehi _6045__83 (.L_HI(net83));
 sg13g2_tiehi _6154__84 (.L_HI(net84));
 sg13g2_tiehi _6044__85 (.L_HI(net85));
 sg13g2_tiehi _6203__86 (.L_HI(net86));
 sg13g2_tiehi _6043__87 (.L_HI(net87));
 sg13g2_tiehi _6153__88 (.L_HI(net88));
 sg13g2_tiehi _6042__89 (.L_HI(net89));
 sg13g2_tiehi _6229__90 (.L_HI(net90));
 sg13g2_tiehi _6041__91 (.L_HI(net91));
 sg13g2_tiehi _6152__92 (.L_HI(net92));
 sg13g2_tiehi _6040__93 (.L_HI(net93));
 sg13g2_tiehi _6087__94 (.L_HI(net94));
 sg13g2_tiehi _6106__95 (.L_HI(net95));
 sg13g2_tiehi _6107__96 (.L_HI(net96));
 sg13g2_tiehi _6202__97 (.L_HI(net97));
 sg13g2_tiehi _6039__98 (.L_HI(net98));
 sg13g2_tiehi _6038__99 (.L_HI(net99));
 sg13g2_tiehi _6035__100 (.L_HI(net100));
 sg13g2_tiehi _6034__101 (.L_HI(net101));
 sg13g2_tiehi _6033__102 (.L_HI(net102));
 sg13g2_tiehi _6032__103 (.L_HI(net103));
 sg13g2_tiehi _6151__104 (.L_HI(net104));
 sg13g2_tiehi _6031__105 (.L_HI(net105));
 sg13g2_tiehi _6217__106 (.L_HI(net106));
 sg13g2_tiehi _6030__107 (.L_HI(net107));
 sg13g2_tiehi _6150__108 (.L_HI(net108));
 sg13g2_tiehi _6029__109 (.L_HI(net109));
 sg13g2_tiehi _6201__110 (.L_HI(net110));
 sg13g2_tiehi _6028__111 (.L_HI(net111));
 sg13g2_tiehi _6149__112 (.L_HI(net112));
 sg13g2_tiehi _6027__113 (.L_HI(net113));
 sg13g2_tiehi _6224__114 (.L_HI(net114));
 sg13g2_tiehi _6026__115 (.L_HI(net115));
 sg13g2_tiehi _6148__116 (.L_HI(net116));
 sg13g2_tiehi _6025__117 (.L_HI(net117));
 sg13g2_tiehi _6200__118 (.L_HI(net118));
 sg13g2_tiehi _6024__119 (.L_HI(net119));
 sg13g2_tiehi _6147__120 (.L_HI(net120));
 sg13g2_tiehi _6023__121 (.L_HI(net121));
 sg13g2_tiehi _6216__122 (.L_HI(net122));
 sg13g2_tiehi _6022__123 (.L_HI(net123));
 sg13g2_tiehi _6021__124 (.L_HI(net124));
 sg13g2_tiehi _6146__125 (.L_HI(net125));
 sg13g2_tiehi _6020__126 (.L_HI(net126));
 sg13g2_tiehi _6019__127 (.L_HI(net127));
 sg13g2_tiehi _6018__128 (.L_HI(net128));
 sg13g2_tiehi _6017__129 (.L_HI(net129));
 sg13g2_tiehi _6016__130 (.L_HI(net130));
 sg13g2_tiehi _6015__131 (.L_HI(net131));
 sg13g2_tiehi _6014__132 (.L_HI(net132));
 sg13g2_tiehi _6013__133 (.L_HI(net133));
 sg13g2_tiehi _6012__134 (.L_HI(net134));
 sg13g2_tiehi _6011__135 (.L_HI(net135));
 sg13g2_tiehi _6010__136 (.L_HI(net136));
 sg13g2_tiehi _6199__137 (.L_HI(net137));
 sg13g2_tiehi _6145__138 (.L_HI(net138));
 sg13g2_tiehi _6228__139 (.L_HI(net139));
 sg13g2_tiehi _6144__140 (.L_HI(net140));
 sg13g2_tiehi _6198__141 (.L_HI(net141));
 sg13g2_tiehi _6143__142 (.L_HI(net142));
 sg13g2_tiehi _6215__143 (.L_HI(net143));
 sg13g2_tiehi _6142__144 (.L_HI(net144));
 sg13g2_tiehi _6197__145 (.L_HI(net145));
 sg13g2_tiehi _6141__146 (.L_HI(net146));
 sg13g2_tiehi _6223__147 (.L_HI(net147));
 sg13g2_tiehi _6140__148 (.L_HI(net148));
 sg13g2_tiehi _6196__149 (.L_HI(net149));
 sg13g2_tiehi _6139__150 (.L_HI(net150));
 sg13g2_tiehi _6214__151 (.L_HI(net151));
 sg13g2_tiehi _6138__152 (.L_HI(net152));
 sg13g2_tiehi _6195__153 (.L_HI(net153));
 sg13g2_tiehi _6137__154 (.L_HI(net154));
 sg13g2_tiehi _6227__155 (.L_HI(net155));
 sg13g2_tiehi _6136__156 (.L_HI(net156));
 sg13g2_tiehi _6194__157 (.L_HI(net157));
 sg13g2_tiehi _6135__158 (.L_HI(net158));
 sg13g2_tiehi _6213__159 (.L_HI(net159));
 sg13g2_tiehi _6134__160 (.L_HI(net160));
 sg13g2_tiehi _6193__161 (.L_HI(net161));
 sg13g2_tiehi _6133__162 (.L_HI(net162));
 sg13g2_tiehi _6192__163 (.L_HI(net163));
 sg13g2_tiehi _6132__164 (.L_HI(net164));
 sg13g2_tiehi _6191__165 (.L_HI(net165));
 sg13g2_tiehi _6131__166 (.L_HI(net166));
 sg13g2_tiehi _6190__167 (.L_HI(net167));
 sg13g2_tiehi _6130__168 (.L_HI(net168));
 sg13g2_tiehi _6189__169 (.L_HI(net169));
 sg13g2_tiehi _6129__170 (.L_HI(net170));
 sg13g2_tiehi _6188__171 (.L_HI(net171));
 sg13g2_tiehi _6128__172 (.L_HI(net172));
 sg13g2_tiehi _6187__173 (.L_HI(net173));
 sg13g2_tiehi _6127__174 (.L_HI(net174));
 sg13g2_tiehi _6222__175 (.L_HI(net175));
 sg13g2_tiehi _6126__176 (.L_HI(net176));
 sg13g2_tiehi _6186__177 (.L_HI(net177));
 sg13g2_tiehi _6125__178 (.L_HI(net178));
 sg13g2_tiehi _6212__179 (.L_HI(net179));
 sg13g2_tiehi _6124__180 (.L_HI(net180));
 sg13g2_tiehi _6185__181 (.L_HI(net181));
 sg13g2_tiehi _6123__182 (.L_HI(net182));
 sg13g2_tiehi _6230__183 (.L_HI(net183));
 sg13g2_tiehi _6122__184 (.L_HI(net184));
 sg13g2_tiehi _6184__185 (.L_HI(net185));
 sg13g2_tiehi _6121__186 (.L_HI(net186));
 sg13g2_tiehi _6211__187 (.L_HI(net187));
 sg13g2_tiehi _6120__188 (.L_HI(net188));
 sg13g2_tiehi _6183__189 (.L_HI(net189));
 sg13g2_tiehi _6119__190 (.L_HI(net190));
 sg13g2_tiehi _6221__191 (.L_HI(net191));
 sg13g2_tiehi _6118__192 (.L_HI(net192));
 sg13g2_tiehi _6182__193 (.L_HI(net193));
 sg13g2_tiehi _6117__194 (.L_HI(net194));
 sg13g2_tiehi _6210__195 (.L_HI(net195));
 sg13g2_tiehi _6116__196 (.L_HI(net196));
 sg13g2_tiehi _6181__197 (.L_HI(net197));
 sg13g2_tiehi _6115__198 (.L_HI(net198));
 sg13g2_tiehi _6226__199 (.L_HI(net199));
 sg13g2_tiehi _6114__200 (.L_HI(net200));
 sg13g2_tiehi _6180__201 (.L_HI(net201));
 sg13g2_tiehi _6113__202 (.L_HI(net202));
 sg13g2_tiehi _6209__203 (.L_HI(net203));
 sg13g2_tiehi _6112__204 (.L_HI(net204));
 sg13g2_tiehi _6179__205 (.L_HI(net205));
 sg13g2_tiehi _6111__206 (.L_HI(net206));
 sg13g2_tiehi _6220__207 (.L_HI(net207));
 sg13g2_tiehi _6110__208 (.L_HI(net208));
 sg13g2_tiehi _6109__209 (.L_HI(net209));
 sg13g2_tiehi _6105__210 (.L_HI(net210));
 sg13g2_tiehi _6104__211 (.L_HI(net211));
 sg13g2_tiehi _6103__212 (.L_HI(net212));
 sg13g2_tiehi _6102__213 (.L_HI(net213));
 sg13g2_tiehi _6101__214 (.L_HI(net214));
 sg13g2_tiehi _6100__215 (.L_HI(net215));
 sg13g2_tiehi _6178__216 (.L_HI(net216));
 sg13g2_tiehi _6099__217 (.L_HI(net217));
 sg13g2_tiehi _6177__218 (.L_HI(net218));
 sg13g2_tiehi _6098__219 (.L_HI(net219));
 sg13g2_tiehi _6176__220 (.L_HI(net220));
 sg13g2_tiehi _6097__221 (.L_HI(net221));
 sg13g2_tiehi _6175__222 (.L_HI(net222));
 sg13g2_tiehi _6096__223 (.L_HI(net223));
 sg13g2_tiehi _6174__224 (.L_HI(net224));
 sg13g2_tiehi _6095__225 (.L_HI(net225));
 sg13g2_tiehi _6173__226 (.L_HI(net226));
 sg13g2_tiehi _6094__227 (.L_HI(net227));
 sg13g2_tiehi _6172__228 (.L_HI(net228));
 sg13g2_tiehi _6093__229 (.L_HI(net229));
 sg13g2_tiehi _6171__230 (.L_HI(net230));
 sg13g2_tiehi tt_um_htfab_bouncy_capsule_231 (.L_HI(net231));
 sg13g2_tiehi tt_um_htfab_bouncy_capsule_232 (.L_HI(net232));
 sg13g2_tiehi tt_um_htfab_bouncy_capsule_233 (.L_HI(net233));
 sg13g2_tiehi tt_um_htfab_bouncy_capsule_234 (.L_HI(net234));
 sg13g2_tiehi tt_um_htfab_bouncy_capsule_235 (.L_HI(net235));
 sg13g2_tiehi tt_um_htfab_bouncy_capsule_236 (.L_HI(net236));
 sg13g2_tiehi tt_um_htfab_bouncy_capsule_237 (.L_HI(net237));
 sg13g2_tiehi tt_um_htfab_bouncy_capsule_238 (.L_HI(net238));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_2 _6461_ (.A(pdm_out),
    .X(uio_out[0]));
 sg13g2_buf_2 _6462_ (.A(pdm_out),
    .X(uio_out[1]));
 sg13g2_buf_2 _6463_ (.A(pdm_out),
    .X(uio_out[2]));
 sg13g2_buf_2 _6464_ (.A(pdm_out),
    .X(uio_out[3]));
 sg13g2_buf_2 _6465_ (.A(pdm_out),
    .X(uio_out[4]));
 sg13g2_buf_2 _6466_ (.A(pdm_out),
    .X(uio_out[5]));
 sg13g2_buf_2 _6467_ (.A(pdm_out),
    .X(uio_out[6]));
 sg13g2_buf_2 _6468_ (.A(pdm_out),
    .X(uio_out[7]));
 sg13g2_buf_1 _6469_ (.A(\i_vga_beam.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _6470_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout813 (.A(_2201_),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(net815),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(_0375_),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(net817),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(_0374_),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(net819),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(_0526_),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(net821),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_0526_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(_0526_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(net825),
    .X(net823));
 sg13g2_buf_1 fanout824 (.A(net825),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(_0525_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_0373_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_2778_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_0534_),
    .X(net828));
 sg13g2_buf_4 fanout829 (.X(net829),
    .A(_0524_));
 sg13g2_buf_2 fanout830 (.A(net831),
    .X(net830));
 sg13g2_buf_4 fanout831 (.X(net831),
    .A(_0505_));
 sg13g2_buf_2 fanout832 (.A(net833),
    .X(net832));
 sg13g2_buf_4 fanout833 (.X(net833),
    .A(_0504_));
 sg13g2_buf_1 fanout834 (.A(_0504_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(net836),
    .X(net835));
 sg13g2_buf_4 fanout836 (.X(net836),
    .A(_0471_));
 sg13g2_buf_2 fanout837 (.A(net838),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_0395_),
    .X(net838));
 sg13g2_buf_4 fanout839 (.X(net839),
    .A(_0395_));
 sg13g2_buf_2 fanout840 (.A(_0395_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(net842),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(net846),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(net846),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(net846),
    .X(net844));
 sg13g2_buf_4 fanout845 (.X(net845),
    .A(net846));
 sg13g2_buf_2 fanout846 (.A(_0394_),
    .X(net846));
 sg13g2_buf_4 fanout847 (.X(net847),
    .A(_0393_));
 sg13g2_buf_4 fanout848 (.X(net848),
    .A(_0483_));
 sg13g2_buf_2 fanout849 (.A(net858),
    .X(net849));
 sg13g2_buf_1 fanout850 (.A(net858),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(net852),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(net858),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(net857),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(net856),
    .X(net854));
 sg13g2_buf_1 fanout855 (.A(net856),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(net857),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(net858),
    .X(net857));
 sg13g2_buf_1 fanout858 (.A(_0472_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_0469_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(net864),
    .X(net860));
 sg13g2_buf_4 fanout861 (.X(net861),
    .A(net862));
 sg13g2_buf_2 fanout862 (.A(net864),
    .X(net862));
 sg13g2_buf_4 fanout863 (.X(net863),
    .A(net864));
 sg13g2_buf_2 fanout864 (.A(_0450_),
    .X(net864));
 sg13g2_buf_4 fanout865 (.X(net865),
    .A(net866));
 sg13g2_buf_4 fanout866 (.X(net866),
    .A(_0449_));
 sg13g2_buf_4 fanout867 (.X(net867),
    .A(_0411_));
 sg13g2_buf_4 fanout868 (.X(net868),
    .A(_1106_));
 sg13g2_buf_2 fanout869 (.A(net870),
    .X(net869));
 sg13g2_buf_1 fanout870 (.A(net871),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_1834_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_2035_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_2033_),
    .X(net873));
 sg13g2_buf_4 fanout874 (.X(net874),
    .A(_2648_));
 sg13g2_buf_4 fanout875 (.X(net875),
    .A(net876));
 sg13g2_buf_2 fanout876 (.A(_2648_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(net878),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(net879),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(net881),
    .X(net879));
 sg13g2_buf_4 fanout880 (.X(net880),
    .A(net881));
 sg13g2_buf_2 fanout881 (.A(_2647_),
    .X(net881));
 sg13g2_buf_4 fanout882 (.X(net882),
    .A(_0859_));
 sg13g2_buf_4 fanout883 (.X(net883),
    .A(_0857_));
 sg13g2_buf_4 fanout884 (.X(net884),
    .A(net885));
 sg13g2_buf_4 fanout885 (.X(net885),
    .A(_0342_));
 sg13g2_buf_2 fanout886 (.A(net888),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(net888),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(net890),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(net890),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_2758_),
    .X(net890));
 sg13g2_buf_4 fanout891 (.X(net891),
    .A(net893));
 sg13g2_buf_2 fanout892 (.A(net893),
    .X(net892));
 sg13g2_buf_4 fanout893 (.X(net893),
    .A(_2757_));
 sg13g2_buf_4 fanout894 (.X(net894),
    .A(net895));
 sg13g2_buf_2 fanout895 (.A(_2696_),
    .X(net895));
 sg13g2_buf_4 fanout896 (.X(net896),
    .A(net897));
 sg13g2_buf_4 fanout897 (.X(net897),
    .A(_2774_));
 sg13g2_buf_4 fanout898 (.X(net898),
    .A(_2569_));
 sg13g2_buf_4 fanout899 (.X(net899),
    .A(_2566_));
 sg13g2_buf_2 fanout900 (.A(net901),
    .X(net900));
 sg13g2_buf_4 fanout901 (.X(net901),
    .A(net902));
 sg13g2_buf_4 fanout902 (.X(net902),
    .A(_2681_));
 sg13g2_buf_2 fanout903 (.A(net904),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(net905),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(_2680_),
    .X(net905));
 sg13g2_buf_4 fanout906 (.X(net906),
    .A(_2680_));
 sg13g2_buf_4 fanout907 (.X(net907),
    .A(_1000_));
 sg13g2_buf_2 fanout908 (.A(_1000_),
    .X(net908));
 sg13g2_buf_4 fanout909 (.X(net909),
    .A(_2530_));
 sg13g2_buf_2 fanout910 (.A(_2041_),
    .X(net910));
 sg13g2_buf_1 fanout911 (.A(_2041_),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(net913),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(_1272_),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(_1272_),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_1032_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_1027_),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(net919),
    .X(net917));
 sg13g2_buf_1 fanout918 (.A(net919),
    .X(net918));
 sg13g2_buf_1 fanout919 (.A(net920),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_2600_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_1525_),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(_1499_),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(_1499_),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(_1498_),
    .X(net924));
 sg13g2_buf_1 fanout925 (.A(_1498_),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(net927),
    .X(net926));
 sg13g2_buf_1 fanout927 (.A(net928),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(_2598_),
    .X(net928));
 sg13g2_buf_4 fanout929 (.X(net929),
    .A(_2092_));
 sg13g2_buf_2 fanout930 (.A(net931),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(net933),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(net933),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(_2091_),
    .X(net933));
 sg13g2_buf_4 fanout934 (.X(net934),
    .A(_2030_));
 sg13g2_buf_4 fanout935 (.X(net935),
    .A(net936));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(_2698_));
 sg13g2_buf_4 fanout937 (.X(net937),
    .A(_2698_));
 sg13g2_buf_4 fanout938 (.X(net938),
    .A(net939));
 sg13g2_buf_2 fanout939 (.A(_2697_),
    .X(net939));
 sg13g2_buf_4 fanout940 (.X(net940),
    .A(net941));
 sg13g2_buf_2 fanout941 (.A(net944),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(net943),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(net944),
    .X(net943));
 sg13g2_buf_4 fanout944 (.X(net944),
    .A(_2697_));
 sg13g2_buf_4 fanout945 (.X(net945),
    .A(_2029_));
 sg13g2_buf_2 fanout946 (.A(net947),
    .X(net946));
 sg13g2_buf_4 fanout947 (.X(net947),
    .A(_1628_));
 sg13g2_buf_4 fanout948 (.X(net948),
    .A(_1628_));
 sg13g2_buf_2 fanout949 (.A(_1510_),
    .X(net949));
 sg13g2_buf_4 fanout950 (.X(net950),
    .A(_1495_));
 sg13g2_buf_2 fanout951 (.A(_1495_),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(net953),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_1494_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_2492_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(_2489_),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_2488_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_2487_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(net959),
    .X(net958));
 sg13g2_buf_1 fanout959 (.A(_2486_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(net961),
    .X(net960));
 sg13g2_buf_1 fanout961 (.A(_2485_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(net963),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_2484_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(net965),
    .X(net964));
 sg13g2_buf_1 fanout965 (.A(_2481_),
    .X(net965));
 sg13g2_buf_4 fanout966 (.X(net966),
    .A(net967));
 sg13g2_buf_2 fanout967 (.A(_2478_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_2478_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_2478_),
    .X(net969));
 sg13g2_buf_4 fanout970 (.X(net970),
    .A(net971));
 sg13g2_buf_4 fanout971 (.X(net971),
    .A(_2477_));
 sg13g2_buf_4 fanout972 (.X(net972),
    .A(net975));
 sg13g2_buf_2 fanout973 (.A(net975),
    .X(net973));
 sg13g2_buf_4 fanout974 (.X(net974),
    .A(net975));
 sg13g2_buf_4 fanout975 (.X(net975),
    .A(_2477_));
 sg13g2_buf_4 fanout976 (.X(net976),
    .A(net979));
 sg13g2_buf_4 fanout977 (.X(net977),
    .A(net979));
 sg13g2_buf_1 fanout978 (.A(net979),
    .X(net978));
 sg13g2_buf_4 fanout979 (.X(net979),
    .A(net982));
 sg13g2_buf_2 fanout980 (.A(net982),
    .X(net980));
 sg13g2_buf_4 fanout981 (.X(net981),
    .A(net982));
 sg13g2_buf_4 fanout982 (.X(net982),
    .A(_2476_));
 sg13g2_buf_4 fanout983 (.X(net983),
    .A(net984));
 sg13g2_buf_4 fanout984 (.X(net984),
    .A(_2475_));
 sg13g2_buf_4 fanout985 (.X(net985),
    .A(net988));
 sg13g2_buf_4 fanout986 (.X(net986),
    .A(net988));
 sg13g2_buf_1 fanout987 (.A(net988),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(net989),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(net990),
    .X(net989));
 sg13g2_buf_4 fanout990 (.X(net990),
    .A(_2475_));
 sg13g2_buf_2 fanout991 (.A(net992),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(net993),
    .X(net992));
 sg13g2_buf_4 fanout993 (.X(net993),
    .A(_2391_));
 sg13g2_buf_4 fanout994 (.X(net994),
    .A(_2375_));
 sg13g2_buf_2 fanout995 (.A(net997),
    .X(net995));
 sg13g2_buf_1 fanout996 (.A(net997),
    .X(net996));
 sg13g2_buf_4 fanout997 (.X(net997),
    .A(net512));
 sg13g2_buf_4 fanout998 (.X(net998),
    .A(\i_collision.i_coll_table.in[5] ));
 sg13g2_buf_2 fanout999 (.A(\i_collision.i_coll_table.in[5] ),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(net1001),
    .X(net1000));
 sg13g2_buf_1 fanout1001 (.A(net1002),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(net539),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(net1004),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(net1005),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(\i_collision.i_coll_table.in[4] ),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(net1008),
    .X(net1006));
 sg13g2_buf_1 fanout1007 (.A(net1008),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(\i_resonator.v[15] ),
    .X(net1008));
 sg13g2_buf_4 fanout1009 (.X(net1009),
    .A(\i_resonator.v[15] ));
 sg13g2_buf_4 fanout1010 (.X(net1010),
    .A(\i_resonator.v[15] ));
 sg13g2_buf_4 fanout1011 (.X(net1011),
    .A(net540));
 sg13g2_buf_4 fanout1012 (.X(net1012),
    .A(net542));
 sg13g2_buf_4 fanout1013 (.X(net1013),
    .A(net536));
 sg13g2_buf_2 fanout1014 (.A(\i_delta_sigma.sample[9] ),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(net1016),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(net1017),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(net1018),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(\i_delta_sigma.sample[11] ),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(net483),
    .X(net1019));
 sg13g2_buf_4 fanout1020 (.X(net1020),
    .A(net543));
 sg13g2_buf_4 fanout1021 (.X(net1021),
    .A(net1022));
 sg13g2_buf_2 fanout1022 (.A(\i_collision.i_coll_table.in[1] ),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(net1024),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(\i_collision.i_coll_table.in[1] ),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(net1026),
    .X(net1025));
 sg13g2_buf_1 fanout1026 (.A(net1027),
    .X(net1026));
 sg13g2_buf_4 fanout1027 (.X(net1027),
    .A(net544));
 sg13g2_buf_2 fanout1028 (.A(net1029),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(net1030),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(net522),
    .X(net1030));
 sg13g2_buf_4 fanout1031 (.X(net1031),
    .A(net549));
 sg13g2_buf_4 fanout1032 (.X(net1032),
    .A(net547));
 sg13g2_buf_2 fanout1033 (.A(net1034),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(net420),
    .X(net1034));
 sg13g2_buf_4 fanout1035 (.X(net1035),
    .A(\i_collision.rotate ));
 sg13g2_buf_1 fanout1036 (.A(\i_collision.rotate ),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(net1038),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_buf_1 fanout1039 (.A(net1042),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(net1042),
    .X(net1040));
 sg13g2_buf_1 fanout1041 (.A(net1042),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(\i_kinematics.update ),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(\i_kinematics.update ),
    .X(net1043));
 sg13g2_buf_1 fanout1044 (.A(net1045),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(\i_kinematics.update ),
    .X(net1045));
 sg13g2_buf_4 fanout1046 (.X(net1046),
    .A(net1048));
 sg13g2_buf_4 fanout1047 (.X(net1047),
    .A(net1048));
 sg13g2_buf_2 fanout1048 (.A(\i_orchestrator.update_resonator ),
    .X(net1048));
 sg13g2_buf_4 fanout1049 (.X(net1049),
    .A(net303));
 sg13g2_buf_1 fanout1050 (.A(\i_collision.i_coll_table.in[0] ),
    .X(net1050));
 sg13g2_buf_4 fanout1051 (.X(net1051),
    .A(\i_capsule.tf_y[9] ));
 sg13g2_buf_2 fanout1052 (.A(\i_orchestrator.vga_y[5] ),
    .X(net1052));
 sg13g2_buf_4 fanout1053 (.X(net1053),
    .A(\i_orchestrator.vga_y[4] ));
 sg13g2_buf_2 fanout1054 (.A(net446),
    .X(net1054));
 sg13g2_buf_4 fanout1055 (.X(net1055),
    .A(\i_orchestrator.vga_y[3] ));
 sg13g2_buf_2 fanout1056 (.A(net533),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(net1058),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(net541),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(net553),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(net337),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(net464),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(net491),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(_2028_),
    .X(net1063));
 sg13g2_buf_1 fanout1064 (.A(_2028_),
    .X(net1064));
 sg13g2_buf_4 fanout1065 (.X(net1065),
    .A(_1629_));
 sg13g2_buf_2 fanout1066 (.A(net1067),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_4 fanout1068 (.X(net1068),
    .A(net1069));
 sg13g2_buf_4 fanout1069 (.X(net1069),
    .A(_2431_));
 sg13g2_buf_4 fanout1070 (.X(net1070),
    .A(_2431_));
 sg13g2_buf_4 fanout1071 (.X(net1071),
    .A(net1073));
 sg13g2_buf_2 fanout1072 (.A(net1073),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(rst_n),
    .X(net1073));
 sg13g2_buf_4 fanout1074 (.X(net1074),
    .A(net1078));
 sg13g2_buf_2 fanout1075 (.A(net1076),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(net1077),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(net1078),
    .X(net1077));
 sg13g2_buf_4 fanout1078 (.X(net1078),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[2]));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tiehi _6092__9 (.L_HI(net9));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_0_clk));
 sg13g2_inv_8 clkload6 (.A(clknet_leaf_33_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_34_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_1_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_2_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_3_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_24_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_27_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_28_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_23_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_4_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_7_clk));
 sg13g2_inv_8 clkload17 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_6_clk));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_10_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_17_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_11_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0071_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0072_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0115_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold4 (.A(\i_orchestrator.sample_counter[9] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0132_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0074_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0010_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0137_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0005_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0238_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0073_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold12 (.A(_1126_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold13 (.A(\i_kinematics.phi[0] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_kinematics.center_y_lo[0] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0178_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold16 (.A(\i_kinematics.center_x_lo[0] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0180_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold18 (.A(\collision_impact[0] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0168_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_orchestrator.tension[2] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold21 (.A(_2310_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold22 (.A(\i_orchestrator.tension[3] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0240_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold24 (.A(\collision_impact[1] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0169_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold26 (.A(\i_transform.track_x[3] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0226_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold28 (.A(\i_orchestrator.lfsr[3] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0121_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i_orchestrator.lfsr[5] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0122_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_orchestrator.lfsr[2] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold33 (.A(\i_orchestrator.lfsr[1] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold34 (.A(\i_orchestrator.sample_counter[3] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0231_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold36 (.A(\i_orchestrator.sample_counter[7] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold37 (.A(_1922_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0235_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold39 (.A(\i_orchestrator.tension[1] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold40 (.A(_2306_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold41 (.A(\i_orchestrator.lfsr[7] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0124_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold43 (.A(\i_orchestrator.sample_counter[8] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0236_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0004_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold46 (.A(_1308_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold47 (.A(\i_transform.image_x[0] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0218_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0066_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0247_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0069_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold52 (.A(_2037_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0282_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold54 (.A(\i_orchestrator.lfsr[6] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold55 (.A(\i_transform.track_y[9] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold56 (.A(_1486_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold57 (.A(\color_entropy[0] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold58 (.A(\center_y[9] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold59 (.A(\i_transform.track_y[3] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0101_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold61 (.A(\i_transform.track_x[9] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold62 (.A(_1986_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold63 (.A(\i_orchestrator.sample_counter[2] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold64 (.A(_1912_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold65 (.A(\i_collision.i_coll_table.in[0] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold66 (.A(\center_x[9] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold67 (.A(\i_kinematics.phi[1] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold68 (.A(\color_entropy[1] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold69 (.A(\i_orchestrator.vga_x[6] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold70 (.A(_1006_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold71 (.A(\i_transform.track_y[0] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0098_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold73 (.A(\i_transform.image_y[0] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0213_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold75 (.A(\i_transform.image_y[4] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold76 (.A(\i_transform.track_y[4] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold77 (.A(_1169_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0102_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold79 (.A(\center_y[2] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0100_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold81 (.A(\i_orchestrator.sample_counter[6] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_transform.image_y[3] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold83 (.A(\i_transform.image_x[1] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold84 (.A(\i_orchestrator.hit_right ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold85 (.A(_1932_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0239_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold87 (.A(\i_orchestrator.vga_y[3] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold88 (.A(\i_orchestrator.vga_x[0] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold89 (.A(_1001_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0076_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold91 (.A(\capsule_color[0] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0241_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold93 (.A(\i_resonator.v[0] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0266_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold95 (.A(\i_kinematics.phi[2] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold96 (.A(\i_orchestrator.sample_counter[5] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold97 (.A(_1920_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold98 (.A(\i_transform.image_y[1] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_orchestrator.vga_x[9] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold100 (.A(\i_orchestrator.hit_bottom ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0043_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold102 (.A(_1954_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0245_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold104 (.A(\i_transform.image_x[3] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold105 (.A(_1885_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold106 (.A(\i_transform.image_x[5] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0152_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold108 (.A(\i_orchestrator.vga_x[2] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold109 (.A(_1002_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold110 (.A(\i_orchestrator.hit_priority[1] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold111 (.A(_1275_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0116_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold113 (.A(\i_transform.track_x[0] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0223_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0011_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold116 (.A(_1320_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold117 (.A(_1321_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_delta_sigma.sample[0] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0254_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold120 (.A(\i_colors.capsule_color[5] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0246_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold122 (.A(\i_kinematics.center_x_lo[1] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0181_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold124 (.A(\i_kinematics.center_y_lo[1] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0179_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0054_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold127 (.A(\i_orchestrator.hit_left ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold128 (.A(\i_delta_sigma.acc[4] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold129 (.A(_1340_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0142_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold131 (.A(\i_kinematics.phi[10] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold132 (.A(\i_transform.track_y[5] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0163_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold134 (.A(\i_collision.vy[0] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold135 (.A(\i_orchestrator.sample_counter[0] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold136 (.A(_1310_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0229_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold138 (.A(\i_orchestrator.sample_counter[4] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold139 (.A(\i_transform.image_y[2] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold140 (.A(\i_delta_sigma.acc[8] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold141 (.A(_1358_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0146_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold143 (.A(\i_orchestrator.hit_top ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold144 (.A(\i_orchestrator.vga_y[9] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold145 (.A(_1149_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0097_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold147 (.A(\i_collision.vx[0] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0175_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold149 (.A(\center_y[2] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold150 (.A(\i_resonator.counter[3] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_transform.image_x[4] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold152 (.A(\center_y[8] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold153 (.A(orient),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0086_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold155 (.A(\i_colors.capsule_color[4] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold156 (.A(_1990_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0252_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold158 (.A(\i_transform.track_y[8] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0166_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold160 (.A(\i_resonator.v[4] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold161 (.A(\i_orchestrator.vga_y[7] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold162 (.A(_1145_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold163 (.A(\i_transform.track_x[4] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0227_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold165 (.A(\i_resonator.v[1] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold166 (.A(_2171_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold167 (.A(\i_resonator.v[6] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold168 (.A(\center_y[3] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold169 (.A(\i_bitmap.in[3] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold170 (.A(_1412_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold171 (.A(\i_delta_sigma.acc[3] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold172 (.A(_1335_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0141_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold174 (.A(\i_transform.image_y[5] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold175 (.A(\capsule_color[1] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold176 (.A(_1944_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold177 (.A(bitmap_pixel),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0287_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold179 (.A(\i_orchestrator.vga_x[8] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold180 (.A(_1009_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0083_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold182 (.A(\i_collision.update ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold183 (.A(\i_resonator.v[3] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold184 (.A(\i_resonator.v[2] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold185 (.A(\i_colors.channel[1] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0002_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold187 (.A(\capsule_color[3] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold188 (.A(\i_orchestrator.trigger_debounce ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0114_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold190 (.A(\i_orchestrator.vga_y[6] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0094_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold192 (.A(\i_resonator.v[5] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold193 (.A(\i_bitmap.in[11] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold194 (.A(\i_colors.channel[0] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0003_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold196 (.A(\i_delta_sigma.acc[0] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold197 (.A(\center_x[2] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold198 (.A(\i_transform.image_x[2] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold199 (.A(\center_y[1] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold200 (.A(\i_delta_sigma.sample[2] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold201 (.A(_2051_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold202 (.A(\i_bitmap.in[6] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold203 (.A(\center_x[4] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0196_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold205 (.A(\center_x[5] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0197_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold207 (.A(\i_transform.track_y[1] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold208 (.A(\i_orchestrator.vga_y[4] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold209 (.A(\center_y[7] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0189_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold211 (.A(\i_colors.channel[2] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold212 (.A(handle_impact),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold213 (.A(\center_y[6] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0188_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold215 (.A(\i_transform.track_x[2] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold216 (.A(_1903_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold217 (.A(\i_transform.track_x[7] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold218 (.A(_1975_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold219 (.A(\i_resonator.v[7] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold220 (.A(\i_kinematics.phi[6] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold221 (.A(\center_y[0] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold222 (.A(\i_bitmap.in[5] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold223 (.A(\center_y[4] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0186_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold225 (.A(\i_orchestrator.vga_x[3] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold226 (.A(\i_orchestrator.vga_x[7] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold227 (.A(\center_y[5] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold228 (.A(\i_resonator.v[9] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold229 (.A(\i_transform.track_x[8] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold230 (.A(_1980_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold231 (.A(\center_x[8] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold232 (.A(\i_orchestrator.vga_y[8] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold233 (.A(\i_transform.track_x[1] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0224_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold235 (.A(\i_delta_sigma.acc[9] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold236 (.A(_1363_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold237 (.A(\i_delta_sigma.acc[1] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold238 (.A(\i_orchestrator.hit_priority[0] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold239 (.A(\center_x[6] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0198_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold241 (.A(\center_x[7] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0199_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold243 (.A(\i_orchestrator.vga_y[0] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold244 (.A(\i_bitmap.in[10] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold245 (.A(\capsule_color[2] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold246 (.A(\i_transform.track_y[6] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0164_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold248 (.A(\i_orchestrator.trigger_resonator[0] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold249 (.A(_2063_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold250 (.A(\i_delta_sigma.sample[3] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold251 (.A(\i_transform.track_y[7] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold252 (.A(\i_delta_sigma.sample[1] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold253 (.A(\i_orchestrator.vga_x[5] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold254 (.A(\i_kinematics.phi[7] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold255 (.A(\i_bitmap.in[4] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold256 (.A(\i_kinematics.phi[5] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold257 (.A(\i_orchestrator.vga_x[4] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold258 (.A(\i_delta_sigma.acc[5] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold259 (.A(\center_x[0] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold260 (.A(\i_capsule.tf_y[8] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold261 (.A(\i_collision.vx[1] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0176_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold263 (.A(\i_capsule.tf_y[7] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold264 (.A(\i_bitmap.in[2] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold265 (.A(\i_bitmap.in[12] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold266 (.A(\i_bitmap.in[0] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold267 (.A(\i_delta_sigma.acc[7] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold268 (.A(_1355_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0145_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold270 (.A(\center_x[3] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0195_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold272 (.A(\i_orchestrator.trigger_resonator[1] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold273 (.A(_2059_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold274 (.A(\i_collision.i_coll_table.in[3] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0290_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold276 (.A(\i_kinematics.phi[4] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold277 (.A(\i_delta_sigma.sample[7] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold278 (.A(\i_collision.vy[1] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold279 (.A(\i_resonator.v[8] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold280 (.A(\i_kinematics.phi[3] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold281 (.A(\i_orchestrator.trigger_resonator[1] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold282 (.A(\i_delta_sigma.acc[6] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold283 (.A(\center_x[1] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold284 (.A(\i_collision.vy[2] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0174_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold286 (.A(\i_delta_sigma.acc[13] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold287 (.A(\i_transform.track_x[6] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0248_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold289 (.A(\i_bitmap.in[8] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold290 (.A(\i_delta_sigma.sample[8] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold291 (.A(\i_bitmap.in[9] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold292 (.A(\i_delta_sigma.acc[2] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold293 (.A(\i_delta_sigma.acc[10] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold294 (.A(\i_capsule.tf_x[8] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold295 (.A(\i_orchestrator.vga_y[2] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold296 (.A(\i_delta_sigma.sample[6] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold297 (.A(\i_orchestrator.update_transform ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold298 (.A(\i_delta_sigma.sample[10] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold299 (.A(\i_resonator.v[11] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold300 (.A(\i_orchestrator.vga_x[4] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold301 (.A(\i_collision.i_coll_table.in[5] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold302 (.A(\i_resonator.v[13] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold303 (.A(\i_orchestrator.vga_y[1] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold304 (.A(\i_resonator.v[10] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold305 (.A(\i_collision.phi[1] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold306 (.A(\i_collision.vx[2] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0177_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold308 (.A(\i_resonator.v[12] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold309 (.A(\i_bitmap.in[1] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold310 (.A(\i_bitmap.in[7] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold311 (.A(\i_capsule.tf_x[9] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold312 (.A(\i_resonator.v[14] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold313 (.A(\i_capsule.tf_x[0] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold314 (.A(\i_delta_sigma.sample[1] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold315 (.A(\i_orchestrator.vga_y[0] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold316 (.A(\i_orchestrator.vga_x[3] ),
    .X(net554));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_fill_1 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_89 ();
 sg13g2_decap_8 FILLER_0_96 ();
 sg13g2_decap_8 FILLER_0_103 ();
 sg13g2_decap_8 FILLER_0_110 ();
 sg13g2_decap_8 FILLER_0_117 ();
 sg13g2_decap_8 FILLER_0_124 ();
 sg13g2_fill_2 FILLER_0_131 ();
 sg13g2_fill_1 FILLER_0_133 ();
 sg13g2_decap_4 FILLER_0_186 ();
 sg13g2_fill_1 FILLER_0_190 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_fill_2 FILLER_0_208 ();
 sg13g2_decap_8 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_221 ();
 sg13g2_decap_8 FILLER_0_228 ();
 sg13g2_decap_8 FILLER_0_235 ();
 sg13g2_decap_4 FILLER_0_242 ();
 sg13g2_decap_4 FILLER_0_250 ();
 sg13g2_fill_2 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_260 ();
 sg13g2_decap_8 FILLER_0_267 ();
 sg13g2_decap_8 FILLER_0_274 ();
 sg13g2_decap_8 FILLER_0_281 ();
 sg13g2_decap_8 FILLER_0_288 ();
 sg13g2_decap_8 FILLER_0_295 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_309 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_4 FILLER_1_96 ();
 sg13g2_fill_1 FILLER_1_116 ();
 sg13g2_fill_2 FILLER_1_186 ();
 sg13g2_fill_1 FILLER_1_198 ();
 sg13g2_fill_2 FILLER_1_229 ();
 sg13g2_fill_1 FILLER_1_231 ();
 sg13g2_fill_1 FILLER_1_251 ();
 sg13g2_fill_2 FILLER_1_258 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_fill_2 FILLER_2_70 ();
 sg13g2_fill_1 FILLER_2_142 ();
 sg13g2_fill_2 FILLER_2_148 ();
 sg13g2_fill_1 FILLER_2_219 ();
 sg13g2_fill_2 FILLER_2_245 ();
 sg13g2_fill_1 FILLER_2_247 ();
 sg13g2_fill_2 FILLER_2_254 ();
 sg13g2_fill_2 FILLER_2_264 ();
 sg13g2_fill_2 FILLER_2_276 ();
 sg13g2_decap_8 FILLER_2_288 ();
 sg13g2_decap_8 FILLER_2_295 ();
 sg13g2_decap_8 FILLER_2_302 ();
 sg13g2_decap_8 FILLER_2_309 ();
 sg13g2_decap_8 FILLER_2_316 ();
 sg13g2_decap_8 FILLER_2_323 ();
 sg13g2_decap_8 FILLER_2_330 ();
 sg13g2_decap_8 FILLER_2_337 ();
 sg13g2_decap_8 FILLER_2_344 ();
 sg13g2_decap_8 FILLER_2_351 ();
 sg13g2_decap_8 FILLER_2_358 ();
 sg13g2_decap_8 FILLER_2_365 ();
 sg13g2_decap_8 FILLER_2_372 ();
 sg13g2_decap_8 FILLER_2_379 ();
 sg13g2_decap_8 FILLER_2_386 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_4 FILLER_3_42 ();
 sg13g2_fill_1 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_fill_1 FILLER_3_63 ();
 sg13g2_fill_1 FILLER_3_109 ();
 sg13g2_fill_1 FILLER_3_153 ();
 sg13g2_fill_2 FILLER_3_174 ();
 sg13g2_fill_1 FILLER_3_176 ();
 sg13g2_fill_1 FILLER_3_210 ();
 sg13g2_fill_1 FILLER_3_226 ();
 sg13g2_fill_1 FILLER_3_265 ();
 sg13g2_decap_8 FILLER_3_295 ();
 sg13g2_decap_8 FILLER_3_302 ();
 sg13g2_decap_8 FILLER_3_309 ();
 sg13g2_decap_8 FILLER_3_316 ();
 sg13g2_decap_8 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_330 ();
 sg13g2_decap_8 FILLER_3_337 ();
 sg13g2_decap_8 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_351 ();
 sg13g2_decap_8 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_fill_2 FILLER_4_14 ();
 sg13g2_fill_1 FILLER_4_16 ();
 sg13g2_fill_2 FILLER_4_69 ();
 sg13g2_fill_1 FILLER_4_71 ();
 sg13g2_fill_2 FILLER_4_87 ();
 sg13g2_fill_1 FILLER_4_89 ();
 sg13g2_fill_2 FILLER_4_95 ();
 sg13g2_fill_1 FILLER_4_97 ();
 sg13g2_fill_2 FILLER_4_108 ();
 sg13g2_fill_1 FILLER_4_150 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_4 FILLER_4_217 ();
 sg13g2_fill_1 FILLER_4_221 ();
 sg13g2_fill_1 FILLER_4_260 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_4 FILLER_5_14 ();
 sg13g2_fill_2 FILLER_5_18 ();
 sg13g2_fill_1 FILLER_5_33 ();
 sg13g2_fill_1 FILLER_5_39 ();
 sg13g2_fill_1 FILLER_5_89 ();
 sg13g2_fill_2 FILLER_5_95 ();
 sg13g2_fill_1 FILLER_5_97 ();
 sg13g2_fill_2 FILLER_5_107 ();
 sg13g2_fill_1 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_fill_1 FILLER_5_157 ();
 sg13g2_fill_1 FILLER_5_173 ();
 sg13g2_fill_2 FILLER_5_182 ();
 sg13g2_fill_1 FILLER_5_184 ();
 sg13g2_decap_4 FILLER_5_190 ();
 sg13g2_fill_1 FILLER_5_194 ();
 sg13g2_decap_8 FILLER_5_198 ();
 sg13g2_decap_8 FILLER_5_205 ();
 sg13g2_decap_4 FILLER_5_212 ();
 sg13g2_fill_1 FILLER_5_216 ();
 sg13g2_fill_1 FILLER_5_222 ();
 sg13g2_fill_1 FILLER_5_236 ();
 sg13g2_decap_4 FILLER_5_254 ();
 sg13g2_fill_2 FILLER_5_267 ();
 sg13g2_fill_1 FILLER_5_269 ();
 sg13g2_decap_8 FILLER_5_285 ();
 sg13g2_decap_8 FILLER_5_292 ();
 sg13g2_decap_8 FILLER_5_299 ();
 sg13g2_decap_8 FILLER_5_306 ();
 sg13g2_decap_8 FILLER_5_313 ();
 sg13g2_decap_8 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_327 ();
 sg13g2_decap_8 FILLER_5_334 ();
 sg13g2_decap_8 FILLER_5_341 ();
 sg13g2_decap_8 FILLER_5_348 ();
 sg13g2_decap_8 FILLER_5_355 ();
 sg13g2_decap_8 FILLER_5_362 ();
 sg13g2_decap_8 FILLER_5_369 ();
 sg13g2_decap_8 FILLER_5_376 ();
 sg13g2_decap_8 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_390 ();
 sg13g2_decap_8 FILLER_5_397 ();
 sg13g2_decap_4 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_fill_2 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_28 ();
 sg13g2_fill_1 FILLER_6_34 ();
 sg13g2_fill_1 FILLER_6_57 ();
 sg13g2_fill_2 FILLER_6_83 ();
 sg13g2_fill_2 FILLER_6_94 ();
 sg13g2_fill_2 FILLER_6_106 ();
 sg13g2_fill_1 FILLER_6_108 ();
 sg13g2_decap_4 FILLER_6_142 ();
 sg13g2_fill_1 FILLER_6_146 ();
 sg13g2_decap_8 FILLER_6_170 ();
 sg13g2_decap_8 FILLER_6_177 ();
 sg13g2_decap_8 FILLER_6_184 ();
 sg13g2_decap_8 FILLER_6_191 ();
 sg13g2_decap_8 FILLER_6_198 ();
 sg13g2_fill_2 FILLER_6_205 ();
 sg13g2_fill_1 FILLER_6_207 ();
 sg13g2_decap_4 FILLER_6_213 ();
 sg13g2_decap_8 FILLER_6_230 ();
 sg13g2_fill_1 FILLER_6_237 ();
 sg13g2_fill_1 FILLER_6_242 ();
 sg13g2_decap_8 FILLER_6_283 ();
 sg13g2_decap_8 FILLER_6_290 ();
 sg13g2_decap_8 FILLER_6_297 ();
 sg13g2_decap_8 FILLER_6_304 ();
 sg13g2_decap_8 FILLER_6_311 ();
 sg13g2_decap_8 FILLER_6_318 ();
 sg13g2_decap_8 FILLER_6_325 ();
 sg13g2_decap_8 FILLER_6_332 ();
 sg13g2_decap_8 FILLER_6_339 ();
 sg13g2_decap_8 FILLER_6_346 ();
 sg13g2_decap_8 FILLER_6_353 ();
 sg13g2_decap_8 FILLER_6_360 ();
 sg13g2_decap_8 FILLER_6_367 ();
 sg13g2_decap_8 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_381 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_decap_8 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_4 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_11 ();
 sg13g2_fill_2 FILLER_7_42 ();
 sg13g2_fill_2 FILLER_7_49 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_73 ();
 sg13g2_fill_1 FILLER_7_80 ();
 sg13g2_fill_1 FILLER_7_85 ();
 sg13g2_fill_2 FILLER_7_142 ();
 sg13g2_decap_8 FILLER_7_170 ();
 sg13g2_fill_2 FILLER_7_177 ();
 sg13g2_fill_1 FILLER_7_179 ();
 sg13g2_fill_2 FILLER_7_185 ();
 sg13g2_fill_1 FILLER_7_223 ();
 sg13g2_fill_2 FILLER_7_233 ();
 sg13g2_fill_1 FILLER_7_247 ();
 sg13g2_decap_8 FILLER_7_291 ();
 sg13g2_decap_8 FILLER_7_298 ();
 sg13g2_decap_8 FILLER_7_305 ();
 sg13g2_decap_8 FILLER_7_312 ();
 sg13g2_decap_8 FILLER_7_319 ();
 sg13g2_decap_8 FILLER_7_326 ();
 sg13g2_decap_8 FILLER_7_333 ();
 sg13g2_decap_8 FILLER_7_340 ();
 sg13g2_decap_8 FILLER_7_347 ();
 sg13g2_decap_8 FILLER_7_354 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_fill_2 FILLER_8_26 ();
 sg13g2_fill_1 FILLER_8_48 ();
 sg13g2_fill_2 FILLER_8_74 ();
 sg13g2_fill_1 FILLER_8_76 ();
 sg13g2_fill_2 FILLER_8_104 ();
 sg13g2_fill_1 FILLER_8_106 ();
 sg13g2_fill_2 FILLER_8_113 ();
 sg13g2_fill_2 FILLER_8_133 ();
 sg13g2_fill_2 FILLER_8_164 ();
 sg13g2_fill_1 FILLER_8_166 ();
 sg13g2_decap_4 FILLER_8_187 ();
 sg13g2_fill_1 FILLER_8_196 ();
 sg13g2_fill_1 FILLER_8_209 ();
 sg13g2_decap_4 FILLER_8_213 ();
 sg13g2_decap_4 FILLER_8_233 ();
 sg13g2_fill_1 FILLER_8_237 ();
 sg13g2_fill_2 FILLER_8_267 ();
 sg13g2_fill_1 FILLER_8_269 ();
 sg13g2_decap_8 FILLER_8_275 ();
 sg13g2_decap_8 FILLER_8_282 ();
 sg13g2_fill_1 FILLER_8_289 ();
 sg13g2_decap_8 FILLER_8_295 ();
 sg13g2_decap_8 FILLER_8_302 ();
 sg13g2_decap_8 FILLER_8_309 ();
 sg13g2_decap_8 FILLER_8_316 ();
 sg13g2_decap_8 FILLER_8_323 ();
 sg13g2_decap_8 FILLER_8_330 ();
 sg13g2_decap_8 FILLER_8_337 ();
 sg13g2_decap_8 FILLER_8_344 ();
 sg13g2_decap_8 FILLER_8_351 ();
 sg13g2_decap_8 FILLER_8_358 ();
 sg13g2_decap_8 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_35 ();
 sg13g2_fill_2 FILLER_9_87 ();
 sg13g2_fill_1 FILLER_9_89 ();
 sg13g2_fill_2 FILLER_9_170 ();
 sg13g2_fill_1 FILLER_9_198 ();
 sg13g2_fill_2 FILLER_9_211 ();
 sg13g2_decap_8 FILLER_9_249 ();
 sg13g2_decap_4 FILLER_9_261 ();
 sg13g2_fill_1 FILLER_9_265 ();
 sg13g2_decap_4 FILLER_9_271 ();
 sg13g2_decap_8 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_316 ();
 sg13g2_decap_8 FILLER_9_323 ();
 sg13g2_decap_8 FILLER_9_330 ();
 sg13g2_decap_8 FILLER_9_337 ();
 sg13g2_decap_8 FILLER_9_344 ();
 sg13g2_decap_8 FILLER_9_351 ();
 sg13g2_decap_8 FILLER_9_358 ();
 sg13g2_decap_8 FILLER_9_365 ();
 sg13g2_decap_8 FILLER_9_372 ();
 sg13g2_decap_8 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_21 ();
 sg13g2_fill_1 FILLER_10_23 ();
 sg13g2_decap_8 FILLER_10_38 ();
 sg13g2_fill_2 FILLER_10_45 ();
 sg13g2_fill_1 FILLER_10_51 ();
 sg13g2_fill_1 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_fill_2 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_4 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_120 ();
 sg13g2_decap_8 FILLER_10_127 ();
 sg13g2_fill_2 FILLER_10_134 ();
 sg13g2_fill_1 FILLER_10_136 ();
 sg13g2_fill_1 FILLER_10_154 ();
 sg13g2_fill_2 FILLER_10_171 ();
 sg13g2_fill_1 FILLER_10_173 ();
 sg13g2_fill_2 FILLER_10_208 ();
 sg13g2_fill_1 FILLER_10_210 ();
 sg13g2_fill_2 FILLER_10_216 ();
 sg13g2_fill_1 FILLER_10_243 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_fill_2 FILLER_10_270 ();
 sg13g2_fill_2 FILLER_10_302 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_decap_4 FILLER_10_320 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_40 ();
 sg13g2_decap_8 FILLER_11_47 ();
 sg13g2_fill_2 FILLER_11_54 ();
 sg13g2_fill_1 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_62 ();
 sg13g2_fill_1 FILLER_11_93 ();
 sg13g2_fill_1 FILLER_11_103 ();
 sg13g2_decap_4 FILLER_11_114 ();
 sg13g2_decap_8 FILLER_11_138 ();
 sg13g2_decap_4 FILLER_11_145 ();
 sg13g2_fill_1 FILLER_11_149 ();
 sg13g2_decap_4 FILLER_11_155 ();
 sg13g2_fill_2 FILLER_11_159 ();
 sg13g2_fill_2 FILLER_11_196 ();
 sg13g2_fill_1 FILLER_11_198 ();
 sg13g2_fill_1 FILLER_11_225 ();
 sg13g2_fill_1 FILLER_11_236 ();
 sg13g2_fill_2 FILLER_11_283 ();
 sg13g2_fill_1 FILLER_11_285 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_fill_2 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_fill_2 FILLER_11_360 ();
 sg13g2_fill_1 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_8 FILLER_11_393 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_fill_1 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_45 ();
 sg13g2_fill_2 FILLER_12_82 ();
 sg13g2_fill_1 FILLER_12_84 ();
 sg13g2_fill_2 FILLER_12_93 ();
 sg13g2_fill_1 FILLER_12_95 ();
 sg13g2_fill_1 FILLER_12_119 ();
 sg13g2_fill_2 FILLER_12_136 ();
 sg13g2_fill_1 FILLER_12_138 ();
 sg13g2_decap_8 FILLER_12_183 ();
 sg13g2_fill_2 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_218 ();
 sg13g2_decap_8 FILLER_12_225 ();
 sg13g2_fill_2 FILLER_12_232 ();
 sg13g2_fill_2 FILLER_12_283 ();
 sg13g2_fill_1 FILLER_12_285 ();
 sg13g2_fill_1 FILLER_12_317 ();
 sg13g2_fill_2 FILLER_12_339 ();
 sg13g2_fill_1 FILLER_12_352 ();
 sg13g2_decap_4 FILLER_12_386 ();
 sg13g2_fill_2 FILLER_12_390 ();
 sg13g2_fill_2 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_13_69 ();
 sg13g2_fill_1 FILLER_13_71 ();
 sg13g2_fill_1 FILLER_13_107 ();
 sg13g2_fill_2 FILLER_13_118 ();
 sg13g2_fill_1 FILLER_13_120 ();
 sg13g2_decap_8 FILLER_13_137 ();
 sg13g2_decap_4 FILLER_13_144 ();
 sg13g2_fill_1 FILLER_13_151 ();
 sg13g2_decap_4 FILLER_13_161 ();
 sg13g2_fill_2 FILLER_13_165 ();
 sg13g2_decap_8 FILLER_13_171 ();
 sg13g2_decap_4 FILLER_13_178 ();
 sg13g2_fill_1 FILLER_13_182 ();
 sg13g2_fill_2 FILLER_13_206 ();
 sg13g2_fill_1 FILLER_13_208 ();
 sg13g2_decap_4 FILLER_13_213 ();
 sg13g2_fill_2 FILLER_13_217 ();
 sg13g2_fill_2 FILLER_13_223 ();
 sg13g2_decap_4 FILLER_13_236 ();
 sg13g2_fill_2 FILLER_13_240 ();
 sg13g2_fill_1 FILLER_13_251 ();
 sg13g2_fill_1 FILLER_13_288 ();
 sg13g2_fill_1 FILLER_13_367 ();
 sg13g2_fill_1 FILLER_13_378 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_4 ();
 sg13g2_fill_2 FILLER_14_63 ();
 sg13g2_fill_1 FILLER_14_77 ();
 sg13g2_fill_2 FILLER_14_102 ();
 sg13g2_fill_2 FILLER_14_117 ();
 sg13g2_fill_1 FILLER_14_119 ();
 sg13g2_fill_2 FILLER_14_137 ();
 sg13g2_fill_1 FILLER_14_147 ();
 sg13g2_fill_2 FILLER_14_156 ();
 sg13g2_fill_2 FILLER_14_211 ();
 sg13g2_decap_8 FILLER_14_247 ();
 sg13g2_fill_2 FILLER_14_254 ();
 sg13g2_fill_1 FILLER_14_359 ();
 sg13g2_fill_1 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_4 FILLER_15_14 ();
 sg13g2_fill_2 FILLER_15_22 ();
 sg13g2_fill_1 FILLER_15_24 ();
 sg13g2_fill_2 FILLER_15_29 ();
 sg13g2_fill_1 FILLER_15_31 ();
 sg13g2_decap_8 FILLER_15_41 ();
 sg13g2_fill_2 FILLER_15_48 ();
 sg13g2_fill_2 FILLER_15_59 ();
 sg13g2_decap_8 FILLER_15_65 ();
 sg13g2_decap_8 FILLER_15_72 ();
 sg13g2_decap_8 FILLER_15_79 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_fill_2 FILLER_15_98 ();
 sg13g2_fill_1 FILLER_15_129 ();
 sg13g2_fill_2 FILLER_15_180 ();
 sg13g2_fill_1 FILLER_15_182 ();
 sg13g2_fill_2 FILLER_15_192 ();
 sg13g2_fill_1 FILLER_15_194 ();
 sg13g2_fill_1 FILLER_15_261 ();
 sg13g2_fill_2 FILLER_15_295 ();
 sg13g2_fill_1 FILLER_15_297 ();
 sg13g2_fill_1 FILLER_15_316 ();
 sg13g2_fill_2 FILLER_15_391 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_4 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_50 ();
 sg13g2_decap_8 FILLER_16_57 ();
 sg13g2_fill_2 FILLER_16_69 ();
 sg13g2_fill_2 FILLER_16_75 ();
 sg13g2_fill_1 FILLER_16_77 ();
 sg13g2_fill_2 FILLER_16_83 ();
 sg13g2_fill_1 FILLER_16_85 ();
 sg13g2_decap_8 FILLER_16_95 ();
 sg13g2_decap_4 FILLER_16_102 ();
 sg13g2_decap_8 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_117 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_fill_2 FILLER_16_125 ();
 sg13g2_fill_1 FILLER_16_127 ();
 sg13g2_decap_8 FILLER_16_145 ();
 sg13g2_decap_4 FILLER_16_152 ();
 sg13g2_fill_2 FILLER_16_156 ();
 sg13g2_fill_1 FILLER_16_171 ();
 sg13g2_decap_4 FILLER_16_225 ();
 sg13g2_decap_4 FILLER_16_261 ();
 sg13g2_decap_4 FILLER_16_277 ();
 sg13g2_fill_2 FILLER_16_281 ();
 sg13g2_decap_4 FILLER_16_287 ();
 sg13g2_fill_1 FILLER_16_291 ();
 sg13g2_fill_2 FILLER_16_309 ();
 sg13g2_fill_1 FILLER_16_311 ();
 sg13g2_fill_1 FILLER_16_335 ();
 sg13g2_fill_1 FILLER_16_349 ();
 sg13g2_fill_1 FILLER_16_372 ();
 sg13g2_fill_2 FILLER_16_385 ();
 sg13g2_fill_1 FILLER_17_26 ();
 sg13g2_fill_1 FILLER_17_47 ();
 sg13g2_fill_1 FILLER_17_64 ();
 sg13g2_fill_2 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_4 FILLER_17_112 ();
 sg13g2_fill_2 FILLER_17_116 ();
 sg13g2_fill_1 FILLER_17_126 ();
 sg13g2_fill_1 FILLER_17_132 ();
 sg13g2_fill_1 FILLER_17_164 ();
 sg13g2_fill_2 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_211 ();
 sg13g2_decap_8 FILLER_17_218 ();
 sg13g2_decap_8 FILLER_17_225 ();
 sg13g2_fill_1 FILLER_17_232 ();
 sg13g2_fill_2 FILLER_17_254 ();
 sg13g2_fill_1 FILLER_17_256 ();
 sg13g2_decap_8 FILLER_17_262 ();
 sg13g2_decap_8 FILLER_17_269 ();
 sg13g2_fill_2 FILLER_17_276 ();
 sg13g2_fill_1 FILLER_17_278 ();
 sg13g2_fill_2 FILLER_17_288 ();
 sg13g2_fill_2 FILLER_17_300 ();
 sg13g2_fill_1 FILLER_17_302 ();
 sg13g2_fill_1 FILLER_17_350 ();
 sg13g2_fill_1 FILLER_17_390 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_fill_1 FILLER_18_117 ();
 sg13g2_fill_2 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_128 ();
 sg13g2_fill_2 FILLER_18_137 ();
 sg13g2_fill_1 FILLER_18_163 ();
 sg13g2_fill_1 FILLER_18_195 ();
 sg13g2_fill_2 FILLER_18_220 ();
 sg13g2_fill_2 FILLER_18_234 ();
 sg13g2_fill_1 FILLER_18_236 ();
 sg13g2_fill_2 FILLER_18_266 ();
 sg13g2_fill_2 FILLER_18_325 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_fill_2 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_374 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_8 ();
 sg13g2_fill_2 FILLER_19_51 ();
 sg13g2_fill_1 FILLER_19_53 ();
 sg13g2_fill_2 FILLER_19_61 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_124 ();
 sg13g2_fill_2 FILLER_19_133 ();
 sg13g2_fill_1 FILLER_19_160 ();
 sg13g2_fill_2 FILLER_19_175 ();
 sg13g2_fill_1 FILLER_19_177 ();
 sg13g2_fill_2 FILLER_19_197 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_fill_2 FILLER_19_205 ();
 sg13g2_fill_2 FILLER_19_242 ();
 sg13g2_decap_8 FILLER_19_253 ();
 sg13g2_decap_4 FILLER_19_265 ();
 sg13g2_fill_1 FILLER_19_274 ();
 sg13g2_fill_1 FILLER_19_296 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_fill_2 FILLER_19_313 ();
 sg13g2_fill_2 FILLER_19_339 ();
 sg13g2_fill_2 FILLER_19_368 ();
 sg13g2_fill_1 FILLER_19_370 ();
 sg13g2_fill_2 FILLER_19_376 ();
 sg13g2_fill_1 FILLER_19_378 ();
 sg13g2_fill_2 FILLER_19_389 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_45 ();
 sg13g2_decap_8 FILLER_20_55 ();
 sg13g2_decap_4 FILLER_20_80 ();
 sg13g2_fill_2 FILLER_20_84 ();
 sg13g2_decap_4 FILLER_20_89 ();
 sg13g2_fill_2 FILLER_20_93 ();
 sg13g2_fill_1 FILLER_20_103 ();
 sg13g2_fill_2 FILLER_20_111 ();
 sg13g2_fill_1 FILLER_20_113 ();
 sg13g2_fill_2 FILLER_20_124 ();
 sg13g2_fill_2 FILLER_20_173 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_fill_1 FILLER_20_205 ();
 sg13g2_fill_2 FILLER_20_261 ();
 sg13g2_fill_1 FILLER_20_263 ();
 sg13g2_fill_1 FILLER_20_295 ();
 sg13g2_fill_2 FILLER_20_313 ();
 sg13g2_fill_2 FILLER_20_320 ();
 sg13g2_fill_2 FILLER_20_342 ();
 sg13g2_fill_2 FILLER_20_369 ();
 sg13g2_fill_2 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_14 ();
 sg13g2_decap_4 FILLER_21_34 ();
 sg13g2_decap_4 FILLER_21_50 ();
 sg13g2_fill_2 FILLER_21_62 ();
 sg13g2_decap_8 FILLER_21_87 ();
 sg13g2_decap_8 FILLER_21_94 ();
 sg13g2_decap_8 FILLER_21_101 ();
 sg13g2_decap_8 FILLER_21_108 ();
 sg13g2_decap_4 FILLER_21_115 ();
 sg13g2_fill_1 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_125 ();
 sg13g2_decap_4 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_136 ();
 sg13g2_fill_2 FILLER_21_180 ();
 sg13g2_fill_2 FILLER_21_195 ();
 sg13g2_fill_2 FILLER_21_229 ();
 sg13g2_fill_2 FILLER_21_271 ();
 sg13g2_fill_1 FILLER_21_342 ();
 sg13g2_decap_4 FILLER_21_351 ();
 sg13g2_fill_2 FILLER_21_371 ();
 sg13g2_fill_1 FILLER_21_373 ();
 sg13g2_fill_2 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_fill_2 FILLER_22_21 ();
 sg13g2_fill_1 FILLER_22_23 ();
 sg13g2_decap_4 FILLER_22_29 ();
 sg13g2_fill_1 FILLER_22_33 ();
 sg13g2_fill_1 FILLER_22_65 ();
 sg13g2_fill_1 FILLER_22_83 ();
 sg13g2_fill_1 FILLER_22_112 ();
 sg13g2_fill_1 FILLER_22_118 ();
 sg13g2_decap_8 FILLER_22_132 ();
 sg13g2_decap_4 FILLER_22_139 ();
 sg13g2_fill_2 FILLER_22_143 ();
 sg13g2_fill_1 FILLER_22_150 ();
 sg13g2_fill_2 FILLER_22_168 ();
 sg13g2_fill_1 FILLER_22_170 ();
 sg13g2_fill_2 FILLER_22_176 ();
 sg13g2_fill_1 FILLER_22_222 ();
 sg13g2_fill_1 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_281 ();
 sg13g2_fill_1 FILLER_22_336 ();
 sg13g2_decap_4 FILLER_22_346 ();
 sg13g2_decap_8 FILLER_22_355 ();
 sg13g2_fill_1 FILLER_22_362 ();
 sg13g2_fill_1 FILLER_22_386 ();
 sg13g2_fill_1 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_26 ();
 sg13g2_decap_8 FILLER_23_33 ();
 sg13g2_fill_2 FILLER_23_40 ();
 sg13g2_fill_1 FILLER_23_42 ();
 sg13g2_fill_2 FILLER_23_109 ();
 sg13g2_fill_1 FILLER_23_111 ();
 sg13g2_fill_1 FILLER_23_128 ();
 sg13g2_fill_2 FILLER_23_156 ();
 sg13g2_fill_2 FILLER_23_181 ();
 sg13g2_decap_4 FILLER_23_197 ();
 sg13g2_fill_1 FILLER_23_201 ();
 sg13g2_fill_1 FILLER_23_289 ();
 sg13g2_fill_2 FILLER_23_316 ();
 sg13g2_decap_4 FILLER_23_351 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_23 ();
 sg13g2_decap_8 FILLER_24_41 ();
 sg13g2_fill_2 FILLER_24_48 ();
 sg13g2_decap_4 FILLER_24_59 ();
 sg13g2_fill_2 FILLER_24_73 ();
 sg13g2_fill_1 FILLER_24_86 ();
 sg13g2_fill_1 FILLER_24_117 ();
 sg13g2_fill_2 FILLER_24_129 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_fill_2 FILLER_24_243 ();
 sg13g2_fill_2 FILLER_24_266 ();
 sg13g2_fill_1 FILLER_24_268 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_fill_1 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_25_54 ();
 sg13g2_decap_8 FILLER_25_61 ();
 sg13g2_decap_8 FILLER_25_68 ();
 sg13g2_decap_8 FILLER_25_80 ();
 sg13g2_fill_2 FILLER_25_87 ();
 sg13g2_fill_2 FILLER_25_129 ();
 sg13g2_fill_2 FILLER_25_135 ();
 sg13g2_fill_1 FILLER_25_150 ();
 sg13g2_fill_2 FILLER_25_173 ();
 sg13g2_decap_4 FILLER_25_214 ();
 sg13g2_fill_1 FILLER_25_218 ();
 sg13g2_decap_8 FILLER_25_232 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_fill_2 FILLER_25_259 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_fill_2 FILLER_25_274 ();
 sg13g2_fill_1 FILLER_25_276 ();
 sg13g2_decap_4 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_317 ();
 sg13g2_decap_4 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_decap_4 FILLER_25_337 ();
 sg13g2_fill_2 FILLER_25_341 ();
 sg13g2_fill_2 FILLER_25_371 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_4 ();
 sg13g2_fill_2 FILLER_26_55 ();
 sg13g2_fill_1 FILLER_26_57 ();
 sg13g2_fill_1 FILLER_26_67 ();
 sg13g2_decap_4 FILLER_26_76 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_fill_1 FILLER_26_130 ();
 sg13g2_fill_1 FILLER_26_140 ();
 sg13g2_fill_1 FILLER_26_149 ();
 sg13g2_decap_4 FILLER_26_155 ();
 sg13g2_fill_1 FILLER_26_159 ();
 sg13g2_decap_4 FILLER_26_164 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_4 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_decap_4 FILLER_26_228 ();
 sg13g2_fill_1 FILLER_26_232 ();
 sg13g2_fill_2 FILLER_26_290 ();
 sg13g2_decap_4 FILLER_26_304 ();
 sg13g2_fill_1 FILLER_26_308 ();
 sg13g2_fill_2 FILLER_26_318 ();
 sg13g2_fill_1 FILLER_26_320 ();
 sg13g2_decap_8 FILLER_26_338 ();
 sg13g2_decap_8 FILLER_26_345 ();
 sg13g2_decap_4 FILLER_26_356 ();
 sg13g2_fill_2 FILLER_26_360 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_14 ();
 sg13g2_fill_1 FILLER_27_43 ();
 sg13g2_fill_2 FILLER_27_103 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_decap_8 FILLER_27_172 ();
 sg13g2_fill_1 FILLER_27_179 ();
 sg13g2_fill_2 FILLER_27_185 ();
 sg13g2_fill_1 FILLER_27_243 ();
 sg13g2_decap_4 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_266 ();
 sg13g2_fill_2 FILLER_27_296 ();
 sg13g2_fill_1 FILLER_27_336 ();
 sg13g2_fill_2 FILLER_27_362 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_18 ();
 sg13g2_fill_2 FILLER_28_40 ();
 sg13g2_fill_1 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_102 ();
 sg13g2_fill_1 FILLER_28_144 ();
 sg13g2_decap_4 FILLER_28_175 ();
 sg13g2_fill_1 FILLER_28_179 ();
 sg13g2_fill_1 FILLER_28_193 ();
 sg13g2_fill_2 FILLER_28_216 ();
 sg13g2_fill_1 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_227 ();
 sg13g2_fill_2 FILLER_28_233 ();
 sg13g2_fill_1 FILLER_28_250 ();
 sg13g2_fill_1 FILLER_28_264 ();
 sg13g2_decap_4 FILLER_28_333 ();
 sg13g2_fill_2 FILLER_28_337 ();
 sg13g2_fill_2 FILLER_28_356 ();
 sg13g2_fill_1 FILLER_28_358 ();
 sg13g2_fill_2 FILLER_28_376 ();
 sg13g2_fill_1 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_14 ();
 sg13g2_fill_1 FILLER_29_16 ();
 sg13g2_fill_1 FILLER_29_34 ();
 sg13g2_fill_1 FILLER_29_40 ();
 sg13g2_fill_2 FILLER_29_46 ();
 sg13g2_fill_1 FILLER_29_48 ();
 sg13g2_fill_2 FILLER_29_70 ();
 sg13g2_fill_1 FILLER_29_81 ();
 sg13g2_fill_2 FILLER_29_92 ();
 sg13g2_fill_2 FILLER_29_129 ();
 sg13g2_fill_2 FILLER_29_144 ();
 sg13g2_fill_1 FILLER_29_146 ();
 sg13g2_fill_1 FILLER_29_153 ();
 sg13g2_fill_2 FILLER_29_170 ();
 sg13g2_fill_1 FILLER_29_198 ();
 sg13g2_decap_4 FILLER_29_225 ();
 sg13g2_fill_1 FILLER_29_229 ();
 sg13g2_fill_2 FILLER_29_316 ();
 sg13g2_fill_1 FILLER_29_318 ();
 sg13g2_fill_2 FILLER_29_336 ();
 sg13g2_fill_2 FILLER_29_359 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_50 ();
 sg13g2_fill_1 FILLER_30_52 ();
 sg13g2_decap_8 FILLER_30_85 ();
 sg13g2_fill_1 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_fill_2 FILLER_30_144 ();
 sg13g2_fill_2 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_222 ();
 sg13g2_decap_8 FILLER_30_229 ();
 sg13g2_fill_2 FILLER_30_236 ();
 sg13g2_fill_1 FILLER_30_238 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_fill_1 FILLER_30_273 ();
 sg13g2_fill_2 FILLER_30_283 ();
 sg13g2_fill_2 FILLER_30_305 ();
 sg13g2_fill_1 FILLER_30_328 ();
 sg13g2_fill_1 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_22 ();
 sg13g2_fill_2 FILLER_31_42 ();
 sg13g2_fill_1 FILLER_31_60 ();
 sg13g2_decap_4 FILLER_31_66 ();
 sg13g2_fill_2 FILLER_31_70 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_fill_2 FILLER_31_81 ();
 sg13g2_fill_1 FILLER_31_83 ();
 sg13g2_decap_8 FILLER_31_94 ();
 sg13g2_decap_4 FILLER_31_109 ();
 sg13g2_fill_2 FILLER_31_113 ();
 sg13g2_fill_2 FILLER_31_146 ();
 sg13g2_fill_2 FILLER_31_159 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_214 ();
 sg13g2_decap_4 FILLER_31_352 ();
 sg13g2_fill_1 FILLER_31_356 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_16 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_fill_2 FILLER_32_62 ();
 sg13g2_fill_1 FILLER_32_64 ();
 sg13g2_fill_1 FILLER_32_79 ();
 sg13g2_fill_2 FILLER_32_92 ();
 sg13g2_decap_8 FILLER_32_99 ();
 sg13g2_fill_2 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_108 ();
 sg13g2_fill_2 FILLER_32_118 ();
 sg13g2_fill_2 FILLER_32_132 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_fill_1 FILLER_32_143 ();
 sg13g2_fill_1 FILLER_32_189 ();
 sg13g2_fill_2 FILLER_32_267 ();
 sg13g2_fill_1 FILLER_32_304 ();
 sg13g2_fill_2 FILLER_32_354 ();
 sg13g2_fill_2 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_18 ();
 sg13g2_fill_1 FILLER_33_45 ();
 sg13g2_fill_1 FILLER_33_70 ();
 sg13g2_decap_4 FILLER_33_96 ();
 sg13g2_fill_2 FILLER_33_100 ();
 sg13g2_fill_2 FILLER_33_128 ();
 sg13g2_decap_4 FILLER_33_135 ();
 sg13g2_decap_8 FILLER_33_211 ();
 sg13g2_fill_2 FILLER_33_218 ();
 sg13g2_fill_1 FILLER_33_268 ();
 sg13g2_fill_2 FILLER_33_278 ();
 sg13g2_fill_1 FILLER_33_280 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_fill_1 FILLER_33_333 ();
 sg13g2_fill_2 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_357 ();
 sg13g2_fill_2 FILLER_33_376 ();
 sg13g2_fill_2 FILLER_33_383 ();
 sg13g2_fill_1 FILLER_33_385 ();
 sg13g2_fill_2 FILLER_33_391 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_28 ();
 sg13g2_decap_4 FILLER_34_34 ();
 sg13g2_fill_1 FILLER_34_50 ();
 sg13g2_fill_1 FILLER_34_92 ();
 sg13g2_fill_2 FILLER_34_107 ();
 sg13g2_decap_4 FILLER_34_118 ();
 sg13g2_decap_8 FILLER_34_131 ();
 sg13g2_fill_1 FILLER_34_145 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_fill_1 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_296 ();
 sg13g2_fill_1 FILLER_34_348 ();
 sg13g2_fill_1 FILLER_34_374 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_fill_1 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_37 ();
 sg13g2_fill_2 FILLER_35_59 ();
 sg13g2_fill_1 FILLER_35_61 ();
 sg13g2_fill_2 FILLER_35_71 ();
 sg13g2_fill_2 FILLER_35_90 ();
 sg13g2_fill_2 FILLER_35_100 ();
 sg13g2_decap_8 FILLER_35_113 ();
 sg13g2_fill_2 FILLER_35_124 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_fill_2 FILLER_35_152 ();
 sg13g2_fill_1 FILLER_35_154 ();
 sg13g2_fill_2 FILLER_35_168 ();
 sg13g2_fill_1 FILLER_35_196 ();
 sg13g2_fill_2 FILLER_35_206 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_fill_1 FILLER_35_222 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_fill_1 FILLER_35_305 ();
 sg13g2_decap_8 FILLER_35_352 ();
 sg13g2_decap_8 FILLER_35_359 ();
 sg13g2_decap_4 FILLER_35_366 ();
 sg13g2_fill_2 FILLER_35_370 ();
 sg13g2_fill_2 FILLER_35_384 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_28 ();
 sg13g2_fill_2 FILLER_36_32 ();
 sg13g2_decap_4 FILLER_36_65 ();
 sg13g2_decap_4 FILLER_36_76 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_4 FILLER_36_106 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_143 ();
 sg13g2_fill_1 FILLER_36_162 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_309 ();
 sg13g2_fill_2 FILLER_36_345 ();
 sg13g2_fill_1 FILLER_36_347 ();
 sg13g2_fill_1 FILLER_36_352 ();
 sg13g2_fill_2 FILLER_36_358 ();
 sg13g2_fill_1 FILLER_36_360 ();
 sg13g2_fill_2 FILLER_36_389 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_53 ();
 sg13g2_decap_8 FILLER_37_58 ();
 sg13g2_fill_1 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_79 ();
 sg13g2_fill_2 FILLER_37_86 ();
 sg13g2_fill_2 FILLER_37_96 ();
 sg13g2_fill_2 FILLER_37_110 ();
 sg13g2_fill_1 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_155 ();
 sg13g2_fill_2 FILLER_37_166 ();
 sg13g2_fill_1 FILLER_37_208 ();
 sg13g2_fill_2 FILLER_37_223 ();
 sg13g2_fill_1 FILLER_37_225 ();
 sg13g2_decap_8 FILLER_37_243 ();
 sg13g2_fill_2 FILLER_37_250 ();
 sg13g2_fill_2 FILLER_37_257 ();
 sg13g2_decap_4 FILLER_37_285 ();
 sg13g2_fill_2 FILLER_37_289 ();
 sg13g2_fill_1 FILLER_37_336 ();
 sg13g2_fill_2 FILLER_37_396 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_4 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_32 ();
 sg13g2_decap_4 FILLER_38_38 ();
 sg13g2_fill_1 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_48 ();
 sg13g2_decap_4 FILLER_38_81 ();
 sg13g2_fill_2 FILLER_38_85 ();
 sg13g2_fill_2 FILLER_38_95 ();
 sg13g2_fill_1 FILLER_38_113 ();
 sg13g2_fill_2 FILLER_38_150 ();
 sg13g2_fill_1 FILLER_38_152 ();
 sg13g2_fill_2 FILLER_38_170 ();
 sg13g2_fill_2 FILLER_38_204 ();
 sg13g2_fill_2 FILLER_38_219 ();
 sg13g2_fill_1 FILLER_38_226 ();
 sg13g2_decap_4 FILLER_38_256 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_4 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_305 ();
 sg13g2_fill_2 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_4 FILLER_39_49 ();
 sg13g2_fill_2 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_123 ();
 sg13g2_decap_4 FILLER_39_130 ();
 sg13g2_fill_1 FILLER_39_134 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_fill_2 FILLER_39_147 ();
 sg13g2_fill_1 FILLER_39_149 ();
 sg13g2_fill_1 FILLER_39_154 ();
 sg13g2_fill_2 FILLER_39_189 ();
 sg13g2_fill_2 FILLER_39_246 ();
 sg13g2_fill_1 FILLER_39_248 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_fill_1 FILLER_39_308 ();
 sg13g2_fill_1 FILLER_39_382 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_fill_2 FILLER_40_21 ();
 sg13g2_fill_1 FILLER_40_37 ();
 sg13g2_fill_2 FILLER_40_53 ();
 sg13g2_fill_1 FILLER_40_62 ();
 sg13g2_fill_2 FILLER_40_114 ();
 sg13g2_fill_2 FILLER_40_124 ();
 sg13g2_decap_4 FILLER_40_155 ();
 sg13g2_fill_1 FILLER_40_159 ();
 sg13g2_fill_2 FILLER_40_181 ();
 sg13g2_decap_4 FILLER_40_207 ();
 sg13g2_fill_2 FILLER_40_225 ();
 sg13g2_fill_1 FILLER_40_239 ();
 sg13g2_fill_2 FILLER_40_254 ();
 sg13g2_fill_2 FILLER_40_282 ();
 sg13g2_decap_8 FILLER_40_310 ();
 sg13g2_decap_4 FILLER_40_317 ();
 sg13g2_fill_1 FILLER_40_321 ();
 sg13g2_decap_4 FILLER_40_349 ();
 sg13g2_fill_1 FILLER_40_353 ();
 sg13g2_fill_2 FILLER_40_370 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_fill_2 FILLER_41_25 ();
 sg13g2_fill_1 FILLER_41_27 ();
 sg13g2_fill_1 FILLER_41_44 ();
 sg13g2_fill_2 FILLER_41_57 ();
 sg13g2_fill_1 FILLER_41_59 ();
 sg13g2_fill_2 FILLER_41_68 ();
 sg13g2_fill_1 FILLER_41_70 ();
 sg13g2_fill_1 FILLER_41_80 ();
 sg13g2_fill_1 FILLER_41_86 ();
 sg13g2_fill_2 FILLER_41_92 ();
 sg13g2_fill_1 FILLER_41_94 ();
 sg13g2_decap_8 FILLER_41_106 ();
 sg13g2_decap_4 FILLER_41_113 ();
 sg13g2_fill_1 FILLER_41_117 ();
 sg13g2_fill_1 FILLER_41_135 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_fill_1 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_193 ();
 sg13g2_decap_4 FILLER_41_205 ();
 sg13g2_fill_1 FILLER_41_209 ();
 sg13g2_fill_2 FILLER_41_241 ();
 sg13g2_fill_1 FILLER_41_243 ();
 sg13g2_fill_2 FILLER_41_285 ();
 sg13g2_fill_1 FILLER_41_309 ();
 sg13g2_fill_2 FILLER_41_354 ();
 sg13g2_fill_1 FILLER_41_356 ();
 sg13g2_decap_4 FILLER_41_370 ();
 sg13g2_fill_2 FILLER_41_374 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_23 ();
 sg13g2_fill_2 FILLER_42_30 ();
 sg13g2_fill_1 FILLER_42_45 ();
 sg13g2_decap_4 FILLER_42_51 ();
 sg13g2_fill_1 FILLER_42_55 ();
 sg13g2_fill_2 FILLER_42_72 ();
 sg13g2_fill_1 FILLER_42_74 ();
 sg13g2_fill_2 FILLER_42_96 ();
 sg13g2_fill_1 FILLER_42_107 ();
 sg13g2_fill_1 FILLER_42_123 ();
 sg13g2_decap_4 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_205 ();
 sg13g2_fill_2 FILLER_42_212 ();
 sg13g2_fill_1 FILLER_42_214 ();
 sg13g2_fill_1 FILLER_42_241 ();
 sg13g2_fill_1 FILLER_42_270 ();
 sg13g2_decap_4 FILLER_42_310 ();
 sg13g2_fill_1 FILLER_42_314 ();
 sg13g2_decap_4 FILLER_42_340 ();
 sg13g2_fill_1 FILLER_42_344 ();
 sg13g2_fill_2 FILLER_42_351 ();
 sg13g2_decap_8 FILLER_42_367 ();
 sg13g2_decap_8 FILLER_42_383 ();
 sg13g2_fill_2 FILLER_42_390 ();
 sg13g2_fill_1 FILLER_42_392 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_9 ();
 sg13g2_decap_8 FILLER_43_15 ();
 sg13g2_decap_4 FILLER_43_22 ();
 sg13g2_fill_2 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_4 FILLER_43_63 ();
 sg13g2_fill_1 FILLER_43_67 ();
 sg13g2_fill_2 FILLER_43_99 ();
 sg13g2_fill_1 FILLER_43_101 ();
 sg13g2_fill_2 FILLER_43_163 ();
 sg13g2_fill_1 FILLER_43_171 ();
 sg13g2_fill_1 FILLER_43_177 ();
 sg13g2_fill_1 FILLER_43_186 ();
 sg13g2_fill_1 FILLER_43_221 ();
 sg13g2_fill_2 FILLER_43_261 ();
 sg13g2_fill_1 FILLER_43_272 ();
 sg13g2_fill_1 FILLER_43_281 ();
 sg13g2_fill_1 FILLER_43_286 ();
 sg13g2_fill_1 FILLER_43_313 ();
 sg13g2_fill_1 FILLER_43_323 ();
 sg13g2_fill_1 FILLER_43_329 ();
 sg13g2_fill_2 FILLER_43_343 ();
 sg13g2_fill_2 FILLER_43_350 ();
 sg13g2_fill_1 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_400 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_15 ();
 sg13g2_fill_1 FILLER_44_17 ();
 sg13g2_decap_4 FILLER_44_43 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_fill_2 FILLER_44_77 ();
 sg13g2_fill_1 FILLER_44_83 ();
 sg13g2_decap_4 FILLER_44_88 ();
 sg13g2_fill_1 FILLER_44_92 ();
 sg13g2_decap_4 FILLER_44_97 ();
 sg13g2_fill_1 FILLER_44_101 ();
 sg13g2_fill_2 FILLER_44_139 ();
 sg13g2_decap_8 FILLER_44_165 ();
 sg13g2_fill_2 FILLER_44_172 ();
 sg13g2_fill_2 FILLER_44_202 ();
 sg13g2_fill_1 FILLER_44_209 ();
 sg13g2_fill_1 FILLER_44_230 ();
 sg13g2_fill_2 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_278 ();
 sg13g2_decap_8 FILLER_44_285 ();
 sg13g2_fill_1 FILLER_44_292 ();
 sg13g2_fill_1 FILLER_44_320 ();
 sg13g2_fill_1 FILLER_44_356 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_4 ();
 sg13g2_fill_2 FILLER_45_27 ();
 sg13g2_fill_1 FILLER_45_29 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_fill_1 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_117 ();
 sg13g2_fill_2 FILLER_45_136 ();
 sg13g2_fill_1 FILLER_45_138 ();
 sg13g2_decap_8 FILLER_45_144 ();
 sg13g2_fill_1 FILLER_45_151 ();
 sg13g2_fill_2 FILLER_45_157 ();
 sg13g2_decap_4 FILLER_45_162 ();
 sg13g2_fill_2 FILLER_45_177 ();
 sg13g2_fill_1 FILLER_45_179 ();
 sg13g2_fill_1 FILLER_45_212 ();
 sg13g2_fill_2 FILLER_45_225 ();
 sg13g2_fill_2 FILLER_45_333 ();
 sg13g2_fill_1 FILLER_45_357 ();
 sg13g2_fill_2 FILLER_45_371 ();
 sg13g2_fill_1 FILLER_45_373 ();
 sg13g2_fill_1 FILLER_45_382 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_27 ();
 sg13g2_fill_2 FILLER_46_50 ();
 sg13g2_fill_1 FILLER_46_52 ();
 sg13g2_decap_4 FILLER_46_70 ();
 sg13g2_fill_1 FILLER_46_100 ();
 sg13g2_decap_8 FILLER_46_113 ();
 sg13g2_fill_2 FILLER_46_120 ();
 sg13g2_fill_2 FILLER_46_135 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_4 FILLER_46_189 ();
 sg13g2_fill_1 FILLER_46_205 ();
 sg13g2_fill_2 FILLER_46_211 ();
 sg13g2_fill_1 FILLER_46_223 ();
 sg13g2_decap_4 FILLER_46_250 ();
 sg13g2_fill_1 FILLER_46_283 ();
 sg13g2_fill_2 FILLER_46_308 ();
 sg13g2_fill_2 FILLER_46_324 ();
 sg13g2_fill_2 FILLER_46_381 ();
 sg13g2_fill_1 FILLER_46_383 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_7 ();
 sg13g2_fill_1 FILLER_47_9 ();
 sg13g2_fill_1 FILLER_47_19 ();
 sg13g2_fill_1 FILLER_47_33 ();
 sg13g2_fill_2 FILLER_47_54 ();
 sg13g2_decap_4 FILLER_47_81 ();
 sg13g2_fill_1 FILLER_47_89 ();
 sg13g2_fill_2 FILLER_47_105 ();
 sg13g2_decap_4 FILLER_47_120 ();
 sg13g2_fill_2 FILLER_47_124 ();
 sg13g2_fill_2 FILLER_47_145 ();
 sg13g2_fill_2 FILLER_47_155 ();
 sg13g2_decap_8 FILLER_47_187 ();
 sg13g2_decap_4 FILLER_47_194 ();
 sg13g2_fill_2 FILLER_47_198 ();
 sg13g2_fill_2 FILLER_47_209 ();
 sg13g2_fill_2 FILLER_47_229 ();
 sg13g2_fill_1 FILLER_47_231 ();
 sg13g2_fill_2 FILLER_47_236 ();
 sg13g2_fill_2 FILLER_47_258 ();
 sg13g2_fill_1 FILLER_47_296 ();
 sg13g2_fill_2 FILLER_47_336 ();
 sg13g2_fill_2 FILLER_47_349 ();
 sg13g2_fill_2 FILLER_47_354 ();
 sg13g2_fill_2 FILLER_47_372 ();
 sg13g2_fill_1 FILLER_47_374 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_4 ();
 sg13g2_fill_1 FILLER_48_21 ();
 sg13g2_fill_2 FILLER_48_32 ();
 sg13g2_decap_8 FILLER_48_82 ();
 sg13g2_decap_4 FILLER_48_89 ();
 sg13g2_fill_1 FILLER_48_93 ();
 sg13g2_fill_2 FILLER_48_104 ();
 sg13g2_decap_8 FILLER_48_123 ();
 sg13g2_decap_8 FILLER_48_130 ();
 sg13g2_fill_1 FILLER_48_151 ();
 sg13g2_fill_2 FILLER_48_192 ();
 sg13g2_fill_2 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_4 FILLER_48_224 ();
 sg13g2_fill_1 FILLER_48_228 ();
 sg13g2_decap_4 FILLER_48_241 ();
 sg13g2_fill_1 FILLER_48_245 ();
 sg13g2_fill_1 FILLER_48_253 ();
 sg13g2_decap_8 FILLER_48_262 ();
 sg13g2_fill_2 FILLER_48_269 ();
 sg13g2_fill_2 FILLER_48_295 ();
 sg13g2_decap_8 FILLER_48_345 ();
 sg13g2_fill_1 FILLER_48_352 ();
 sg13g2_decap_4 FILLER_48_356 ();
 sg13g2_fill_1 FILLER_48_360 ();
 sg13g2_fill_1 FILLER_48_366 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_27 ();
 sg13g2_decap_8 FILLER_49_78 ();
 sg13g2_fill_1 FILLER_49_85 ();
 sg13g2_fill_2 FILLER_49_138 ();
 sg13g2_fill_2 FILLER_49_152 ();
 sg13g2_fill_1 FILLER_49_154 ();
 sg13g2_decap_4 FILLER_49_159 ();
 sg13g2_fill_1 FILLER_49_176 ();
 sg13g2_decap_4 FILLER_49_181 ();
 sg13g2_fill_2 FILLER_49_185 ();
 sg13g2_decap_8 FILLER_49_213 ();
 sg13g2_decap_8 FILLER_49_220 ();
 sg13g2_fill_2 FILLER_49_246 ();
 sg13g2_fill_2 FILLER_49_265 ();
 sg13g2_decap_8 FILLER_49_351 ();
 sg13g2_fill_2 FILLER_49_391 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_2 ();
 sg13g2_fill_1 FILLER_50_25 ();
 sg13g2_fill_2 FILLER_50_35 ();
 sg13g2_fill_1 FILLER_50_37 ();
 sg13g2_fill_2 FILLER_50_43 ();
 sg13g2_fill_2 FILLER_50_69 ();
 sg13g2_fill_1 FILLER_50_71 ();
 sg13g2_fill_2 FILLER_50_77 ();
 sg13g2_fill_1 FILLER_50_79 ();
 sg13g2_fill_1 FILLER_50_109 ();
 sg13g2_fill_2 FILLER_50_127 ();
 sg13g2_decap_8 FILLER_50_156 ();
 sg13g2_decap_8 FILLER_50_163 ();
 sg13g2_fill_2 FILLER_50_170 ();
 sg13g2_decap_4 FILLER_50_181 ();
 sg13g2_fill_1 FILLER_50_185 ();
 sg13g2_fill_2 FILLER_50_220 ();
 sg13g2_decap_4 FILLER_50_232 ();
 sg13g2_fill_2 FILLER_50_241 ();
 sg13g2_fill_2 FILLER_50_251 ();
 sg13g2_fill_2 FILLER_50_272 ();
 sg13g2_fill_1 FILLER_50_274 ();
 sg13g2_fill_2 FILLER_50_332 ();
 sg13g2_fill_2 FILLER_50_392 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_7 ();
 sg13g2_fill_1 FILLER_51_9 ();
 sg13g2_fill_2 FILLER_51_14 ();
 sg13g2_fill_1 FILLER_51_16 ();
 sg13g2_fill_1 FILLER_51_22 ();
 sg13g2_fill_1 FILLER_51_33 ();
 sg13g2_fill_2 FILLER_51_58 ();
 sg13g2_fill_1 FILLER_51_73 ();
 sg13g2_fill_2 FILLER_51_113 ();
 sg13g2_fill_1 FILLER_51_115 ();
 sg13g2_fill_2 FILLER_51_144 ();
 sg13g2_fill_1 FILLER_51_151 ();
 sg13g2_fill_2 FILLER_51_192 ();
 sg13g2_fill_1 FILLER_51_194 ();
 sg13g2_fill_2 FILLER_51_271 ();
 sg13g2_fill_2 FILLER_51_316 ();
 sg13g2_fill_1 FILLER_51_318 ();
 sg13g2_fill_1 FILLER_51_374 ();
 sg13g2_fill_1 FILLER_51_388 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_13 ();
 sg13g2_fill_1 FILLER_52_15 ();
 sg13g2_fill_2 FILLER_52_27 ();
 sg13g2_fill_1 FILLER_52_29 ();
 sg13g2_fill_1 FILLER_52_72 ();
 sg13g2_fill_1 FILLER_52_79 ();
 sg13g2_fill_2 FILLER_52_119 ();
 sg13g2_fill_2 FILLER_52_191 ();
 sg13g2_fill_1 FILLER_52_193 ();
 sg13g2_fill_1 FILLER_52_220 ();
 sg13g2_fill_1 FILLER_52_230 ();
 sg13g2_fill_2 FILLER_52_259 ();
 sg13g2_fill_1 FILLER_52_261 ();
 sg13g2_fill_2 FILLER_52_291 ();
 sg13g2_fill_1 FILLER_52_350 ();
 sg13g2_fill_1 FILLER_52_376 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_46 ();
 sg13g2_fill_1 FILLER_53_48 ();
 sg13g2_fill_2 FILLER_53_54 ();
 sg13g2_fill_2 FILLER_53_71 ();
 sg13g2_fill_1 FILLER_53_73 ();
 sg13g2_fill_2 FILLER_53_103 ();
 sg13g2_fill_2 FILLER_53_114 ();
 sg13g2_decap_4 FILLER_53_132 ();
 sg13g2_fill_1 FILLER_53_166 ();
 sg13g2_fill_2 FILLER_53_193 ();
 sg13g2_fill_1 FILLER_53_195 ();
 sg13g2_fill_2 FILLER_53_234 ();
 sg13g2_decap_4 FILLER_53_244 ();
 sg13g2_fill_2 FILLER_53_248 ();
 sg13g2_fill_1 FILLER_53_254 ();
 sg13g2_fill_2 FILLER_53_263 ();
 sg13g2_fill_1 FILLER_53_265 ();
 sg13g2_fill_2 FILLER_53_284 ();
 sg13g2_fill_1 FILLER_53_290 ();
 sg13g2_fill_2 FILLER_53_335 ();
 sg13g2_fill_1 FILLER_53_370 ();
 sg13g2_fill_2 FILLER_53_397 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_7 ();
 sg13g2_fill_1 FILLER_54_9 ();
 sg13g2_fill_2 FILLER_54_71 ();
 sg13g2_fill_1 FILLER_54_73 ();
 sg13g2_decap_8 FILLER_54_85 ();
 sg13g2_decap_8 FILLER_54_92 ();
 sg13g2_decap_8 FILLER_54_99 ();
 sg13g2_decap_8 FILLER_54_106 ();
 sg13g2_decap_4 FILLER_54_113 ();
 sg13g2_fill_1 FILLER_54_117 ();
 sg13g2_fill_2 FILLER_54_126 ();
 sg13g2_decap_4 FILLER_54_137 ();
 sg13g2_fill_2 FILLER_54_141 ();
 sg13g2_decap_4 FILLER_54_156 ();
 sg13g2_fill_2 FILLER_54_160 ();
 sg13g2_fill_2 FILLER_54_172 ();
 sg13g2_fill_1 FILLER_54_182 ();
 sg13g2_fill_2 FILLER_54_207 ();
 sg13g2_fill_2 FILLER_54_235 ();
 sg13g2_fill_1 FILLER_54_237 ();
 sg13g2_fill_2 FILLER_54_276 ();
 sg13g2_fill_1 FILLER_54_278 ();
 sg13g2_decap_4 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_13 ();
 sg13g2_fill_2 FILLER_55_19 ();
 sg13g2_fill_1 FILLER_55_21 ();
 sg13g2_fill_2 FILLER_55_26 ();
 sg13g2_fill_2 FILLER_55_41 ();
 sg13g2_fill_1 FILLER_55_54 ();
 sg13g2_decap_8 FILLER_55_59 ();
 sg13g2_fill_1 FILLER_55_66 ();
 sg13g2_fill_2 FILLER_55_81 ();
 sg13g2_decap_4 FILLER_55_87 ();
 sg13g2_fill_2 FILLER_55_91 ();
 sg13g2_fill_2 FILLER_55_134 ();
 sg13g2_fill_1 FILLER_55_136 ();
 sg13g2_decap_4 FILLER_55_142 ();
 sg13g2_fill_1 FILLER_55_167 ();
 sg13g2_decap_8 FILLER_55_182 ();
 sg13g2_decap_4 FILLER_55_189 ();
 sg13g2_fill_2 FILLER_55_193 ();
 sg13g2_fill_1 FILLER_55_263 ();
 sg13g2_fill_2 FILLER_55_281 ();
 sg13g2_fill_1 FILLER_55_360 ();
 sg13g2_fill_1 FILLER_55_366 ();
 sg13g2_fill_1 FILLER_55_382 ();
 sg13g2_fill_2 FILLER_56_16 ();
 sg13g2_fill_1 FILLER_56_18 ();
 sg13g2_fill_2 FILLER_56_24 ();
 sg13g2_fill_1 FILLER_56_26 ();
 sg13g2_fill_1 FILLER_56_62 ();
 sg13g2_fill_1 FILLER_56_93 ();
 sg13g2_fill_2 FILLER_56_128 ();
 sg13g2_fill_1 FILLER_56_142 ();
 sg13g2_fill_1 FILLER_56_174 ();
 sg13g2_fill_2 FILLER_56_184 ();
 sg13g2_fill_2 FILLER_56_210 ();
 sg13g2_fill_1 FILLER_56_212 ();
 sg13g2_fill_2 FILLER_56_218 ();
 sg13g2_fill_2 FILLER_56_239 ();
 sg13g2_fill_1 FILLER_56_241 ();
 sg13g2_fill_1 FILLER_56_247 ();
 sg13g2_decap_4 FILLER_56_252 ();
 sg13g2_decap_8 FILLER_56_274 ();
 sg13g2_fill_2 FILLER_56_281 ();
 sg13g2_fill_1 FILLER_56_283 ();
 sg13g2_fill_2 FILLER_56_317 ();
 sg13g2_fill_1 FILLER_56_328 ();
 sg13g2_fill_2 FILLER_56_353 ();
 sg13g2_fill_1 FILLER_56_355 ();
 sg13g2_fill_1 FILLER_56_382 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_decap_4 FILLER_57_24 ();
 sg13g2_fill_1 FILLER_57_28 ();
 sg13g2_fill_2 FILLER_57_33 ();
 sg13g2_fill_1 FILLER_57_35 ();
 sg13g2_fill_2 FILLER_57_78 ();
 sg13g2_fill_1 FILLER_57_94 ();
 sg13g2_fill_1 FILLER_57_106 ();
 sg13g2_fill_2 FILLER_57_131 ();
 sg13g2_fill_1 FILLER_57_133 ();
 sg13g2_fill_2 FILLER_57_175 ();
 sg13g2_fill_1 FILLER_57_177 ();
 sg13g2_fill_2 FILLER_57_198 ();
 sg13g2_fill_1 FILLER_57_249 ();
 sg13g2_fill_1 FILLER_57_270 ();
 sg13g2_fill_1 FILLER_57_279 ();
 sg13g2_fill_1 FILLER_57_358 ();
 sg13g2_fill_1 FILLER_57_368 ();
 sg13g2_fill_1 FILLER_57_397 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_21 ();
 sg13g2_fill_1 FILLER_58_32 ();
 sg13g2_decap_8 FILLER_58_38 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_fill_2 FILLER_58_56 ();
 sg13g2_decap_4 FILLER_58_64 ();
 sg13g2_fill_2 FILLER_58_68 ();
 sg13g2_decap_8 FILLER_58_74 ();
 sg13g2_fill_2 FILLER_58_81 ();
 sg13g2_decap_4 FILLER_58_108 ();
 sg13g2_fill_2 FILLER_58_112 ();
 sg13g2_fill_1 FILLER_58_144 ();
 sg13g2_decap_8 FILLER_58_154 ();
 sg13g2_fill_2 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_fill_2 FILLER_58_289 ();
 sg13g2_fill_1 FILLER_58_357 ();
 sg13g2_fill_2 FILLER_58_373 ();
 sg13g2_fill_2 FILLER_58_389 ();
 sg13g2_fill_1 FILLER_58_391 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_16 ();
 sg13g2_fill_1 FILLER_59_18 ();
 sg13g2_fill_2 FILLER_59_24 ();
 sg13g2_fill_2 FILLER_59_31 ();
 sg13g2_fill_1 FILLER_59_33 ();
 sg13g2_fill_1 FILLER_59_56 ();
 sg13g2_fill_1 FILLER_59_62 ();
 sg13g2_decap_4 FILLER_59_77 ();
 sg13g2_fill_1 FILLER_59_81 ();
 sg13g2_fill_2 FILLER_59_92 ();
 sg13g2_decap_8 FILLER_59_99 ();
 sg13g2_decap_8 FILLER_59_106 ();
 sg13g2_decap_8 FILLER_59_113 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_decap_8 FILLER_59_140 ();
 sg13g2_decap_4 FILLER_59_147 ();
 sg13g2_fill_1 FILLER_59_151 ();
 sg13g2_fill_1 FILLER_59_165 ();
 sg13g2_fill_2 FILLER_59_182 ();
 sg13g2_fill_1 FILLER_59_184 ();
 sg13g2_fill_2 FILLER_59_220 ();
 sg13g2_fill_2 FILLER_59_231 ();
 sg13g2_decap_4 FILLER_59_268 ();
 sg13g2_fill_1 FILLER_59_272 ();
 sg13g2_fill_1 FILLER_59_282 ();
 sg13g2_fill_1 FILLER_59_297 ();
 sg13g2_fill_2 FILLER_59_352 ();
 sg13g2_fill_1 FILLER_59_354 ();
 sg13g2_fill_2 FILLER_59_381 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_2 ();
 sg13g2_fill_2 FILLER_60_18 ();
 sg13g2_fill_1 FILLER_60_20 ();
 sg13g2_fill_2 FILLER_60_32 ();
 sg13g2_fill_1 FILLER_60_34 ();
 sg13g2_fill_1 FILLER_60_80 ();
 sg13g2_decap_4 FILLER_60_98 ();
 sg13g2_fill_1 FILLER_60_102 ();
 sg13g2_fill_2 FILLER_60_116 ();
 sg13g2_fill_2 FILLER_60_154 ();
 sg13g2_decap_8 FILLER_60_183 ();
 sg13g2_fill_2 FILLER_60_190 ();
 sg13g2_fill_1 FILLER_60_192 ();
 sg13g2_decap_8 FILLER_60_211 ();
 sg13g2_fill_1 FILLER_60_218 ();
 sg13g2_fill_2 FILLER_60_223 ();
 sg13g2_fill_1 FILLER_60_331 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_24 ();
 sg13g2_fill_2 FILLER_61_105 ();
 sg13g2_decap_4 FILLER_61_123 ();
 sg13g2_decap_4 FILLER_61_132 ();
 sg13g2_fill_1 FILLER_61_136 ();
 sg13g2_decap_4 FILLER_61_141 ();
 sg13g2_fill_2 FILLER_61_145 ();
 sg13g2_fill_1 FILLER_61_157 ();
 sg13g2_fill_1 FILLER_61_171 ();
 sg13g2_decap_4 FILLER_61_185 ();
 sg13g2_decap_8 FILLER_61_200 ();
 sg13g2_fill_2 FILLER_61_211 ();
 sg13g2_decap_4 FILLER_61_223 ();
 sg13g2_fill_2 FILLER_61_240 ();
 sg13g2_fill_2 FILLER_61_268 ();
 sg13g2_fill_1 FILLER_61_270 ();
 sg13g2_fill_2 FILLER_61_302 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_7 ();
 sg13g2_fill_2 FILLER_62_30 ();
 sg13g2_fill_2 FILLER_62_47 ();
 sg13g2_decap_4 FILLER_62_64 ();
 sg13g2_fill_2 FILLER_62_68 ();
 sg13g2_decap_8 FILLER_62_100 ();
 sg13g2_decap_4 FILLER_62_107 ();
 sg13g2_fill_2 FILLER_62_131 ();
 sg13g2_fill_1 FILLER_62_147 ();
 sg13g2_decap_4 FILLER_62_189 ();
 sg13g2_fill_2 FILLER_62_244 ();
 sg13g2_fill_1 FILLER_62_246 ();
 sg13g2_fill_1 FILLER_62_265 ();
 sg13g2_fill_1 FILLER_62_297 ();
 sg13g2_fill_1 FILLER_62_327 ();
 sg13g2_fill_1 FILLER_62_365 ();
 sg13g2_fill_2 FILLER_62_370 ();
 sg13g2_fill_2 FILLER_62_382 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_7 ();
 sg13g2_decap_4 FILLER_63_29 ();
 sg13g2_fill_2 FILLER_63_33 ();
 sg13g2_fill_1 FILLER_63_49 ();
 sg13g2_fill_2 FILLER_63_55 ();
 sg13g2_fill_1 FILLER_63_57 ();
 sg13g2_decap_4 FILLER_63_62 ();
 sg13g2_fill_2 FILLER_63_66 ();
 sg13g2_decap_8 FILLER_63_73 ();
 sg13g2_decap_4 FILLER_63_80 ();
 sg13g2_fill_1 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_89 ();
 sg13g2_decap_8 FILLER_63_96 ();
 sg13g2_fill_1 FILLER_63_103 ();
 sg13g2_decap_8 FILLER_63_107 ();
 sg13g2_fill_1 FILLER_63_118 ();
 sg13g2_fill_1 FILLER_63_141 ();
 sg13g2_fill_1 FILLER_63_166 ();
 sg13g2_fill_2 FILLER_63_184 ();
 sg13g2_decap_4 FILLER_63_242 ();
 sg13g2_fill_2 FILLER_63_246 ();
 sg13g2_decap_4 FILLER_63_274 ();
 sg13g2_fill_2 FILLER_63_324 ();
 sg13g2_fill_2 FILLER_63_334 ();
 sg13g2_fill_1 FILLER_63_355 ();
 sg13g2_fill_1 FILLER_63_369 ();
 sg13g2_fill_2 FILLER_63_396 ();
 sg13g2_fill_1 FILLER_63_398 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_18 ();
 sg13g2_fill_2 FILLER_64_25 ();
 sg13g2_fill_1 FILLER_64_27 ();
 sg13g2_fill_2 FILLER_64_56 ();
 sg13g2_fill_1 FILLER_64_58 ();
 sg13g2_fill_2 FILLER_64_74 ();
 sg13g2_fill_1 FILLER_64_76 ();
 sg13g2_fill_1 FILLER_64_96 ();
 sg13g2_fill_2 FILLER_64_138 ();
 sg13g2_decap_8 FILLER_64_158 ();
 sg13g2_decap_4 FILLER_64_165 ();
 sg13g2_decap_4 FILLER_64_173 ();
 sg13g2_fill_2 FILLER_64_177 ();
 sg13g2_fill_1 FILLER_64_201 ();
 sg13g2_fill_2 FILLER_64_272 ();
 sg13g2_fill_2 FILLER_64_286 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_23 ();
 sg13g2_fill_1 FILLER_65_25 ();
 sg13g2_fill_2 FILLER_65_40 ();
 sg13g2_fill_1 FILLER_65_42 ();
 sg13g2_fill_2 FILLER_65_49 ();
 sg13g2_fill_2 FILLER_65_62 ();
 sg13g2_decap_4 FILLER_65_77 ();
 sg13g2_fill_2 FILLER_65_144 ();
 sg13g2_fill_2 FILLER_65_150 ();
 sg13g2_fill_2 FILLER_65_169 ();
 sg13g2_fill_1 FILLER_65_171 ();
 sg13g2_fill_2 FILLER_65_186 ();
 sg13g2_fill_2 FILLER_65_223 ();
 sg13g2_fill_2 FILLER_65_256 ();
 sg13g2_fill_1 FILLER_65_258 ();
 sg13g2_fill_1 FILLER_65_285 ();
 sg13g2_fill_2 FILLER_65_341 ();
 sg13g2_fill_2 FILLER_65_393 ();
 sg13g2_fill_1 FILLER_65_395 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_2 ();
 sg13g2_decap_4 FILLER_66_48 ();
 sg13g2_fill_1 FILLER_66_82 ();
 sg13g2_fill_1 FILLER_66_97 ();
 sg13g2_fill_1 FILLER_66_124 ();
 sg13g2_fill_1 FILLER_66_149 ();
 sg13g2_fill_2 FILLER_66_202 ();
 sg13g2_fill_2 FILLER_66_239 ();
 sg13g2_fill_1 FILLER_66_290 ();
 sg13g2_fill_1 FILLER_66_331 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_4 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_4 ();
 sg13g2_fill_2 FILLER_67_47 ();
 sg13g2_fill_1 FILLER_67_49 ();
 sg13g2_fill_1 FILLER_67_64 ();
 sg13g2_fill_2 FILLER_67_70 ();
 sg13g2_fill_2 FILLER_67_81 ();
 sg13g2_decap_8 FILLER_67_87 ();
 sg13g2_decap_4 FILLER_67_94 ();
 sg13g2_fill_2 FILLER_67_105 ();
 sg13g2_fill_1 FILLER_67_107 ();
 sg13g2_fill_1 FILLER_67_113 ();
 sg13g2_fill_2 FILLER_67_138 ();
 sg13g2_fill_1 FILLER_67_156 ();
 sg13g2_fill_1 FILLER_67_175 ();
 sg13g2_fill_2 FILLER_67_249 ();
 sg13g2_fill_2 FILLER_67_327 ();
 sg13g2_fill_1 FILLER_67_334 ();
 sg13g2_fill_1 FILLER_67_358 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_19 ();
 sg13g2_decap_8 FILLER_68_36 ();
 sg13g2_decap_8 FILLER_68_43 ();
 sg13g2_fill_2 FILLER_68_70 ();
 sg13g2_fill_2 FILLER_68_78 ();
 sg13g2_decap_8 FILLER_68_85 ();
 sg13g2_decap_8 FILLER_68_92 ();
 sg13g2_fill_2 FILLER_68_99 ();
 sg13g2_fill_2 FILLER_68_106 ();
 sg13g2_fill_1 FILLER_68_108 ();
 sg13g2_fill_1 FILLER_68_117 ();
 sg13g2_fill_2 FILLER_68_139 ();
 sg13g2_fill_1 FILLER_68_185 ();
 sg13g2_fill_2 FILLER_68_208 ();
 sg13g2_fill_1 FILLER_68_210 ();
 sg13g2_fill_1 FILLER_68_217 ();
 sg13g2_fill_1 FILLER_68_227 ();
 sg13g2_fill_2 FILLER_68_233 ();
 sg13g2_fill_1 FILLER_68_235 ();
 sg13g2_fill_2 FILLER_68_254 ();
 sg13g2_fill_2 FILLER_68_267 ();
 sg13g2_fill_1 FILLER_68_269 ();
 sg13g2_fill_2 FILLER_68_337 ();
 sg13g2_fill_1 FILLER_68_339 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_23 ();
 sg13g2_fill_1 FILLER_69_25 ();
 sg13g2_fill_2 FILLER_69_31 ();
 sg13g2_fill_2 FILLER_69_48 ();
 sg13g2_fill_2 FILLER_69_63 ();
 sg13g2_fill_2 FILLER_69_78 ();
 sg13g2_decap_4 FILLER_69_88 ();
 sg13g2_fill_2 FILLER_69_92 ();
 sg13g2_fill_1 FILLER_69_103 ();
 sg13g2_fill_1 FILLER_69_108 ();
 sg13g2_fill_1 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_123 ();
 sg13g2_fill_1 FILLER_69_130 ();
 sg13g2_decap_4 FILLER_69_139 ();
 sg13g2_decap_8 FILLER_69_152 ();
 sg13g2_fill_2 FILLER_69_172 ();
 sg13g2_fill_1 FILLER_69_191 ();
 sg13g2_fill_2 FILLER_69_207 ();
 sg13g2_fill_2 FILLER_69_231 ();
 sg13g2_fill_1 FILLER_69_233 ();
 sg13g2_fill_2 FILLER_69_244 ();
 sg13g2_fill_1 FILLER_69_281 ();
 sg13g2_fill_1 FILLER_69_287 ();
 sg13g2_fill_1 FILLER_69_309 ();
 sg13g2_fill_2 FILLER_69_322 ();
 sg13g2_fill_1 FILLER_69_363 ();
 sg13g2_fill_2 FILLER_70_16 ();
 sg13g2_fill_2 FILLER_70_33 ();
 sg13g2_fill_1 FILLER_70_35 ();
 sg13g2_fill_2 FILLER_70_49 ();
 sg13g2_fill_2 FILLER_70_94 ();
 sg13g2_fill_1 FILLER_70_96 ();
 sg13g2_decap_8 FILLER_70_129 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_fill_1 FILLER_70_147 ();
 sg13g2_fill_2 FILLER_70_176 ();
 sg13g2_fill_1 FILLER_70_178 ();
 sg13g2_fill_1 FILLER_70_197 ();
 sg13g2_fill_1 FILLER_70_215 ();
 sg13g2_fill_1 FILLER_70_231 ();
 sg13g2_fill_1 FILLER_70_250 ();
 sg13g2_fill_1 FILLER_70_255 ();
 sg13g2_fill_1 FILLER_70_260 ();
 sg13g2_fill_2 FILLER_70_278 ();
 sg13g2_fill_1 FILLER_70_307 ();
 sg13g2_fill_1 FILLER_70_354 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_fill_2 FILLER_71_70 ();
 sg13g2_fill_1 FILLER_71_72 ();
 sg13g2_fill_2 FILLER_71_133 ();
 sg13g2_fill_2 FILLER_71_140 ();
 sg13g2_fill_1 FILLER_71_150 ();
 sg13g2_fill_2 FILLER_71_174 ();
 sg13g2_fill_1 FILLER_71_193 ();
 sg13g2_fill_2 FILLER_71_214 ();
 sg13g2_fill_1 FILLER_71_216 ();
 sg13g2_fill_2 FILLER_71_339 ();
 sg13g2_fill_2 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_72_2 ();
 sg13g2_fill_1 FILLER_72_58 ();
 sg13g2_fill_2 FILLER_72_68 ();
 sg13g2_fill_2 FILLER_72_75 ();
 sg13g2_fill_1 FILLER_72_77 ();
 sg13g2_fill_1 FILLER_72_83 ();
 sg13g2_fill_2 FILLER_72_121 ();
 sg13g2_fill_1 FILLER_72_123 ();
 sg13g2_fill_1 FILLER_72_151 ();
 sg13g2_fill_1 FILLER_72_302 ();
 sg13g2_fill_2 FILLER_72_352 ();
 sg13g2_fill_2 FILLER_72_398 ();
 sg13g2_decap_4 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_4 ();
 sg13g2_fill_2 FILLER_73_31 ();
 sg13g2_fill_1 FILLER_73_33 ();
 sg13g2_fill_2 FILLER_73_49 ();
 sg13g2_decap_4 FILLER_73_55 ();
 sg13g2_fill_2 FILLER_73_59 ();
 sg13g2_decap_4 FILLER_73_66 ();
 sg13g2_decap_8 FILLER_73_79 ();
 sg13g2_decap_4 FILLER_73_86 ();
 sg13g2_fill_2 FILLER_73_90 ();
 sg13g2_fill_2 FILLER_73_127 ();
 sg13g2_fill_1 FILLER_73_129 ();
 sg13g2_decap_4 FILLER_73_135 ();
 sg13g2_fill_2 FILLER_73_139 ();
 sg13g2_fill_2 FILLER_73_144 ();
 sg13g2_fill_1 FILLER_73_151 ();
 sg13g2_fill_2 FILLER_73_155 ();
 sg13g2_fill_1 FILLER_73_157 ();
 sg13g2_fill_2 FILLER_73_185 ();
 sg13g2_fill_2 FILLER_73_337 ();
 sg13g2_fill_1 FILLER_73_353 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_30 ();
 sg13g2_fill_1 FILLER_74_37 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_fill_2 FILLER_74_56 ();
 sg13g2_fill_1 FILLER_74_58 ();
 sg13g2_fill_2 FILLER_74_67 ();
 sg13g2_decap_8 FILLER_74_81 ();
 sg13g2_decap_4 FILLER_74_88 ();
 sg13g2_fill_1 FILLER_74_92 ();
 sg13g2_decap_4 FILLER_74_106 ();
 sg13g2_fill_2 FILLER_74_110 ();
 sg13g2_decap_8 FILLER_74_120 ();
 sg13g2_decap_8 FILLER_74_127 ();
 sg13g2_decap_8 FILLER_74_134 ();
 sg13g2_fill_1 FILLER_74_141 ();
 sg13g2_decap_8 FILLER_74_152 ();
 sg13g2_decap_8 FILLER_74_159 ();
 sg13g2_decap_4 FILLER_74_178 ();
 sg13g2_fill_1 FILLER_74_230 ();
 sg13g2_fill_2 FILLER_74_257 ();
 sg13g2_fill_2 FILLER_74_327 ();
 sg13g2_fill_1 FILLER_74_339 ();
 sg13g2_fill_2 FILLER_74_350 ();
 sg13g2_fill_1 FILLER_74_371 ();
 sg13g2_fill_2 FILLER_74_381 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_4 FILLER_75_7 ();
 sg13g2_fill_1 FILLER_75_11 ();
 sg13g2_fill_1 FILLER_75_42 ();
 sg13g2_fill_1 FILLER_75_52 ();
 sg13g2_fill_1 FILLER_75_71 ();
 sg13g2_fill_2 FILLER_75_92 ();
 sg13g2_fill_1 FILLER_75_94 ();
 sg13g2_fill_2 FILLER_75_110 ();
 sg13g2_fill_1 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_123 ();
 sg13g2_fill_1 FILLER_75_130 ();
 sg13g2_fill_2 FILLER_75_152 ();
 sg13g2_fill_1 FILLER_75_159 ();
 sg13g2_fill_1 FILLER_75_188 ();
 sg13g2_fill_2 FILLER_75_216 ();
 sg13g2_fill_1 FILLER_75_218 ();
 sg13g2_fill_1 FILLER_75_247 ();
 sg13g2_fill_2 FILLER_75_262 ();
 sg13g2_fill_1 FILLER_75_296 ();
 sg13g2_fill_1 FILLER_75_310 ();
 sg13g2_fill_1 FILLER_75_348 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_fill_1 FILLER_76_59 ();
 sg13g2_fill_2 FILLER_76_84 ();
 sg13g2_fill_2 FILLER_76_101 ();
 sg13g2_fill_1 FILLER_76_129 ();
 sg13g2_fill_2 FILLER_76_179 ();
 sg13g2_fill_2 FILLER_76_210 ();
 sg13g2_fill_2 FILLER_76_226 ();
 sg13g2_fill_2 FILLER_76_302 ();
 sg13g2_fill_2 FILLER_76_323 ();
 sg13g2_fill_1 FILLER_76_334 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_fill_1 FILLER_77_132 ();
 sg13g2_fill_2 FILLER_77_185 ();
 sg13g2_fill_1 FILLER_77_187 ();
 sg13g2_fill_2 FILLER_77_203 ();
 sg13g2_fill_1 FILLER_77_231 ();
 sg13g2_fill_1 FILLER_77_293 ();
 sg13g2_fill_1 FILLER_77_330 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_fill_2 FILLER_78_28 ();
 sg13g2_fill_2 FILLER_78_35 ();
 sg13g2_fill_2 FILLER_78_54 ();
 sg13g2_fill_2 FILLER_78_80 ();
 sg13g2_fill_2 FILLER_78_136 ();
 sg13g2_fill_1 FILLER_78_209 ();
 sg13g2_fill_2 FILLER_78_389 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_4 FILLER_79_42 ();
 sg13g2_fill_2 FILLER_79_59 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_fill_2 FILLER_79_84 ();
 sg13g2_fill_1 FILLER_79_86 ();
 sg13g2_fill_2 FILLER_79_100 ();
 sg13g2_fill_1 FILLER_79_102 ();
 sg13g2_fill_2 FILLER_79_108 ();
 sg13g2_fill_1 FILLER_79_110 ();
 sg13g2_decap_8 FILLER_79_125 ();
 sg13g2_fill_2 FILLER_79_169 ();
 sg13g2_fill_1 FILLER_79_171 ();
 sg13g2_fill_1 FILLER_79_198 ();
 sg13g2_fill_2 FILLER_79_375 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_fill_2 FILLER_80_100 ();
 sg13g2_fill_2 FILLER_80_110 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_8 FILLER_80_123 ();
 sg13g2_decap_8 FILLER_80_130 ();
 sg13g2_decap_8 FILLER_80_137 ();
 sg13g2_fill_2 FILLER_80_144 ();
 sg13g2_decap_8 FILLER_80_154 ();
 sg13g2_decap_8 FILLER_80_161 ();
 sg13g2_fill_1 FILLER_80_168 ();
 sg13g2_fill_1 FILLER_80_256 ();
 sg13g2_fill_2 FILLER_80_299 ();
 sg13g2_fill_1 FILLER_80_301 ();
 sg13g2_fill_2 FILLER_80_365 ();
 assign uio_oe[0] = net231;
 assign uio_oe[1] = net232;
 assign uio_oe[2] = net233;
 assign uio_oe[3] = net234;
 assign uio_oe[4] = net235;
 assign uio_oe[5] = net236;
 assign uio_oe[6] = net237;
 assign uio_oe[7] = net238;
endmodule

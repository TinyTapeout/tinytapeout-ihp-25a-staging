module tt_um_betz_morse_keyer (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire \main.aux_dah_o ;
 wire \main.aux_dit_o ;
 wire \main.aux_morse_o ;
 wire \main.buzzer_o ;
 wire \main.code_dah ;
 wire \main.code_dit ;
 wire \main.dah_r ;
 wire \main.db0.cnt[0] ;
 wire \main.db0.cnt[10] ;
 wire \main.db0.cnt[11] ;
 wire \main.db0.cnt[12] ;
 wire \main.db0.cnt[13] ;
 wire \main.db0.cnt[1] ;
 wire \main.db0.cnt[2] ;
 wire \main.db0.cnt[3] ;
 wire \main.db0.cnt[4] ;
 wire \main.db0.cnt[5] ;
 wire \main.db0.cnt[6] ;
 wire \main.db0.cnt[7] ;
 wire \main.db0.cnt[8] ;
 wire \main.db0.cnt[9] ;
 wire \main.db0.sig_o ;
 wire \main.db0.sig_r[0] ;
 wire \main.db0.sig_r[1] ;
 wire \main.db0.sig_r[2] ;
 wire \main.db1.cnt[0] ;
 wire \main.db1.cnt[10] ;
 wire \main.db1.cnt[11] ;
 wire \main.db1.cnt[12] ;
 wire \main.db1.cnt[13] ;
 wire \main.db1.cnt[1] ;
 wire \main.db1.cnt[2] ;
 wire \main.db1.cnt[3] ;
 wire \main.db1.cnt[4] ;
 wire \main.db1.cnt[5] ;
 wire \main.db1.cnt[6] ;
 wire \main.db1.cnt[7] ;
 wire \main.db1.cnt[8] ;
 wire \main.db1.cnt[9] ;
 wire \main.db1.sig_r[0] ;
 wire \main.db1.sig_r[1] ;
 wire \main.db1.sig_r[2] ;
 wire \main.display.data[0] ;
 wire \main.display.data[1] ;
 wire \main.display.data[2] ;
 wire \main.display.data[3] ;
 wire \main.display.data[4] ;
 wire \main.display.data[5] ;
 wire \main.display.mask[0] ;
 wire \main.display.mask[1] ;
 wire \main.display.mask[2] ;
 wire \main.display.mask[3] ;
 wire \main.display.mask[4] ;
 wire \main.display.mask[5] ;
 wire \main.display.strobe_i ;
 wire \main.dit_pulse ;
 wire \main.dit_timer.clk128 ;
 wire \main.dit_timer.clk16 ;
 wire \main.dit_timer.clk2 ;
 wire \main.dit_timer.clk256 ;
 wire \main.dit_timer.clk32 ;
 wire \main.dit_timer.clk4 ;
 wire \main.dit_timer.clk512 ;
 wire \main.dit_timer.clk64 ;
 wire \main.dit_timer.clk8 ;
 wire \main.dit_timer.div1.in_r ;
 wire \main.dit_timer.div2.in_r ;
 wire \main.dit_timer.div3.in_r ;
 wire \main.dit_timer.div4.in_r ;
 wire \main.dit_timer.div5.in_r ;
 wire \main.dit_timer.div6.in_r ;
 wire \main.dit_timer.div7.in_r ;
 wire \main.dit_timer.div8.in_r ;
 wire \main.dit_timer.last_clk512 ;
 wire \main.dit_timer.morse_i ;
 wire \main.dit_timer.pause_count[0] ;
 wire \main.dit_timer.pause_count[1] ;
 wire \main.dit_timer.pause_count[2] ;
 wire \main.dit_timer.pause_count[3] ;
 wire \main.dit_timer.pause_count[4] ;
 wire \main.dit_timer.pause_count[5] ;
 wire \main.dit_timer.timer[0] ;
 wire \main.dit_timer.timer[10] ;
 wire \main.dit_timer.timer[11] ;
 wire \main.dit_timer.timer[1] ;
 wire \main.dit_timer.timer[2] ;
 wire \main.dit_timer.timer[3] ;
 wire \main.dit_timer.timer[4] ;
 wire \main.dit_timer.timer[5] ;
 wire \main.dit_timer.timer[6] ;
 wire \main.dit_timer.timer[7] ;
 wire \main.dit_timer.timer[8] ;
 wire \main.dit_timer.timer[9] ;
 wire \main.dit_timer.timer_en ;
 wire \main.encoder.high_ct[0] ;
 wire \main.encoder.high_ct[1] ;
 wire \main.encoder.low_ct[0] ;
 wire \main.encoder.low_ct[1] ;
 wire \main.encoder.low_ct[2] ;
 wire \main.encoder.low_ct[3] ;
 wire \main.encoder.low_ct[4] ;
 wire \main.encoder.low_ct[5] ;
 wire \main.iambic_morse ;
 wire \main.keyer.current_state[0] ;
 wire \main.keyer.current_state[1] ;
 wire \main.keyer.current_state[2] ;
 wire \main.keyer.current_state[3] ;
 wire \main.keyer.current_state[4] ;
 wire \main.keyer.current_state[5] ;
 wire \main.keyer.current_state[6] ;
 wire \main.keyer.current_state[7] ;
 wire \main.keyer.current_state[8] ;
 wire \main.keyer.dah_count[0] ;
 wire \main.keyer.dah_count[1] ;
 wire net10;
 wire net11;
 wire net25;
 wire net26;
 wire net27;
 wire clknet_0_clk;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;

 sg13g2_inv_1 _0659_ (.Y(_0119_),
    .A(net88));
 sg13g2_inv_1 _0660_ (.Y(_0120_),
    .A(net192));
 sg13g2_inv_1 _0661_ (.Y(_0121_),
    .A(net225));
 sg13g2_inv_2 _0662_ (.Y(_0122_),
    .A(net133));
 sg13g2_inv_2 _0663_ (.Y(_0123_),
    .A(net125));
 sg13g2_inv_1 _0664_ (.Y(_0124_),
    .A(net96));
 sg13g2_inv_1 _0665_ (.Y(_0125_),
    .A(net99));
 sg13g2_inv_1 _0666_ (.Y(_0126_),
    .A(net118));
 sg13g2_inv_1 _0667_ (.Y(_0127_),
    .A(net147));
 sg13g2_inv_2 _0668_ (.Y(_0128_),
    .A(net134));
 sg13g2_inv_2 _0669_ (.Y(_0129_),
    .A(net156));
 sg13g2_inv_1 _0670_ (.Y(_0130_),
    .A(net94));
 sg13g2_inv_1 _0671_ (.Y(_0131_),
    .A(net104));
 sg13g2_inv_1 _0672_ (.Y(_0132_),
    .A(net218));
 sg13g2_inv_1 _0673_ (.Y(_0133_),
    .A(net106));
 sg13g2_inv_1 _0674_ (.Y(_0134_),
    .A(net263));
 sg13g2_inv_1 _0675_ (.Y(_0135_),
    .A(\main.dit_timer.pause_count[1] ));
 sg13g2_inv_1 _0676_ (.Y(_0136_),
    .A(net67));
 sg13g2_inv_1 _0677_ (.Y(_0137_),
    .A(\main.dit_timer.pause_count[3] ));
 sg13g2_inv_1 _0678_ (.Y(_0138_),
    .A(net73));
 sg13g2_inv_1 _0679_ (.Y(_0139_),
    .A(\main.display.mask[4] ));
 sg13g2_inv_1 _0680_ (.Y(_0140_),
    .A(net194));
 sg13g2_inv_1 _0681_ (.Y(_0141_),
    .A(net188));
 sg13g2_inv_1 _0682_ (.Y(_0142_),
    .A(net186));
 sg13g2_inv_1 _0683_ (.Y(_0143_),
    .A(net182));
 sg13g2_inv_1 _0684_ (.Y(_0144_),
    .A(net180));
 sg13g2_inv_1 _0685_ (.Y(_0145_),
    .A(net176));
 sg13g2_inv_1 _0686_ (.Y(_0146_),
    .A(net232));
 sg13g2_inv_1 _0687_ (.Y(_0147_),
    .A(net161));
 sg13g2_inv_1 _0688_ (.Y(_0148_),
    .A(net274));
 sg13g2_inv_2 _0689_ (.Y(_0149_),
    .A(net195));
 sg13g2_inv_1 _0690_ (.Y(_0150_),
    .A(net141));
 sg13g2_inv_1 _0691_ (.Y(_0151_),
    .A(net154));
 sg13g2_inv_1 _0692_ (.Y(_0152_),
    .A(net149));
 sg13g2_inv_1 _0693_ (.Y(_0153_),
    .A(net219));
 sg13g2_inv_1 _0694_ (.Y(_0154_),
    .A(net127));
 sg13g2_inv_1 _0695_ (.Y(_0155_),
    .A(net144));
 sg13g2_inv_1 _0696_ (.Y(_0156_),
    .A(net229));
 sg13g2_nand2_1 _0697_ (.Y(_0157_),
    .A(net190),
    .B(net122));
 sg13g2_a21oi_1 _0698_ (.A1(net190),
    .A2(net122),
    .Y(_0158_),
    .B1(net70));
 sg13g2_inv_1 _0699_ (.Y(_0159_),
    .A(_0158_));
 sg13g2_nand2_1 _0700_ (.Y(_0160_),
    .A(net191),
    .B(net140));
 sg13g2_o21ai_1 _0701_ (.B1(_0160_),
    .Y(_0161_),
    .A1(net132),
    .A2(_0158_));
 sg13g2_o21ai_1 _0702_ (.B1(net87),
    .Y(_0162_),
    .A1(net175),
    .A2(_0157_));
 sg13g2_nand2_1 _0703_ (.Y(_0032_),
    .A(_0161_),
    .B(_0162_));
 sg13g2_nor2b_1 _0704_ (.A(net1),
    .B_N(\main.db0.sig_o ),
    .Y(_0163_));
 sg13g2_a21oi_2 _0705_ (.B1(_0163_),
    .Y(_0164_),
    .A2(net1),
    .A1(net124));
 sg13g2_inv_2 _0706_ (.Y(\main.dit_timer.morse_i ),
    .A(_0164_));
 sg13g2_nand2_1 _0707_ (.Y(_0165_),
    .A(net87),
    .B(net2));
 sg13g2_and2_1 _0708_ (.A(net117),
    .B(net191),
    .X(_0166_));
 sg13g2_nand2_1 _0709_ (.Y(_0167_),
    .A(net120),
    .B(_0165_));
 sg13g2_a22oi_1 _0710_ (.Y(_0168_),
    .B1(net175),
    .B2(_0159_),
    .A2(\main.keyer.current_state[5] ),
    .A1(net191));
 sg13g2_o21ai_1 _0711_ (.B1(_0168_),
    .Y(_0003_),
    .A1(_0166_),
    .A2(_0167_));
 sg13g2_nand3_1 _0712_ (.B(net175),
    .C(net122),
    .A(net2),
    .Y(_0169_));
 sg13g2_nor2_1 _0713_ (.A(net190),
    .B(net151),
    .Y(_0170_));
 sg13g2_a22oi_1 _0714_ (.Y(_0004_),
    .B1(_0169_),
    .B2(_0170_),
    .A2(_0126_),
    .A1(net190));
 sg13g2_a21oi_1 _0715_ (.A1(net87),
    .A2(net2),
    .Y(_0171_),
    .B1(net91));
 sg13g2_nor2_2 _0716_ (.A(\main.keyer.current_state[4] ),
    .B(net91),
    .Y(_0172_));
 sg13g2_nor3_1 _0717_ (.A(_0166_),
    .B(_0171_),
    .C(net92),
    .Y(_0002_));
 sg13g2_nand3_1 _0718_ (.B(net175),
    .C(\main.keyer.current_state[8] ),
    .A(net2),
    .Y(_0173_));
 sg13g2_a21oi_1 _0719_ (.A1(_0126_),
    .A2(_0173_),
    .Y(_0006_),
    .B1(net190));
 sg13g2_nor2b_1 _0720_ (.A(net191),
    .B_N(net140),
    .Y(_0174_));
 sg13g2_a22oi_1 _0721_ (.Y(_0175_),
    .B1(_0174_),
    .B2(_0165_),
    .A2(_0166_),
    .A1(net120));
 sg13g2_inv_1 _0722_ (.Y(_0001_),
    .A(_0175_));
 sg13g2_a21oi_1 _0723_ (.A1(net2),
    .A2(net175),
    .Y(_0176_),
    .B1(net190));
 sg13g2_a22oi_1 _0724_ (.Y(_0177_),
    .B1(_0176_),
    .B2(net122),
    .A2(\main.keyer.current_state[8] ),
    .A1(net190));
 sg13g2_inv_1 _0725_ (.Y(_0005_),
    .A(net123));
 sg13g2_nand2_1 _0726_ (.Y(_0178_),
    .A(net91),
    .B(_0166_));
 sg13g2_a21oi_1 _0727_ (.A1(net87),
    .A2(\main.keyer.current_state[2] ),
    .Y(_0179_),
    .B1(net129));
 sg13g2_inv_1 _0728_ (.Y(_0180_),
    .A(_0179_));
 sg13g2_o21ai_1 _0729_ (.B1(_0120_),
    .Y(_0181_),
    .A1(net2),
    .A2(net129));
 sg13g2_o21ai_1 _0730_ (.B1(_0178_),
    .Y(_0000_),
    .A1(net130),
    .A2(_0181_));
 sg13g2_nand3_1 _0731_ (.B(_0132_),
    .C(net92),
    .A(_0126_),
    .Y(_0008_));
 sg13g2_nand2_1 _0732_ (.Y(_0182_),
    .A(\main.db0.sig_o ),
    .B(net70));
 sg13g2_a22oi_1 _0733_ (.Y(_0183_),
    .B1(_0180_),
    .B2(net190),
    .A2(_0176_),
    .A1(\main.keyer.current_state[8] ));
 sg13g2_o21ai_1 _0734_ (.B1(_0183_),
    .Y(_0007_),
    .A1(net175),
    .A2(net71));
 sg13g2_nor2b_2 _0735_ (.A(net85),
    .B_N(\main.dit_timer.morse_i ),
    .Y(_0184_));
 sg13g2_nand2b_2 _0736_ (.Y(_0185_),
    .B(\main.dit_timer.morse_i ),
    .A_N(net85));
 sg13g2_nand3_1 _0737_ (.B(\main.dit_timer.timer[0] ),
    .C(net101),
    .A(\main.dit_timer.timer[1] ),
    .Y(_0186_));
 sg13g2_and4_2 _0738_ (.A(\main.dit_timer.timer[1] ),
    .B(\main.dit_timer.timer[0] ),
    .C(\main.dit_timer.timer[3] ),
    .D(\main.dit_timer.timer[2] ),
    .X(_0187_));
 sg13g2_and2_1 _0739_ (.A(\main.dit_timer.timer[5] ),
    .B(\main.dit_timer.timer[4] ),
    .X(_0188_));
 sg13g2_and2_1 _0740_ (.A(_0187_),
    .B(_0188_),
    .X(_0189_));
 sg13g2_and4_1 _0741_ (.A(net109),
    .B(net160),
    .C(_0187_),
    .D(_0188_),
    .X(_0190_));
 sg13g2_nand4_1 _0742_ (.B(net160),
    .C(_0187_),
    .A(net109),
    .Y(_0191_),
    .D(_0188_));
 sg13g2_xor2_1 _0743_ (.B(net223),
    .A(net6),
    .X(_0192_));
 sg13g2_xor2_1 _0744_ (.B(\main.dit_timer.timer[10] ),
    .A(net5),
    .X(_0193_));
 sg13g2_xor2_1 _0745_ (.B(net112),
    .A(net4),
    .X(_0194_));
 sg13g2_xor2_1 _0746_ (.B(net269),
    .A(net3),
    .X(_0195_));
 sg13g2_nor4_2 _0747_ (.A(_0192_),
    .B(_0193_),
    .C(_0194_),
    .Y(_0196_),
    .D(_0195_));
 sg13g2_nand2_1 _0748_ (.Y(_0197_),
    .A(_0190_),
    .B(net270));
 sg13g2_nor2_1 _0749_ (.A(_0184_),
    .B(_0197_),
    .Y(_0009_));
 sg13g2_nand3_1 _0750_ (.B(_0190_),
    .C(_0196_),
    .A(_0164_),
    .Y(_0198_));
 sg13g2_or2_1 _0751_ (.X(_0199_),
    .B(\main.dit_timer.morse_i ),
    .A(\main.dit_timer.timer_en ));
 sg13g2_o21ai_1 _0752_ (.B1(_0185_),
    .Y(_0200_),
    .A1(_0134_),
    .A2(_0198_));
 sg13g2_nor2b_1 _0753_ (.A(_0200_),
    .B_N(_0199_),
    .Y(_0010_));
 sg13g2_nand2_1 _0754_ (.Y(_0201_),
    .A(net85),
    .B(_0164_));
 sg13g2_and3_1 _0755_ (.X(_0020_),
    .A(net85),
    .B(net58),
    .C(_0164_));
 sg13g2_nor2_1 _0756_ (.A(net58),
    .B(_0201_),
    .Y(_0021_));
 sg13g2_a22oi_1 _0757_ (.Y(_0202_),
    .B1(_0184_),
    .B2(net103),
    .A2(net231),
    .A1(net192));
 sg13g2_nand2_1 _0758_ (.Y(_0022_),
    .A(_0201_),
    .B(_0202_));
 sg13g2_nor2_1 _0759_ (.A(_0026_),
    .B(_0164_),
    .Y(\main.buzzer_o ));
 sg13g2_nor2_2 _0760_ (.A(net174),
    .B(\main.dit_timer.morse_i ),
    .Y(_0203_));
 sg13g2_a21oi_1 _0761_ (.A1(net174),
    .A2(_0133_),
    .Y(_0033_),
    .B1(_0203_));
 sg13g2_nor2b_1 _0762_ (.A(net192),
    .B_N(net58),
    .Y(_0204_));
 sg13g2_a21oi_1 _0763_ (.A1(net192),
    .A2(net106),
    .Y(_0205_),
    .B1(_0204_));
 sg13g2_nor2_1 _0764_ (.A(_0203_),
    .B(_0205_),
    .Y(_0034_));
 sg13g2_nor2b_1 _0765_ (.A(\main.dit_timer.div8.in_r ),
    .B_N(net34),
    .Y(_0206_));
 sg13g2_mux2_1 _0766_ (.A0(net38),
    .A1(net46),
    .S(_0206_),
    .X(_0035_));
 sg13g2_nor2_2 _0767_ (.A(\main.code_dit ),
    .B(net267),
    .Y(_0207_));
 sg13g2_nor2_2 _0768_ (.A(_0149_),
    .B(_0207_),
    .Y(_0208_));
 sg13g2_nand2_1 _0769_ (.Y(_0209_),
    .A(net195),
    .B(_0207_));
 sg13g2_o21ai_1 _0770_ (.B1(net170),
    .Y(_0210_),
    .A1(\main.display.mask[0] ),
    .A2(net138));
 sg13g2_inv_1 _0771_ (.Y(_0036_),
    .A(net139));
 sg13g2_a22oi_1 _0772_ (.Y(_0211_),
    .B1(_0208_),
    .B2(net221),
    .A2(_0149_),
    .A1(net145));
 sg13g2_inv_1 _0773_ (.Y(_0037_),
    .A(net222));
 sg13g2_a22oi_1 _0774_ (.Y(_0212_),
    .B1(_0208_),
    .B2(net145),
    .A2(_0149_),
    .A1(net136));
 sg13g2_inv_1 _0775_ (.Y(_0038_),
    .A(net146));
 sg13g2_a22oi_1 _0776_ (.Y(_0213_),
    .B1(net171),
    .B2(net136),
    .A2(_0149_),
    .A1(\main.display.mask[3] ));
 sg13g2_inv_1 _0777_ (.Y(_0039_),
    .A(net137));
 sg13g2_a22oi_1 _0778_ (.Y(_0214_),
    .B1(net171),
    .B2(net152),
    .A2(_0149_),
    .A1(\main.display.mask[4] ));
 sg13g2_inv_1 _0779_ (.Y(_0040_),
    .A(net153));
 sg13g2_a22oi_1 _0780_ (.Y(_0215_),
    .B1(net171),
    .B2(net243),
    .A2(_0149_),
    .A1(net193));
 sg13g2_inv_1 _0781_ (.Y(_0041_),
    .A(_0215_));
 sg13g2_nand2_2 _0782_ (.Y(_0216_),
    .A(_0185_),
    .B(_0197_));
 sg13g2_nor2b_1 _0783_ (.A(\main.dit_timer.last_clk512 ),
    .B_N(\main.dit_timer.clk512 ),
    .Y(_0217_));
 sg13g2_o21ai_1 _0784_ (.B1(_0217_),
    .Y(_0218_),
    .A1(\main.dit_timer.timer_en ),
    .A2(\main.dit_timer.morse_i ));
 sg13g2_a221oi_1 _0785_ (.B2(_0217_),
    .C1(_0184_),
    .B1(_0199_),
    .A1(_0190_),
    .Y(_0219_),
    .A2(_0196_));
 sg13g2_nand2_1 _0786_ (.Y(_0220_),
    .A(net234),
    .B(_0219_));
 sg13g2_or2_2 _0787_ (.X(_0221_),
    .B(_0219_),
    .A(_0184_));
 sg13g2_o21ai_1 _0788_ (.B1(_0220_),
    .Y(_0042_),
    .A1(net234),
    .A2(_0221_));
 sg13g2_xnor2_1 _0789_ (.Y(_0222_),
    .A(net158),
    .B(\main.dit_timer.timer[0] ));
 sg13g2_nand2_1 _0790_ (.Y(_0223_),
    .A(net158),
    .B(_0219_));
 sg13g2_o21ai_1 _0791_ (.B1(_0223_),
    .Y(_0043_),
    .A1(_0221_),
    .A2(_0222_));
 sg13g2_a21o_1 _0792_ (.A2(\main.dit_timer.timer[0] ),
    .A1(\main.dit_timer.timer[1] ),
    .B1(net101),
    .X(_0224_));
 sg13g2_nand2_1 _0793_ (.Y(_0225_),
    .A(_0186_),
    .B(_0224_));
 sg13g2_nand2_1 _0794_ (.Y(_0226_),
    .A(net101),
    .B(_0219_));
 sg13g2_o21ai_1 _0795_ (.B1(_0226_),
    .Y(_0044_),
    .A1(_0221_),
    .A2(_0225_));
 sg13g2_xor2_1 _0796_ (.B(_0186_),
    .A(net107),
    .X(_0227_));
 sg13g2_nand2_1 _0797_ (.Y(_0228_),
    .A(net107),
    .B(_0219_));
 sg13g2_o21ai_1 _0798_ (.B1(_0228_),
    .Y(_0045_),
    .A1(_0221_),
    .A2(_0227_));
 sg13g2_nor2_1 _0799_ (.A(_0026_),
    .B(_0187_),
    .Y(_0229_));
 sg13g2_and2_1 _0800_ (.A(_0026_),
    .B(_0187_),
    .X(_0230_));
 sg13g2_nor3_1 _0801_ (.A(_0218_),
    .B(_0229_),
    .C(_0230_),
    .Y(_0231_));
 sg13g2_nor2b_1 _0802_ (.A(net115),
    .B_N(_0218_),
    .Y(_0232_));
 sg13g2_nor3_1 _0803_ (.A(_0216_),
    .B(_0231_),
    .C(_0232_),
    .Y(_0046_));
 sg13g2_a21oi_1 _0804_ (.A1(net115),
    .A2(_0187_),
    .Y(_0233_),
    .B1(net131));
 sg13g2_nor3_1 _0805_ (.A(_0189_),
    .B(_0221_),
    .C(_0233_),
    .Y(_0234_));
 sg13g2_a21o_1 _0806_ (.A2(_0219_),
    .A1(net131),
    .B1(_0234_),
    .X(_0047_));
 sg13g2_xnor2_1 _0807_ (.Y(_0235_),
    .A(net160),
    .B(_0189_));
 sg13g2_nand2_1 _0808_ (.Y(_0236_),
    .A(net160),
    .B(_0219_));
 sg13g2_o21ai_1 _0809_ (.B1(_0236_),
    .Y(_0048_),
    .A1(_0221_),
    .A2(_0235_));
 sg13g2_a21oi_1 _0810_ (.A1(\main.dit_timer.timer[6] ),
    .A2(_0189_),
    .Y(_0237_),
    .B1(net109));
 sg13g2_or2_1 _0811_ (.X(_0238_),
    .B(_0237_),
    .A(_0190_));
 sg13g2_nand2_1 _0812_ (.Y(_0239_),
    .A(net109),
    .B(_0219_));
 sg13g2_o21ai_1 _0813_ (.B1(_0239_),
    .Y(_0049_),
    .A1(_0221_),
    .A2(_0238_));
 sg13g2_nor2_1 _0814_ (.A(_0191_),
    .B(_0218_),
    .Y(_0240_));
 sg13g2_xnor2_1 _0815_ (.Y(_0241_),
    .A(net241),
    .B(_0240_));
 sg13g2_nor2_1 _0816_ (.A(_0216_),
    .B(_0241_),
    .Y(_0050_));
 sg13g2_a21oi_1 _0817_ (.A1(\main.dit_timer.timer[8] ),
    .A2(_0240_),
    .Y(_0242_),
    .B1(net112));
 sg13g2_nand2_1 _0818_ (.Y(_0243_),
    .A(\main.dit_timer.timer[8] ),
    .B(net112));
 sg13g2_nor3_2 _0819_ (.A(_0191_),
    .B(_0218_),
    .C(_0243_),
    .Y(_0244_));
 sg13g2_nor3_1 _0820_ (.A(_0216_),
    .B(net113),
    .C(_0244_),
    .Y(_0051_));
 sg13g2_or2_1 _0821_ (.X(_0245_),
    .B(_0244_),
    .A(net273));
 sg13g2_nand2_1 _0822_ (.Y(_0246_),
    .A(net273),
    .B(_0244_));
 sg13g2_and4_1 _0823_ (.A(_0185_),
    .B(_0197_),
    .C(_0245_),
    .D(_0246_),
    .X(_0052_));
 sg13g2_xor2_1 _0824_ (.B(_0246_),
    .A(net223),
    .X(_0247_));
 sg13g2_nor2_1 _0825_ (.A(_0216_),
    .B(net224),
    .Y(_0053_));
 sg13g2_nand2_1 _0826_ (.Y(_0248_),
    .A(net98),
    .B(\main.dit_timer.morse_i ));
 sg13g2_nand2_2 _0827_ (.Y(_0249_),
    .A(_0198_),
    .B(_0248_));
 sg13g2_a21oi_2 _0828_ (.B1(_0184_),
    .Y(_0250_),
    .A2(_0248_),
    .A1(_0198_));
 sg13g2_mux2_1 _0829_ (.A0(net60),
    .A1(_0185_),
    .S(_0249_),
    .X(_0054_));
 sg13g2_nand2_1 _0830_ (.Y(_0251_),
    .A(net60),
    .B(_0250_));
 sg13g2_o21ai_1 _0831_ (.B1(net61),
    .Y(_0055_),
    .A1(_0135_),
    .A2(_0249_));
 sg13g2_nand2_1 _0832_ (.Y(_0252_),
    .A(net82),
    .B(_0250_));
 sg13g2_o21ai_1 _0833_ (.B1(net83),
    .Y(_0056_),
    .A1(_0136_),
    .A2(_0249_));
 sg13g2_nand2_1 _0834_ (.Y(_0253_),
    .A(net67),
    .B(_0250_));
 sg13g2_o21ai_1 _0835_ (.B1(net68),
    .Y(_0057_),
    .A1(_0137_),
    .A2(_0249_));
 sg13g2_nand2_1 _0836_ (.Y(_0254_),
    .A(net79),
    .B(_0250_));
 sg13g2_o21ai_1 _0837_ (.B1(net80),
    .Y(_0058_),
    .A1(_0138_),
    .A2(_0249_));
 sg13g2_nand2_1 _0838_ (.Y(_0255_),
    .A(net73),
    .B(_0250_));
 sg13g2_o21ai_1 _0839_ (.B1(net74),
    .Y(_0059_),
    .A1(_0134_),
    .A2(_0249_));
 sg13g2_nor2b_1 _0840_ (.A(\main.dit_timer.div1.in_r ),
    .B_N(net31),
    .Y(_0256_));
 sg13g2_mux2_1 _0841_ (.A0(net39),
    .A1(net54),
    .S(_0256_),
    .X(_0060_));
 sg13g2_nor2b_1 _0842_ (.A(\main.dit_timer.div2.in_r ),
    .B_N(net39),
    .Y(_0257_));
 sg13g2_mux2_1 _0843_ (.A0(net33),
    .A1(net48),
    .S(_0257_),
    .X(_0061_));
 sg13g2_nor2b_1 _0844_ (.A(\main.dit_timer.div3.in_r ),
    .B_N(net33),
    .Y(_0258_));
 sg13g2_mux2_1 _0845_ (.A0(net32),
    .A1(net44),
    .S(_0258_),
    .X(_0062_));
 sg13g2_nor2b_1 _0846_ (.A(\main.dit_timer.div4.in_r ),
    .B_N(net32),
    .Y(_0259_));
 sg13g2_mux2_1 _0847_ (.A0(net37),
    .A1(net56),
    .S(_0259_),
    .X(_0063_));
 sg13g2_nor2b_1 _0848_ (.A(\main.dit_timer.div5.in_r ),
    .B_N(net37),
    .Y(_0260_));
 sg13g2_mux2_1 _0849_ (.A0(net35),
    .A1(net52),
    .S(_0260_),
    .X(_0064_));
 sg13g2_nor2b_1 _0850_ (.A(\main.dit_timer.div6.in_r ),
    .B_N(net35),
    .Y(_0261_));
 sg13g2_mux2_1 _0851_ (.A0(net30),
    .A1(net42),
    .S(_0261_),
    .X(_0065_));
 sg13g2_nor2b_1 _0852_ (.A(\main.dit_timer.div7.in_r ),
    .B_N(net30),
    .Y(_0262_));
 sg13g2_mux2_1 _0853_ (.A0(net34),
    .A1(net50),
    .S(_0262_),
    .X(_0066_));
 sg13g2_o21ai_1 _0854_ (.B1(net171),
    .Y(_0263_),
    .A1(net267),
    .A2(net194));
 sg13g2_o21ai_1 _0855_ (.B1(net268),
    .Y(_0067_),
    .A1(_0141_),
    .A2(net195));
 sg13g2_o21ai_1 _0856_ (.B1(net171),
    .Y(_0264_),
    .A1(net194),
    .A2(net188));
 sg13g2_o21ai_1 _0857_ (.B1(_0264_),
    .Y(_0068_),
    .A1(_0142_),
    .A2(net195));
 sg13g2_o21ai_1 _0858_ (.B1(net171),
    .Y(_0265_),
    .A1(net194),
    .A2(net186));
 sg13g2_o21ai_1 _0859_ (.B1(_0265_),
    .Y(_0069_),
    .A1(_0143_),
    .A2(net195));
 sg13g2_o21ai_1 _0860_ (.B1(net171),
    .Y(_0266_),
    .A1(net194),
    .A2(net182));
 sg13g2_o21ai_1 _0861_ (.B1(net272),
    .Y(_0070_),
    .A1(net173),
    .A2(net195));
 sg13g2_o21ai_1 _0862_ (.B1(net171),
    .Y(_0267_),
    .A1(net193),
    .A2(net180));
 sg13g2_o21ai_1 _0863_ (.B1(_0267_),
    .Y(_0071_),
    .A1(_0145_),
    .A2(net195));
 sg13g2_o21ai_1 _0864_ (.B1(_0208_),
    .Y(_0268_),
    .A1(net193),
    .A2(net176));
 sg13g2_o21ai_1 _0865_ (.B1(_0268_),
    .Y(_0072_),
    .A1(_0148_),
    .A2(net195));
 sg13g2_or2_1 _0866_ (.X(_0269_),
    .B(\main.db1.cnt[3] ),
    .A(\main.db1.cnt[2] ));
 sg13g2_nor2b_1 _0867_ (.A(\main.db1.cnt[5] ),
    .B_N(\main.db1.cnt[4] ),
    .Y(_0270_));
 sg13g2_nand2b_1 _0868_ (.Y(_0271_),
    .B(_0023_),
    .A_N(\main.db1.cnt[6] ));
 sg13g2_a21oi_1 _0869_ (.A1(_0269_),
    .A2(_0270_),
    .Y(_0272_),
    .B1(_0271_));
 sg13g2_o21ai_1 _0870_ (.B1(_0122_),
    .Y(_0273_),
    .A1(_0123_),
    .A2(_0272_));
 sg13g2_a21oi_1 _0871_ (.A1(\main.db1.cnt[9] ),
    .A2(_0273_),
    .Y(_0274_),
    .B1(net225));
 sg13g2_a21o_2 _0872_ (.A2(_0273_),
    .A1(\main.db1.cnt[9] ),
    .B1(\main.db1.cnt[10] ),
    .X(_0275_));
 sg13g2_or2_2 _0873_ (.X(_0276_),
    .B(\main.db1.sig_r[1] ),
    .A(\main.db1.sig_r[2] ));
 sg13g2_nand2_2 _0874_ (.Y(_0277_),
    .A(net143),
    .B(net41));
 sg13g2_nand2_1 _0875_ (.Y(_0278_),
    .A(_0276_),
    .B(_0277_));
 sg13g2_and4_2 _0876_ (.A(\main.db1.cnt[13] ),
    .B(\main.db1.cnt[12] ),
    .C(\main.db1.cnt[11] ),
    .D(net168),
    .X(_0279_));
 sg13g2_nand4_1 _0877_ (.B(\main.db1.cnt[12] ),
    .C(\main.db1.cnt[11] ),
    .A(\main.db1.cnt[13] ),
    .Y(_0280_),
    .D(net168));
 sg13g2_nor2_1 _0878_ (.A(net164),
    .B(net166),
    .Y(_0281_));
 sg13g2_nand2_1 _0879_ (.Y(_0282_),
    .A(_0275_),
    .B(_0279_));
 sg13g2_o21ai_1 _0880_ (.B1(\main.db1.cnt[0] ),
    .Y(_0283_),
    .A1(net164),
    .A2(net166));
 sg13g2_a22oi_1 _0881_ (.Y(_0284_),
    .B1(_0279_),
    .B2(_0275_),
    .A2(_0277_),
    .A1(_0276_));
 sg13g2_mux2_1 _0882_ (.A0(_0284_),
    .A1(_0281_),
    .S(net260),
    .X(_0073_));
 sg13g2_nand2_1 _0883_ (.Y(_0285_),
    .A(\main.db1.cnt[0] ),
    .B(net232));
 sg13g2_nand2_1 _0884_ (.Y(_0286_),
    .A(net168),
    .B(_0285_));
 sg13g2_o21ai_1 _0885_ (.B1(_0286_),
    .Y(_0287_),
    .A1(net164),
    .A2(net166));
 sg13g2_a22oi_1 _0886_ (.Y(_0074_),
    .B1(_0286_),
    .B2(_0282_),
    .A2(_0283_),
    .A1(_0146_));
 sg13g2_or2_1 _0887_ (.X(_0288_),
    .B(_0285_),
    .A(net227));
 sg13g2_a221oi_1 _0888_ (.B2(_0275_),
    .C1(_0288_),
    .B1(_0279_),
    .A1(_0276_),
    .Y(_0289_),
    .A2(_0277_));
 sg13g2_a21o_1 _0889_ (.A2(_0287_),
    .A1(net227),
    .B1(_0289_),
    .X(_0075_));
 sg13g2_and3_1 _0890_ (.X(_0290_),
    .A(\main.db1.cnt[2] ),
    .B(\main.db1.cnt[0] ),
    .C(\main.db1.cnt[1] ));
 sg13g2_and4_1 _0891_ (.A(\main.db1.cnt[2] ),
    .B(net99),
    .C(\main.db1.cnt[0] ),
    .D(\main.db1.cnt[1] ),
    .X(_0291_));
 sg13g2_a21o_1 _0892_ (.A2(_0277_),
    .A1(_0276_),
    .B1(_0291_),
    .X(_0292_));
 sg13g2_o21ai_1 _0893_ (.B1(_0292_),
    .Y(_0293_),
    .A1(net164),
    .A2(net166));
 sg13g2_o21ai_1 _0894_ (.B1(_0290_),
    .Y(_0294_),
    .A1(_0274_),
    .A2(_0280_));
 sg13g2_a22oi_1 _0895_ (.Y(_0076_),
    .B1(_0294_),
    .B2(_0125_),
    .A2(_0292_),
    .A1(net162));
 sg13g2_nand2b_1 _0896_ (.Y(_0295_),
    .B(_0291_),
    .A_N(net235));
 sg13g2_a221oi_1 _0897_ (.B2(_0275_),
    .C1(_0295_),
    .B1(_0279_),
    .A1(_0276_),
    .Y(_0296_),
    .A2(_0277_));
 sg13g2_a21o_1 _0898_ (.A2(_0293_),
    .A1(net235),
    .B1(_0296_),
    .X(_0077_));
 sg13g2_and3_1 _0899_ (.X(_0297_),
    .A(\main.db1.cnt[5] ),
    .B(_0275_),
    .C(_0279_));
 sg13g2_and2_1 _0900_ (.A(\main.db1.cnt[4] ),
    .B(_0291_),
    .X(_0298_));
 sg13g2_xnor2_1 _0901_ (.Y(_0299_),
    .A(net257),
    .B(_0298_));
 sg13g2_a21o_1 _0902_ (.A2(_0299_),
    .A1(_0284_),
    .B1(_0297_),
    .X(_0078_));
 sg13g2_and2_1 _0903_ (.A(\main.db1.cnt[5] ),
    .B(_0298_),
    .X(_0300_));
 sg13g2_nand4_1 _0904_ (.B(\main.db1.cnt[5] ),
    .C(\main.db1.cnt[4] ),
    .A(net96),
    .Y(_0301_),
    .D(_0291_));
 sg13g2_nand2_1 _0905_ (.Y(_0302_),
    .A(net168),
    .B(_0301_));
 sg13g2_o21ai_1 _0906_ (.B1(_0302_),
    .Y(_0303_),
    .A1(net164),
    .A2(net166));
 sg13g2_o21ai_1 _0907_ (.B1(_0300_),
    .Y(_0304_),
    .A1(net164),
    .A2(net166));
 sg13g2_a22oi_1 _0908_ (.Y(_0079_),
    .B1(_0304_),
    .B2(_0124_),
    .A2(_0302_),
    .A1(net162));
 sg13g2_nand2b_1 _0909_ (.Y(_0305_),
    .B(_0123_),
    .A_N(_0301_));
 sg13g2_a221oi_1 _0910_ (.B2(_0275_),
    .C1(_0305_),
    .B1(_0279_),
    .A1(_0276_),
    .Y(_0306_),
    .A2(_0277_));
 sg13g2_a21o_1 _0911_ (.A2(_0303_),
    .A1(net125),
    .B1(_0306_),
    .X(_0080_));
 sg13g2_nor2_1 _0912_ (.A(_0123_),
    .B(_0301_),
    .Y(_0307_));
 sg13g2_nor3_2 _0913_ (.A(_0122_),
    .B(_0123_),
    .C(_0301_),
    .Y(_0308_));
 sg13g2_or3_1 _0914_ (.A(_0122_),
    .B(_0123_),
    .C(_0301_),
    .X(_0309_));
 sg13g2_nand2_1 _0915_ (.Y(_0310_),
    .A(net168),
    .B(_0309_));
 sg13g2_o21ai_1 _0916_ (.B1(_0310_),
    .Y(_0311_),
    .A1(net164),
    .A2(net166));
 sg13g2_o21ai_1 _0917_ (.B1(_0307_),
    .Y(_0312_),
    .A1(net164),
    .A2(net166));
 sg13g2_a22oi_1 _0918_ (.Y(_0081_),
    .B1(_0312_),
    .B2(_0122_),
    .A2(_0310_),
    .A1(net162));
 sg13g2_nand2b_1 _0919_ (.Y(_0313_),
    .B(_0308_),
    .A_N(net253));
 sg13g2_a221oi_1 _0920_ (.B2(_0275_),
    .C1(_0313_),
    .B1(_0279_),
    .A1(_0276_),
    .Y(_0314_),
    .A2(_0277_));
 sg13g2_a21o_1 _0921_ (.A2(_0311_),
    .A1(net253),
    .B1(_0314_),
    .X(_0082_));
 sg13g2_and2_1 _0922_ (.A(\main.db1.cnt[9] ),
    .B(_0308_),
    .X(_0315_));
 sg13g2_nand3_1 _0923_ (.B(\main.db1.cnt[9] ),
    .C(_0308_),
    .A(net225),
    .Y(_0316_));
 sg13g2_nand2_1 _0924_ (.Y(_0317_),
    .A(net168),
    .B(_0316_));
 sg13g2_o21ai_1 _0925_ (.B1(_0315_),
    .Y(_0318_),
    .A1(_0274_),
    .A2(_0280_));
 sg13g2_a22oi_1 _0926_ (.Y(_0083_),
    .B1(_0318_),
    .B2(_0121_),
    .A2(_0317_),
    .A1(net162));
 sg13g2_nor2b_1 _0927_ (.A(net249),
    .B_N(_0316_),
    .Y(_0319_));
 sg13g2_nand3_1 _0928_ (.B(net225),
    .C(\main.db1.cnt[9] ),
    .A(net249),
    .Y(_0320_));
 sg13g2_nor4_2 _0929_ (.A(_0122_),
    .B(_0123_),
    .C(_0301_),
    .Y(_0321_),
    .D(_0320_));
 sg13g2_o21ai_1 _0930_ (.B1(net168),
    .Y(_0322_),
    .A1(_0309_),
    .A2(_0320_));
 sg13g2_o21ai_1 _0931_ (.B1(net162),
    .Y(_0084_),
    .A1(net250),
    .A2(_0322_));
 sg13g2_and2_1 _0932_ (.A(net265),
    .B(_0321_),
    .X(_0323_));
 sg13g2_o21ai_1 _0933_ (.B1(net168),
    .Y(_0324_),
    .A1(net265),
    .A2(_0321_));
 sg13g2_o21ai_1 _0934_ (.B1(net162),
    .Y(_0085_),
    .A1(_0323_),
    .A2(_0324_));
 sg13g2_nor2_1 _0935_ (.A(net244),
    .B(_0323_),
    .Y(_0325_));
 sg13g2_nand3_1 _0936_ (.B(\main.db1.cnt[12] ),
    .C(_0321_),
    .A(net244),
    .Y(_0326_));
 sg13g2_nand2_1 _0937_ (.Y(_0327_),
    .A(_0278_),
    .B(_0326_));
 sg13g2_o21ai_1 _0938_ (.B1(net162),
    .Y(_0086_),
    .A1(net245),
    .A2(_0327_));
 sg13g2_nor2b_1 _0939_ (.A(_0028_),
    .B_N(net186),
    .Y(_0328_));
 sg13g2_nor2_2 _0940_ (.A(net188),
    .B(net185),
    .Y(_0329_));
 sg13g2_or2_1 _0941_ (.X(_0330_),
    .B(net185),
    .A(net188));
 sg13g2_o21ai_1 _0942_ (.B1(net178),
    .Y(_0331_),
    .A1(net188),
    .A2(net185));
 sg13g2_or2_1 _0943_ (.X(_0332_),
    .B(_0331_),
    .A(_0328_));
 sg13g2_nor2b_1 _0944_ (.A(net184),
    .B_N(net187),
    .Y(_0333_));
 sg13g2_nand2b_1 _0945_ (.Y(_0334_),
    .B(net187),
    .A_N(net183));
 sg13g2_nor2b_2 _0946_ (.A(net188),
    .B_N(net185),
    .Y(_0335_));
 sg13g2_nand2b_2 _0947_ (.Y(_0336_),
    .B(net185),
    .A_N(net189));
 sg13g2_a21oi_1 _0948_ (.A1(net184),
    .A2(_0336_),
    .Y(_0337_),
    .B1(_0333_));
 sg13g2_nor2_1 _0949_ (.A(net182),
    .B(_0329_),
    .Y(_0338_));
 sg13g2_mux2_1 _0950_ (.A0(_0329_),
    .A1(_0335_),
    .S(net181),
    .X(_0339_));
 sg13g2_nor2_1 _0951_ (.A(net178),
    .B(_0339_),
    .Y(_0340_));
 sg13g2_o21ai_1 _0952_ (.B1(_0332_),
    .Y(_0341_),
    .A1(net178),
    .A2(_0339_));
 sg13g2_nand2_1 _0953_ (.Y(_0342_),
    .A(\main.display.mask[0] ),
    .B(\main.display.mask[1] ));
 sg13g2_and3_1 _0954_ (.X(_0343_),
    .A(\main.display.mask[0] ),
    .B(\main.display.mask[1] ),
    .C(\main.display.mask[2] ));
 sg13g2_nand4_1 _0955_ (.B(\main.display.mask[1] ),
    .C(\main.display.mask[2] ),
    .A(\main.display.mask[0] ),
    .Y(_0344_),
    .D(\main.display.mask[3] ));
 sg13g2_nor3_1 _0956_ (.A(_0139_),
    .B(net193),
    .C(_0344_),
    .Y(_0345_));
 sg13g2_nor4_2 _0957_ (.A(_0139_),
    .B(net194),
    .C(\main.display.data[5] ),
    .Y(_0346_),
    .D(_0344_));
 sg13g2_nand2_1 _0958_ (.Y(_0347_),
    .A(net188),
    .B(net186));
 sg13g2_nor2_1 _0959_ (.A(net186),
    .B(net183),
    .Y(_0348_));
 sg13g2_or2_2 _0960_ (.X(_0349_),
    .B(net183),
    .A(net187));
 sg13g2_nor2_1 _0961_ (.A(net183),
    .B(net172),
    .Y(_0350_));
 sg13g2_nor2b_2 _0962_ (.A(net185),
    .B_N(net189),
    .Y(_0351_));
 sg13g2_nand2b_2 _0963_ (.Y(_0352_),
    .B(net189),
    .A_N(net185));
 sg13g2_nor2_1 _0964_ (.A(_0141_),
    .B(net178),
    .Y(_0353_));
 sg13g2_nand2b_2 _0965_ (.Y(_0354_),
    .B(net189),
    .A_N(net180));
 sg13g2_a21oi_1 _0966_ (.A1(_0349_),
    .A2(_0354_),
    .Y(_0355_),
    .B1(_0351_));
 sg13g2_o21ai_1 _0967_ (.B1(_0346_),
    .Y(_0356_),
    .A1(net177),
    .A2(_0355_));
 sg13g2_a21oi_1 _0968_ (.A1(net177),
    .A2(_0341_),
    .Y(_0357_),
    .B1(_0356_));
 sg13g2_nor3_2 _0969_ (.A(_0139_),
    .B(_0140_),
    .C(_0344_),
    .Y(_0358_));
 sg13g2_nand4_1 _0970_ (.B(\main.display.mask[4] ),
    .C(net193),
    .A(\main.display.mask[3] ),
    .Y(_0359_),
    .D(_0343_));
 sg13g2_nor2_1 _0971_ (.A(net183),
    .B(net173),
    .Y(_0360_));
 sg13g2_nand2b_1 _0972_ (.Y(_0361_),
    .B(net179),
    .A_N(net184));
 sg13g2_nand2b_1 _0973_ (.Y(_0362_),
    .B(net176),
    .A_N(\main.display.data[5] ));
 sg13g2_nor2_1 _0974_ (.A(_0336_),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_nor3_2 _0975_ (.A(_0336_),
    .B(_0361_),
    .C(_0362_),
    .Y(_0364_));
 sg13g2_nor2_2 _0976_ (.A(net176),
    .B(\main.display.data[5] ),
    .Y(_0365_));
 sg13g2_nand2b_2 _0977_ (.Y(_0366_),
    .B(net181),
    .A_N(net185));
 sg13g2_and4_1 _0978_ (.A(net184),
    .B(net179),
    .C(_0329_),
    .D(_0365_),
    .X(_0367_));
 sg13g2_nor2_1 _0979_ (.A(_0364_),
    .B(_0367_),
    .Y(_0368_));
 sg13g2_nand3_1 _0980_ (.B(\main.display.data[5] ),
    .C(_0360_),
    .A(net176),
    .Y(_0369_));
 sg13g2_o21ai_1 _0981_ (.B1(_0368_),
    .Y(_0370_),
    .A1(_0330_),
    .A2(_0369_));
 sg13g2_nand2_2 _0982_ (.Y(_0371_),
    .A(net189),
    .B(net180));
 sg13g2_nor3_1 _0983_ (.A(\main.display.data[4] ),
    .B(_0366_),
    .C(_0371_),
    .Y(_0372_));
 sg13g2_nand2b_2 _0984_ (.Y(_0373_),
    .B(\main.display.data[5] ),
    .A_N(net176));
 sg13g2_nor3_1 _0985_ (.A(_0366_),
    .B(_0371_),
    .C(_0373_),
    .Y(_0374_));
 sg13g2_nor3_1 _0986_ (.A(_0336_),
    .B(_0361_),
    .C(_0373_),
    .Y(_0375_));
 sg13g2_or2_1 _0987_ (.X(_0376_),
    .B(_0375_),
    .A(_0374_));
 sg13g2_o21ai_1 _0988_ (.B1(_0358_),
    .Y(_0377_),
    .A1(_0370_),
    .A2(_0376_));
 sg13g2_nor3_1 _0989_ (.A(\main.display.mask[3] ),
    .B(\main.display.mask[4] ),
    .C(net193),
    .Y(_0378_));
 sg13g2_or4_1 _0990_ (.A(\main.display.mask[2] ),
    .B(\main.display.mask[3] ),
    .C(\main.display.mask[4] ),
    .D(net193),
    .X(_0379_));
 sg13g2_nand2b_1 _0991_ (.Y(_0380_),
    .B(\main.display.mask[0] ),
    .A_N(\main.display.mask[1] ));
 sg13g2_or3_1 _0992_ (.A(net180),
    .B(net176),
    .C(\main.display.data[5] ),
    .X(_0381_));
 sg13g2_nor4_2 _0993_ (.A(_0349_),
    .B(_0379_),
    .C(_0380_),
    .Y(_0382_),
    .D(_0381_));
 sg13g2_a21oi_1 _0994_ (.A1(_0141_),
    .A2(_0382_),
    .Y(_0383_),
    .B1(net169));
 sg13g2_nor2_2 _0995_ (.A(net183),
    .B(net179),
    .Y(_0384_));
 sg13g2_nor4_2 _0996_ (.A(net183),
    .B(_0342_),
    .C(_0379_),
    .Y(_0385_),
    .D(_0381_));
 sg13g2_inv_1 _0997_ (.Y(_0386_),
    .A(_0385_));
 sg13g2_nor2_1 _0998_ (.A(_0335_),
    .B(_0386_),
    .Y(_0387_));
 sg13g2_nor2_2 _0999_ (.A(_0143_),
    .B(_0351_),
    .Y(_0388_));
 sg13g2_nand4_1 _1000_ (.B(_0343_),
    .C(_0365_),
    .A(net173),
    .Y(_0389_),
    .D(_0378_));
 sg13g2_a21o_1 _1001_ (.A2(_0388_),
    .A1(_0336_),
    .B1(_0389_),
    .X(_0390_));
 sg13g2_nor3_2 _1002_ (.A(\main.display.mask[4] ),
    .B(net193),
    .C(_0344_),
    .Y(_0391_));
 sg13g2_nand2b_1 _1003_ (.Y(_0392_),
    .B(net181),
    .A_N(_0029_));
 sg13g2_nor2_1 _1004_ (.A(_0143_),
    .B(net180),
    .Y(_0393_));
 sg13g2_o21ai_1 _1005_ (.B1(net173),
    .Y(_0394_),
    .A1(net181),
    .A2(_0336_));
 sg13g2_inv_1 _1006_ (.Y(_0395_),
    .A(_0394_));
 sg13g2_o21ai_1 _1007_ (.B1(_0383_),
    .Y(_0396_),
    .A1(_0338_),
    .A2(_0390_));
 sg13g2_nand2_2 _1008_ (.Y(_0397_),
    .A(_0365_),
    .B(_0391_));
 sg13g2_a221oi_1 _1009_ (.B2(_0395_),
    .C1(_0397_),
    .B1(_0392_),
    .A1(net178),
    .Y(_0398_),
    .A2(_0366_));
 sg13g2_nor4_2 _1010_ (.A(_0357_),
    .B(_0387_),
    .C(_0396_),
    .Y(_0399_),
    .D(_0398_));
 sg13g2_a22oi_1 _1011_ (.Y(_0087_),
    .B1(_0377_),
    .B2(_0399_),
    .A2(net170),
    .A1(_0150_));
 sg13g2_and2_1 _1012_ (.A(net177),
    .B(_0332_),
    .X(_0400_));
 sg13g2_mux2_1 _1013_ (.A0(net188),
    .A1(_0347_),
    .S(net182),
    .X(_0401_));
 sg13g2_a21oi_1 _1014_ (.A1(net178),
    .A2(_0401_),
    .Y(_0402_),
    .B1(net177));
 sg13g2_a22oi_1 _1015_ (.Y(_0403_),
    .B1(_0393_),
    .B2(_0347_),
    .A2(_0384_),
    .A1(_0030_));
 sg13g2_a22oi_1 _1016_ (.Y(_0404_),
    .B1(_0402_),
    .B2(_0403_),
    .A2(_0400_),
    .A1(_0394_));
 sg13g2_nand2b_1 _1017_ (.Y(_0405_),
    .B(_0346_),
    .A_N(_0404_));
 sg13g2_nand2_1 _1018_ (.Y(_0406_),
    .A(_0363_),
    .B(_0384_));
 sg13g2_nor3_1 _1019_ (.A(_0334_),
    .B(_0371_),
    .C(_0373_),
    .Y(_0407_));
 sg13g2_nor4_1 _1020_ (.A(_0364_),
    .B(_0367_),
    .C(_0374_),
    .D(_0407_),
    .Y(_0408_));
 sg13g2_a21oi_1 _1021_ (.A1(_0406_),
    .A2(_0408_),
    .Y(_0409_),
    .B1(_0359_));
 sg13g2_xnor2_1 _1022_ (.Y(_0410_),
    .A(net173),
    .B(_0337_));
 sg13g2_and4_1 _1023_ (.A(_0365_),
    .B(_0391_),
    .C(_0401_),
    .D(_0410_),
    .X(_0411_));
 sg13g2_a21oi_1 _1024_ (.A1(_0351_),
    .A2(_0385_),
    .Y(_0412_),
    .B1(net170));
 sg13g2_a21oi_2 _1025_ (.B1(net183),
    .Y(_0413_),
    .A2(net187),
    .A1(net189));
 sg13g2_a21o_1 _1026_ (.A2(net172),
    .A1(net184),
    .B1(_0413_),
    .X(_0414_));
 sg13g2_o21ai_1 _1027_ (.B1(_0412_),
    .Y(_0415_),
    .A1(_0389_),
    .A2(_0414_));
 sg13g2_nor3_1 _1028_ (.A(_0409_),
    .B(_0411_),
    .C(_0415_),
    .Y(_0416_));
 sg13g2_a22oi_1 _1029_ (.Y(_0088_),
    .B1(_0405_),
    .B2(_0416_),
    .A2(net170),
    .A1(_0151_));
 sg13g2_nor2_1 _1030_ (.A(net184),
    .B(_0335_),
    .Y(_0417_));
 sg13g2_o21ai_1 _1031_ (.B1(net173),
    .Y(_0418_),
    .A1(net182),
    .A2(_0335_));
 sg13g2_o21ai_1 _1032_ (.B1(net173),
    .Y(_0419_),
    .A1(net181),
    .A2(net172));
 sg13g2_a22oi_1 _1033_ (.Y(_0420_),
    .B1(_0419_),
    .B2(_0400_),
    .A2(_0418_),
    .A1(_0402_));
 sg13g2_nand2b_1 _1034_ (.Y(_0421_),
    .B(_0346_),
    .A_N(_0420_));
 sg13g2_nor4_1 _1035_ (.A(_0145_),
    .B(_0148_),
    .C(_0334_),
    .D(_0354_),
    .Y(_0422_));
 sg13g2_nor4_1 _1036_ (.A(_0364_),
    .B(_0374_),
    .C(_0375_),
    .D(_0422_),
    .Y(_0423_));
 sg13g2_nor2_1 _1037_ (.A(_0359_),
    .B(_0423_),
    .Y(_0424_));
 sg13g2_xnor2_1 _1038_ (.Y(_0425_),
    .A(_0354_),
    .B(_0388_));
 sg13g2_nor3_1 _1039_ (.A(_0335_),
    .B(_0397_),
    .C(_0425_),
    .Y(_0426_));
 sg13g2_a21oi_1 _1040_ (.A1(net172),
    .A2(_0385_),
    .Y(_0427_),
    .B1(net169));
 sg13g2_o21ai_1 _1041_ (.B1(_0427_),
    .Y(_0428_),
    .A1(_0333_),
    .A2(_0389_));
 sg13g2_nor3_1 _1042_ (.A(_0424_),
    .B(_0426_),
    .C(_0428_),
    .Y(_0429_));
 sg13g2_a22oi_1 _1043_ (.Y(_0089_),
    .B1(_0421_),
    .B2(_0429_),
    .A2(net170),
    .A1(_0152_));
 sg13g2_o21ai_1 _1044_ (.B1(net178),
    .Y(_0430_),
    .A1(_0028_),
    .A2(_0351_));
 sg13g2_o21ai_1 _1045_ (.B1(_0430_),
    .Y(_0431_),
    .A1(net178),
    .A2(_0337_));
 sg13g2_a21oi_1 _1046_ (.A1(net177),
    .A2(_0431_),
    .Y(_0432_),
    .B1(_0356_));
 sg13g2_o21ai_1 _1047_ (.B1(_0358_),
    .Y(_0433_),
    .A1(_0370_),
    .A2(_0372_));
 sg13g2_o21ai_1 _1048_ (.B1(_0366_),
    .Y(_0434_),
    .A1(_0333_),
    .A2(_0353_));
 sg13g2_a221oi_1 _1049_ (.B2(net172),
    .C1(_0397_),
    .B1(_0434_),
    .A1(_0352_),
    .Y(_0435_),
    .A2(_0384_));
 sg13g2_nor2_2 _1050_ (.A(net169),
    .B(_0382_),
    .Y(_0436_));
 sg13g2_inv_1 _1051_ (.Y(_0437_),
    .A(_0436_));
 sg13g2_nor2_1 _1052_ (.A(_0388_),
    .B(_0417_),
    .Y(_0438_));
 sg13g2_o21ai_1 _1053_ (.B1(_0436_),
    .Y(_0439_),
    .A1(_0389_),
    .A2(_0438_));
 sg13g2_nor3_1 _1054_ (.A(_0432_),
    .B(_0435_),
    .C(_0439_),
    .Y(_0440_));
 sg13g2_a22oi_1 _1055_ (.Y(_0090_),
    .B1(_0433_),
    .B2(_0440_),
    .A2(net169),
    .A1(_0153_));
 sg13g2_nand2_1 _1056_ (.Y(_0441_),
    .A(net177),
    .B(_0430_));
 sg13g2_a21oi_1 _1057_ (.A1(_0141_),
    .A2(_0366_),
    .Y(_0442_),
    .B1(net179));
 sg13g2_nor2_1 _1058_ (.A(net173),
    .B(_0336_),
    .Y(_0443_));
 sg13g2_nor3_1 _1059_ (.A(_0441_),
    .B(_0442_),
    .C(_0443_),
    .Y(_0444_));
 sg13g2_nand2_1 _1060_ (.Y(_0445_),
    .A(_0328_),
    .B(_0353_));
 sg13g2_a221oi_1 _1061_ (.B2(_0445_),
    .C1(\main.display.data[4] ),
    .B1(_0361_),
    .A1(net179),
    .Y(_0446_),
    .A2(net172));
 sg13g2_o21ai_1 _1062_ (.B1(_0346_),
    .Y(_0447_),
    .A1(_0444_),
    .A2(_0446_));
 sg13g2_a21oi_1 _1063_ (.A1(_0352_),
    .A2(_0417_),
    .Y(_0448_),
    .B1(_0389_));
 sg13g2_nand2_1 _1064_ (.Y(_0449_),
    .A(_0358_),
    .B(_0364_));
 sg13g2_o21ai_1 _1065_ (.B1(_0354_),
    .Y(_0450_),
    .A1(_0331_),
    .A2(_0413_));
 sg13g2_o21ai_1 _1066_ (.B1(_0449_),
    .Y(_0451_),
    .A1(_0397_),
    .A2(_0450_));
 sg13g2_nor4_1 _1067_ (.A(_0385_),
    .B(_0437_),
    .C(_0448_),
    .D(_0451_),
    .Y(_0452_));
 sg13g2_a22oi_1 _1068_ (.Y(_0091_),
    .B1(_0447_),
    .B2(_0452_),
    .A2(net169),
    .A1(_0154_));
 sg13g2_nand3_1 _1069_ (.B(_0348_),
    .C(_0371_),
    .A(_0145_),
    .Y(_0453_));
 sg13g2_o21ai_1 _1070_ (.B1(_0453_),
    .Y(_0454_),
    .A1(_0340_),
    .A2(_0441_));
 sg13g2_nand2_1 _1071_ (.Y(_0455_),
    .A(_0346_),
    .B(_0454_));
 sg13g2_a21oi_1 _1072_ (.A1(net172),
    .A2(_0413_),
    .Y(_0456_),
    .B1(_0390_));
 sg13g2_o21ai_1 _1073_ (.B1(_0436_),
    .Y(_0457_),
    .A1(_0352_),
    .A2(_0386_));
 sg13g2_nor2_1 _1074_ (.A(_0360_),
    .B(_0393_),
    .Y(_0458_));
 sg13g2_and3_1 _1075_ (.X(_0459_),
    .A(_0358_),
    .B(_0363_),
    .C(_0458_));
 sg13g2_a21o_1 _1076_ (.A2(_0413_),
    .A1(net172),
    .B1(_0388_),
    .X(_0460_));
 sg13g2_a221oi_1 _1077_ (.B2(net179),
    .C1(_0397_),
    .B1(_0460_),
    .A1(_0349_),
    .Y(_0461_),
    .A2(_0353_));
 sg13g2_nor4_1 _1078_ (.A(_0456_),
    .B(_0457_),
    .C(_0459_),
    .D(_0461_),
    .Y(_0462_));
 sg13g2_a22oi_1 _1079_ (.Y(_0092_),
    .B1(_0455_),
    .B2(_0462_),
    .A2(net169),
    .A1(_0155_));
 sg13g2_a21o_1 _1080_ (.A2(_0458_),
    .A1(_0347_),
    .B1(_0145_),
    .X(_0463_));
 sg13g2_nor3_1 _1081_ (.A(_0142_),
    .B(net180),
    .C(_0030_),
    .Y(_0464_));
 sg13g2_or4_1 _1082_ (.A(net177),
    .B(_0348_),
    .C(_0360_),
    .D(_0464_),
    .X(_0465_));
 sg13g2_nand4_1 _1083_ (.B(_0371_),
    .C(_0463_),
    .A(_0346_),
    .Y(_0466_),
    .D(_0465_));
 sg13g2_nor2_1 _1084_ (.A(net181),
    .B(_0029_),
    .Y(_0467_));
 sg13g2_a21oi_1 _1085_ (.A1(net181),
    .A2(_0336_),
    .Y(_0468_),
    .B1(_0467_));
 sg13g2_nor2_1 _1086_ (.A(_0389_),
    .B(_0468_),
    .Y(_0469_));
 sg13g2_o21ai_1 _1087_ (.B1(_0436_),
    .Y(_0470_),
    .A1(_0329_),
    .A2(_0386_));
 sg13g2_xnor2_1 _1088_ (.Y(_0471_),
    .A(net181),
    .B(_0351_));
 sg13g2_nor2_1 _1089_ (.A(_0144_),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_nor3_1 _1090_ (.A(_0397_),
    .B(_0442_),
    .C(_0472_),
    .Y(_0473_));
 sg13g2_nor3_1 _1091_ (.A(_0349_),
    .B(_0354_),
    .C(_0373_),
    .Y(_0474_));
 sg13g2_nor3_1 _1092_ (.A(_0364_),
    .B(_0367_),
    .C(_0474_),
    .Y(_0475_));
 sg13g2_nor2_1 _1093_ (.A(_0359_),
    .B(_0475_),
    .Y(_0476_));
 sg13g2_nor4_1 _1094_ (.A(_0469_),
    .B(_0470_),
    .C(_0473_),
    .D(_0476_),
    .Y(_0477_));
 sg13g2_a22oi_1 _1095_ (.Y(_0093_),
    .B1(_0466_),
    .B2(_0477_),
    .A2(net169),
    .A1(_0156_));
 sg13g2_nor2_1 _1096_ (.A(_0028_),
    .B(_0352_),
    .Y(_0478_));
 sg13g2_a22oi_1 _1097_ (.Y(_0479_),
    .B1(_0391_),
    .B2(_0478_),
    .A2(_0350_),
    .A1(_0345_));
 sg13g2_or4_1 _1098_ (.A(net176),
    .B(\main.display.data[5] ),
    .C(_0027_),
    .D(_0479_),
    .X(_0480_));
 sg13g2_nor3_1 _1099_ (.A(_0354_),
    .B(_0362_),
    .C(_0366_),
    .Y(_0481_));
 sg13g2_nor3_1 _1100_ (.A(_0407_),
    .B(_0422_),
    .C(_0481_),
    .Y(_0482_));
 sg13g2_o21ai_1 _1101_ (.B1(_0480_),
    .Y(_0483_),
    .A1(_0359_),
    .A2(_0482_));
 sg13g2_mux2_1 _1102_ (.A0(_0483_),
    .A1(net237),
    .S(net169),
    .X(_0094_));
 sg13g2_a21oi_1 _1103_ (.A1(_0119_),
    .A2(_0120_),
    .Y(_0095_),
    .B1(net92));
 sg13g2_nor2_1 _1104_ (.A(net88),
    .B(_0120_),
    .Y(_0484_));
 sg13g2_nor2_1 _1105_ (.A(\main.keyer.dah_count[1] ),
    .B(net191),
    .Y(_0485_));
 sg13g2_nor3_1 _1106_ (.A(_0172_),
    .B(net89),
    .C(_0485_),
    .Y(_0096_));
 sg13g2_or2_1 _1107_ (.X(_0486_),
    .B(\main.db0.cnt[3] ),
    .A(\main.db0.cnt[2] ));
 sg13g2_nor2b_1 _1108_ (.A(\main.db0.cnt[5] ),
    .B_N(\main.db0.cnt[4] ),
    .Y(_0487_));
 sg13g2_nand2b_1 _1109_ (.Y(_0488_),
    .B(_0024_),
    .A_N(\main.db0.cnt[6] ));
 sg13g2_a21oi_1 _1110_ (.A1(_0486_),
    .A2(_0487_),
    .Y(_0489_),
    .B1(_0488_));
 sg13g2_o21ai_1 _1111_ (.B1(_0128_),
    .Y(_0490_),
    .A1(_0129_),
    .A2(_0489_));
 sg13g2_a21oi_1 _1112_ (.A1(\main.db0.cnt[9] ),
    .A2(_0490_),
    .Y(_0491_),
    .B1(net147));
 sg13g2_a21o_2 _1113_ (.A2(_0490_),
    .A1(\main.db0.cnt[9] ),
    .B1(\main.db0.cnt[10] ),
    .X(_0492_));
 sg13g2_or2_2 _1114_ (.X(_0493_),
    .B(\main.db0.sig_r[1] ),
    .A(\main.db0.sig_r[2] ));
 sg13g2_nand2_2 _1115_ (.Y(_0494_),
    .A(net242),
    .B(net36));
 sg13g2_nand2_1 _1116_ (.Y(_0495_),
    .A(_0493_),
    .B(_0494_));
 sg13g2_and4_2 _1117_ (.A(\main.db0.cnt[13] ),
    .B(\main.db0.cnt[12] ),
    .C(\main.db0.cnt[11] ),
    .D(net167),
    .X(_0496_));
 sg13g2_nand4_1 _1118_ (.B(\main.db0.cnt[12] ),
    .C(\main.db0.cnt[11] ),
    .A(\main.db0.cnt[13] ),
    .Y(_0497_),
    .D(net167));
 sg13g2_nor2_1 _1119_ (.A(net163),
    .B(net165),
    .Y(_0498_));
 sg13g2_nand2_2 _1120_ (.Y(_0499_),
    .A(_0492_),
    .B(_0496_));
 sg13g2_o21ai_1 _1121_ (.B1(\main.db0.cnt[0] ),
    .Y(_0500_),
    .A1(_0491_),
    .A2(_0497_));
 sg13g2_a22oi_1 _1122_ (.Y(_0501_),
    .B1(_0496_),
    .B2(_0492_),
    .A2(_0494_),
    .A1(_0493_));
 sg13g2_mux2_1 _1123_ (.A0(_0501_),
    .A1(_0498_),
    .S(net259),
    .X(_0097_));
 sg13g2_nand2_1 _1124_ (.Y(_0502_),
    .A(\main.db0.cnt[0] ),
    .B(net161));
 sg13g2_nand2_1 _1125_ (.Y(_0503_),
    .A(_0495_),
    .B(_0502_));
 sg13g2_o21ai_1 _1126_ (.B1(_0503_),
    .Y(_0504_),
    .A1(net163),
    .A2(net165));
 sg13g2_a22oi_1 _1127_ (.Y(_0098_),
    .B1(_0503_),
    .B2(_0499_),
    .A2(_0500_),
    .A1(_0147_));
 sg13g2_or2_1 _1128_ (.X(_0505_),
    .B(_0502_),
    .A(net216));
 sg13g2_a221oi_1 _1129_ (.B2(_0492_),
    .C1(_0505_),
    .B1(_0496_),
    .A1(_0493_),
    .Y(_0506_),
    .A2(_0494_));
 sg13g2_a21o_1 _1130_ (.A2(_0504_),
    .A1(net216),
    .B1(_0506_),
    .X(_0099_));
 sg13g2_and3_1 _1131_ (.X(_0507_),
    .A(\main.db0.cnt[2] ),
    .B(\main.db0.cnt[0] ),
    .C(\main.db0.cnt[1] ));
 sg13g2_and4_1 _1132_ (.A(\main.db0.cnt[2] ),
    .B(net104),
    .C(\main.db0.cnt[0] ),
    .D(\main.db0.cnt[1] ),
    .X(_0508_));
 sg13g2_a21o_1 _1133_ (.A2(_0494_),
    .A1(_0493_),
    .B1(_0508_),
    .X(_0509_));
 sg13g2_o21ai_1 _1134_ (.B1(_0509_),
    .Y(_0510_),
    .A1(_0491_),
    .A2(_0497_));
 sg13g2_o21ai_1 _1135_ (.B1(_0507_),
    .Y(_0511_),
    .A1(net163),
    .A2(net165));
 sg13g2_a22oi_1 _1136_ (.Y(_0100_),
    .B1(_0511_),
    .B2(_0131_),
    .A2(_0509_),
    .A1(_0499_));
 sg13g2_nand2b_1 _1137_ (.Y(_0512_),
    .B(_0508_),
    .A_N(net239));
 sg13g2_a221oi_1 _1138_ (.B2(_0492_),
    .C1(_0512_),
    .B1(_0496_),
    .A1(_0493_),
    .Y(_0513_),
    .A2(_0494_));
 sg13g2_a21o_1 _1139_ (.A2(_0510_),
    .A1(net239),
    .B1(_0513_),
    .X(_0101_));
 sg13g2_and3_1 _1140_ (.X(_0514_),
    .A(\main.db0.cnt[5] ),
    .B(_0492_),
    .C(_0496_));
 sg13g2_and2_1 _1141_ (.A(\main.db0.cnt[4] ),
    .B(_0508_),
    .X(_0515_));
 sg13g2_xnor2_1 _1142_ (.Y(_0516_),
    .A(net261),
    .B(_0515_));
 sg13g2_a21o_1 _1143_ (.A2(_0516_),
    .A1(_0501_),
    .B1(_0514_),
    .X(_0102_));
 sg13g2_and2_1 _1144_ (.A(\main.db0.cnt[5] ),
    .B(_0515_),
    .X(_0517_));
 sg13g2_nand4_1 _1145_ (.B(\main.db0.cnt[5] ),
    .C(\main.db0.cnt[4] ),
    .A(net94),
    .Y(_0518_),
    .D(_0508_));
 sg13g2_nand2_1 _1146_ (.Y(_0519_),
    .A(net167),
    .B(_0518_));
 sg13g2_o21ai_1 _1147_ (.B1(_0519_),
    .Y(_0520_),
    .A1(net163),
    .A2(net165));
 sg13g2_o21ai_1 _1148_ (.B1(_0517_),
    .Y(_0521_),
    .A1(net163),
    .A2(net165));
 sg13g2_a22oi_1 _1149_ (.Y(_0103_),
    .B1(_0521_),
    .B2(_0130_),
    .A2(_0519_),
    .A1(_0499_));
 sg13g2_nand2b_1 _1150_ (.Y(_0522_),
    .B(_0129_),
    .A_N(_0518_));
 sg13g2_a221oi_1 _1151_ (.B2(_0492_),
    .C1(_0522_),
    .B1(_0496_),
    .A1(_0493_),
    .Y(_0523_),
    .A2(_0494_));
 sg13g2_a21o_1 _1152_ (.A2(_0520_),
    .A1(net156),
    .B1(_0523_),
    .X(_0104_));
 sg13g2_nor2_1 _1153_ (.A(_0129_),
    .B(_0518_),
    .Y(_0524_));
 sg13g2_nor3_2 _1154_ (.A(_0128_),
    .B(_0129_),
    .C(_0518_),
    .Y(_0525_));
 sg13g2_or3_1 _1155_ (.A(_0128_),
    .B(_0129_),
    .C(_0518_),
    .X(_0526_));
 sg13g2_nand2_1 _1156_ (.Y(_0527_),
    .A(net167),
    .B(_0526_));
 sg13g2_o21ai_1 _1157_ (.B1(_0527_),
    .Y(_0528_),
    .A1(net163),
    .A2(net165));
 sg13g2_o21ai_1 _1158_ (.B1(_0524_),
    .Y(_0529_),
    .A1(net163),
    .A2(net165));
 sg13g2_a22oi_1 _1159_ (.Y(_0105_),
    .B1(_0529_),
    .B2(_0128_),
    .A2(_0527_),
    .A1(_0499_));
 sg13g2_nand2b_1 _1160_ (.Y(_0530_),
    .B(_0525_),
    .A_N(net251));
 sg13g2_a221oi_1 _1161_ (.B2(_0492_),
    .C1(_0530_),
    .B1(_0496_),
    .A1(_0493_),
    .Y(_0531_),
    .A2(_0494_));
 sg13g2_a21o_1 _1162_ (.A2(_0528_),
    .A1(net251),
    .B1(_0531_),
    .X(_0106_));
 sg13g2_and2_1 _1163_ (.A(\main.db0.cnt[9] ),
    .B(_0525_),
    .X(_0532_));
 sg13g2_nand3_1 _1164_ (.B(\main.db0.cnt[9] ),
    .C(_0525_),
    .A(net147),
    .Y(_0533_));
 sg13g2_nand2_1 _1165_ (.Y(_0534_),
    .A(net167),
    .B(_0533_));
 sg13g2_o21ai_1 _1166_ (.B1(_0532_),
    .Y(_0535_),
    .A1(net163),
    .A2(net165));
 sg13g2_a22oi_1 _1167_ (.Y(_0107_),
    .B1(_0535_),
    .B2(_0127_),
    .A2(_0534_),
    .A1(_0499_));
 sg13g2_nor2b_1 _1168_ (.A(net247),
    .B_N(_0533_),
    .Y(_0536_));
 sg13g2_nand3_1 _1169_ (.B(net147),
    .C(net278),
    .A(net247),
    .Y(_0537_));
 sg13g2_nor4_2 _1170_ (.A(_0128_),
    .B(_0129_),
    .C(_0518_),
    .Y(_0538_),
    .D(_0537_));
 sg13g2_o21ai_1 _1171_ (.B1(net167),
    .Y(_0539_),
    .A1(_0526_),
    .A2(_0537_));
 sg13g2_o21ai_1 _1172_ (.B1(_0499_),
    .Y(_0108_),
    .A1(net248),
    .A2(_0539_));
 sg13g2_and2_1 _1173_ (.A(net266),
    .B(_0538_),
    .X(_0540_));
 sg13g2_o21ai_1 _1174_ (.B1(net167),
    .Y(_0541_),
    .A1(net266),
    .A2(_0538_));
 sg13g2_o21ai_1 _1175_ (.B1(_0499_),
    .Y(_0109_),
    .A1(_0540_),
    .A2(_0541_));
 sg13g2_nor2_1 _1176_ (.A(net254),
    .B(_0540_),
    .Y(_0542_));
 sg13g2_nand3_1 _1177_ (.B(\main.db0.cnt[12] ),
    .C(_0538_),
    .A(net254),
    .Y(_0543_));
 sg13g2_nand2_1 _1178_ (.Y(_0544_),
    .A(net167),
    .B(_0543_));
 sg13g2_o21ai_1 _1179_ (.B1(_0499_),
    .Y(_0110_),
    .A1(net255),
    .A2(_0544_));
 sg13g2_mux2_1 _1180_ (.A0(net143),
    .A1(net175),
    .S(net162),
    .X(_0111_));
 sg13g2_mux2_1 _1181_ (.A0(net87),
    .A1(net242),
    .S(_0498_),
    .X(_0112_));
 sg13g2_a21o_1 _1182_ (.A2(net63),
    .A1(net174),
    .B1(_0203_),
    .X(_0113_));
 sg13g2_a22oi_1 _1183_ (.Y(_0545_),
    .B1(_0203_),
    .B2(net63),
    .A2(\main.encoder.low_ct[1] ),
    .A1(net174));
 sg13g2_inv_1 _1184_ (.Y(_0114_),
    .A(net64));
 sg13g2_a22oi_1 _1185_ (.Y(_0546_),
    .B1(_0203_),
    .B2(net103),
    .A2(net76),
    .A1(net174));
 sg13g2_inv_1 _1186_ (.Y(_0115_),
    .A(_0546_));
 sg13g2_a22oi_1 _1187_ (.Y(_0547_),
    .B1(_0203_),
    .B2(net76),
    .A2(\main.encoder.low_ct[3] ),
    .A1(net174));
 sg13g2_inv_1 _1188_ (.Y(_0116_),
    .A(net77));
 sg13g2_a22oi_1 _1189_ (.Y(_0548_),
    .B1(_0203_),
    .B2(net78),
    .A2(net65),
    .A1(net174));
 sg13g2_inv_1 _1190_ (.Y(_0117_),
    .A(_0548_));
 sg13g2_a22oi_1 _1191_ (.Y(_0549_),
    .B1(_0203_),
    .B2(net65),
    .A2(\main.encoder.low_ct[5] ),
    .A1(net174));
 sg13g2_inv_1 _1192_ (.Y(_0118_),
    .A(net66));
 sg13g2_dfrbp_1 _1193_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net210),
    .D(_0032_),
    .Q_N(\main.keyer.current_state[0] ),
    .Q(_0031_));
 sg13g2_dfrbp_1 _1194_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net207),
    .D(_0000_),
    .Q_N(_0629_),
    .Q(\main.keyer.current_state[1] ));
 sg13g2_dfrbp_1 _1195_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net207),
    .D(_0001_),
    .Q_N(_0630_),
    .Q(\main.keyer.current_state[2] ));
 sg13g2_dfrbp_1 _1196_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net212),
    .D(_0002_),
    .Q_N(_0631_),
    .Q(\main.keyer.current_state[3] ));
 sg13g2_dfrbp_1 _1197_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net212),
    .D(net121),
    .Q_N(_0632_),
    .Q(\main.keyer.current_state[4] ));
 sg13g2_dfrbp_1 _1198_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net211),
    .D(_0004_),
    .Q_N(_0633_),
    .Q(\main.keyer.current_state[5] ));
 sg13g2_dfrbp_1 _1199_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net210),
    .D(_0005_),
    .Q_N(_0634_),
    .Q(\main.keyer.current_state[6] ));
 sg13g2_dfrbp_1 _1200_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net211),
    .D(net119),
    .Q_N(_0635_),
    .Q(\main.keyer.current_state[7] ));
 sg13g2_dfrbp_1 _1201_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net210),
    .D(net72),
    .Q_N(_0636_),
    .Q(\main.keyer.current_state[8] ));
 sg13g2_dfrbp_1 _1202_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net201),
    .D(net59),
    .Q_N(_0628_),
    .Q(\main.code_dit ));
 sg13g2_dfrbp_1 _1203_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net210),
    .D(_0033_),
    .Q_N(_0627_),
    .Q(\main.encoder.high_ct[0] ));
 sg13g2_dfrbp_1 _1204_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net210),
    .D(_0034_),
    .Q_N(_0637_),
    .Q(\main.encoder.high_ct[1] ));
 sg13g2_dfrbp_1 _1205_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net201),
    .D(net86),
    .Q_N(_0626_),
    .Q(\main.code_dah ));
 sg13g2_dfrbp_1 _1206_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net201),
    .D(net47),
    .Q_N(_0019_),
    .Q(\main.dit_timer.clk512 ));
 sg13g2_dfrbp_1 _1207_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net201),
    .D(_0022_),
    .Q_N(_0625_),
    .Q(\main.display.strobe_i ));
 sg13g2_dfrbp_1 _1208_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net198),
    .D(_0036_),
    .Q_N(_0624_),
    .Q(\main.display.mask[0] ));
 sg13g2_dfrbp_1 _1209_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net196),
    .D(_0037_),
    .Q_N(_0623_),
    .Q(\main.display.mask[1] ));
 sg13g2_dfrbp_1 _1210_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net196),
    .D(_0038_),
    .Q_N(_0622_),
    .Q(\main.display.mask[2] ));
 sg13g2_dfrbp_1 _1211_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net196),
    .D(_0039_),
    .Q_N(_0621_),
    .Q(\main.display.mask[3] ));
 sg13g2_dfrbp_1 _1212_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net196),
    .D(_0040_),
    .Q_N(_0620_),
    .Q(\main.display.mask[4] ));
 sg13g2_dfrbp_1 _1213_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net196),
    .D(_0041_),
    .Q_N(_0638_),
    .Q(\main.display.mask[5] ));
 sg13g2_dfrbp_1 _1214_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net17),
    .D(net38),
    .Q_N(_0619_),
    .Q(\main.dit_timer.last_clk512 ));
 sg13g2_dfrbp_1 _1215_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net211),
    .D(_0042_),
    .Q_N(_0618_),
    .Q(\main.dit_timer.timer[0] ));
 sg13g2_dfrbp_1 _1216_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net211),
    .D(net159),
    .Q_N(_0617_),
    .Q(\main.dit_timer.timer[1] ));
 sg13g2_dfrbp_1 _1217_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net211),
    .D(net102),
    .Q_N(_0616_),
    .Q(\main.dit_timer.timer[2] ));
 sg13g2_dfrbp_1 _1218_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net212),
    .D(net108),
    .Q_N(_0615_),
    .Q(\main.dit_timer.timer[3] ));
 sg13g2_dfrbp_1 _1219_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net213),
    .D(net116),
    .Q_N(_0026_),
    .Q(\main.dit_timer.timer[4] ));
 sg13g2_dfrbp_1 _1220_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net212),
    .D(_0047_),
    .Q_N(_0614_),
    .Q(\main.dit_timer.timer[5] ));
 sg13g2_dfrbp_1 _1221_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net212),
    .D(_0048_),
    .Q_N(_0613_),
    .Q(\main.dit_timer.timer[6] ));
 sg13g2_dfrbp_1 _1222_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net212),
    .D(net110),
    .Q_N(_0612_),
    .Q(\main.dit_timer.timer[7] ));
 sg13g2_dfrbp_1 _1223_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net212),
    .D(_0050_),
    .Q_N(_0611_),
    .Q(\main.dit_timer.timer[8] ));
 sg13g2_dfrbp_1 _1224_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net213),
    .D(net114),
    .Q_N(_0610_),
    .Q(\main.dit_timer.timer[9] ));
 sg13g2_dfrbp_1 _1225_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net213),
    .D(_0052_),
    .Q_N(_0609_),
    .Q(\main.dit_timer.timer[10] ));
 sg13g2_dfrbp_1 _1226_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net213),
    .D(_0053_),
    .Q_N(_0639_),
    .Q(\main.dit_timer.timer[11] ));
 sg13g2_dfrbp_1 _1227_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net209),
    .D(net264),
    .Q_N(_0640_),
    .Q(\main.dit_timer.timer_en ));
 sg13g2_dfrbp_1 _1228_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net211),
    .D(_0009_),
    .Q_N(_0641_),
    .Q(\main.dit_pulse ));
 sg13g2_dfrbp_1 _1229_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net196),
    .D(net28),
    .Q_N(_0011_),
    .Q(\main.dit_timer.clk2 ));
 sg13g2_dfrbp_1 _1230_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net209),
    .D(_0054_),
    .Q_N(_0608_),
    .Q(\main.dit_timer.pause_count[0] ));
 sg13g2_dfrbp_1 _1231_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net209),
    .D(net62),
    .Q_N(_0607_),
    .Q(\main.dit_timer.pause_count[1] ));
 sg13g2_dfrbp_1 _1232_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net209),
    .D(net84),
    .Q_N(_0606_),
    .Q(\main.dit_timer.pause_count[2] ));
 sg13g2_dfrbp_1 _1233_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net209),
    .D(net69),
    .Q_N(_0605_),
    .Q(\main.dit_timer.pause_count[3] ));
 sg13g2_dfrbp_1 _1234_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net209),
    .D(net81),
    .Q_N(_0604_),
    .Q(\main.dit_timer.pause_count[4] ));
 sg13g2_dfrbp_1 _1235_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net209),
    .D(net75),
    .Q_N(_0642_),
    .Q(\main.dit_timer.pause_count[5] ));
 sg13g2_dfrbp_1 _1236_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net196),
    .D(net31),
    .Q_N(_0603_),
    .Q(\main.dit_timer.div1.in_r ));
 sg13g2_dfrbp_1 _1237_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net196),
    .D(net55),
    .Q_N(_0012_),
    .Q(\main.dit_timer.clk4 ));
 sg13g2_dfrbp_1 _1238_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net197),
    .D(net39),
    .Q_N(_0602_),
    .Q(\main.dit_timer.div2.in_r ));
 sg13g2_dfrbp_1 _1239_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net197),
    .D(net49),
    .Q_N(_0013_),
    .Q(\main.dit_timer.clk8 ));
 sg13g2_dfrbp_1 _1240_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net197),
    .D(net33),
    .Q_N(_0601_),
    .Q(\main.dit_timer.div3.in_r ));
 sg13g2_dfrbp_1 _1241_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net197),
    .D(net45),
    .Q_N(_0014_),
    .Q(\main.dit_timer.clk16 ));
 sg13g2_dfrbp_1 _1242_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net197),
    .D(net32),
    .Q_N(_0600_),
    .Q(\main.dit_timer.div4.in_r ));
 sg13g2_dfrbp_1 _1243_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net197),
    .D(net57),
    .Q_N(_0015_),
    .Q(\main.dit_timer.clk32 ));
 sg13g2_dfrbp_1 _1244_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net197),
    .D(net37),
    .Q_N(_0599_),
    .Q(\main.dit_timer.div5.in_r ));
 sg13g2_dfrbp_1 _1245_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net200),
    .D(net53),
    .Q_N(_0016_),
    .Q(\main.dit_timer.clk64 ));
 sg13g2_dfrbp_1 _1246_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net199),
    .D(net35),
    .Q_N(_0598_),
    .Q(\main.dit_timer.div6.in_r ));
 sg13g2_dfrbp_1 _1247_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net199),
    .D(net43),
    .Q_N(_0017_),
    .Q(\main.dit_timer.clk128 ));
 sg13g2_dfrbp_1 _1248_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net199),
    .D(net30),
    .Q_N(_0597_),
    .Q(\main.dit_timer.div7.in_r ));
 sg13g2_dfrbp_1 _1249_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net199),
    .D(net51),
    .Q_N(_0018_),
    .Q(\main.dit_timer.clk256 ));
 sg13g2_dfrbp_1 _1250_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net198),
    .D(net34),
    .Q_N(_0596_),
    .Q(\main.dit_timer.div8.in_r ));
 sg13g2_dfrbp_1 _1251_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net203),
    .D(_0067_),
    .Q_N(_0030_),
    .Q(\main.display.data[0] ));
 sg13g2_dfrbp_1 _1252_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net203),
    .D(_0068_),
    .Q_N(_0029_),
    .Q(\main.display.data[1] ));
 sg13g2_dfrbp_1 _1253_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net203),
    .D(_0069_),
    .Q_N(_0028_),
    .Q(\main.display.data[2] ));
 sg13g2_dfrbp_1 _1254_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net203),
    .D(_0070_),
    .Q_N(_0027_),
    .Q(\main.display.data[3] ));
 sg13g2_dfrbp_1 _1255_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net201),
    .D(_0071_),
    .Q_N(_0595_),
    .Q(\main.display.data[4] ));
 sg13g2_dfrbp_1 _1256_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net201),
    .D(net275),
    .Q_N(_0594_),
    .Q(\main.display.data[5] ));
 sg13g2_dfrbp_1 _1257_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net205),
    .D(_0073_),
    .Q_N(_0593_),
    .Q(\main.db1.cnt[0] ));
 sg13g2_dfrbp_1 _1258_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net204),
    .D(net233),
    .Q_N(_0592_),
    .Q(\main.db1.cnt[1] ));
 sg13g2_dfrbp_1 _1259_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net204),
    .D(net228),
    .Q_N(_0591_),
    .Q(\main.db1.cnt[2] ));
 sg13g2_dfrbp_1 _1260_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net198),
    .D(net100),
    .Q_N(_0590_),
    .Q(\main.db1.cnt[3] ));
 sg13g2_dfrbp_1 _1261_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net199),
    .D(net236),
    .Q_N(_0589_),
    .Q(\main.db1.cnt[4] ));
 sg13g2_dfrbp_1 _1262_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net198),
    .D(net258),
    .Q_N(_0023_),
    .Q(\main.db1.cnt[5] ));
 sg13g2_dfrbp_1 _1263_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net198),
    .D(net97),
    .Q_N(_0588_),
    .Q(\main.db1.cnt[6] ));
 sg13g2_dfrbp_1 _1264_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net198),
    .D(net126),
    .Q_N(_0587_),
    .Q(\main.db1.cnt[7] ));
 sg13g2_dfrbp_1 _1265_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net198),
    .D(_0081_),
    .Q_N(_0586_),
    .Q(\main.db1.cnt[8] ));
 sg13g2_dfrbp_1 _1266_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net198),
    .D(_0082_),
    .Q_N(_0585_),
    .Q(\main.db1.cnt[9] ));
 sg13g2_dfrbp_1 _1267_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net204),
    .D(net226),
    .Q_N(_0584_),
    .Q(\main.db1.cnt[10] ));
 sg13g2_dfrbp_1 _1268_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net204),
    .D(_0084_),
    .Q_N(_0583_),
    .Q(\main.db1.cnt[11] ));
 sg13g2_dfrbp_1 _1269_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net204),
    .D(_0085_),
    .Q_N(_0582_),
    .Q(\main.db1.cnt[12] ));
 sg13g2_dfrbp_1 _1270_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net204),
    .D(net246),
    .Q_N(_0581_),
    .Q(\main.db1.cnt[13] ));
 sg13g2_dfrbp_1 _1271_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net202),
    .D(net142),
    .Q_N(_0580_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1272_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net202),
    .D(net155),
    .Q_N(_0579_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1273_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net201),
    .D(net150),
    .Q_N(_0578_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1274_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net201),
    .D(net220),
    .Q_N(_0577_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1275_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net202),
    .D(net128),
    .Q_N(_0576_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1276_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net203),
    .D(_0092_),
    .Q_N(_0575_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1277_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net203),
    .D(net230),
    .Q_N(_0574_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1278_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net202),
    .D(net238),
    .Q_N(_0643_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _1279_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net22),
    .D(_0008_),
    .Q_N(_0573_),
    .Q(\main.iambic_morse ));
 sg13g2_dfrbp_1 _1280_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net21),
    .D(net93),
    .Q_N(_0572_),
    .Q(\main.keyer.dah_count[0] ));
 sg13g2_dfrbp_1 _1281_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net19),
    .D(net90),
    .Q_N(_0644_),
    .Q(\main.keyer.dah_count[1] ));
 sg13g2_dfrbp_1 _1282_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net209),
    .D(net8),
    .Q_N(_0645_),
    .Q(\main.db1.sig_r[0] ));
 sg13g2_dfrbp_1 _1283_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net204),
    .D(net40),
    .Q_N(_0646_),
    .Q(\main.db1.sig_r[1] ));
 sg13g2_dfrbp_1 _1284_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net205),
    .D(net41),
    .Q_N(_0571_),
    .Q(\main.db1.sig_r[2] ));
 sg13g2_dfrbp_1 _1285_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net207),
    .D(_0097_),
    .Q_N(_0570_),
    .Q(\main.db0.cnt[0] ));
 sg13g2_dfrbp_1 _1286_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net206),
    .D(net215),
    .Q_N(_0569_),
    .Q(\main.db0.cnt[1] ));
 sg13g2_dfrbp_1 _1287_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net207),
    .D(net217),
    .Q_N(_0568_),
    .Q(\main.db0.cnt[2] ));
 sg13g2_dfrbp_1 _1288_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net207),
    .D(net105),
    .Q_N(_0567_),
    .Q(\main.db0.cnt[3] ));
 sg13g2_dfrbp_1 _1289_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net207),
    .D(net240),
    .Q_N(_0566_),
    .Q(\main.db0.cnt[4] ));
 sg13g2_dfrbp_1 _1290_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net207),
    .D(net262),
    .Q_N(_0024_),
    .Q(\main.db0.cnt[5] ));
 sg13g2_dfrbp_1 _1291_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net208),
    .D(net95),
    .Q_N(_0565_),
    .Q(\main.db0.cnt[6] ));
 sg13g2_dfrbp_1 _1292_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net206),
    .D(net157),
    .Q_N(_0564_),
    .Q(\main.db0.cnt[7] ));
 sg13g2_dfrbp_1 _1293_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net206),
    .D(net135),
    .Q_N(_0563_),
    .Q(\main.db0.cnt[8] ));
 sg13g2_dfrbp_1 _1294_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net206),
    .D(net252),
    .Q_N(_0562_),
    .Q(\main.db0.cnt[9] ));
 sg13g2_dfrbp_1 _1295_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net206),
    .D(net148),
    .Q_N(_0561_),
    .Q(\main.db0.cnt[10] ));
 sg13g2_dfrbp_1 _1296_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net206),
    .D(_0108_),
    .Q_N(_0560_),
    .Q(\main.db0.cnt[11] ));
 sg13g2_dfrbp_1 _1297_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net206),
    .D(_0109_),
    .Q_N(_0559_),
    .Q(\main.db0.cnt[12] ));
 sg13g2_dfrbp_1 _1298_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net206),
    .D(net256),
    .Q_N(_0558_),
    .Q(\main.db0.cnt[13] ));
 sg13g2_dfrbp_1 _1299_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net205),
    .D(_0111_),
    .Q_N(_0647_),
    .Q(\main.dah_r ));
 sg13g2_dfrbp_1 _1300_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net211),
    .D(net7),
    .Q_N(_0648_),
    .Q(\main.db0.sig_r[0] ));
 sg13g2_dfrbp_1 _1301_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net211),
    .D(net29),
    .Q_N(_0649_),
    .Q(\main.db0.sig_r[1] ));
 sg13g2_dfrbp_1 _1302_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net207),
    .D(net36),
    .Q_N(_0557_),
    .Q(\main.db0.sig_r[2] ));
 sg13g2_dfrbp_1 _1303_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net208),
    .D(_0112_),
    .Q_N(_0650_),
    .Q(\main.db0.sig_o ));
 sg13g2_dfrbp_1 _1304_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net23),
    .D(\main.dit_timer.morse_i ),
    .Q_N(_0025_),
    .Q(\main.aux_morse_o ));
 sg13g2_dfrbp_1 _1305_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net20),
    .D(net175),
    .Q_N(_0651_),
    .Q(\main.aux_dah_o ));
 sg13g2_dfrbp_1 _1306_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net18),
    .D(net87),
    .Q_N(_0556_),
    .Q(\main.aux_dit_o ));
 sg13g2_dfrbp_1 _1307_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net210),
    .D(_0113_),
    .Q_N(_0555_),
    .Q(\main.encoder.low_ct[0] ));
 sg13g2_dfrbp_1 _1308_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net210),
    .D(_0114_),
    .Q_N(_0554_),
    .Q(\main.encoder.low_ct[1] ));
 sg13g2_dfrbp_1 _1309_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net205),
    .D(_0115_),
    .Q_N(_0553_),
    .Q(\main.encoder.low_ct[2] ));
 sg13g2_dfrbp_1 _1310_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net205),
    .D(_0116_),
    .Q_N(_0552_),
    .Q(\main.encoder.low_ct[3] ));
 sg13g2_dfrbp_1 _1311_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net204),
    .D(_0117_),
    .Q_N(_0551_),
    .Q(\main.encoder.low_ct[4] ));
 sg13g2_dfrbp_1 _1312_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net210),
    .D(_0118_),
    .Q_N(_0550_),
    .Q(\main.encoder.low_ct[5] ));
 sg13g2_tiehi _1306__18 (.L_HI(net18));
 sg13g2_tiehi _1281__19 (.L_HI(net19));
 sg13g2_tiehi _1305__20 (.L_HI(net20));
 sg13g2_tiehi _1280__21 (.L_HI(net21));
 sg13g2_tiehi _1279__22 (.L_HI(net22));
 sg13g2_tiehi _1304__23 (.L_HI(net23));
 sg13g2_tiehi tt_um_betz_morse_keyer_24 (.L_HI(net24));
 sg13g2_tiehi tt_um_betz_morse_keyer_25 (.L_HI(net25));
 sg13g2_tiehi tt_um_betz_morse_keyer_26 (.L_HI(net26));
 sg13g2_tiehi tt_um_betz_morse_keyer_27 (.L_HI(net27));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_betz_morse_keyer_10 (.L_LO(net10));
 sg13g2_tielo tt_um_betz_morse_keyer_11 (.L_LO(net11));
 sg13g2_tielo tt_um_betz_morse_keyer_12 (.L_LO(net12));
 sg13g2_tielo tt_um_betz_morse_keyer_13 (.L_LO(net13));
 sg13g2_tielo tt_um_betz_morse_keyer_14 (.L_LO(net14));
 sg13g2_tielo tt_um_betz_morse_keyer_15 (.L_LO(net15));
 sg13g2_tielo tt_um_betz_morse_keyer_16 (.L_LO(net16));
 sg13g2_tiehi _1214__17 (.L_HI(net17));
 sg13g2_buf_1 _1332_ (.A(\main.aux_dit_o ),
    .X(uio_out[2]));
 sg13g2_buf_2 _1333_ (.A(\main.aux_dah_o ),
    .X(uio_out[3]));
 sg13g2_buf_1 _1334_ (.A(\main.aux_morse_o ),
    .X(uio_out[4]));
 sg13g2_buf_2 _1335_ (.A(\main.buzzer_o ),
    .X(uio_out[5]));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(_0282_));
 sg13g2_buf_2 fanout163 (.A(_0491_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_0274_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_0497_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_0280_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_0495_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_0278_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(net170),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_0209_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_0208_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_0330_),
    .X(net172));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(_0144_));
 sg13g2_buf_2 fanout174 (.A(_0120_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(net132),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(net177),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(\main.display.data[4] ),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(net179),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(net180),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(net277),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(net182),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(net276),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(\main.display.data[2] ),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(\main.display.data[2] ),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(net187),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(\main.display.data[1] ),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(net189),
    .X(net188));
 sg13g2_buf_4 fanout189 (.X(net189),
    .A(\main.display.data[0] ));
 sg13g2_buf_2 fanout190 (.A(net192),
    .X(net190));
 sg13g2_buf_1 fanout191 (.A(net192),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(net111),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(net194),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(net271),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(net138),
    .X(net195));
 sg13g2_buf_4 fanout196 (.X(net196),
    .A(net197));
 sg13g2_buf_4 fanout197 (.X(net197),
    .A(net200));
 sg13g2_buf_4 fanout198 (.X(net198),
    .A(net200));
 sg13g2_buf_2 fanout199 (.A(net200),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(rst_n),
    .X(net200));
 sg13g2_buf_4 fanout201 (.X(net201),
    .A(net203));
 sg13g2_buf_2 fanout202 (.A(net203),
    .X(net202));
 sg13g2_buf_4 fanout203 (.X(net203),
    .A(rst_n));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(net214));
 sg13g2_buf_2 fanout205 (.A(net214),
    .X(net205));
 sg13g2_buf_4 fanout206 (.X(net206),
    .A(net208));
 sg13g2_buf_4 fanout207 (.X(net207),
    .A(net208));
 sg13g2_buf_2 fanout208 (.A(net214),
    .X(net208));
 sg13g2_buf_4 fanout209 (.X(net209),
    .A(net213));
 sg13g2_buf_4 fanout210 (.X(net210),
    .A(net213));
 sg13g2_buf_4 fanout211 (.X(net211),
    .A(net212));
 sg13g2_buf_4 fanout212 (.X(net212),
    .A(net213));
 sg13g2_buf_4 fanout213 (.X(net213),
    .A(net214));
 sg13g2_buf_2 fanout214 (.A(rst_n),
    .X(net214));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[0]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_tielo tt_um_betz_morse_keyer_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0011_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold2 (.A(\main.db0.sig_r[0] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold3 (.A(\main.dit_timer.clk128 ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold4 (.A(\main.dit_timer.clk2 ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold5 (.A(\main.dit_timer.clk16 ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold6 (.A(\main.dit_timer.clk8 ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold7 (.A(\main.dit_timer.clk256 ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold8 (.A(\main.dit_timer.clk64 ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold9 (.A(\main.db0.sig_r[1] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold10 (.A(\main.dit_timer.clk32 ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold11 (.A(\main.dit_timer.clk512 ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold12 (.A(\main.dit_timer.clk4 ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold13 (.A(\main.db1.sig_r[0] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold14 (.A(\main.db1.sig_r[1] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0017_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0065_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0014_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0062_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0019_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0035_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0013_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0061_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0018_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0066_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0016_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0064_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0012_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0060_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0015_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0063_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold31 (.A(\main.encoder.high_ct[1] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0021_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold33 (.A(\main.dit_timer.pause_count[0] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0251_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0055_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold36 (.A(\main.encoder.low_ct[0] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0545_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold38 (.A(\main.encoder.low_ct[4] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0549_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold40 (.A(\main.dit_timer.pause_count[2] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0253_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0057_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold43 (.A(\main.keyer.current_state[0] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0182_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0007_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold46 (.A(\main.dit_timer.pause_count[4] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0255_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0059_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold49 (.A(\main.encoder.low_ct[2] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0547_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold51 (.A(\main.encoder.low_ct[3] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold52 (.A(\main.dit_timer.pause_count[3] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0254_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0058_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold55 (.A(\main.dit_timer.pause_count[1] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0252_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0056_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold58 (.A(\main.aux_morse_o ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0020_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold60 (.A(\main.db0.sig_o ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold61 (.A(\main.keyer.dah_count[0] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0484_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0096_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold64 (.A(\main.keyer.current_state[3] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0172_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0095_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold67 (.A(\main.db0.cnt[6] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0103_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold69 (.A(\main.db1.cnt[6] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0079_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0025_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold72 (.A(\main.db1.cnt[3] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0076_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold74 (.A(\main.dit_timer.timer[2] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0044_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold76 (.A(\main.encoder.low_ct[1] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold77 (.A(\main.db0.cnt[3] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0100_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold79 (.A(\main.encoder.high_ct[0] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold80 (.A(\main.dit_timer.timer[3] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0045_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold82 (.A(\main.dit_timer.timer[7] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0049_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold84 (.A(\main.dit_pulse ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold85 (.A(\main.dit_timer.timer[9] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0242_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0051_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold88 (.A(\main.dit_timer.timer[4] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0046_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold90 (.A(\main.keyer.dah_count[1] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold91 (.A(\main.keyer.current_state[7] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0006_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold93 (.A(\main.keyer.current_state[4] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0003_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold95 (.A(\main.keyer.current_state[6] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0177_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold97 (.A(\main.iambic_morse ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold98 (.A(\main.db1.cnt[7] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0080_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold100 (.A(uo_out[4]),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0091_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold102 (.A(\main.keyer.current_state[1] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0179_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold104 (.A(\main.dit_timer.timer[5] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold105 (.A(\main.dah_r ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold106 (.A(\main.db1.cnt[8] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold107 (.A(\main.db0.cnt[8] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0105_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold109 (.A(\main.display.mask[2] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0213_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold111 (.A(\main.display.strobe_i ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0210_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold113 (.A(\main.keyer.current_state[2] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold114 (.A(uo_out[0]),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0087_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold116 (.A(\main.db1.sig_r[2] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold117 (.A(uo_out[5]),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold118 (.A(\main.display.mask[1] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0212_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold120 (.A(\main.db0.cnt[10] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0107_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold122 (.A(uo_out[2]),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0089_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold124 (.A(\main.keyer.current_state[5] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold125 (.A(\main.display.mask[3] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0214_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold127 (.A(uo_out[1]),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0088_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold129 (.A(\main.db0.cnt[7] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0104_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold131 (.A(\main.dit_timer.timer[1] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0043_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold133 (.A(\main.dit_timer.timer[6] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold134 (.A(\main.db0.cnt[1] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0098_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold136 (.A(\main.db0.cnt[2] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0099_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold138 (.A(\main.keyer.current_state[8] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold139 (.A(uo_out[3]),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0090_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold141 (.A(\main.display.mask[0] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0211_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold143 (.A(\main.dit_timer.timer[11] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0247_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold145 (.A(\main.db1.cnt[10] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0083_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold147 (.A(\main.db1.cnt[2] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0075_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold149 (.A(uo_out[6]),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0093_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold151 (.A(\main.encoder.low_ct[5] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold152 (.A(\main.db1.cnt[1] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0074_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold154 (.A(\main.dit_timer.timer[0] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold155 (.A(\main.db1.cnt[4] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0077_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold157 (.A(uo_out[7]),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0094_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold159 (.A(\main.db0.cnt[4] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0101_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold161 (.A(\main.dit_timer.timer[8] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold162 (.A(\main.db0.sig_r[2] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold163 (.A(\main.display.mask[4] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold164 (.A(\main.db1.cnt[13] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0325_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0086_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold167 (.A(\main.db0.cnt[11] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0536_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold169 (.A(\main.db1.cnt[11] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0319_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold171 (.A(\main.db0.cnt[9] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0106_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold173 (.A(\main.db1.cnt[9] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold174 (.A(\main.db0.cnt[13] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0542_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0110_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0023_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0078_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold179 (.A(\main.db0.cnt[0] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold180 (.A(\main.db1.cnt[0] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0024_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0102_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold183 (.A(\main.dit_timer.pause_count[5] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0010_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold185 (.A(\main.db1.cnt[12] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold186 (.A(\main.db0.cnt[12] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold187 (.A(\main.code_dah ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0263_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold189 (.A(\main.dit_timer.timer[8] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0196_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold191 (.A(\main.display.mask[5] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0266_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold193 (.A(\main.dit_timer.timer[10] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold194 (.A(\main.display.data[5] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0072_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold196 (.A(\main.display.data[2] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold197 (.A(\main.display.data[3] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold198 (.A(\main.db0.cnt[9] ),
    .X(net278));
 sg13g2_antennanp ANTENNA_1 (.A(_0050_));
 sg13g2_antennanp ANTENNA_2 (.A(net7));
 sg13g2_antennanp ANTENNA_3 (.A(_0050_));
 sg13g2_antennanp ANTENNA_4 (.A(net7));
 sg13g2_antennanp ANTENNA_5 (.A(_0050_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_4 FILLER_7_368 ();
 sg13g2_fill_2 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_387 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_4 FILLER_8_336 ();
 sg13g2_fill_1 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_345 ();
 sg13g2_fill_2 FILLER_8_352 ();
 sg13g2_fill_1 FILLER_8_354 ();
 sg13g2_fill_1 FILLER_8_392 ();
 sg13g2_fill_1 FILLER_8_403 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_fill_1 FILLER_9_329 ();
 sg13g2_fill_2 FILLER_9_380 ();
 sg13g2_fill_1 FILLER_9_404 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_fill_1 FILLER_10_308 ();
 sg13g2_fill_1 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_4 FILLER_11_308 ();
 sg13g2_fill_1 FILLER_11_312 ();
 sg13g2_fill_1 FILLER_11_348 ();
 sg13g2_fill_2 FILLER_11_360 ();
 sg13g2_fill_1 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_4 FILLER_12_238 ();
 sg13g2_fill_2 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_248 ();
 sg13g2_decap_8 FILLER_12_255 ();
 sg13g2_decap_8 FILLER_12_262 ();
 sg13g2_decap_8 FILLER_12_269 ();
 sg13g2_decap_8 FILLER_12_276 ();
 sg13g2_decap_8 FILLER_12_283 ();
 sg13g2_decap_8 FILLER_12_290 ();
 sg13g2_decap_4 FILLER_12_297 ();
 sg13g2_fill_1 FILLER_12_301 ();
 sg13g2_fill_1 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_4 FILLER_13_224 ();
 sg13g2_fill_2 FILLER_13_228 ();
 sg13g2_fill_2 FILLER_13_240 ();
 sg13g2_fill_1 FILLER_13_242 ();
 sg13g2_fill_2 FILLER_13_273 ();
 sg13g2_fill_1 FILLER_13_275 ();
 sg13g2_decap_8 FILLER_13_281 ();
 sg13g2_decap_8 FILLER_13_288 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_fill_1 FILLER_14_175 ();
 sg13g2_decap_4 FILLER_14_180 ();
 sg13g2_fill_1 FILLER_14_184 ();
 sg13g2_fill_1 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_195 ();
 sg13g2_decap_8 FILLER_14_202 ();
 sg13g2_decap_8 FILLER_14_209 ();
 sg13g2_decap_8 FILLER_14_216 ();
 sg13g2_fill_1 FILLER_14_339 ();
 sg13g2_fill_2 FILLER_14_354 ();
 sg13g2_fill_2 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_fill_2 FILLER_15_168 ();
 sg13g2_fill_1 FILLER_15_179 ();
 sg13g2_fill_1 FILLER_15_185 ();
 sg13g2_fill_2 FILLER_15_212 ();
 sg13g2_fill_1 FILLER_15_236 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_4 FILLER_16_154 ();
 sg13g2_fill_1 FILLER_16_158 ();
 sg13g2_decap_4 FILLER_16_226 ();
 sg13g2_fill_2 FILLER_16_230 ();
 sg13g2_fill_1 FILLER_16_242 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_fill_2 FILLER_16_277 ();
 sg13g2_fill_1 FILLER_16_279 ();
 sg13g2_fill_1 FILLER_16_361 ();
 sg13g2_fill_1 FILLER_16_367 ();
 sg13g2_fill_2 FILLER_16_396 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_4 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_260 ();
 sg13g2_fill_1 FILLER_17_262 ();
 sg13g2_fill_2 FILLER_17_284 ();
 sg13g2_fill_1 FILLER_17_286 ();
 sg13g2_fill_1 FILLER_17_368 ();
 sg13g2_fill_1 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_fill_1 FILLER_18_161 ();
 sg13g2_decap_4 FILLER_18_167 ();
 sg13g2_fill_2 FILLER_18_171 ();
 sg13g2_fill_1 FILLER_18_182 ();
 sg13g2_fill_2 FILLER_18_213 ();
 sg13g2_decap_8 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_230 ();
 sg13g2_fill_2 FILLER_18_236 ();
 sg13g2_fill_1 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_4 FILLER_19_84 ();
 sg13g2_fill_2 FILLER_19_88 ();
 sg13g2_decap_4 FILLER_19_131 ();
 sg13g2_decap_8 FILLER_19_149 ();
 sg13g2_fill_2 FILLER_19_156 ();
 sg13g2_fill_1 FILLER_19_158 ();
 sg13g2_fill_1 FILLER_19_215 ();
 sg13g2_fill_2 FILLER_19_233 ();
 sg13g2_fill_1 FILLER_19_235 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_fill_2 FILLER_19_275 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_4 FILLER_20_84 ();
 sg13g2_fill_2 FILLER_20_88 ();
 sg13g2_fill_1 FILLER_20_134 ();
 sg13g2_fill_2 FILLER_20_161 ();
 sg13g2_fill_1 FILLER_20_163 ();
 sg13g2_fill_1 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_277 ();
 sg13g2_fill_1 FILLER_20_297 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_4 FILLER_21_77 ();
 sg13g2_fill_2 FILLER_21_81 ();
 sg13g2_fill_1 FILLER_21_114 ();
 sg13g2_decap_4 FILLER_21_124 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_170 ();
 sg13g2_fill_1 FILLER_21_216 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_fill_1 FILLER_21_275 ();
 sg13g2_fill_2 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_4 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_55 ();
 sg13g2_decap_4 FILLER_22_62 ();
 sg13g2_fill_2 FILLER_22_66 ();
 sg13g2_fill_2 FILLER_22_87 ();
 sg13g2_fill_2 FILLER_22_113 ();
 sg13g2_fill_1 FILLER_22_259 ();
 sg13g2_fill_2 FILLER_22_350 ();
 sg13g2_fill_1 FILLER_22_352 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_2 FILLER_23_61 ();
 sg13g2_fill_1 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_116 ();
 sg13g2_fill_1 FILLER_23_148 ();
 sg13g2_fill_2 FILLER_23_184 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_fill_2 FILLER_23_283 ();
 sg13g2_fill_1 FILLER_23_319 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_fill_2 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_4 FILLER_24_42 ();
 sg13g2_decap_4 FILLER_24_77 ();
 sg13g2_fill_2 FILLER_24_174 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_236 ();
 sg13g2_fill_1 FILLER_24_269 ();
 sg13g2_fill_1 FILLER_24_339 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_4 FILLER_25_68 ();
 sg13g2_fill_1 FILLER_25_106 ();
 sg13g2_fill_1 FILLER_25_183 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_fill_1 FILLER_25_340 ();
 sg13g2_fill_1 FILLER_25_352 ();
 sg13g2_fill_2 FILLER_25_372 ();
 sg13g2_fill_1 FILLER_25_393 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_4 FILLER_26_49 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_fill_2 FILLER_26_99 ();
 sg13g2_fill_1 FILLER_26_110 ();
 sg13g2_fill_1 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_142 ();
 sg13g2_fill_2 FILLER_26_209 ();
 sg13g2_fill_2 FILLER_26_237 ();
 sg13g2_decap_4 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_4 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_60 ();
 sg13g2_decap_4 FILLER_27_75 ();
 sg13g2_fill_1 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_141 ();
 sg13g2_fill_1 FILLER_27_154 ();
 sg13g2_fill_2 FILLER_27_189 ();
 sg13g2_fill_2 FILLER_27_229 ();
 sg13g2_fill_2 FILLER_27_239 ();
 sg13g2_fill_1 FILLER_27_241 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_fill_2 FILLER_27_319 ();
 sg13g2_fill_1 FILLER_27_340 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_4 FILLER_28_127 ();
 sg13g2_fill_2 FILLER_28_161 ();
 sg13g2_fill_2 FILLER_28_233 ();
 sg13g2_fill_1 FILLER_28_235 ();
 sg13g2_fill_1 FILLER_28_276 ();
 sg13g2_fill_1 FILLER_28_286 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_4 FILLER_29_56 ();
 sg13g2_fill_2 FILLER_29_60 ();
 sg13g2_fill_2 FILLER_29_99 ();
 sg13g2_fill_1 FILLER_29_136 ();
 sg13g2_fill_2 FILLER_29_186 ();
 sg13g2_fill_1 FILLER_29_278 ();
 sg13g2_fill_2 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_373 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_fill_2 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_74 ();
 sg13g2_fill_1 FILLER_30_114 ();
 sg13g2_decap_4 FILLER_30_125 ();
 sg13g2_fill_1 FILLER_30_134 ();
 sg13g2_fill_1 FILLER_30_154 ();
 sg13g2_fill_1 FILLER_30_316 ();
 sg13g2_fill_1 FILLER_30_334 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_4 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_53 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_fill_2 FILLER_31_112 ();
 sg13g2_fill_1 FILLER_31_125 ();
 sg13g2_fill_1 FILLER_31_148 ();
 sg13g2_fill_1 FILLER_31_188 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_201 ();
 sg13g2_fill_1 FILLER_31_263 ();
 sg13g2_fill_2 FILLER_31_289 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_71 ();
 sg13g2_fill_2 FILLER_32_75 ();
 sg13g2_fill_1 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_170 ();
 sg13g2_fill_1 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_188 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_fill_1 FILLER_32_250 ();
 sg13g2_fill_1 FILLER_32_349 ();
 sg13g2_fill_1 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_fill_2 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_30 ();
 sg13g2_decap_4 FILLER_33_70 ();
 sg13g2_fill_1 FILLER_33_90 ();
 sg13g2_fill_1 FILLER_33_104 ();
 sg13g2_fill_1 FILLER_33_132 ();
 sg13g2_fill_2 FILLER_33_260 ();
 sg13g2_fill_2 FILLER_33_271 ();
 sg13g2_fill_2 FILLER_33_327 ();
 sg13g2_fill_2 FILLER_33_334 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_fill_2 FILLER_34_56 ();
 sg13g2_fill_2 FILLER_34_65 ();
 sg13g2_fill_1 FILLER_34_73 ();
 sg13g2_fill_2 FILLER_34_81 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_fill_1 FILLER_34_99 ();
 sg13g2_fill_2 FILLER_34_109 ();
 sg13g2_fill_1 FILLER_34_138 ();
 sg13g2_fill_1 FILLER_34_149 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_194 ();
 sg13g2_fill_1 FILLER_34_215 ();
 sg13g2_fill_1 FILLER_34_259 ();
 sg13g2_fill_2 FILLER_34_296 ();
 sg13g2_fill_1 FILLER_34_312 ();
 sg13g2_fill_2 FILLER_34_362 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_4 FILLER_35_42 ();
 sg13g2_fill_2 FILLER_35_46 ();
 sg13g2_fill_1 FILLER_35_72 ();
 sg13g2_fill_1 FILLER_35_95 ();
 sg13g2_fill_1 FILLER_35_106 ();
 sg13g2_fill_1 FILLER_35_125 ();
 sg13g2_fill_2 FILLER_35_158 ();
 sg13g2_fill_1 FILLER_35_181 ();
 sg13g2_fill_2 FILLER_35_259 ();
 sg13g2_fill_1 FILLER_35_367 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_71 ();
 sg13g2_fill_1 FILLER_36_121 ();
 sg13g2_fill_1 FILLER_36_268 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_340 ();
 sg13g2_fill_2 FILLER_36_376 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_4 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_53 ();
 sg13g2_fill_2 FILLER_37_87 ();
 sg13g2_fill_2 FILLER_37_114 ();
 sg13g2_fill_1 FILLER_37_228 ();
 sg13g2_fill_1 FILLER_37_257 ();
 sg13g2_fill_1 FILLER_37_312 ();
 sg13g2_fill_2 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_44 ();
 sg13g2_fill_2 FILLER_38_77 ();
 sg13g2_fill_1 FILLER_38_109 ();
 sg13g2_fill_2 FILLER_38_139 ();
 sg13g2_fill_2 FILLER_38_219 ();
 sg13g2_fill_2 FILLER_38_270 ();
 sg13g2_fill_2 FILLER_38_349 ();
 sg13g2_fill_2 FILLER_38_377 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net24;
 assign uio_oe[3] = net25;
 assign uio_oe[4] = net26;
 assign uio_oe[5] = net27;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[0] = net13;
 assign uio_out[1] = net14;
 assign uio_out[6] = net15;
 assign uio_out[7] = net16;
endmodule

module tt_um_gregac_tiny_nn (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire clknet_leaf_0_clk;
 wire \u_tiny_nn_top.core_accumulate_result[0] ;
 wire \u_tiny_nn_top.core_accumulate_result[10] ;
 wire \u_tiny_nn_top.core_accumulate_result[11] ;
 wire \u_tiny_nn_top.core_accumulate_result[12] ;
 wire \u_tiny_nn_top.core_accumulate_result[13] ;
 wire \u_tiny_nn_top.core_accumulate_result[14] ;
 wire \u_tiny_nn_top.core_accumulate_result[15] ;
 wire \u_tiny_nn_top.core_accumulate_result[1] ;
 wire \u_tiny_nn_top.core_accumulate_result[2] ;
 wire \u_tiny_nn_top.core_accumulate_result[3] ;
 wire \u_tiny_nn_top.core_accumulate_result[4] ;
 wire \u_tiny_nn_top.core_accumulate_result[5] ;
 wire \u_tiny_nn_top.core_accumulate_result[6] ;
 wire \u_tiny_nn_top.core_accumulate_result[7] ;
 wire \u_tiny_nn_top.core_accumulate_result[8] ;
 wire \u_tiny_nn_top.core_accumulate_result[9] ;
 wire \u_tiny_nn_top.core_mul_add_op_b_en ;
 wire \u_tiny_nn_top.counter_q[0] ;
 wire \u_tiny_nn_top.counter_q[1] ;
 wire \u_tiny_nn_top.counter_q[2] ;
 wire \u_tiny_nn_top.counter_q[3] ;
 wire \u_tiny_nn_top.counter_q[4] ;
 wire \u_tiny_nn_top.counter_q[5] ;
 wire \u_tiny_nn_top.counter_q[6] ;
 wire \u_tiny_nn_top.counter_q[7] ;
 wire \u_tiny_nn_top.data_i_q[0] ;
 wire \u_tiny_nn_top.data_i_q[10] ;
 wire \u_tiny_nn_top.data_i_q[11] ;
 wire \u_tiny_nn_top.data_i_q[12] ;
 wire \u_tiny_nn_top.data_i_q[13] ;
 wire \u_tiny_nn_top.data_i_q[14] ;
 wire \u_tiny_nn_top.data_i_q[15] ;
 wire \u_tiny_nn_top.data_i_q[1] ;
 wire \u_tiny_nn_top.data_i_q[2] ;
 wire \u_tiny_nn_top.data_i_q[3] ;
 wire \u_tiny_nn_top.data_i_q[4] ;
 wire \u_tiny_nn_top.data_i_q[5] ;
 wire \u_tiny_nn_top.data_i_q[6] ;
 wire \u_tiny_nn_top.data_i_q[7] ;
 wire \u_tiny_nn_top.data_i_q[8] ;
 wire \u_tiny_nn_top.data_i_q[9] ;
 wire \u_tiny_nn_top.max_val_q[0] ;
 wire \u_tiny_nn_top.max_val_q[10] ;
 wire \u_tiny_nn_top.max_val_q[11] ;
 wire \u_tiny_nn_top.max_val_q[12] ;
 wire \u_tiny_nn_top.max_val_q[13] ;
 wire \u_tiny_nn_top.max_val_q[14] ;
 wire \u_tiny_nn_top.max_val_q[15] ;
 wire \u_tiny_nn_top.max_val_q[1] ;
 wire \u_tiny_nn_top.max_val_q[2] ;
 wire \u_tiny_nn_top.max_val_q[3] ;
 wire \u_tiny_nn_top.max_val_q[4] ;
 wire \u_tiny_nn_top.max_val_q[5] ;
 wire \u_tiny_nn_top.max_val_q[6] ;
 wire \u_tiny_nn_top.max_val_q[7] ;
 wire \u_tiny_nn_top.max_val_q[8] ;
 wire \u_tiny_nn_top.max_val_q[9] ;
 wire \u_tiny_nn_top.max_val_skid_q[0] ;
 wire \u_tiny_nn_top.max_val_skid_q[1] ;
 wire \u_tiny_nn_top.max_val_skid_q[2] ;
 wire \u_tiny_nn_top.max_val_skid_q[3] ;
 wire \u_tiny_nn_top.max_val_skid_q[4] ;
 wire \u_tiny_nn_top.max_val_skid_q[5] ;
 wire \u_tiny_nn_top.max_val_skid_q[6] ;
 wire \u_tiny_nn_top.max_val_skid_q[7] ;
 wire \u_tiny_nn_top.param_write_q[0] ;
 wire \u_tiny_nn_top.param_write_q[1] ;
 wire \u_tiny_nn_top.param_write_q[2] ;
 wire \u_tiny_nn_top.param_write_q[3] ;
 wire \u_tiny_nn_top.param_write_q[4] ;
 wire \u_tiny_nn_top.param_write_q[5] ;
 wire \u_tiny_nn_top.param_write_q[6] ;
 wire \u_tiny_nn_top.param_write_q[7] ;
 wire \u_tiny_nn_top.phase_q ;
 wire \u_tiny_nn_top.relu_q ;
 wire \u_tiny_nn_top.start_count_q[0] ;
 wire \u_tiny_nn_top.start_count_q[1] ;
 wire \u_tiny_nn_top.start_count_q[2] ;
 wire \u_tiny_nn_top.start_count_q[3] ;
 wire \u_tiny_nn_top.start_count_q[4] ;
 wire \u_tiny_nn_top.start_count_q[5] ;
 wire \u_tiny_nn_top.start_count_q[6] ;
 wire \u_tiny_nn_top.start_count_q[7] ;
 wire \u_tiny_nn_top.state_q[0] ;
 wire \u_tiny_nn_top.state_q[10] ;
 wire \u_tiny_nn_top.state_q[12] ;
 wire \u_tiny_nn_top.state_q[13] ;
 wire \u_tiny_nn_top.state_q[14] ;
 wire \u_tiny_nn_top.state_q[15] ;
 wire \u_tiny_nn_top.state_q[16] ;
 wire \u_tiny_nn_top.state_q[17] ;
 wire \u_tiny_nn_top.state_q[1] ;
 wire \u_tiny_nn_top.state_q[2] ;
 wire \u_tiny_nn_top.state_q[3] ;
 wire \u_tiny_nn_top.state_q[4] ;
 wire \u_tiny_nn_top.state_q[5] ;
 wire \u_tiny_nn_top.state_q[6] ;
 wire \u_tiny_nn_top.state_q[7] ;
 wire \u_tiny_nn_top.state_q[8] ;
 wire \u_tiny_nn_top.state_q[9] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][0] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][10] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][11] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][12] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][13] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][14] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][15] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][1] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][2] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][3] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][4] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][5] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][6] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][7] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][8] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[0][9] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][0] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][10] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][11] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][12] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][13] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][14] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][15] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][1] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][2] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][3] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][4] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][5] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][6] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][7] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][8] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_0_q[1][9] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][0] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][10] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][11] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][12] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][13] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][14] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][15] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][1] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][2] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][3] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][4] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][5] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][6] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][7] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][8] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[0][9] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][0] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][10] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][11] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][12] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][13] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][14] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][15] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][1] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][2] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][3] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][4] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][5] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][6] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][7] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][8] ;
 wire \u_tiny_nn_top.u_core.accumulate_level_1_q[1][9] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[0] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[10] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[11] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[12] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[13] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[14] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[15] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[1] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[2] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[3] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[4] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[5] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[6] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[7] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[8] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[9] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[0] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[10] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[11] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[12] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[13] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[14] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[15] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[1] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[2] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[3] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[4] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[5] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[6] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[7] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[8] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[9] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[0] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[10] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[11] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[12] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[13] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[14] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[15] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[1] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[2] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[3] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[4] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[5] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[6] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[7] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[8] ;
 wire \u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[9] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][0] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][10] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][11] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][12] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][13] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][14] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][15] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][1] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][2] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][3] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][4] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][5] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][6] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][7] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][8] ;
 wire \u_tiny_nn_top.u_core.mul_add_op_a_q[1][9] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][0] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][10] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][11] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][12] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][13] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][14] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][15] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][1] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][2] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][3] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][4] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][5] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][6] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][7] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][8] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[0][9] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][0] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][10] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][11] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][12] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][13] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][14] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][15] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][1] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][2] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][3] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][4] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][5] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][6] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][7] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][8] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[1][9] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][0] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][10] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][11] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][12] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][13] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][14] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][15] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][1] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][2] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][3] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][4] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][5] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][6] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][7] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][8] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[2][9] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][0] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][10] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][11] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][12] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][13] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][14] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][15] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][1] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][2] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][3] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][4] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][5] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][6] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][7] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][8] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[3][9] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][0] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][10] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][11] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][12] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][13] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][14] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][15] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][1] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][2] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][3] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][4] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][5] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][6] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][7] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][8] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[4][9] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][0] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][10] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][11] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][12] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][13] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][14] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][15] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][1] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][2] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][3] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][4] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][5] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][6] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][7] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][8] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[5][9] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][0] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][10] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][11] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][12] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][13] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][14] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][15] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][1] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][2] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][3] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][4] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][5] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][6] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][7] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][8] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[6][9] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][0] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][10] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][11] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][12] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][13] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][14] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][15] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][1] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][2] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][3] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][4] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][5] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][6] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][7] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][8] ;
 wire \u_tiny_nn_top.u_core.mul_val_op_q[7][9] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][0] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][10] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][11] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][12] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][13] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][14] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][15] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][1] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][2] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][3] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][4] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][5] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][6] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][7] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][8] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[0][9] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][0] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][10] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][11] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][12] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][13] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][14] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][15] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][1] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][2] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][3] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][4] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][5] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][6] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][7] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][8] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[1][9] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][0] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][10] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][11] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][12] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][13] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][14] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][15] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][1] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][2] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][3] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][4] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][5] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][6] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][7] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][8] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[2][9] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][0] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][10] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][11] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][12] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][13] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][14] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][15] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][1] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][2] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][3] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][4] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][5] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][6] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][7] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][8] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[3][9] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][0] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][10] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][11] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][12] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][13] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][14] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][15] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][1] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][2] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][3] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][4] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][5] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][6] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][7] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][8] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[4][9] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][0] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][10] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][11] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][12] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][13] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][14] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][15] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][1] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][2] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][3] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][4] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][5] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][6] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][7] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][8] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[5][9] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][0] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][10] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][11] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][12] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][13] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][14] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][15] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][1] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][2] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][3] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][4] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][5] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][6] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][7] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][8] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[6][9] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][0] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][10] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][11] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][12] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][13] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][14] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][15] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][1] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][2] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][3] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][4] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][5] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][6] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][7] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][8] ;
 wire \u_tiny_nn_top.u_core.param_val_op_q[7][9] ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;

 sg13g2_inv_1 _06099_ (.Y(_00638_),
    .A(net1827));
 sg13g2_inv_1 _06100_ (.Y(_00639_),
    .A(\u_tiny_nn_top.data_i_q[13] ));
 sg13g2_inv_1 _06101_ (.Y(_00640_),
    .A(net1828));
 sg13g2_inv_1 _06102_ (.Y(_00641_),
    .A(\u_tiny_nn_top.data_i_q[11] ));
 sg13g2_inv_2 _06103_ (.Y(_00642_),
    .A(\u_tiny_nn_top.data_i_q[10] ));
 sg13g2_inv_2 _06104_ (.Y(_00643_),
    .A(\u_tiny_nn_top.data_i_q[9] ));
 sg13g2_inv_2 _06105_ (.Y(_00644_),
    .A(net1831));
 sg13g2_inv_2 _06106_ (.Y(_00645_),
    .A(\u_tiny_nn_top.data_i_q[2] ));
 sg13g2_inv_2 _06107_ (.Y(_00646_),
    .A(\u_tiny_nn_top.data_i_q[0] ));
 sg13g2_inv_1 _06108_ (.Y(_00647_),
    .A(net1802));
 sg13g2_inv_1 _06109_ (.Y(_00648_),
    .A(net1809));
 sg13g2_inv_1 _06110_ (.Y(_00649_),
    .A(net1813));
 sg13g2_inv_1 _06111_ (.Y(_00650_),
    .A(net1818));
 sg13g2_inv_1 _06112_ (.Y(_00651_),
    .A(net1822));
 sg13g2_inv_1 _06113_ (.Y(_00652_),
    .A(net674));
 sg13g2_inv_1 _06114_ (.Y(_00653_),
    .A(net1855));
 sg13g2_inv_1 _06115_ (.Y(_00654_),
    .A(net1031));
 sg13g2_inv_2 _06116_ (.Y(_00655_),
    .A(net1103));
 sg13g2_inv_1 _06117_ (.Y(_00656_),
    .A(net1797));
 sg13g2_inv_1 _06118_ (.Y(_00657_),
    .A(\u_tiny_nn_top.state_q[15] ));
 sg13g2_inv_1 _06119_ (.Y(_00658_),
    .A(\u_tiny_nn_top.state_q[3] ));
 sg13g2_inv_1 _06120_ (.Y(_00659_),
    .A(net1788));
 sg13g2_inv_2 _06121_ (.Y(_00660_),
    .A(net1793));
 sg13g2_inv_1 _06122_ (.Y(_00661_),
    .A(net1789));
 sg13g2_inv_1 _06123_ (.Y(_00662_),
    .A(net491));
 sg13g2_inv_1 _06124_ (.Y(_00663_),
    .A(net1015));
 sg13g2_inv_1 _06125_ (.Y(_00664_),
    .A(\u_tiny_nn_top.max_val_q[3] ));
 sg13g2_inv_1 _06126_ (.Y(_00665_),
    .A(\u_tiny_nn_top.max_val_q[2] ));
 sg13g2_inv_1 _06127_ (.Y(_00666_),
    .A(\u_tiny_nn_top.max_val_q[5] ));
 sg13g2_inv_1 _06128_ (.Y(_00667_),
    .A(net1001));
 sg13g2_inv_1 _06129_ (.Y(_00668_),
    .A(\u_tiny_nn_top.max_val_q[8] ));
 sg13g2_inv_1 _06130_ (.Y(_00669_),
    .A(\u_tiny_nn_top.max_val_q[9] ));
 sg13g2_inv_1 _06131_ (.Y(_00670_),
    .A(\u_tiny_nn_top.max_val_q[13] ));
 sg13g2_inv_1 _06132_ (.Y(_00671_),
    .A(\u_tiny_nn_top.max_val_q[12] ));
 sg13g2_inv_1 _06133_ (.Y(_00672_),
    .A(_00017_));
 sg13g2_inv_1 _06134_ (.Y(_00673_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][15] ));
 sg13g2_inv_1 _06135_ (.Y(_00674_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][13] ));
 sg13g2_inv_2 _06136_ (.Y(_00675_),
    .A(_00019_));
 sg13g2_inv_2 _06137_ (.Y(_00676_),
    .A(net1102));
 sg13g2_inv_1 _06138_ (.Y(_00677_),
    .A(net1047));
 sg13g2_inv_1 _06139_ (.Y(_00678_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][13] ));
 sg13g2_inv_1 _06140_ (.Y(_00679_),
    .A(_00038_));
 sg13g2_inv_1 _06141_ (.Y(_00680_),
    .A(_00037_));
 sg13g2_inv_1 _06142_ (.Y(_00681_),
    .A(_00042_));
 sg13g2_inv_1 _06143_ (.Y(_00682_),
    .A(_00041_));
 sg13g2_inv_1 _06144_ (.Y(_00683_),
    .A(\u_tiny_nn_top.u_core.mul_val_op_q[2][0] ));
 sg13g2_inv_1 _06145_ (.Y(_00684_),
    .A(net892));
 sg13g2_inv_1 _06146_ (.Y(_00685_),
    .A(_00046_));
 sg13g2_inv_1 _06147_ (.Y(_00686_),
    .A(_00045_));
 sg13g2_inv_1 _06148_ (.Y(_00687_),
    .A(_00048_));
 sg13g2_inv_1 _06149_ (.Y(_00688_),
    .A(_00047_));
 sg13g2_inv_1 _06150_ (.Y(_00689_),
    .A(_00050_));
 sg13g2_inv_1 _06151_ (.Y(_00690_),
    .A(_00049_));
 sg13g2_inv_1 _06152_ (.Y(_00691_),
    .A(_00054_));
 sg13g2_inv_1 _06153_ (.Y(_00692_),
    .A(_00053_));
 sg13g2_inv_1 _06154_ (.Y(_00693_),
    .A(_00056_));
 sg13g2_inv_1 _06155_ (.Y(_00694_),
    .A(_00055_));
 sg13g2_inv_1 _06156_ (.Y(_00695_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[15] ));
 sg13g2_inv_1 _06157_ (.Y(_00696_),
    .A(net1084));
 sg13g2_inv_1 _06158_ (.Y(_00697_),
    .A(net1075));
 sg13g2_inv_1 _06159_ (.Y(_00698_),
    .A(net997));
 sg13g2_inv_1 _06160_ (.Y(_00699_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[12] ));
 sg13g2_inv_1 _06161_ (.Y(_00700_),
    .A(net1069));
 sg13g2_inv_2 _06162_ (.Y(_00701_),
    .A(net1005));
 sg13g2_inv_2 _06163_ (.Y(_00702_),
    .A(net1017));
 sg13g2_inv_2 _06164_ (.Y(_00703_),
    .A(_00072_));
 sg13g2_inv_1 _06165_ (.Y(_00704_),
    .A(_00075_));
 sg13g2_inv_1 _06166_ (.Y(_00705_),
    .A(net820));
 sg13g2_inv_1 _06167_ (.Y(_00706_),
    .A(net786));
 sg13g2_inv_1 _06168_ (.Y(_00707_),
    .A(net823));
 sg13g2_inv_1 _06169_ (.Y(_00708_),
    .A(net795));
 sg13g2_inv_1 _06170_ (.Y(_00709_),
    .A(net1100));
 sg13g2_inv_1 _06171_ (.Y(_00710_),
    .A(net691));
 sg13g2_inv_1 _06172_ (.Y(_00711_),
    .A(net832));
 sg13g2_inv_1 _06173_ (.Y(_00712_),
    .A(net815));
 sg13g2_inv_1 _06174_ (.Y(_00713_),
    .A(net811));
 sg13g2_inv_1 _06175_ (.Y(_00714_),
    .A(net841));
 sg13g2_inv_1 _06176_ (.Y(_00715_),
    .A(net771));
 sg13g2_inv_1 _06177_ (.Y(_00716_),
    .A(net794));
 sg13g2_inv_1 _06178_ (.Y(_00717_),
    .A(net956));
 sg13g2_inv_1 _06179_ (.Y(_00718_),
    .A(net887));
 sg13g2_inv_1 _06180_ (.Y(_00719_),
    .A(net734));
 sg13g2_inv_1 _06181_ (.Y(_00720_),
    .A(net798));
 sg13g2_inv_1 _06182_ (.Y(_00721_),
    .A(net930));
 sg13g2_inv_1 _06183_ (.Y(_00722_),
    .A(_00113_));
 sg13g2_inv_1 _06184_ (.Y(_00723_),
    .A(net1801));
 sg13g2_inv_1 _06185_ (.Y(_00724_),
    .A(net949));
 sg13g2_inv_1 _06186_ (.Y(_00725_),
    .A(net932));
 sg13g2_inv_1 _06187_ (.Y(_00726_),
    .A(net988));
 sg13g2_inv_1 _06188_ (.Y(_00727_),
    .A(net966));
 sg13g2_inv_1 _06189_ (.Y(_00728_),
    .A(net945));
 sg13g2_inv_1 _06190_ (.Y(_00729_),
    .A(net964));
 sg13g2_inv_1 _06191_ (.Y(_00730_),
    .A(net965));
 sg13g2_inv_1 _06192_ (.Y(_00731_),
    .A(net1034));
 sg13g2_inv_1 _06193_ (.Y(_00732_),
    .A(net1013));
 sg13g2_inv_1 _06194_ (.Y(_00733_),
    .A(net1049));
 sg13g2_inv_1 _06195_ (.Y(_00734_),
    .A(net1104));
 sg13g2_inv_1 _06196_ (.Y(_00735_),
    .A(net1111));
 sg13g2_inv_1 _06197_ (.Y(_00736_),
    .A(net1093));
 sg13g2_inv_1 _06198_ (.Y(_00737_),
    .A(net1071));
 sg13g2_inv_1 _06199_ (.Y(_00738_),
    .A(net1079));
 sg13g2_inv_2 _06200_ (.Y(_00739_),
    .A(net1073));
 sg13g2_inv_1 _06201_ (.Y(_00740_),
    .A(net942));
 sg13g2_inv_1 _06202_ (.Y(_00741_),
    .A(net943));
 sg13g2_inv_1 _06203_ (.Y(_00742_),
    .A(net962));
 sg13g2_inv_1 _06204_ (.Y(_00743_),
    .A(net959));
 sg13g2_inv_1 _06205_ (.Y(_00744_),
    .A(net928));
 sg13g2_inv_1 _06206_ (.Y(_00745_),
    .A(net952));
 sg13g2_inv_1 _06207_ (.Y(_00746_),
    .A(net979));
 sg13g2_inv_1 _06208_ (.Y(_00747_),
    .A(net1012));
 sg13g2_inv_1 _06209_ (.Y(_00748_),
    .A(net1083));
 sg13g2_inv_1 _06210_ (.Y(_00749_),
    .A(net1041));
 sg13g2_inv_1 _06211_ (.Y(_00750_),
    .A(net1106));
 sg13g2_inv_1 _06212_ (.Y(_00751_),
    .A(net1107));
 sg13g2_inv_1 _06213_ (.Y(_00752_),
    .A(net1108));
 sg13g2_inv_2 _06214_ (.Y(_00753_),
    .A(net1063));
 sg13g2_inv_2 _06215_ (.Y(_00754_),
    .A(net1085));
 sg13g2_inv_2 _06216_ (.Y(_00755_),
    .A(net1086));
 sg13g2_inv_1 _06217_ (.Y(_00756_),
    .A(_00119_));
 sg13g2_inv_1 _06218_ (.Y(_00757_),
    .A(_00138_));
 sg13g2_inv_1 _06219_ (.Y(_00758_),
    .A(_00137_));
 sg13g2_inv_1 _06220_ (.Y(_00759_),
    .A(_00140_));
 sg13g2_inv_1 _06221_ (.Y(_00760_),
    .A(_00139_));
 sg13g2_inv_1 _06222_ (.Y(_00761_),
    .A(net1052));
 sg13g2_inv_1 _06223_ (.Y(_00762_),
    .A(net1022));
 sg13g2_inv_1 _06224_ (.Y(_00763_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][13] ));
 sg13g2_inv_1 _06225_ (.Y(_00764_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][3] ));
 sg13g2_inv_1 _06226_ (.Y(_00765_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][2] ));
 sg13g2_inv_1 _06227_ (.Y(_00766_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][5] ));
 sg13g2_inv_1 _06228_ (.Y(_00767_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][4] ));
 sg13g2_inv_1 _06229_ (.Y(_00768_),
    .A(_00142_));
 sg13g2_inv_1 _06230_ (.Y(_00769_),
    .A(net1109));
 sg13g2_inv_1 _06231_ (.Y(_00770_),
    .A(net1044));
 sg13g2_inv_1 _06232_ (.Y(_00771_),
    .A(_00150_));
 sg13g2_inv_1 _06233_ (.Y(_00772_),
    .A(_00149_));
 sg13g2_inv_1 _06234_ (.Y(_00773_),
    .A(_00154_));
 sg13g2_inv_1 _06235_ (.Y(_00774_),
    .A(net903));
 sg13g2_nor4_2 _06236_ (.A(\u_tiny_nn_top.counter_q[4] ),
    .B(\u_tiny_nn_top.counter_q[5] ),
    .C(\u_tiny_nn_top.counter_q[7] ),
    .Y(_00775_),
    .D(\u_tiny_nn_top.counter_q[6] ));
 sg13g2_or4_2 _06237_ (.A(\u_tiny_nn_top.counter_q[4] ),
    .B(\u_tiny_nn_top.counter_q[5] ),
    .C(\u_tiny_nn_top.counter_q[7] ),
    .D(\u_tiny_nn_top.counter_q[6] ),
    .X(_00776_));
 sg13g2_nor2_1 _06238_ (.A(net1857),
    .B(net1855),
    .Y(_00777_));
 sg13g2_nor3_1 _06239_ (.A(net1857),
    .B(net1856),
    .C(\u_tiny_nn_top.counter_q[2] ),
    .Y(_00778_));
 sg13g2_or2_2 _06240_ (.X(_00779_),
    .B(\u_tiny_nn_top.counter_q[3] ),
    .A(\u_tiny_nn_top.counter_q[2] ));
 sg13g2_nor4_2 _06241_ (.A(net1860),
    .B(net1855),
    .C(\u_tiny_nn_top.counter_q[2] ),
    .Y(_00780_),
    .D(\u_tiny_nn_top.counter_q[3] ));
 sg13g2_or4_2 _06242_ (.A(net1860),
    .B(net1856),
    .C(\u_tiny_nn_top.counter_q[2] ),
    .D(\u_tiny_nn_top.counter_q[3] ),
    .X(_00781_));
 sg13g2_nor2_1 _06243_ (.A(_00776_),
    .B(_00781_),
    .Y(_00782_));
 sg13g2_nand2_1 _06244_ (.Y(_00783_),
    .A(_00775_),
    .B(_00780_));
 sg13g2_nand2b_2 _06245_ (.Y(_00784_),
    .B(net1855),
    .A_N(net1860));
 sg13g2_nor2_1 _06246_ (.A(_00776_),
    .B(_00779_),
    .Y(_00785_));
 sg13g2_nor3_2 _06247_ (.A(_00776_),
    .B(_00779_),
    .C(_00784_),
    .Y(_00786_));
 sg13g2_nor2_1 _06248_ (.A(\u_tiny_nn_top.state_q[4] ),
    .B(\u_tiny_nn_top.state_q[14] ),
    .Y(_00787_));
 sg13g2_or2_1 _06249_ (.X(_00788_),
    .B(\u_tiny_nn_top.state_q[14] ),
    .A(\u_tiny_nn_top.state_q[4] ));
 sg13g2_o21ai_1 _06250_ (.B1(net1765),
    .Y(_00789_),
    .A1(\u_tiny_nn_top.state_q[3] ),
    .A2(\u_tiny_nn_top.state_q[6] ));
 sg13g2_nor2_1 _06251_ (.A(\u_tiny_nn_top.state_q[14] ),
    .B(\u_tiny_nn_top.state_q[10] ),
    .Y(_00790_));
 sg13g2_o21ai_1 _06252_ (.B1(_00790_),
    .Y(_00791_),
    .A1(_00786_),
    .A2(_00789_));
 sg13g2_nor3_2 _06253_ (.A(net1824),
    .B(net1827),
    .C(\u_tiny_nn_top.data_i_q[13] ),
    .Y(_00792_));
 sg13g2_nand2_1 _06254_ (.Y(_00793_),
    .A(net1828),
    .B(_00792_));
 sg13g2_nor2_1 _06255_ (.A(net1781),
    .B(net1780),
    .Y(_00794_));
 sg13g2_and3_2 _06256_ (.X(_00795_),
    .A(net1824),
    .B(net1114),
    .C(_00794_));
 sg13g2_nor3_2 _06257_ (.A(net1824),
    .B(net1827),
    .C(net1781),
    .Y(_00796_));
 sg13g2_nor3_2 _06258_ (.A(net1824),
    .B(net1784),
    .C(\u_tiny_nn_top.data_i_q[13] ),
    .Y(_00797_));
 sg13g2_nor4_2 _06259_ (.A(_00660_),
    .B(_00795_),
    .C(_00796_),
    .Y(_00798_),
    .D(_00797_));
 sg13g2_a21oi_1 _06260_ (.A1(net1828),
    .A2(_00792_),
    .Y(_00799_),
    .B1(_00660_));
 sg13g2_nand2_1 _06261_ (.Y(_00800_),
    .A(net1793),
    .B(_00793_));
 sg13g2_nand2_1 _06262_ (.Y(_00801_),
    .A(\u_tiny_nn_top.state_q[13] ),
    .B(net1740));
 sg13g2_nor3_1 _06263_ (.A(\u_tiny_nn_top.data_i_q[11] ),
    .B(\u_tiny_nn_top.data_i_q[10] ),
    .C(\u_tiny_nn_top.data_i_q[9] ),
    .Y(_00802_));
 sg13g2_inv_1 _06264_ (.Y(_00803_),
    .A(_00802_));
 sg13g2_nor4_2 _06265_ (.A(net1777),
    .B(net1776),
    .C(net1774),
    .Y(_00804_),
    .D(_00644_));
 sg13g2_nand3_1 _06266_ (.B(_00795_),
    .C(_00803_),
    .A(\u_tiny_nn_top.state_q[0] ),
    .Y(_00805_));
 sg13g2_o21ai_1 _06267_ (.B1(_00801_),
    .Y(_00806_),
    .A1(_00804_),
    .A2(_00805_));
 sg13g2_nor2_1 _06268_ (.A(net1830),
    .B(_00803_),
    .Y(_00807_));
 sg13g2_nand2_1 _06269_ (.Y(_00808_),
    .A(_00795_),
    .B(_00807_));
 sg13g2_nand2_1 _06270_ (.Y(_00809_),
    .A(net1830),
    .B(_00795_));
 sg13g2_nand2_1 _06271_ (.Y(_00810_),
    .A(_00795_),
    .B(_00804_));
 sg13g2_a221oi_1 _06272_ (.B2(\u_tiny_nn_top.state_q[17] ),
    .C1(_00806_),
    .B1(_00810_),
    .A1(\u_tiny_nn_top.state_q[8] ),
    .Y(_00811_),
    .A2(_00808_));
 sg13g2_a221oi_1 _06273_ (.B2(_00798_),
    .C1(net1003),
    .B1(_00793_),
    .A1(net1740),
    .Y(_00812_),
    .A2(_00791_));
 sg13g2_and2_1 _06274_ (.A(_00811_),
    .B(_00812_),
    .X(_00187_));
 sg13g2_xnor2_1 _06275_ (.Y(_00813_),
    .A(\u_tiny_nn_top.counter_q[7] ),
    .B(\u_tiny_nn_top.start_count_q[7] ));
 sg13g2_xnor2_1 _06276_ (.Y(_00814_),
    .A(net1856),
    .B(\u_tiny_nn_top.start_count_q[1] ));
 sg13g2_xor2_1 _06277_ (.B(\u_tiny_nn_top.start_count_q[0] ),
    .A(net1857),
    .X(_00815_));
 sg13g2_xnor2_1 _06278_ (.Y(_00816_),
    .A(\u_tiny_nn_top.counter_q[3] ),
    .B(\u_tiny_nn_top.start_count_q[3] ));
 sg13g2_xnor2_1 _06279_ (.Y(_00817_),
    .A(\u_tiny_nn_top.counter_q[2] ),
    .B(\u_tiny_nn_top.start_count_q[2] ));
 sg13g2_xnor2_1 _06280_ (.Y(_00818_),
    .A(\u_tiny_nn_top.counter_q[5] ),
    .B(\u_tiny_nn_top.start_count_q[5] ));
 sg13g2_xnor2_1 _06281_ (.Y(_00819_),
    .A(\u_tiny_nn_top.counter_q[6] ),
    .B(\u_tiny_nn_top.start_count_q[6] ));
 sg13g2_xnor2_1 _06282_ (.Y(_00820_),
    .A(\u_tiny_nn_top.counter_q[4] ),
    .B(\u_tiny_nn_top.start_count_q[4] ));
 sg13g2_nand4_1 _06283_ (.B(_00814_),
    .C(_00819_),
    .A(_00813_),
    .Y(_00821_),
    .D(_00820_));
 sg13g2_nand3_1 _06284_ (.B(_00817_),
    .C(_00818_),
    .A(_00816_),
    .Y(_00822_));
 sg13g2_nor3_2 _06285_ (.A(_00815_),
    .B(_00821_),
    .C(_00822_),
    .Y(_00823_));
 sg13g2_nand2b_1 _06286_ (.Y(_00824_),
    .B(net918),
    .A_N(_00823_));
 sg13g2_nor2_1 _06287_ (.A(\u_tiny_nn_top.state_q[15] ),
    .B(net1790),
    .Y(_00825_));
 sg13g2_or2_2 _06288_ (.X(_00826_),
    .B(net1790),
    .A(\u_tiny_nn_top.state_q[15] ));
 sg13g2_a21oi_1 _06289_ (.A1(_00097_),
    .A2(net1730),
    .Y(_00827_),
    .B1(net1763));
 sg13g2_nand2_2 _06290_ (.Y(_00828_),
    .A(\u_tiny_nn_top.state_q[12] ),
    .B(net1736));
 sg13g2_nand2b_2 _06291_ (.Y(_00829_),
    .B(_00828_),
    .A_N(\u_tiny_nn_top.state_q[7] ));
 sg13g2_nand2_1 _06292_ (.Y(_00830_),
    .A(\u_tiny_nn_top.max_val_skid_q[7] ),
    .B(_00829_));
 sg13g2_nor2_1 _06293_ (.A(\u_tiny_nn_top.state_q[6] ),
    .B(\u_tiny_nn_top.state_q[10] ),
    .Y(_00831_));
 sg13g2_nor3_2 _06294_ (.A(\u_tiny_nn_top.state_q[3] ),
    .B(\u_tiny_nn_top.state_q[6] ),
    .C(\u_tiny_nn_top.state_q[10] ),
    .Y(_00832_));
 sg13g2_nand2_2 _06295_ (.Y(_00833_),
    .A(_00658_),
    .B(_00831_));
 sg13g2_nor3_2 _06296_ (.A(net1788),
    .B(\u_tiny_nn_top.state_q[17] ),
    .C(\u_tiny_nn_top.state_q[8] ),
    .Y(_00834_));
 sg13g2_inv_1 _06297_ (.Y(_00835_),
    .A(_00834_));
 sg13g2_nor3_2 _06298_ (.A(net1788),
    .B(\u_tiny_nn_top.state_q[8] ),
    .C(_00833_),
    .Y(_00836_));
 sg13g2_nand2_2 _06299_ (.Y(_00837_),
    .A(_00832_),
    .B(_00834_));
 sg13g2_nor2_1 _06300_ (.A(\u_tiny_nn_top.state_q[12] ),
    .B(\u_tiny_nn_top.state_q[15] ),
    .Y(_00838_));
 sg13g2_nor2_2 _06301_ (.A(\u_tiny_nn_top.state_q[12] ),
    .B(_00826_),
    .Y(_00839_));
 sg13g2_nand2_2 _06302_ (.Y(_00840_),
    .A(_00655_),
    .B(net1763));
 sg13g2_nor4_2 _06303_ (.A(\u_tiny_nn_top.state_q[7] ),
    .B(net1764),
    .C(_00837_),
    .Y(_00841_),
    .D(_00840_));
 sg13g2_o21ai_1 _06304_ (.B1(_00788_),
    .Y(_00842_),
    .A1(net1852),
    .A2(net798));
 sg13g2_a21oi_1 _06305_ (.A1(net1852),
    .A2(_00721_),
    .Y(_00843_),
    .B1(_00842_));
 sg13g2_nand2_1 _06306_ (.Y(_00844_),
    .A(net1858),
    .B(\u_tiny_nn_top.state_q[8] ));
 sg13g2_a221oi_1 _06307_ (.B2(net1859),
    .C1(_00843_),
    .B1(\u_tiny_nn_top.state_q[8] ),
    .A1(\u_tiny_nn_top.counter_q[7] ),
    .Y(_00845_),
    .A2(net1788));
 sg13g2_nor2b_1 _06308_ (.A(net1859),
    .B_N(net918),
    .Y(_00846_));
 sg13g2_a21oi_1 _06309_ (.A1(net1859),
    .A2(_00097_),
    .Y(_00847_),
    .B1(_00846_));
 sg13g2_a21oi_1 _06310_ (.A1(_00833_),
    .A2(_00847_),
    .Y(_00848_),
    .B1(_00841_));
 sg13g2_nand3_1 _06311_ (.B(_00845_),
    .C(_00848_),
    .A(_00830_),
    .Y(_00849_));
 sg13g2_xnor2_1 _06312_ (.Y(_00850_),
    .A(net1823),
    .B(\u_tiny_nn_top.max_val_q[15] ));
 sg13g2_nor2_1 _06313_ (.A(net1783),
    .B(\u_tiny_nn_top.max_val_q[14] ),
    .Y(_00851_));
 sg13g2_a22oi_1 _06314_ (.Y(_00852_),
    .B1(\u_tiny_nn_top.max_val_q[10] ),
    .B2(net1776),
    .A2(\u_tiny_nn_top.max_val_q[9] ),
    .A1(net1774));
 sg13g2_a22oi_1 _06315_ (.Y(_00853_),
    .B1(_00669_),
    .B2(\u_tiny_nn_top.data_i_q[9] ),
    .A2(_00668_),
    .A1(net1830));
 sg13g2_nand2b_1 _06316_ (.Y(_00854_),
    .B(\u_tiny_nn_top.max_val_q[7] ),
    .A_N(net1833));
 sg13g2_o21ai_1 _06317_ (.B1(_00854_),
    .Y(_00855_),
    .A1(net1830),
    .A2(_00668_));
 sg13g2_nand2_1 _06318_ (.Y(_00856_),
    .A(_00853_),
    .B(_00855_));
 sg13g2_and2_1 _06319_ (.A(_00852_),
    .B(_00856_),
    .X(_00857_));
 sg13g2_a22oi_1 _06320_ (.Y(_00858_),
    .B1(_00671_),
    .B2(net1829),
    .A2(_00670_),
    .A1(\u_tiny_nn_top.data_i_q[13] ));
 sg13g2_nand2b_1 _06321_ (.Y(_00859_),
    .B(\u_tiny_nn_top.data_i_q[11] ),
    .A_N(\u_tiny_nn_top.max_val_q[11] ));
 sg13g2_nand2b_1 _06322_ (.Y(_00860_),
    .B(\u_tiny_nn_top.data_i_q[10] ),
    .A_N(\u_tiny_nn_top.max_val_q[10] ));
 sg13g2_nand2_1 _06323_ (.Y(_00861_),
    .A(_00859_),
    .B(_00860_));
 sg13g2_nand3_1 _06324_ (.B(_00859_),
    .C(_00860_),
    .A(_00858_),
    .Y(_00862_));
 sg13g2_a22oi_1 _06325_ (.Y(_00863_),
    .B1(\u_tiny_nn_top.max_val_q[14] ),
    .B2(net1783),
    .A2(\u_tiny_nn_top.max_val_q[13] ),
    .A1(net1782));
 sg13g2_a22oi_1 _06326_ (.Y(_00864_),
    .B1(\u_tiny_nn_top.max_val_q[12] ),
    .B2(net1779),
    .A2(\u_tiny_nn_top.max_val_q[11] ),
    .A1(net1777));
 sg13g2_o21ai_1 _06327_ (.B1(_00864_),
    .Y(_00865_),
    .A1(_00857_),
    .A2(_00861_));
 sg13g2_nand2_1 _06328_ (.Y(_00866_),
    .A(_00858_),
    .B(_00865_));
 sg13g2_a21oi_1 _06329_ (.A1(_00863_),
    .A2(_00866_),
    .Y(_00867_),
    .B1(_00851_));
 sg13g2_nand2b_1 _06330_ (.Y(_00868_),
    .B(\u_tiny_nn_top.max_val_q[6] ),
    .A_N(net1838));
 sg13g2_o21ai_1 _06331_ (.B1(_00868_),
    .Y(_00869_),
    .A1(net1840),
    .A2(_00666_));
 sg13g2_a22oi_1 _06332_ (.Y(_00870_),
    .B1(_00667_),
    .B2(net1843),
    .A2(_00666_),
    .A1(net1840));
 sg13g2_a22oi_1 _06333_ (.Y(_00871_),
    .B1(_00665_),
    .B2(\u_tiny_nn_top.data_i_q[2] ),
    .A2(_00664_),
    .A1(net1847));
 sg13g2_nor2_1 _06334_ (.A(net1847),
    .B(_00664_),
    .Y(_00872_));
 sg13g2_a21oi_1 _06335_ (.A1(net1771),
    .A2(\u_tiny_nn_top.max_val_q[2] ),
    .Y(_00873_),
    .B1(_00872_));
 sg13g2_and2_1 _06336_ (.A(_00871_),
    .B(_00873_),
    .X(_00874_));
 sg13g2_xor2_1 _06337_ (.B(\u_tiny_nn_top.max_val_q[1] ),
    .A(net1849),
    .X(_00875_));
 sg13g2_a21oi_1 _06338_ (.A1(net1769),
    .A2(\u_tiny_nn_top.max_val_q[0] ),
    .Y(_00876_),
    .B1(_00875_));
 sg13g2_a21oi_1 _06339_ (.A1(net1849),
    .A2(_00663_),
    .Y(_00877_),
    .B1(_00876_));
 sg13g2_nand2b_1 _06340_ (.Y(_00878_),
    .B(_00874_),
    .A_N(_00877_));
 sg13g2_o21ai_1 _06341_ (.B1(_00878_),
    .Y(_00879_),
    .A1(_00871_),
    .A2(_00872_));
 sg13g2_nand2b_1 _06342_ (.Y(_00880_),
    .B(\u_tiny_nn_top.max_val_q[4] ),
    .A_N(net1843));
 sg13g2_nand2b_1 _06343_ (.Y(_00881_),
    .B(\u_tiny_nn_top.data_i_q[0] ),
    .A_N(\u_tiny_nn_top.max_val_q[0] ));
 sg13g2_nand3_1 _06344_ (.B(_00876_),
    .C(_00881_),
    .A(_00874_),
    .Y(_00882_));
 sg13g2_nand3_1 _06345_ (.B(_00880_),
    .C(_00882_),
    .A(_00879_),
    .Y(_00883_));
 sg13g2_a21oi_1 _06346_ (.A1(_00870_),
    .A2(_00883_),
    .Y(_00884_),
    .B1(_00869_));
 sg13g2_nor2b_1 _06347_ (.A(\u_tiny_nn_top.max_val_q[7] ),
    .B_N(net1833),
    .Y(_00885_));
 sg13g2_nor2b_1 _06348_ (.A(\u_tiny_nn_top.max_val_q[6] ),
    .B_N(net1838),
    .Y(_00886_));
 sg13g2_nand4_1 _06349_ (.B(_00853_),
    .C(_00863_),
    .A(_00852_),
    .Y(_00887_),
    .D(_00864_));
 sg13g2_nor4_1 _06350_ (.A(_00851_),
    .B(_00855_),
    .C(_00862_),
    .D(_00885_),
    .Y(_00888_));
 sg13g2_nand2b_1 _06351_ (.Y(_00889_),
    .B(_00888_),
    .A_N(_00887_));
 sg13g2_nor3_1 _06352_ (.A(_00884_),
    .B(_00886_),
    .C(_00889_),
    .Y(_00890_));
 sg13g2_o21ai_1 _06353_ (.B1(_00850_),
    .Y(_00891_),
    .A1(_00867_),
    .A2(_00890_));
 sg13g2_nor3_1 _06354_ (.A(\u_tiny_nn_top.max_val_q[5] ),
    .B(\u_tiny_nn_top.max_val_q[4] ),
    .C(\u_tiny_nn_top.max_val_q[6] ),
    .Y(_00892_));
 sg13g2_nor3_1 _06355_ (.A(\u_tiny_nn_top.max_val_q[1] ),
    .B(\u_tiny_nn_top.max_val_q[0] ),
    .C(\u_tiny_nn_top.max_val_q[3] ),
    .Y(_00893_));
 sg13g2_nand3_1 _06356_ (.B(_00892_),
    .C(_00893_),
    .A(_00665_),
    .Y(_00894_));
 sg13g2_inv_1 _06357_ (.Y(_00895_),
    .A(_00894_));
 sg13g2_nand4_1 _06358_ (.B(\u_tiny_nn_top.max_val_q[13] ),
    .C(\u_tiny_nn_top.max_val_q[12] ),
    .A(\u_tiny_nn_top.max_val_q[11] ),
    .Y(_00896_),
    .D(\u_tiny_nn_top.max_val_q[14] ));
 sg13g2_nand4_1 _06359_ (.B(\u_tiny_nn_top.max_val_q[8] ),
    .C(\u_tiny_nn_top.max_val_q[9] ),
    .A(\u_tiny_nn_top.max_val_q[7] ),
    .Y(_00897_),
    .D(\u_tiny_nn_top.max_val_q[10] ));
 sg13g2_nor2_1 _06360_ (.A(_00896_),
    .B(_00897_),
    .Y(_00898_));
 sg13g2_nor4_1 _06361_ (.A(net1827),
    .B(\u_tiny_nn_top.data_i_q[13] ),
    .C(net1829),
    .D(net1833),
    .Y(_00899_));
 sg13g2_and2_1 _06362_ (.A(_00807_),
    .B(_00899_),
    .X(_00900_));
 sg13g2_or4_1 _06363_ (.A(net1846),
    .B(\u_tiny_nn_top.data_i_q[2] ),
    .C(net1849),
    .D(\u_tiny_nn_top.data_i_q[0] ),
    .X(_00901_));
 sg13g2_nor3_2 _06364_ (.A(net1841),
    .B(net1844),
    .C(_00901_),
    .Y(_00902_));
 sg13g2_nor2_1 _06365_ (.A(net1823),
    .B(net1837),
    .Y(_00903_));
 sg13g2_and2_1 _06366_ (.A(_00900_),
    .B(_00903_),
    .X(_00904_));
 sg13g2_a22oi_1 _06367_ (.Y(_00905_),
    .B1(_00902_),
    .B2(_00904_),
    .A2(_00898_),
    .A1(_00895_));
 sg13g2_and2_1 _06368_ (.A(_00168_),
    .B(_00905_),
    .X(_00906_));
 sg13g2_nand2_1 _06369_ (.Y(_00907_),
    .A(net1823),
    .B(_00867_));
 sg13g2_nand2_1 _06370_ (.Y(_00908_),
    .A(_00905_),
    .B(_00907_));
 sg13g2_nand4_1 _06371_ (.B(net1833),
    .C(_00794_),
    .A(net1827),
    .Y(_00909_),
    .D(_00804_));
 sg13g2_nand3b_1 _06372_ (.B(_00902_),
    .C(net1834),
    .Y(_00910_),
    .A_N(net1837));
 sg13g2_nor2_1 _06373_ (.A(_00909_),
    .B(_00910_),
    .Y(_00911_));
 sg13g2_a221oi_1 _06374_ (.B2(\u_tiny_nn_top.max_val_q[15] ),
    .C1(_00911_),
    .B1(_00908_),
    .A1(_00891_),
    .Y(_00912_),
    .A2(_00906_));
 sg13g2_and2_1 _06375_ (.A(_00850_),
    .B(_00880_),
    .X(_00913_));
 sg13g2_nand3b_1 _06376_ (.B(_00870_),
    .C(_00913_),
    .Y(_00914_),
    .A_N(_00869_));
 sg13g2_nor4_1 _06377_ (.A(_00882_),
    .B(_00886_),
    .C(_00889_),
    .D(_00914_),
    .Y(_00915_));
 sg13g2_nand2_1 _06378_ (.Y(_00916_),
    .A(_00017_),
    .B(_00902_));
 sg13g2_nor4_1 _06379_ (.A(\u_tiny_nn_top.max_val_q[11] ),
    .B(\u_tiny_nn_top.max_val_q[13] ),
    .C(\u_tiny_nn_top.max_val_q[12] ),
    .D(\u_tiny_nn_top.max_val_q[14] ),
    .Y(_00917_));
 sg13g2_nor4_1 _06380_ (.A(\u_tiny_nn_top.max_val_q[7] ),
    .B(\u_tiny_nn_top.max_val_q[8] ),
    .C(\u_tiny_nn_top.max_val_q[9] ),
    .D(\u_tiny_nn_top.max_val_q[10] ),
    .Y(_00918_));
 sg13g2_and2_1 _06381_ (.A(_00917_),
    .B(_00918_),
    .X(_00919_));
 sg13g2_o21ai_1 _06382_ (.B1(_00919_),
    .Y(_00920_),
    .A1(\u_tiny_nn_top.max_val_q[15] ),
    .A2(_00894_));
 sg13g2_o21ai_1 _06383_ (.B1(_00900_),
    .Y(_00921_),
    .A1(net1823),
    .A2(_00916_));
 sg13g2_nand2b_1 _06384_ (.Y(_00922_),
    .B(_00911_),
    .A_N(_00168_));
 sg13g2_nor2b_1 _06385_ (.A(_00909_),
    .B_N(_00916_),
    .Y(_00923_));
 sg13g2_a21oi_1 _06386_ (.A1(_00894_),
    .A2(_00898_),
    .Y(_00924_),
    .B1(_00923_));
 sg13g2_nand4_1 _06387_ (.B(_00921_),
    .C(_00922_),
    .A(_00920_),
    .Y(_00925_),
    .D(_00924_));
 sg13g2_or3_1 _06388_ (.A(_00912_),
    .B(_00915_),
    .C(_00925_),
    .X(_00926_));
 sg13g2_nor2_2 _06389_ (.A(_00655_),
    .B(net1736),
    .Y(_00927_));
 sg13g2_nand2_1 _06390_ (.Y(_00928_),
    .A(\u_tiny_nn_top.state_q[12] ),
    .B(net1740));
 sg13g2_mux2_2 _06391_ (.A0(net1833),
    .A1(\u_tiny_nn_top.max_val_q[7] ),
    .S(net1480),
    .X(_00929_));
 sg13g2_a221oi_1 _06392_ (.B2(_00929_),
    .C1(_00849_),
    .B1(_00927_),
    .A1(_00824_),
    .Y(_00186_),
    .A2(_00827_));
 sg13g2_mux2_1 _06393_ (.A0(net1096),
    .A1(_00095_),
    .S(net1730),
    .X(_00930_));
 sg13g2_and2_1 _06394_ (.A(\u_tiny_nn_top.state_q[17] ),
    .B(_00785_),
    .X(_00931_));
 sg13g2_mux2_1 _06395_ (.A0(_00096_),
    .A1(_00095_),
    .S(net1858),
    .X(_00932_));
 sg13g2_nor2_1 _06396_ (.A(net1852),
    .B(net887),
    .Y(_00933_));
 sg13g2_nor2b_1 _06397_ (.A(net734),
    .B_N(net1852),
    .Y(_00934_));
 sg13g2_nor3_2 _06398_ (.A(net1765),
    .B(_00933_),
    .C(_00934_),
    .Y(_00935_));
 sg13g2_nor2b_1 _06399_ (.A(net1860),
    .B_N(\u_tiny_nn_top.state_q[8] ),
    .Y(_00936_));
 sg13g2_a21oi_1 _06400_ (.A1(\u_tiny_nn_top.counter_q[6] ),
    .A2(net1788),
    .Y(_00937_),
    .B1(_00936_));
 sg13g2_o21ai_1 _06401_ (.B1(_00937_),
    .Y(_00938_),
    .A1(_00832_),
    .A2(_00932_));
 sg13g2_a221oi_1 _06402_ (.B2(_00784_),
    .C1(_00938_),
    .B1(_00931_),
    .A1(net852),
    .Y(_00939_),
    .A2(_00829_));
 sg13g2_o21ai_1 _06403_ (.B1(_00939_),
    .Y(_00940_),
    .A1(_00825_),
    .A2(net1097));
 sg13g2_nor2b_1 _06404_ (.A(\u_tiny_nn_top.max_val_q[6] ),
    .B_N(net1478),
    .Y(_00941_));
 sg13g2_nor2_1 _06405_ (.A(net1837),
    .B(net1480),
    .Y(_00942_));
 sg13g2_nor3_2 _06406_ (.A(net1726),
    .B(_00941_),
    .C(_00942_),
    .Y(_00943_));
 sg13g2_nor4_2 _06407_ (.A(_00841_),
    .B(_00935_),
    .C(_00940_),
    .Y(_00185_),
    .D(_00943_));
 sg13g2_mux2_1 _06408_ (.A0(net1067),
    .A1(_00093_),
    .S(net1730),
    .X(_00944_));
 sg13g2_a21o_1 _06409_ (.A2(_00786_),
    .A1(\u_tiny_nn_top.state_q[17] ),
    .B1(_00841_),
    .X(_00945_));
 sg13g2_o21ai_1 _06410_ (.B1(_00788_),
    .Y(_00946_),
    .A1(net1852),
    .A2(net794));
 sg13g2_a21oi_2 _06411_ (.B1(_00946_),
    .Y(_00947_),
    .A2(_00717_),
    .A1(net1852));
 sg13g2_mux2_1 _06412_ (.A0(_00094_),
    .A1(_00093_),
    .S(net1858),
    .X(_00948_));
 sg13g2_a22oi_1 _06413_ (.Y(_00949_),
    .B1(\u_tiny_nn_top.state_q[8] ),
    .B2(net1859),
    .A2(net1788),
    .A1(\u_tiny_nn_top.counter_q[5] ));
 sg13g2_o21ai_1 _06414_ (.B1(_00949_),
    .Y(_00950_),
    .A1(_00832_),
    .A2(_00948_));
 sg13g2_a21oi_1 _06415_ (.A1(net773),
    .A2(_00829_),
    .Y(_00951_),
    .B1(_00950_));
 sg13g2_o21ai_1 _06416_ (.B1(_00951_),
    .Y(_00952_),
    .A1(_00825_),
    .A2(_00944_));
 sg13g2_nor2_1 _06417_ (.A(net1840),
    .B(net1478),
    .Y(_00953_));
 sg13g2_a21oi_1 _06418_ (.A1(_00666_),
    .A2(net1478),
    .Y(_00954_),
    .B1(net1726));
 sg13g2_nor2b_2 _06419_ (.A(_00953_),
    .B_N(_00954_),
    .Y(_00955_));
 sg13g2_nor4_2 _06420_ (.A(_00945_),
    .B(_00947_),
    .C(_00952_),
    .Y(_00184_),
    .D(_00955_));
 sg13g2_nand2_1 _06421_ (.Y(_00956_),
    .A(net1861),
    .B(net1855));
 sg13g2_nand3_1 _06422_ (.B(net1855),
    .C(_00785_),
    .A(net1861),
    .Y(_00957_));
 sg13g2_a21oi_1 _06423_ (.A1(\u_tiny_nn_top.counter_q[4] ),
    .A2(net1788),
    .Y(_00958_),
    .B1(_00936_));
 sg13g2_o21ai_1 _06424_ (.B1(_00958_),
    .Y(_00959_),
    .A1(_00162_),
    .A2(_00957_));
 sg13g2_mux2_1 _06425_ (.A0(_00092_),
    .A1(_00091_),
    .S(net1730),
    .X(_00960_));
 sg13g2_nand2_1 _06426_ (.Y(_00961_),
    .A(net1854),
    .B(\u_tiny_nn_top.core_accumulate_result[12] ));
 sg13g2_o21ai_1 _06427_ (.B1(_00961_),
    .Y(_00962_),
    .A1(net1854),
    .A2(_00714_));
 sg13g2_mux2_1 _06428_ (.A0(_00092_),
    .A1(net1099),
    .S(net1858),
    .X(_00963_));
 sg13g2_a221oi_1 _06429_ (.B2(net1764),
    .C1(_00841_),
    .B1(_00962_),
    .A1(_00835_),
    .Y(_00964_),
    .A2(_00959_));
 sg13g2_o21ai_1 _06430_ (.B1(_00964_),
    .Y(_00965_),
    .A1(net1763),
    .A2(_00960_));
 sg13g2_a21oi_1 _06431_ (.A1(net829),
    .A2(_00829_),
    .Y(_00966_),
    .B1(_00965_));
 sg13g2_o21ai_1 _06432_ (.B1(_00966_),
    .Y(_00967_),
    .A1(_00832_),
    .A2(_00963_));
 sg13g2_nor2_1 _06433_ (.A(net1843),
    .B(net1477),
    .Y(_00968_));
 sg13g2_a21oi_1 _06434_ (.A1(_00667_),
    .A2(net1477),
    .Y(_00969_),
    .B1(_00968_));
 sg13g2_a21oi_1 _06435_ (.A1(_00927_),
    .A2(_00969_),
    .Y(_00183_),
    .B1(_00967_));
 sg13g2_mux2_1 _06436_ (.A0(net1094),
    .A1(_00089_),
    .S(net1730),
    .X(_00970_));
 sg13g2_mux2_1 _06437_ (.A0(_00090_),
    .A1(_00089_),
    .S(net1858),
    .X(_00971_));
 sg13g2_a21oi_1 _06438_ (.A1(net1853),
    .A2(_00713_),
    .Y(_00972_),
    .B1(net1766));
 sg13g2_o21ai_1 _06439_ (.B1(_00972_),
    .Y(_00973_),
    .A1(net1852),
    .A2(net815));
 sg13g2_o21ai_1 _06440_ (.B1(_00973_),
    .Y(_00974_),
    .A1(_00654_),
    .A2(_00659_));
 sg13g2_o21ai_1 _06441_ (.B1(_00844_),
    .Y(_00975_),
    .A1(_00832_),
    .A2(_00971_));
 sg13g2_a221oi_1 _06442_ (.B2(_00956_),
    .C1(_00975_),
    .B1(_00931_),
    .A1(net835),
    .Y(_00976_),
    .A2(_00829_));
 sg13g2_o21ai_1 _06443_ (.B1(_00976_),
    .Y(_00977_),
    .A1(net1763),
    .A2(net1095));
 sg13g2_nor2_1 _06444_ (.A(net1846),
    .B(net1477),
    .Y(_00978_));
 sg13g2_a21oi_1 _06445_ (.A1(_00664_),
    .A2(net1477),
    .Y(_00979_),
    .B1(net1726));
 sg13g2_nor2b_2 _06446_ (.A(_00978_),
    .B_N(_00979_),
    .Y(_00980_));
 sg13g2_nor4_2 _06447_ (.A(_00841_),
    .B(_00974_),
    .C(_00977_),
    .Y(_00182_),
    .D(_00980_));
 sg13g2_nand2b_1 _06448_ (.Y(_00981_),
    .B(net1064),
    .A_N(_00823_));
 sg13g2_a21oi_1 _06449_ (.A1(_00087_),
    .A2(_00823_),
    .Y(_00982_),
    .B1(net1763));
 sg13g2_nor2_1 _06450_ (.A(net1852),
    .B(\u_tiny_nn_top.core_accumulate_result[2] ),
    .Y(_00983_));
 sg13g2_a21oi_1 _06451_ (.A1(net1853),
    .A2(_00711_),
    .Y(_00984_),
    .B1(_00983_));
 sg13g2_mux2_1 _06452_ (.A0(_00088_),
    .A1(_00087_),
    .S(net1859),
    .X(_00985_));
 sg13g2_a22oi_1 _06453_ (.Y(_00986_),
    .B1(net1764),
    .B2(_00984_),
    .A2(\u_tiny_nn_top.state_q[13] ),
    .A1(\u_tiny_nn_top.counter_q[2] ));
 sg13g2_o21ai_1 _06454_ (.B1(_00986_),
    .Y(_00987_),
    .A1(_00832_),
    .A2(_00985_));
 sg13g2_nor4_2 _06455_ (.A(_00841_),
    .B(_00931_),
    .C(_00936_),
    .Y(_00988_),
    .D(_00987_));
 sg13g2_a22oi_1 _06456_ (.Y(_00989_),
    .B1(_00981_),
    .B2(_00982_),
    .A2(_00829_),
    .A1(\u_tiny_nn_top.max_val_skid_q[2] ));
 sg13g2_nor2_1 _06457_ (.A(\u_tiny_nn_top.data_i_q[2] ),
    .B(net1478),
    .Y(_00990_));
 sg13g2_a21oi_1 _06458_ (.A1(_00665_),
    .A2(net1477),
    .Y(_00991_),
    .B1(net1726));
 sg13g2_nand2b_2 _06459_ (.Y(_00992_),
    .B(_00991_),
    .A_N(_00990_));
 sg13g2_and3_1 _06460_ (.X(_00181_),
    .A(_00988_),
    .B(net1065),
    .C(_00992_));
 sg13g2_a21oi_1 _06461_ (.A1(_00085_),
    .A2(net1730),
    .Y(_00993_),
    .B1(net1763));
 sg13g2_o21ai_1 _06462_ (.B1(_00993_),
    .Y(_00994_),
    .A1(_00709_),
    .A2(net1730));
 sg13g2_nor2b_1 _06463_ (.A(\u_tiny_nn_top.core_accumulate_result[9] ),
    .B_N(net1853),
    .Y(_00995_));
 sg13g2_nor2_1 _06464_ (.A(net1853),
    .B(\u_tiny_nn_top.core_accumulate_result[1] ),
    .Y(_00996_));
 sg13g2_nor3_2 _06465_ (.A(net1766),
    .B(_00995_),
    .C(_00996_),
    .Y(_00997_));
 sg13g2_mux2_1 _06466_ (.A0(_00086_),
    .A1(_00085_),
    .S(net1858),
    .X(_00998_));
 sg13g2_a22oi_1 _06467_ (.Y(_00999_),
    .B1(\u_tiny_nn_top.state_q[8] ),
    .B2(net1860),
    .A2(net1788),
    .A1(net1855));
 sg13g2_o21ai_1 _06468_ (.B1(_00999_),
    .Y(_01000_),
    .A1(_00832_),
    .A2(_00998_));
 sg13g2_nor3_1 _06469_ (.A(_00841_),
    .B(_00997_),
    .C(_01000_),
    .Y(_01001_));
 sg13g2_a22oi_1 _06470_ (.Y(_01002_),
    .B1(_00931_),
    .B2(_00653_),
    .A2(_00829_),
    .A1(\u_tiny_nn_top.max_val_skid_q[1] ));
 sg13g2_nand3_1 _06471_ (.B(_01001_),
    .C(_01002_),
    .A(net1101),
    .Y(_01003_));
 sg13g2_nor2_1 _06472_ (.A(net1849),
    .B(net1477),
    .Y(_01004_));
 sg13g2_a21oi_1 _06473_ (.A1(_00663_),
    .A2(net1477),
    .Y(_01005_),
    .B1(_01004_));
 sg13g2_a21oi_1 _06474_ (.A1(_00927_),
    .A2(_01005_),
    .Y(_00180_),
    .B1(_01003_));
 sg13g2_mux2_1 _06475_ (.A0(_00084_),
    .A1(_00083_),
    .S(net1730),
    .X(_01006_));
 sg13g2_nand2b_1 _06476_ (.Y(_01007_),
    .B(net1858),
    .A_N(_00083_));
 sg13g2_o21ai_1 _06477_ (.B1(_01007_),
    .Y(_01008_),
    .A1(net1858),
    .A2(_00084_));
 sg13g2_o21ai_1 _06478_ (.B1(net1764),
    .Y(_01009_),
    .A1(net1853),
    .A2(\u_tiny_nn_top.core_accumulate_result[0] ));
 sg13g2_a21oi_1 _06479_ (.A1(net1853),
    .A2(_00706_),
    .Y(_01010_),
    .B1(_01009_));
 sg13g2_nand2b_1 _06480_ (.Y(_01011_),
    .B(net1857),
    .A_N(_00165_));
 sg13g2_o21ai_1 _06481_ (.B1(_01011_),
    .Y(_01012_),
    .A1(net1857),
    .A2(_00167_));
 sg13g2_a221oi_1 _06482_ (.B2(_00835_),
    .C1(_01010_),
    .B1(_01012_),
    .A1(_00833_),
    .Y(_01013_),
    .A2(_01008_));
 sg13g2_nand2b_1 _06483_ (.Y(_01014_),
    .B(_01013_),
    .A_N(_00945_));
 sg13g2_a21oi_1 _06484_ (.A1(net704),
    .A2(_00829_),
    .Y(_01015_),
    .B1(_01014_));
 sg13g2_o21ai_1 _06485_ (.B1(_01015_),
    .Y(_01016_),
    .A1(net1763),
    .A2(_01006_));
 sg13g2_nor2b_1 _06486_ (.A(net1033),
    .B_N(net1481),
    .Y(_01017_));
 sg13g2_nor2_1 _06487_ (.A(\u_tiny_nn_top.data_i_q[0] ),
    .B(net1481),
    .Y(_01018_));
 sg13g2_nor3_1 _06488_ (.A(net1726),
    .B(_01017_),
    .C(_01018_),
    .Y(_01019_));
 sg13g2_nor2_1 _06489_ (.A(_01016_),
    .B(_01019_),
    .Y(_00179_));
 sg13g2_nand4_1 _06490_ (.B(\u_tiny_nn_top.data_i_q[2] ),
    .C(net1849),
    .A(net1846),
    .Y(_01020_),
    .D(\u_tiny_nn_top.data_i_q[0] ));
 sg13g2_nand4_1 _06491_ (.B(net1837),
    .C(net1841),
    .A(net1834),
    .Y(_01021_),
    .D(net1844));
 sg13g2_nor3_2 _06492_ (.A(_00810_),
    .B(_01020_),
    .C(_01021_),
    .Y(_01022_));
 sg13g2_inv_1 _06493_ (.Y(_01023_),
    .A(net1555));
 sg13g2_nand2_1 _06494_ (.Y(_01024_),
    .A(net993),
    .B(_01023_));
 sg13g2_o21ai_1 _06495_ (.B1(_01024_),
    .Y(_00013_),
    .A1(_00652_),
    .A2(_00656_));
 sg13g2_nand3_1 _06496_ (.B(net1736),
    .C(net1765),
    .A(net989),
    .Y(_01025_));
 sg13g2_nand3_1 _06497_ (.B(_00786_),
    .C(_01022_),
    .A(\u_tiny_nn_top.state_q[15] ),
    .Y(_01026_));
 sg13g2_nand2_1 _06498_ (.Y(_00012_),
    .A(_01025_),
    .B(_01026_));
 sg13g2_nor2b_2 _06499_ (.A(_01022_),
    .B_N(net1791),
    .Y(_01027_));
 sg13g2_nand2_1 _06500_ (.Y(_01028_),
    .A(net1854),
    .B(net1791));
 sg13g2_nor2_1 _06501_ (.A(net976),
    .B(_01027_),
    .Y(_01029_));
 sg13g2_nand2_1 _06502_ (.Y(_00011_),
    .A(_01028_),
    .B(_01029_));
 sg13g2_a21oi_1 _06503_ (.A1(_00660_),
    .A2(net676),
    .Y(_00010_),
    .B1(_00810_));
 sg13g2_a21oi_2 _06504_ (.B1(_00657_),
    .Y(_01030_),
    .A2(net1555),
    .A1(_00786_));
 sg13g2_nand3b_1 _06505_ (.B(_00785_),
    .C(net1861),
    .Y(_01031_),
    .A_N(net1855));
 sg13g2_inv_1 _06506_ (.Y(_01032_),
    .A(_01031_));
 sg13g2_nand2_1 _06507_ (.Y(_01033_),
    .A(_01030_),
    .B(_01031_));
 sg13g2_or2_1 _06508_ (.X(_01034_),
    .B(_01031_),
    .A(_00163_));
 sg13g2_nand3b_1 _06509_ (.B(_01033_),
    .C(_01034_),
    .Y(_00009_),
    .A_N(net884));
 sg13g2_nand2_1 _06510_ (.Y(_01035_),
    .A(\u_tiny_nn_top.state_q[14] ),
    .B(net1736));
 sg13g2_o21ai_1 _06511_ (.B1(_01035_),
    .Y(_00008_),
    .A1(net489),
    .A2(_01023_));
 sg13g2_nor2_2 _06512_ (.A(_00803_),
    .B(_00809_),
    .Y(_01036_));
 sg13g2_nand2_1 _06513_ (.Y(_01037_),
    .A(\u_tiny_nn_top.state_q[0] ),
    .B(_01036_));
 sg13g2_o21ai_1 _06514_ (.B1(_01037_),
    .Y(_00007_),
    .A1(net485),
    .A2(net1740));
 sg13g2_and2_1 _06515_ (.A(net1829),
    .B(_00797_),
    .X(_01038_));
 sg13g2_nand2_1 _06516_ (.Y(_01039_),
    .A(net1793),
    .B(_01038_));
 sg13g2_o21ai_1 _06517_ (.B1(_01039_),
    .Y(_00006_),
    .A1(_00655_),
    .A2(net1555));
 sg13g2_nor2_1 _06518_ (.A(net1768),
    .B(net1555),
    .Y(_01040_));
 sg13g2_nand2_2 _06519_ (.Y(_01041_),
    .A(net1790),
    .B(net1739));
 sg13g2_nor2b_2 _06520_ (.A(_01040_),
    .B_N(_01041_),
    .Y(_01042_));
 sg13g2_nand2b_1 _06521_ (.Y(_00005_),
    .B(_01042_),
    .A_N(net521));
 sg13g2_nand2_1 _06522_ (.Y(_01043_),
    .A(net1791),
    .B(net1555));
 sg13g2_nand3_1 _06523_ (.B(net491),
    .C(net1555),
    .A(net1792),
    .Y(_01044_));
 sg13g2_or4_2 _06524_ (.A(net806),
    .B(_00776_),
    .C(_00779_),
    .D(_00956_),
    .X(_01045_));
 sg13g2_nand2b_1 _06525_ (.Y(_01046_),
    .B(_00956_),
    .A_N(_00777_));
 sg13g2_nand3_1 _06526_ (.B(net1736),
    .C(_00957_),
    .A(\u_tiny_nn_top.state_q[10] ),
    .Y(_01047_));
 sg13g2_nand3_1 _06527_ (.B(_01045_),
    .C(_01047_),
    .A(_01044_),
    .Y(_00004_));
 sg13g2_nor2_2 _06528_ (.A(_00652_),
    .B(net1797),
    .Y(_01048_));
 sg13g2_nand3_1 _06529_ (.B(net1793),
    .C(_00792_),
    .A(net1828),
    .Y(_01049_));
 sg13g2_nand2b_1 _06530_ (.Y(_00016_),
    .B(_01049_),
    .A_N(_01048_));
 sg13g2_a21oi_1 _06531_ (.A1(_00660_),
    .A2(net487),
    .Y(_00015_),
    .B1(_00808_));
 sg13g2_a22oi_1 _06532_ (.Y(_01050_),
    .B1(net1555),
    .B2(net1790),
    .A2(net1765),
    .A1(net983));
 sg13g2_nor2_1 _06533_ (.A(net1739),
    .B(net984),
    .Y(_00014_));
 sg13g2_nand2_2 _06534_ (.Y(_01051_),
    .A(net1779),
    .B(_00797_));
 sg13g2_nor2_1 _06535_ (.A(_00660_),
    .B(_01051_),
    .Y(_00001_));
 sg13g2_nand2_1 _06536_ (.Y(_01052_),
    .A(net1793),
    .B(_00796_));
 sg13g2_nor2_1 _06537_ (.A(net1828),
    .B(_01052_),
    .Y(_00000_));
 sg13g2_nor2_1 _06538_ (.A(net1780),
    .B(_01052_),
    .Y(_00003_));
 sg13g2_nor2_1 _06539_ (.A(_00655_),
    .B(_01023_),
    .Y(_00002_));
 sg13g2_nor2_1 _06540_ (.A(net1830),
    .B(_01052_),
    .Y(_01053_));
 sg13g2_a21oi_1 _06541_ (.A1(_00774_),
    .A2(_01052_),
    .Y(_00188_),
    .B1(_01053_));
 sg13g2_nor3_1 _06542_ (.A(net674),
    .B(net1791),
    .C(net884),
    .Y(_01054_));
 sg13g2_a22oi_1 _06543_ (.Y(_01055_),
    .B1(_01054_),
    .B2(_00660_),
    .A2(_01051_),
    .A1(_00799_));
 sg13g2_nor2b_1 _06544_ (.A(_01051_),
    .B_N(_01054_),
    .Y(_01056_));
 sg13g2_nor2b_2 _06545_ (.A(net1854),
    .B_N(net1791),
    .Y(_01057_));
 sg13g2_a21oi_1 _06546_ (.A1(net1801),
    .A2(_01048_),
    .Y(_01058_),
    .B1(_01057_));
 sg13g2_nand2b_1 _06547_ (.Y(_01059_),
    .B(_01058_),
    .A_N(_01056_));
 sg13g2_mux2_1 _06548_ (.A0(net1864),
    .A1(_01059_),
    .S(_01055_),
    .X(_00189_));
 sg13g2_a21o_2 _06549_ (.A2(_00797_),
    .A1(net1793),
    .B1(_00000_),
    .X(_01060_));
 sg13g2_nor2_1 _06550_ (.A(net839),
    .B(net1554),
    .Y(_01061_));
 sg13g2_a21oi_1 _06551_ (.A1(net1770),
    .A2(net1554),
    .Y(_00190_),
    .B1(_01061_));
 sg13g2_mux2_1 _06552_ (.A0(net784),
    .A1(net1851),
    .S(net1554),
    .X(_00191_));
 sg13g2_nor2_1 _06553_ (.A(net760),
    .B(net1554),
    .Y(_01062_));
 sg13g2_a21oi_1 _06554_ (.A1(net1772),
    .A2(net1554),
    .Y(_00192_),
    .B1(_01062_));
 sg13g2_mux2_1 _06555_ (.A0(net827),
    .A1(\u_tiny_nn_top.data_i_q[3] ),
    .S(net1554),
    .X(_00193_));
 sg13g2_mux2_1 _06556_ (.A0(net759),
    .A1(net1845),
    .S(_01060_),
    .X(_00194_));
 sg13g2_mux2_1 _06557_ (.A0(net761),
    .A1(net1842),
    .S(_01060_),
    .X(_00195_));
 sg13g2_mux2_1 _06558_ (.A0(net799),
    .A1(net1839),
    .S(net1554),
    .X(_00196_));
 sg13g2_mux2_1 _06559_ (.A0(net808),
    .A1(net1836),
    .S(net1554),
    .X(_00197_));
 sg13g2_nor2_2 _06560_ (.A(net1792),
    .B(net1764),
    .Y(_01063_));
 sg13g2_and2_1 _06561_ (.A(_00839_),
    .B(_01063_),
    .X(_01064_));
 sg13g2_nor2_1 _06562_ (.A(net1793),
    .B(_00837_),
    .Y(_01065_));
 sg13g2_a21oi_1 _06563_ (.A1(_01064_),
    .A2(_01065_),
    .Y(_01066_),
    .B1(_00798_));
 sg13g2_nand4_1 _06564_ (.B(_01024_),
    .C(_01028_),
    .A(_00811_),
    .Y(_01067_),
    .D(_01066_));
 sg13g2_and3_2 _06565_ (.X(_01068_),
    .A(_00162_),
    .B(_00836_),
    .C(_01064_));
 sg13g2_nand3_1 _06566_ (.B(_00836_),
    .C(_01064_),
    .A(_00162_),
    .Y(_01069_));
 sg13g2_nor2_2 _06567_ (.A(\u_tiny_nn_top.state_q[4] ),
    .B(net1765),
    .Y(_01070_));
 sg13g2_nor3_1 _06568_ (.A(net1791),
    .B(\u_tiny_nn_top.state_q[17] ),
    .C(_01070_),
    .Y(_01071_));
 sg13g2_nand3b_1 _06569_ (.B(_00099_),
    .C(net1740),
    .Y(_01072_),
    .A_N(\u_tiny_nn_top.state_q[17] ));
 sg13g2_o21ai_1 _06570_ (.B1(_01072_),
    .Y(_01073_),
    .A1(_00099_),
    .A2(net1740));
 sg13g2_nand2_1 _06571_ (.Y(_01074_),
    .A(net1738),
    .B(_00836_));
 sg13g2_o21ai_1 _06572_ (.B1(_01069_),
    .Y(_01075_),
    .A1(net1857),
    .A2(_00836_));
 sg13g2_a21oi_1 _06573_ (.A1(_01043_),
    .A2(_01073_),
    .Y(_01076_),
    .B1(_01071_));
 sg13g2_a221oi_1 _06574_ (.B2(_01042_),
    .C1(net1857),
    .B1(_00838_),
    .A1(net1112),
    .Y(_01077_),
    .A2(net1738));
 sg13g2_nor3_1 _06575_ (.A(_01075_),
    .B(_01076_),
    .C(_01077_),
    .Y(_01078_));
 sg13g2_o21ai_1 _06576_ (.B1(\u_tiny_nn_top.data_i_q[0] ),
    .Y(_01079_),
    .A1(_00795_),
    .A2(_01038_));
 sg13g2_o21ai_1 _06577_ (.B1(_01079_),
    .Y(_01080_),
    .A1(_00797_),
    .A2(_01036_));
 sg13g2_nor2_1 _06578_ (.A(_01069_),
    .B(_01080_),
    .Y(_01081_));
 sg13g2_nor3_1 _06579_ (.A(net1503),
    .B(_01078_),
    .C(_01081_),
    .Y(_01082_));
 sg13g2_a21o_1 _06580_ (.A2(net1503),
    .A1(net1857),
    .B1(_01082_),
    .X(_00198_));
 sg13g2_nand2_1 _06581_ (.Y(_01083_),
    .A(net1856),
    .B(net1503));
 sg13g2_a22oi_1 _06582_ (.Y(_01084_),
    .B1(_01046_),
    .B2(_00840_),
    .A2(net1555),
    .A1(net1790));
 sg13g2_a22oi_1 _06583_ (.Y(_01085_),
    .B1(_01026_),
    .B2(_01084_),
    .A2(net1739),
    .A1(_00102_));
 sg13g2_a21oi_1 _06584_ (.A1(_00164_),
    .A2(net1764),
    .Y(_01086_),
    .B1(net1791));
 sg13g2_nor2_1 _06585_ (.A(net1739),
    .B(_01086_),
    .Y(_01087_));
 sg13g2_o21ai_1 _06586_ (.B1(_01046_),
    .Y(_01088_),
    .A1(_00837_),
    .A2(_01087_));
 sg13g2_nand3_1 _06587_ (.B(_01069_),
    .C(_01088_),
    .A(_01043_),
    .Y(_01089_));
 sg13g2_nor2_1 _06588_ (.A(_01085_),
    .B(_01089_),
    .Y(_01090_));
 sg13g2_a22oi_1 _06589_ (.Y(_01091_),
    .B1(_00803_),
    .B2(_00795_),
    .A2(_00796_),
    .A1(net1829));
 sg13g2_nor2_1 _06590_ (.A(_00101_),
    .B(_00809_),
    .Y(_01092_));
 sg13g2_a21oi_1 _06591_ (.A1(net1849),
    .A2(_01038_),
    .Y(_01093_),
    .B1(_01092_));
 sg13g2_nand4_1 _06592_ (.B(_01068_),
    .C(_01091_),
    .A(_01051_),
    .Y(_01094_),
    .D(_01093_));
 sg13g2_nand2b_1 _06593_ (.Y(_01095_),
    .B(_01094_),
    .A_N(net1503));
 sg13g2_o21ai_1 _06594_ (.B1(_01083_),
    .Y(_00199_),
    .A1(_01090_),
    .A2(_01095_));
 sg13g2_xor2_1 _06595_ (.B(_00777_),
    .A(_00103_),
    .X(_01096_));
 sg13g2_nor2_1 _06596_ (.A(\u_tiny_nn_top.state_q[14] ),
    .B(_01027_),
    .Y(_01097_));
 sg13g2_a21oi_1 _06597_ (.A1(_00103_),
    .A2(net1738),
    .Y(_01098_),
    .B1(_01097_));
 sg13g2_nor2_2 _06598_ (.A(\u_tiny_nn_top.state_q[12] ),
    .B(_01030_),
    .Y(_01099_));
 sg13g2_a22oi_1 _06599_ (.Y(_01100_),
    .B1(_01042_),
    .B2(_01099_),
    .A2(net1738),
    .A1(_00104_));
 sg13g2_nor2_1 _06600_ (.A(_01098_),
    .B(_01100_),
    .Y(_01101_));
 sg13g2_a21oi_1 _06601_ (.A1(net1736),
    .A2(_01096_),
    .Y(_01102_),
    .B1(_01101_));
 sg13g2_a221oi_1 _06602_ (.B2(net1738),
    .C1(_01096_),
    .B1(_00836_),
    .A1(_00832_),
    .Y(_01103_),
    .A2(_00834_));
 sg13g2_nor4_1 _06603_ (.A(\u_tiny_nn_top.state_q[4] ),
    .B(_01068_),
    .C(_01102_),
    .D(_01103_),
    .Y(_01104_));
 sg13g2_or2_2 _06604_ (.X(_01105_),
    .B(_01038_),
    .A(_01036_));
 sg13g2_a21oi_1 _06605_ (.A1(\u_tiny_nn_top.data_i_q[2] ),
    .A2(_01105_),
    .Y(_01106_),
    .B1(_01069_));
 sg13g2_nor3_1 _06606_ (.A(net1503),
    .B(_01104_),
    .C(_01106_),
    .Y(_01107_));
 sg13g2_a21o_1 _06607_ (.A2(net1503),
    .A1(net1048),
    .B1(_01107_),
    .X(_00200_));
 sg13g2_nor2_2 _06608_ (.A(_01027_),
    .B(_01070_),
    .Y(_01108_));
 sg13g2_a21oi_1 _06609_ (.A1(_00105_),
    .A2(net1738),
    .Y(_01109_),
    .B1(_01108_));
 sg13g2_nand2b_1 _06610_ (.Y(_01110_),
    .B(_00840_),
    .A_N(_00106_));
 sg13g2_xor2_1 _06611_ (.B(_00778_),
    .A(_00105_),
    .X(_01111_));
 sg13g2_a22oi_1 _06612_ (.Y(_01112_),
    .B1(_01042_),
    .B2(_01099_),
    .A2(net1738),
    .A1(_00106_));
 sg13g2_a21oi_1 _06613_ (.A1(_00837_),
    .A2(_01074_),
    .Y(_01113_),
    .B1(_01112_));
 sg13g2_a21oi_1 _06614_ (.A1(_01110_),
    .A2(_01111_),
    .Y(_01114_),
    .B1(_01113_));
 sg13g2_a21oi_1 _06615_ (.A1(net1736),
    .A2(_01111_),
    .Y(_01115_),
    .B1(_01068_));
 sg13g2_o21ai_1 _06616_ (.B1(_01115_),
    .Y(_01116_),
    .A1(_01109_),
    .A2(_01114_));
 sg13g2_nand3_1 _06617_ (.B(_01068_),
    .C(_01105_),
    .A(net1848),
    .Y(_01117_));
 sg13g2_nor2b_1 _06618_ (.A(net1503),
    .B_N(_01117_),
    .Y(_01118_));
 sg13g2_a22oi_1 _06619_ (.Y(_00201_),
    .B1(_01116_),
    .B2(_01118_),
    .A2(net1503),
    .A1(_00654_));
 sg13g2_a21oi_1 _06620_ (.A1(\u_tiny_nn_top.state_q[12] ),
    .A2(net1736),
    .Y(_01119_),
    .B1(_01030_));
 sg13g2_nor2_1 _06621_ (.A(_00837_),
    .B(_01040_),
    .Y(_01120_));
 sg13g2_nand3_1 _06622_ (.B(_01119_),
    .C(_01120_),
    .A(_01108_),
    .Y(_01121_));
 sg13g2_nand2_1 _06623_ (.Y(_01122_),
    .A(_01074_),
    .B(_01121_));
 sg13g2_xnor2_1 _06624_ (.Y(_01123_),
    .A(_00107_),
    .B(_00781_));
 sg13g2_nor2_1 _06625_ (.A(_01122_),
    .B(_01123_),
    .Y(_01124_));
 sg13g2_o21ai_1 _06626_ (.B1(net1739),
    .Y(_01125_),
    .A1(_01027_),
    .A2(_01070_));
 sg13g2_nor2_1 _06627_ (.A(_00107_),
    .B(_01125_),
    .Y(_01126_));
 sg13g2_nor3_1 _06628_ (.A(_00108_),
    .B(net1737),
    .C(_00839_),
    .Y(_01127_));
 sg13g2_nor4_1 _06629_ (.A(_01068_),
    .B(_01124_),
    .C(_01126_),
    .D(_01127_),
    .Y(_01128_));
 sg13g2_a21oi_1 _06630_ (.A1(net1845),
    .A2(_01105_),
    .Y(_01129_),
    .B1(_01069_));
 sg13g2_nor3_1 _06631_ (.A(net1504),
    .B(_01128_),
    .C(_01129_),
    .Y(_01130_));
 sg13g2_a21o_1 _06632_ (.A2(net1504),
    .A1(net1053),
    .B1(_01130_),
    .X(_00202_));
 sg13g2_a22oi_1 _06633_ (.Y(_01131_),
    .B1(_01099_),
    .B2(_01120_),
    .A2(_00836_),
    .A1(net1738));
 sg13g2_nor2b_1 _06634_ (.A(_01131_),
    .B_N(_01108_),
    .Y(_01132_));
 sg13g2_nor2_1 _06635_ (.A(\u_tiny_nn_top.counter_q[4] ),
    .B(_00781_),
    .Y(_01133_));
 sg13g2_nor3_1 _06636_ (.A(\u_tiny_nn_top.counter_q[4] ),
    .B(_00109_),
    .C(_00781_),
    .Y(_01134_));
 sg13g2_nand2_1 _06637_ (.Y(_01135_),
    .A(_01074_),
    .B(_01133_));
 sg13g2_a221oi_1 _06638_ (.B2(_00109_),
    .C1(_01132_),
    .B1(_01135_),
    .A1(_01125_),
    .Y(_01136_),
    .A2(_01134_));
 sg13g2_nor3_1 _06639_ (.A(_00110_),
    .B(net1737),
    .C(_00839_),
    .Y(_01137_));
 sg13g2_nor3_1 _06640_ (.A(_01068_),
    .B(_01136_),
    .C(_01137_),
    .Y(_01138_));
 sg13g2_a21oi_1 _06641_ (.A1(net1842),
    .A2(_01105_),
    .Y(_01139_),
    .B1(_01069_));
 sg13g2_nor3_1 _06642_ (.A(net1504),
    .B(_01138_),
    .C(_01139_),
    .Y(_01140_));
 sg13g2_a21o_1 _06643_ (.A2(net1504),
    .A1(net1024),
    .B1(_01140_),
    .X(_00203_));
 sg13g2_nand2b_2 _06644_ (.Y(_01141_),
    .B(_01133_),
    .A_N(\u_tiny_nn_top.counter_q[5] ));
 sg13g2_xor2_1 _06645_ (.B(_01141_),
    .A(_00111_),
    .X(_01142_));
 sg13g2_nand2_1 _06646_ (.Y(_01143_),
    .A(_01131_),
    .B(_01142_));
 sg13g2_nor2_1 _06647_ (.A(_00775_),
    .B(_01141_),
    .Y(_01144_));
 sg13g2_xor2_1 _06648_ (.B(_01144_),
    .A(_00111_),
    .X(_01145_));
 sg13g2_nor3_1 _06649_ (.A(_00112_),
    .B(net1737),
    .C(_00839_),
    .Y(_01146_));
 sg13g2_o21ai_1 _06650_ (.B1(_01069_),
    .Y(_01147_),
    .A1(_01108_),
    .A2(_01145_));
 sg13g2_nor2_1 _06651_ (.A(_01146_),
    .B(_01147_),
    .Y(_01148_));
 sg13g2_a22oi_1 _06652_ (.Y(_01149_),
    .B1(_01038_),
    .B2(_00672_),
    .A2(_01036_),
    .A1(net1837));
 sg13g2_a221oi_1 _06653_ (.B2(_01068_),
    .C1(net1504),
    .B1(_01149_),
    .A1(_01143_),
    .Y(_01150_),
    .A2(_01148_));
 sg13g2_a21o_1 _06654_ (.A2(net1504),
    .A1(net1039),
    .B1(_01150_),
    .X(_00204_));
 sg13g2_nor2_1 _06655_ (.A(\u_tiny_nn_top.counter_q[6] ),
    .B(_01141_),
    .Y(_01151_));
 sg13g2_and2_1 _06656_ (.A(_01125_),
    .B(_01151_),
    .X(_01152_));
 sg13g2_nor3_1 _06657_ (.A(_00113_),
    .B(_01132_),
    .C(_01152_),
    .Y(_01153_));
 sg13g2_nor4_1 _06658_ (.A(\u_tiny_nn_top.counter_q[6] ),
    .B(_00722_),
    .C(_01122_),
    .D(_01141_),
    .Y(_01154_));
 sg13g2_nor3_1 _06659_ (.A(_00114_),
    .B(net1737),
    .C(_00839_),
    .Y(_01155_));
 sg13g2_nor4_1 _06660_ (.A(_01068_),
    .B(_01153_),
    .C(_01154_),
    .D(_01155_),
    .Y(_01156_));
 sg13g2_a21oi_1 _06661_ (.A1(net1836),
    .A2(_01105_),
    .Y(_01157_),
    .B1(_01069_));
 sg13g2_nor3_1 _06662_ (.A(net1504),
    .B(_01156_),
    .C(_01157_),
    .Y(_01158_));
 sg13g2_a21o_1 _06663_ (.A2(net1504),
    .A1(net1008),
    .B1(_01158_),
    .X(_00205_));
 sg13g2_nor2_1 _06664_ (.A(_00662_),
    .B(_01063_),
    .Y(_00206_));
 sg13g2_nand2_1 _06665_ (.Y(_01159_),
    .A(net704),
    .B(net1724));
 sg13g2_mux2_1 _06666_ (.A0(_00644_),
    .A1(_00668_),
    .S(net1479),
    .X(_01160_));
 sg13g2_o21ai_1 _06667_ (.B1(_01159_),
    .Y(_00207_),
    .A1(net1724),
    .A2(_01160_));
 sg13g2_nand2_1 _06668_ (.Y(_01161_),
    .A(net877),
    .B(net1724));
 sg13g2_mux2_1 _06669_ (.A0(net1774),
    .A1(_00669_),
    .S(net1479),
    .X(_01162_));
 sg13g2_o21ai_1 _06670_ (.B1(_01161_),
    .Y(_00208_),
    .A1(net1725),
    .A2(_01162_));
 sg13g2_nand2_1 _06671_ (.Y(_01163_),
    .A(net901),
    .B(net1725));
 sg13g2_nor2b_1 _06672_ (.A(\u_tiny_nn_top.max_val_q[10] ),
    .B_N(net1479),
    .Y(_01164_));
 sg13g2_o21ai_1 _06673_ (.B1(_00927_),
    .Y(_01165_),
    .A1(\u_tiny_nn_top.data_i_q[10] ),
    .A2(net1480));
 sg13g2_o21ai_1 _06674_ (.B1(_01163_),
    .Y(_00209_),
    .A1(_01164_),
    .A2(_01165_));
 sg13g2_nand2_1 _06675_ (.Y(_01166_),
    .A(net835),
    .B(net1725));
 sg13g2_nor2b_1 _06676_ (.A(\u_tiny_nn_top.max_val_q[11] ),
    .B_N(net1479),
    .Y(_01167_));
 sg13g2_o21ai_1 _06677_ (.B1(_00927_),
    .Y(_01168_),
    .A1(\u_tiny_nn_top.data_i_q[11] ),
    .A2(net1480));
 sg13g2_o21ai_1 _06678_ (.B1(_01166_),
    .Y(_00210_),
    .A1(_01167_),
    .A2(_01168_));
 sg13g2_nand2_1 _06679_ (.Y(_01169_),
    .A(net829),
    .B(net1724));
 sg13g2_mux2_1 _06680_ (.A0(net1780),
    .A1(_00671_),
    .S(net1479),
    .X(_01170_));
 sg13g2_o21ai_1 _06681_ (.B1(_01169_),
    .Y(_00211_),
    .A1(net1724),
    .A2(_01170_));
 sg13g2_nand2_1 _06682_ (.Y(_01171_),
    .A(net773),
    .B(net1725));
 sg13g2_mux2_1 _06683_ (.A0(net1781),
    .A1(_00670_),
    .S(net1479),
    .X(_01172_));
 sg13g2_o21ai_1 _06684_ (.B1(_01171_),
    .Y(_00212_),
    .A1(net1724),
    .A2(_01172_));
 sg13g2_nand2_1 _06685_ (.Y(_01173_),
    .A(net852),
    .B(net1724));
 sg13g2_nor2b_1 _06686_ (.A(\u_tiny_nn_top.max_val_q[14] ),
    .B_N(net1479),
    .Y(_01174_));
 sg13g2_o21ai_1 _06687_ (.B1(_00927_),
    .Y(_01175_),
    .A1(net1827),
    .A2(net1480));
 sg13g2_o21ai_1 _06688_ (.B1(_01173_),
    .Y(_00213_),
    .A1(_01174_),
    .A2(_01175_));
 sg13g2_nand2_1 _06689_ (.Y(_01176_),
    .A(net936),
    .B(net1724));
 sg13g2_nor2b_1 _06690_ (.A(\u_tiny_nn_top.max_val_q[15] ),
    .B_N(net1479),
    .Y(_01177_));
 sg13g2_o21ai_1 _06691_ (.B1(_00927_),
    .Y(_01178_),
    .A1(net1823),
    .A2(net1480));
 sg13g2_o21ai_1 _06692_ (.B1(_01176_),
    .Y(_00214_),
    .A1(_01177_),
    .A2(_01178_));
 sg13g2_nor4_1 _06693_ (.A(_00658_),
    .B(_00776_),
    .C(_00779_),
    .D(_00784_),
    .Y(_01179_));
 sg13g2_or4_2 _06694_ (.A(_00658_),
    .B(_00776_),
    .C(_00779_),
    .D(_00784_),
    .X(_01180_));
 sg13g2_a21o_1 _06695_ (.A2(_00658_),
    .A1(_00657_),
    .B1(_01034_),
    .X(_01181_));
 sg13g2_and2_1 _06696_ (.A(_01180_),
    .B(_01181_),
    .X(_01182_));
 sg13g2_nand2_2 _06697_ (.Y(_01183_),
    .A(_01180_),
    .B(_01181_));
 sg13g2_o21ai_1 _06698_ (.B1(net1854),
    .Y(_01184_),
    .A1(\u_tiny_nn_top.state_q[4] ),
    .A2(\u_tiny_nn_top.state_q[14] ));
 sg13g2_nand2b_1 _06699_ (.Y(_01185_),
    .B(_00786_),
    .A_N(_00831_));
 sg13g2_and2_1 _06700_ (.A(_00161_),
    .B(_00831_),
    .X(_01186_));
 sg13g2_a21o_2 _06701_ (.A2(_01185_),
    .A1(_01041_),
    .B1(_01186_),
    .X(_01187_));
 sg13g2_a21oi_2 _06702_ (.B1(_01186_),
    .Y(_01188_),
    .A2(_01185_),
    .A1(_01041_));
 sg13g2_and3_1 _06703_ (.X(_01189_),
    .A(_01182_),
    .B(net1762),
    .C(_01187_));
 sg13g2_or4_1 _06704_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[3] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[2] ),
    .C(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[5] ),
    .D(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[4] ),
    .X(_01190_));
 sg13g2_nor3_1 _06705_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[1] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[0] ),
    .C(_01190_),
    .Y(_01191_));
 sg13g2_nor3_1 _06706_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[12] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[11] ),
    .C(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[14] ),
    .Y(_01192_));
 sg13g2_nor4_1 _06707_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[8] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[7] ),
    .C(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[10] ),
    .D(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[9] ),
    .Y(_01193_));
 sg13g2_nand3_1 _06708_ (.B(_01192_),
    .C(_01193_),
    .A(_00702_),
    .Y(_01194_));
 sg13g2_nand3_1 _06709_ (.B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[11] ),
    .C(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[14] ),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[12] ),
    .Y(_01195_));
 sg13g2_nand4_1 _06710_ (.B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[7] ),
    .C(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[10] ),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[8] ),
    .Y(_01196_),
    .D(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[9] ));
 sg13g2_nor3_1 _06711_ (.A(_00702_),
    .B(_01195_),
    .C(_01196_),
    .Y(_01197_));
 sg13g2_inv_1 _06712_ (.Y(_01198_),
    .A(_01197_));
 sg13g2_a22oi_1 _06713_ (.Y(_01199_),
    .B1(_01194_),
    .B2(_01198_),
    .A2(_01191_),
    .A1(_00071_));
 sg13g2_nor2_1 _06714_ (.A(_00695_),
    .B(_01194_),
    .Y(_01200_));
 sg13g2_o21ai_1 _06715_ (.B1(_00826_),
    .Y(_01201_),
    .A1(_00776_),
    .A2(_00781_));
 sg13g2_nand4_1 _06716_ (.B(_00662_),
    .C(_00775_),
    .A(net1791),
    .Y(_01202_),
    .D(_00780_));
 sg13g2_and4_2 _06717_ (.A(_01045_),
    .B(_01180_),
    .C(_01201_),
    .D(_01202_),
    .X(_01203_));
 sg13g2_nand4_1 _06718_ (.B(_01180_),
    .C(_01201_),
    .A(_01045_),
    .Y(_01204_),
    .D(_01202_));
 sg13g2_nor2_1 _06719_ (.A(net1792),
    .B(\u_tiny_nn_top.state_q[10] ),
    .Y(_01205_));
 sg13g2_nor4_2 _06720_ (.A(\u_tiny_nn_top.state_q[3] ),
    .B(net1792),
    .C(\u_tiny_nn_top.state_q[10] ),
    .Y(_01206_),
    .D(_00826_));
 sg13g2_nand3_1 _06721_ (.B(net1763),
    .C(_01205_),
    .A(_00658_),
    .Y(_01207_));
 sg13g2_nand2_1 _06722_ (.Y(_01208_),
    .A(_01204_),
    .B(_01207_));
 sg13g2_mux2_2 _06723_ (.A0(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][6] ),
    .A1(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][6] ),
    .S(net1672),
    .X(_01209_));
 sg13g2_nand2b_1 _06724_ (.Y(_01210_),
    .B(net1671),
    .A_N(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][5] ));
 sg13g2_o21ai_1 _06725_ (.B1(_01210_),
    .Y(_01211_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][5] ),
    .A2(net1671));
 sg13g2_mux2_1 _06726_ (.A0(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][5] ),
    .A1(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][5] ),
    .S(net1671),
    .X(_01212_));
 sg13g2_nand2b_1 _06727_ (.Y(_01213_),
    .B(net1672),
    .A_N(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][4] ));
 sg13g2_o21ai_1 _06728_ (.B1(_01213_),
    .Y(_01214_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][4] ),
    .A2(net1672));
 sg13g2_nand3b_1 _06729_ (.B(_01211_),
    .C(_01214_),
    .Y(_01215_),
    .A_N(_01209_));
 sg13g2_nand2b_1 _06730_ (.Y(_01216_),
    .B(net1672),
    .A_N(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][3] ));
 sg13g2_o21ai_1 _06731_ (.B1(_01216_),
    .Y(_01217_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][3] ),
    .A2(net1672));
 sg13g2_inv_1 _06732_ (.Y(_01218_),
    .A(_01217_));
 sg13g2_mux2_2 _06733_ (.A0(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][0] ),
    .A1(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][0] ),
    .S(net1672),
    .X(_01219_));
 sg13g2_mux2_2 _06734_ (.A0(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][1] ),
    .A1(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][1] ),
    .S(net1671),
    .X(_01220_));
 sg13g2_nand2b_1 _06735_ (.Y(_01221_),
    .B(net1671),
    .A_N(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][2] ));
 sg13g2_o21ai_1 _06736_ (.B1(_01221_),
    .Y(_01222_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][2] ),
    .A2(net1672));
 sg13g2_inv_1 _06737_ (.Y(_01223_),
    .A(_01222_));
 sg13g2_nand2b_1 _06738_ (.Y(_01224_),
    .B(_01222_),
    .A_N(_01220_));
 sg13g2_nor4_2 _06739_ (.A(_01215_),
    .B(_01218_),
    .C(_01219_),
    .Y(_01225_),
    .D(_01224_));
 sg13g2_nand2b_1 _06740_ (.Y(_01226_),
    .B(net1671),
    .A_N(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][15] ));
 sg13g2_o21ai_1 _06741_ (.B1(_01226_),
    .Y(_01227_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][15] ),
    .A2(net1671));
 sg13g2_mux2_2 _06742_ (.A0(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][15] ),
    .A1(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][15] ),
    .S(net1671),
    .X(_01228_));
 sg13g2_and2_1 _06743_ (.A(_01225_),
    .B(_01227_),
    .X(_01229_));
 sg13g2_a21oi_2 _06744_ (.B1(_00058_),
    .Y(_01230_),
    .A2(_01207_),
    .A1(_01204_));
 sg13g2_nor3_2 _06745_ (.A(_00057_),
    .B(_01203_),
    .C(_01206_),
    .Y(_01231_));
 sg13g2_or2_1 _06746_ (.X(_01232_),
    .B(_01231_),
    .A(_01230_));
 sg13g2_nor2_2 _06747_ (.A(_01230_),
    .B(_01231_),
    .Y(_01233_));
 sg13g2_nor3_2 _06748_ (.A(_00676_),
    .B(_01203_),
    .C(_01206_),
    .Y(_01234_));
 sg13g2_a21oi_2 _06749_ (.B1(_01234_),
    .Y(_01235_),
    .A2(net1673),
    .A1(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][7] ));
 sg13g2_a21o_1 _06750_ (.A2(net1673),
    .A1(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][7] ),
    .B1(_01234_),
    .X(_01236_));
 sg13g2_mux2_2 _06751_ (.A0(_00061_),
    .A1(_00062_),
    .S(net1673),
    .X(_01237_));
 sg13g2_nand3_1 _06752_ (.B(_01204_),
    .C(_01207_),
    .A(_00065_),
    .Y(_01238_));
 sg13g2_o21ai_1 _06753_ (.B1(_00066_),
    .Y(_01239_),
    .A1(_01203_),
    .A2(_01206_));
 sg13g2_and2_2 _06754_ (.A(_01238_),
    .B(_01239_),
    .X(_01240_));
 sg13g2_nand2_1 _06755_ (.Y(_01241_),
    .A(_01238_),
    .B(_01239_));
 sg13g2_nand4_1 _06756_ (.B(_01235_),
    .C(_01237_),
    .A(_01233_),
    .Y(_01242_),
    .D(_01241_));
 sg13g2_nand3_1 _06757_ (.B(_01204_),
    .C(_01207_),
    .A(_00067_),
    .Y(_01243_));
 sg13g2_o21ai_1 _06758_ (.B1(_00068_),
    .Y(_01244_),
    .A1(_01203_),
    .A2(_01206_));
 sg13g2_nand2_2 _06759_ (.Y(_01245_),
    .A(_01243_),
    .B(_01244_));
 sg13g2_a21oi_2 _06760_ (.B1(_00064_),
    .Y(_01246_),
    .A2(_01207_),
    .A1(_01204_));
 sg13g2_nor3_2 _06761_ (.A(_00063_),
    .B(_01203_),
    .C(_01206_),
    .Y(_01247_));
 sg13g2_nor2_2 _06762_ (.A(_01246_),
    .B(_01247_),
    .Y(_01248_));
 sg13g2_mux2_2 _06763_ (.A0(_00059_),
    .A1(_00060_),
    .S(net1673),
    .X(_01249_));
 sg13g2_a21o_1 _06764_ (.A2(_01207_),
    .A1(_01204_),
    .B1(_00070_),
    .X(_01250_));
 sg13g2_nand3b_1 _06765_ (.B(_01204_),
    .C(_01207_),
    .Y(_01251_),
    .A_N(_00069_));
 sg13g2_and2_2 _06766_ (.A(_01250_),
    .B(_01251_),
    .X(_01252_));
 sg13g2_nand4_1 _06767_ (.B(_01248_),
    .C(_01249_),
    .A(_01245_),
    .Y(_01253_),
    .D(_01252_));
 sg13g2_nor2_1 _06768_ (.A(_01242_),
    .B(_01253_),
    .Y(_01254_));
 sg13g2_nor2b_1 _06769_ (.A(_01229_),
    .B_N(_01254_),
    .Y(_01255_));
 sg13g2_nor3_1 _06770_ (.A(_01199_),
    .B(_01200_),
    .C(_01255_),
    .Y(_01256_));
 sg13g2_nor4_1 _06771_ (.A(_01233_),
    .B(_01237_),
    .C(_01245_),
    .D(_01248_),
    .Y(_01257_));
 sg13g2_nor4_1 _06772_ (.A(_01235_),
    .B(_01241_),
    .C(_01249_),
    .D(_01252_),
    .Y(_01258_));
 sg13g2_nand2_1 _06773_ (.Y(_01259_),
    .A(_01257_),
    .B(_01258_));
 sg13g2_inv_1 _06774_ (.Y(_01260_),
    .A(_01259_));
 sg13g2_and2_2 _06775_ (.A(_01256_),
    .B(_01259_),
    .X(_01261_));
 sg13g2_inv_1 _06776_ (.Y(_01262_),
    .A(_01261_));
 sg13g2_a21o_1 _06777_ (.A2(_01256_),
    .A1(_01225_),
    .B1(_01261_),
    .X(_01263_));
 sg13g2_nand2_1 _06778_ (.Y(_01264_),
    .A(_01225_),
    .B(_01260_));
 sg13g2_nand2b_1 _06779_ (.Y(_01265_),
    .B(_01191_),
    .A_N(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[6] ));
 sg13g2_nor2_2 _06780_ (.A(_01198_),
    .B(_01265_),
    .Y(_01266_));
 sg13g2_xnor2_1 _06781_ (.Y(_01267_),
    .A(_00695_),
    .B(_01228_));
 sg13g2_nand4_1 _06782_ (.B(_01260_),
    .C(_01266_),
    .A(_01225_),
    .Y(_01268_),
    .D(_01267_));
 sg13g2_and2_2 _06783_ (.A(_01263_),
    .B(_01268_),
    .X(_01269_));
 sg13g2_nor3_1 _06784_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[15] ),
    .B(_01194_),
    .C(_01265_),
    .Y(_01270_));
 sg13g2_or3_2 _06785_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[15] ),
    .B(_01194_),
    .C(_01265_),
    .X(_01271_));
 sg13g2_xor2_1 _06786_ (.B(_01249_),
    .A(_00080_),
    .X(_01272_));
 sg13g2_inv_1 _06787_ (.Y(_01273_),
    .A(_01272_));
 sg13g2_nand2b_1 _06788_ (.Y(_01274_),
    .B(_01237_),
    .A_N(_00073_));
 sg13g2_xnor2_1 _06789_ (.Y(_01275_),
    .A(_00073_),
    .B(_01237_));
 sg13g2_nand2_1 _06790_ (.Y(_01276_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[8] ),
    .B(_01233_));
 sg13g2_nor2_1 _06791_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[8] ),
    .B(_01233_),
    .Y(_01277_));
 sg13g2_o21ai_1 _06792_ (.B1(_00696_),
    .Y(_01278_),
    .A1(_01230_),
    .A2(_01231_));
 sg13g2_xnor2_1 _06793_ (.Y(_01279_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[8] ),
    .B(_01232_));
 sg13g2_inv_1 _06794_ (.Y(_01280_),
    .A(_01279_));
 sg13g2_xnor2_1 _06795_ (.Y(_01281_),
    .A(_00074_),
    .B(_01235_));
 sg13g2_a21oi_2 _06796_ (.B1(_00703_),
    .Y(_01282_),
    .A2(_01251_),
    .A1(_01250_));
 sg13g2_and3_1 _06797_ (.X(_01283_),
    .A(_00703_),
    .B(_01250_),
    .C(_01251_));
 sg13g2_nor2_1 _06798_ (.A(_01282_),
    .B(_01283_),
    .Y(_01284_));
 sg13g2_a21oi_1 _06799_ (.A1(_01243_),
    .A2(_01244_),
    .Y(_01285_),
    .B1(_00701_));
 sg13g2_and3_1 _06800_ (.X(_01286_),
    .A(_00701_),
    .B(_01243_),
    .C(_01244_));
 sg13g2_nor2_1 _06801_ (.A(_01285_),
    .B(_01286_),
    .Y(_01287_));
 sg13g2_nor4_2 _06802_ (.A(_01282_),
    .B(_01283_),
    .C(_01285_),
    .Y(_01288_),
    .D(_01286_));
 sg13g2_nand3_1 _06803_ (.B(_01238_),
    .C(_01239_),
    .A(_00700_),
    .Y(_01289_));
 sg13g2_o21ai_1 _06804_ (.B1(_00699_),
    .Y(_01290_),
    .A1(_01246_),
    .A2(_01247_));
 sg13g2_and2_1 _06805_ (.A(_01289_),
    .B(_01290_),
    .X(_01291_));
 sg13g2_nor3_1 _06806_ (.A(_00699_),
    .B(_01246_),
    .C(_01247_),
    .Y(_01292_));
 sg13g2_a21oi_1 _06807_ (.A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[11] ),
    .A2(_01241_),
    .Y(_01293_),
    .B1(_01292_));
 sg13g2_and3_1 _06808_ (.X(_01294_),
    .A(_01288_),
    .B(_01291_),
    .C(_01293_));
 sg13g2_nand3_1 _06809_ (.B(_01291_),
    .C(_01293_),
    .A(_01288_),
    .Y(_01295_));
 sg13g2_nor2_1 _06810_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[10] ),
    .B(_01249_),
    .Y(_01296_));
 sg13g2_nand2_1 _06811_ (.Y(_01297_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[10] ),
    .B(_01249_));
 sg13g2_xnor2_1 _06812_ (.Y(_01298_),
    .A(_00697_),
    .B(_01249_));
 sg13g2_nand3_1 _06813_ (.B(_01235_),
    .C(_01278_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[7] ),
    .Y(_01299_));
 sg13g2_nand4_1 _06814_ (.B(_01276_),
    .C(_01298_),
    .A(_01275_),
    .Y(_01300_),
    .D(_01299_));
 sg13g2_nor2_1 _06815_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[9] ),
    .B(_01237_),
    .Y(_01301_));
 sg13g2_a21oi_1 _06816_ (.A1(_01297_),
    .A2(_01301_),
    .Y(_01302_),
    .B1(_01296_));
 sg13g2_a21oi_2 _06817_ (.B1(_01295_),
    .Y(_01303_),
    .A2(_01302_),
    .A1(_01300_));
 sg13g2_a21o_2 _06818_ (.A2(_01302_),
    .A1(_01300_),
    .B1(_01295_),
    .X(_01304_));
 sg13g2_and4_1 _06819_ (.A(_01275_),
    .B(_01279_),
    .C(_01281_),
    .D(_01298_),
    .X(_01305_));
 sg13g2_nand4_1 _06820_ (.B(_01279_),
    .C(_01281_),
    .A(_01275_),
    .Y(_01306_),
    .D(_01298_));
 sg13g2_a21oi_1 _06821_ (.A1(_01289_),
    .A2(_01290_),
    .Y(_01307_),
    .B1(_01292_));
 sg13g2_nor2_1 _06822_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[13] ),
    .B(_01252_),
    .Y(_01308_));
 sg13g2_nor2_1 _06823_ (.A(_00704_),
    .B(_01245_),
    .Y(_01309_));
 sg13g2_a21o_1 _06824_ (.A2(_01308_),
    .A1(_01287_),
    .B1(_01309_),
    .X(_01310_));
 sg13g2_a221oi_1 _06825_ (.B2(_01287_),
    .C1(_01309_),
    .B1(_01308_),
    .A1(_01288_),
    .Y(_01311_),
    .A2(_01307_));
 sg13g2_a221oi_1 _06826_ (.B2(_01288_),
    .C1(_01310_),
    .B1(_01307_),
    .A1(_01294_),
    .Y(_01312_),
    .A2(_01305_));
 sg13g2_o21ai_1 _06827_ (.B1(_01311_),
    .Y(_01313_),
    .A1(_01295_),
    .A2(_01306_));
 sg13g2_nor2_2 _06828_ (.A(_01303_),
    .B(_01313_),
    .Y(_01314_));
 sg13g2_nand2_1 _06829_ (.Y(_01315_),
    .A(_01304_),
    .B(_01312_));
 sg13g2_nand3_1 _06830_ (.B(_01304_),
    .C(_01312_),
    .A(_00074_),
    .Y(_01316_));
 sg13g2_o21ai_1 _06831_ (.B1(_01235_),
    .Y(_01317_),
    .A1(_01303_),
    .A2(_01313_));
 sg13g2_nand2_2 _06832_ (.Y(_01318_),
    .A(_01316_),
    .B(_01317_));
 sg13g2_a21oi_2 _06833_ (.B1(_01281_),
    .Y(_01319_),
    .A2(_01317_),
    .A1(_01316_));
 sg13g2_nand3_1 _06834_ (.B(_01304_),
    .C(_01312_),
    .A(_01232_),
    .Y(_01320_));
 sg13g2_nor3_1 _06835_ (.A(_00077_),
    .B(_01303_),
    .C(_01313_),
    .Y(_01321_));
 sg13g2_o21ai_1 _06836_ (.B1(_01320_),
    .Y(_01322_),
    .A1(_01277_),
    .A2(_01321_));
 sg13g2_o21ai_1 _06837_ (.B1(_01322_),
    .Y(_01323_),
    .A1(_01280_),
    .A2(_01319_));
 sg13g2_nor2_1 _06838_ (.A(_01274_),
    .B(net1495),
    .Y(_01324_));
 sg13g2_a221oi_1 _06839_ (.B2(_01275_),
    .C1(_01324_),
    .B1(_01323_),
    .A1(_01301_),
    .Y(_01325_),
    .A2(net1495));
 sg13g2_nand2b_1 _06840_ (.Y(_01326_),
    .B(_01272_),
    .A_N(_01325_));
 sg13g2_nor2_1 _06841_ (.A(_00082_),
    .B(net1496),
    .Y(_01327_));
 sg13g2_xnor2_1 _06842_ (.Y(_01328_),
    .A(_00082_),
    .B(_01240_));
 sg13g2_o21ai_1 _06843_ (.B1(_01328_),
    .Y(_01329_),
    .A1(_01289_),
    .A2(_01314_));
 sg13g2_nor2_1 _06844_ (.A(_01327_),
    .B(_01329_),
    .Y(_01330_));
 sg13g2_xor2_1 _06845_ (.B(_01248_),
    .A(_00081_),
    .X(_01331_));
 sg13g2_xnor2_1 _06846_ (.Y(_01332_),
    .A(_01330_),
    .B(_01331_));
 sg13g2_xnor2_1 _06847_ (.Y(_01333_),
    .A(_00075_),
    .B(_01245_));
 sg13g2_nand2_1 _06848_ (.Y(_01334_),
    .A(_00702_),
    .B(net1496));
 sg13g2_a22oi_1 _06849_ (.Y(_01335_),
    .B1(_01334_),
    .B2(_01282_),
    .A2(net1496),
    .A1(_01283_));
 sg13g2_xnor2_1 _06850_ (.Y(_01336_),
    .A(_01333_),
    .B(_01335_));
 sg13g2_nand2_1 _06851_ (.Y(_01337_),
    .A(_00080_),
    .B(_01314_));
 sg13g2_nand2b_1 _06852_ (.Y(_01338_),
    .B(net1495),
    .A_N(_01296_));
 sg13g2_a21oi_1 _06853_ (.A1(_01337_),
    .A2(_01338_),
    .Y(_01339_),
    .B1(_01273_));
 sg13g2_xnor2_1 _06854_ (.Y(_01340_),
    .A(_01328_),
    .B(_01339_));
 sg13g2_nor2_1 _06855_ (.A(_01290_),
    .B(_01314_),
    .Y(_01341_));
 sg13g2_o21ai_1 _06856_ (.B1(_01331_),
    .Y(_01342_),
    .A1(_00081_),
    .A2(net1496));
 sg13g2_nor3_1 _06857_ (.A(_01284_),
    .B(_01341_),
    .C(_01342_),
    .Y(_01343_));
 sg13g2_o21ai_1 _06858_ (.B1(_01284_),
    .Y(_01344_),
    .A1(_01341_),
    .A2(_01342_));
 sg13g2_nand2b_1 _06859_ (.Y(_01345_),
    .B(_01344_),
    .A_N(_01343_));
 sg13g2_and4_1 _06860_ (.A(_01332_),
    .B(_01336_),
    .C(_01340_),
    .D(_01345_),
    .X(_01346_));
 sg13g2_nand2_1 _06861_ (.Y(_01347_),
    .A(_01273_),
    .B(_01325_));
 sg13g2_nand3_1 _06862_ (.B(_01346_),
    .C(_01347_),
    .A(_01326_),
    .Y(_01348_));
 sg13g2_inv_1 _06863_ (.Y(_01349_),
    .A(_01348_));
 sg13g2_nand3_1 _06864_ (.B(_01304_),
    .C(_01312_),
    .A(_01228_),
    .Y(_01350_));
 sg13g2_mux2_2 _06865_ (.A0(_00076_),
    .A1(_01227_),
    .S(net1498),
    .X(_01351_));
 sg13g2_o21ai_1 _06866_ (.B1(_01350_),
    .Y(_01352_),
    .A1(_00076_),
    .A2(net1498));
 sg13g2_nand2_2 _06867_ (.Y(_01353_),
    .A(_01349_),
    .B(_01352_));
 sg13g2_nand2_1 _06868_ (.Y(_01354_),
    .A(_00076_),
    .B(net1498));
 sg13g2_o21ai_1 _06869_ (.B1(_01354_),
    .Y(_01355_),
    .A1(_01228_),
    .A2(net1497));
 sg13g2_inv_1 _06870_ (.Y(_01356_),
    .A(_01355_));
 sg13g2_a21oi_2 _06871_ (.B1(_01356_),
    .Y(_01357_),
    .A2(_01352_),
    .A1(_01349_));
 sg13g2_xnor2_1 _06872_ (.Y(_01358_),
    .A(_01353_),
    .B(_01355_));
 sg13g2_xor2_1 _06873_ (.B(_01323_),
    .A(_01275_),
    .X(_01359_));
 sg13g2_xnor2_1 _06874_ (.Y(_01360_),
    .A(_01275_),
    .B(_01323_));
 sg13g2_nor2_1 _06875_ (.A(_01348_),
    .B(net1476),
    .Y(_01361_));
 sg13g2_a21oi_2 _06876_ (.B1(_01348_),
    .Y(_01362_),
    .A2(net1476),
    .A1(_01351_));
 sg13g2_xnor2_1 _06877_ (.Y(_01363_),
    .A(_01279_),
    .B(_01319_));
 sg13g2_xnor2_1 _06878_ (.Y(_01364_),
    .A(_01280_),
    .B(_01319_));
 sg13g2_nor2_1 _06879_ (.A(_01352_),
    .B(_01364_),
    .Y(_01365_));
 sg13g2_xnor2_1 _06880_ (.Y(_01366_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[7] ),
    .B(_01236_));
 sg13g2_xnor2_1 _06881_ (.Y(_01367_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[7] ),
    .B(_01235_));
 sg13g2_nor2_1 _06882_ (.A(_01351_),
    .B(net1529),
    .Y(_01368_));
 sg13g2_mux2_1 _06883_ (.A0(_00079_),
    .A1(_01211_),
    .S(net1498),
    .X(_01369_));
 sg13g2_mux2_1 _06884_ (.A0(_00078_),
    .A1(_01214_),
    .S(net1498),
    .X(_01370_));
 sg13g2_and2_1 _06885_ (.A(_01369_),
    .B(_01370_),
    .X(_01371_));
 sg13g2_mux2_1 _06886_ (.A0(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[3] ),
    .A1(_01218_),
    .S(net1498),
    .X(_01372_));
 sg13g2_nand3_1 _06887_ (.B(_01304_),
    .C(_01312_),
    .A(_01219_),
    .Y(_01373_));
 sg13g2_o21ai_1 _06888_ (.B1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[0] ),
    .Y(_01374_),
    .A1(_01303_),
    .A2(_01313_));
 sg13g2_nand2_1 _06889_ (.Y(_01375_),
    .A(_01373_),
    .B(_01374_));
 sg13g2_nand3_1 _06890_ (.B(_01304_),
    .C(_01312_),
    .A(_01220_),
    .Y(_01376_));
 sg13g2_o21ai_1 _06891_ (.B1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[1] ),
    .Y(_01377_),
    .A1(_01303_),
    .A2(_01313_));
 sg13g2_nand2_1 _06892_ (.Y(_01378_),
    .A(_01376_),
    .B(_01377_));
 sg13g2_and4_1 _06893_ (.A(_01373_),
    .B(_01374_),
    .C(_01376_),
    .D(_01377_),
    .X(_01379_));
 sg13g2_nand4_1 _06894_ (.B(_01374_),
    .C(_01376_),
    .A(_01373_),
    .Y(_01380_),
    .D(_01377_));
 sg13g2_mux2_1 _06895_ (.A0(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[2] ),
    .A1(_01223_),
    .S(net1498),
    .X(_01381_));
 sg13g2_o21ai_1 _06896_ (.B1(_01352_),
    .Y(_01382_),
    .A1(_01380_),
    .A2(_01381_));
 sg13g2_nor3_2 _06897_ (.A(_01372_),
    .B(_01380_),
    .C(_01381_),
    .Y(_01383_));
 sg13g2_nor2_1 _06898_ (.A(_01351_),
    .B(_01383_),
    .Y(_01384_));
 sg13g2_a21oi_2 _06899_ (.B1(_01351_),
    .Y(_01385_),
    .A2(_01383_),
    .A1(_01371_));
 sg13g2_nand2_1 _06900_ (.Y(_01386_),
    .A(_01209_),
    .B(net1497));
 sg13g2_o21ai_1 _06901_ (.B1(_01386_),
    .Y(_01387_),
    .A1(_00071_),
    .A2(net1498));
 sg13g2_a21o_1 _06902_ (.A2(_01387_),
    .A1(_01352_),
    .B1(_01385_),
    .X(_01388_));
 sg13g2_a21oi_1 _06903_ (.A1(_01352_),
    .A2(_01387_),
    .Y(_01389_),
    .B1(_01385_));
 sg13g2_a21oi_1 _06904_ (.A1(net1529),
    .A2(_01389_),
    .Y(_01390_),
    .B1(_01368_));
 sg13g2_a21oi_1 _06905_ (.A1(_01364_),
    .A2(_01390_),
    .Y(_01391_),
    .B1(_01365_));
 sg13g2_o21ai_1 _06906_ (.B1(_01362_),
    .Y(_01392_),
    .A1(net1476),
    .A2(_01391_));
 sg13g2_nand2_1 _06907_ (.Y(_01393_),
    .A(_00071_),
    .B(net1497));
 sg13g2_o21ai_1 _06908_ (.B1(_01393_),
    .Y(_01394_),
    .A1(_01209_),
    .A2(net1499));
 sg13g2_mux2_1 _06909_ (.A0(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[1] ),
    .A1(_01220_),
    .S(net1495),
    .X(_01395_));
 sg13g2_mux2_1 _06910_ (.A0(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[0] ),
    .A1(_01219_),
    .S(net1495),
    .X(_01396_));
 sg13g2_inv_1 _06911_ (.Y(_01397_),
    .A(_01396_));
 sg13g2_nor2_1 _06912_ (.A(_01395_),
    .B(_01396_),
    .Y(_01398_));
 sg13g2_nand2_1 _06913_ (.Y(_01399_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[2] ),
    .B(net1497));
 sg13g2_o21ai_1 _06914_ (.B1(_01399_),
    .Y(_01400_),
    .A1(_01222_),
    .A2(net1497));
 sg13g2_nand2_1 _06915_ (.Y(_01401_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[3] ),
    .B(net1497));
 sg13g2_o21ai_1 _06916_ (.B1(_01401_),
    .Y(_01402_),
    .A1(_01217_),
    .A2(net1497));
 sg13g2_nor2_2 _06917_ (.A(_01355_),
    .B(_01398_),
    .Y(_01403_));
 sg13g2_a21oi_2 _06918_ (.B1(_01403_),
    .Y(_01404_),
    .A2(_01400_),
    .A1(_01356_));
 sg13g2_nand2_1 _06919_ (.Y(_01405_),
    .A(_01356_),
    .B(_01402_));
 sg13g2_mux2_1 _06920_ (.A0(_00078_),
    .A1(_01214_),
    .S(net1495),
    .X(_01406_));
 sg13g2_nand3_1 _06921_ (.B(_01405_),
    .C(_01406_),
    .A(_01404_),
    .Y(_01407_));
 sg13g2_nand2_1 _06922_ (.Y(_01408_),
    .A(_00079_),
    .B(net1497));
 sg13g2_o21ai_1 _06923_ (.B1(_01408_),
    .Y(_01409_),
    .A1(_01212_),
    .A2(net1499));
 sg13g2_and2_1 _06924_ (.A(_01356_),
    .B(_01407_),
    .X(_01410_));
 sg13g2_nor2_1 _06925_ (.A(_01355_),
    .B(_01409_),
    .Y(_01411_));
 sg13g2_nor2_1 _06926_ (.A(_01410_),
    .B(_01411_),
    .Y(_01412_));
 sg13g2_o21ai_1 _06927_ (.B1(_01412_),
    .Y(_01413_),
    .A1(_01355_),
    .A2(_01394_));
 sg13g2_or2_1 _06928_ (.X(_01414_),
    .B(_01413_),
    .A(_01392_));
 sg13g2_xnor2_1 _06929_ (.Y(_01415_),
    .A(_01392_),
    .B(_01413_));
 sg13g2_a21oi_1 _06930_ (.A1(_01370_),
    .A2(_01383_),
    .Y(_01416_),
    .B1(_01351_));
 sg13g2_xnor2_1 _06931_ (.Y(_01417_),
    .A(_01369_),
    .B(_01416_));
 sg13g2_xor2_1 _06932_ (.B(_01416_),
    .A(_01369_),
    .X(_01418_));
 sg13g2_nand2_1 _06933_ (.Y(_01419_),
    .A(_01367_),
    .B(_01417_));
 sg13g2_xnor2_1 _06934_ (.Y(_01420_),
    .A(_01370_),
    .B(_01384_));
 sg13g2_mux2_1 _06935_ (.A0(_01417_),
    .A1(_01420_),
    .S(net1529),
    .X(_01421_));
 sg13g2_xor2_1 _06936_ (.B(_01387_),
    .A(_01385_),
    .X(_01422_));
 sg13g2_xnor2_1 _06937_ (.Y(_01423_),
    .A(_01385_),
    .B(_01387_));
 sg13g2_mux2_1 _06938_ (.A0(_01388_),
    .A1(_01423_),
    .S(net1529),
    .X(_01424_));
 sg13g2_mux4_1 _06939_ (.S0(_01364_),
    .A0(_01389_),
    .A1(_01417_),
    .A2(_01422_),
    .A3(_01420_),
    .S1(net1529),
    .X(_01425_));
 sg13g2_or2_1 _06940_ (.X(_01426_),
    .B(_01425_),
    .A(net1476));
 sg13g2_and2_1 _06941_ (.A(_01362_),
    .B(_01426_),
    .X(_01427_));
 sg13g2_a21o_1 _06942_ (.A2(_01405_),
    .A1(_01404_),
    .B1(_01406_),
    .X(_01428_));
 sg13g2_and2_1 _06943_ (.A(_01407_),
    .B(_01428_),
    .X(_01429_));
 sg13g2_nor2_1 _06944_ (.A(_01427_),
    .B(_01429_),
    .Y(_01430_));
 sg13g2_xnor2_1 _06945_ (.Y(_01431_),
    .A(_01372_),
    .B(_01382_));
 sg13g2_nand2_1 _06946_ (.Y(_01432_),
    .A(_01367_),
    .B(_01431_));
 sg13g2_nand3_1 _06947_ (.B(_01380_),
    .C(_01381_),
    .A(_01352_),
    .Y(_01433_));
 sg13g2_a21o_1 _06948_ (.A2(_01380_),
    .A1(_01352_),
    .B1(_01381_),
    .X(_01434_));
 sg13g2_and2_1 _06949_ (.A(_01433_),
    .B(_01434_),
    .X(_01435_));
 sg13g2_mux2_1 _06950_ (.A0(_01431_),
    .A1(_01435_),
    .S(_01366_),
    .X(_01436_));
 sg13g2_nor2_1 _06951_ (.A(_01359_),
    .B(_01363_),
    .Y(_01437_));
 sg13g2_and2_1 _06952_ (.A(_01436_),
    .B(_01437_),
    .X(_01438_));
 sg13g2_nor2_1 _06953_ (.A(_01359_),
    .B(_01364_),
    .Y(_01439_));
 sg13g2_a21o_1 _06954_ (.A2(_01439_),
    .A1(_01421_),
    .B1(_01438_),
    .X(_01440_));
 sg13g2_a21oi_1 _06955_ (.A1(_01364_),
    .A2(_01424_),
    .Y(_01441_),
    .B1(_01365_));
 sg13g2_nor2_1 _06956_ (.A(_01348_),
    .B(_01360_),
    .Y(_01442_));
 sg13g2_a22oi_1 _06957_ (.Y(_01443_),
    .B1(_01441_),
    .B2(_01442_),
    .A2(_01440_),
    .A1(_01349_));
 sg13g2_xnor2_1 _06958_ (.Y(_01444_),
    .A(_01400_),
    .B(_01403_));
 sg13g2_or2_1 _06959_ (.X(_01445_),
    .B(_01444_),
    .A(_01443_));
 sg13g2_mux2_1 _06960_ (.A0(_01417_),
    .A1(_01422_),
    .S(_01367_),
    .X(_01446_));
 sg13g2_mux4_1 _06961_ (.S0(net1529),
    .A0(_01351_),
    .A1(_01388_),
    .A2(_01423_),
    .A3(_01418_),
    .S1(_01364_),
    .X(_01447_));
 sg13g2_and2_1 _06962_ (.A(net1476),
    .B(_01447_),
    .X(_01448_));
 sg13g2_and2_1 _06963_ (.A(net1529),
    .B(_01431_),
    .X(_01449_));
 sg13g2_a21oi_1 _06964_ (.A1(_01367_),
    .A2(_01420_),
    .Y(_01450_),
    .B1(_01449_));
 sg13g2_a22oi_1 _06965_ (.Y(_01451_),
    .B1(_01376_),
    .B2(_01377_),
    .A2(_01374_),
    .A1(_01373_));
 sg13g2_nor3_1 _06966_ (.A(_01351_),
    .B(_01379_),
    .C(_01451_),
    .Y(_01452_));
 sg13g2_and2_1 _06967_ (.A(_01351_),
    .B(_01378_),
    .X(_01453_));
 sg13g2_nor2_1 _06968_ (.A(_01452_),
    .B(_01453_),
    .Y(_01454_));
 sg13g2_o21ai_1 _06969_ (.B1(net1529),
    .Y(_01455_),
    .A1(_01452_),
    .A2(_01453_));
 sg13g2_nand3_1 _06970_ (.B(_01433_),
    .C(_01434_),
    .A(_01367_),
    .Y(_01456_));
 sg13g2_and2_1 _06971_ (.A(_01455_),
    .B(_01456_),
    .X(_01457_));
 sg13g2_inv_1 _06972_ (.Y(_01458_),
    .A(_01457_));
 sg13g2_nand4_1 _06973_ (.B(_01364_),
    .C(_01455_),
    .A(_01360_),
    .Y(_01459_),
    .D(_01456_));
 sg13g2_nand4_1 _06974_ (.B(_01346_),
    .C(_01347_),
    .A(_01326_),
    .Y(_01460_),
    .D(_01459_));
 sg13g2_a21o_1 _06975_ (.A2(_01450_),
    .A1(_01439_),
    .B1(_01460_),
    .X(_01461_));
 sg13g2_nand2_1 _06976_ (.Y(_01462_),
    .A(_01395_),
    .B(_01396_));
 sg13g2_a22oi_1 _06977_ (.Y(_01463_),
    .B1(_01403_),
    .B2(_01462_),
    .A2(_01395_),
    .A1(_01355_));
 sg13g2_nor3_1 _06978_ (.A(_01448_),
    .B(_01461_),
    .C(_01463_),
    .Y(_01464_));
 sg13g2_o21ai_1 _06979_ (.B1(_01463_),
    .Y(_01465_),
    .A1(_01448_),
    .A2(_01461_));
 sg13g2_nor2b_1 _06980_ (.A(_01464_),
    .B_N(_01465_),
    .Y(_01466_));
 sg13g2_a21oi_1 _06981_ (.A1(_01367_),
    .A2(_01378_),
    .Y(_01467_),
    .B1(_01375_));
 sg13g2_a21oi_1 _06982_ (.A1(_01367_),
    .A2(_01454_),
    .Y(_01468_),
    .B1(_01467_));
 sg13g2_and2_1 _06983_ (.A(_01437_),
    .B(_01468_),
    .X(_01469_));
 sg13g2_a221oi_1 _06984_ (.B2(_01439_),
    .C1(_01469_),
    .B1(_01436_),
    .A1(_01359_),
    .Y(_01470_),
    .A2(_01425_));
 sg13g2_nor3_2 _06985_ (.A(_01348_),
    .B(_01397_),
    .C(_01470_),
    .Y(_01471_));
 sg13g2_a21oi_1 _06986_ (.A1(_01465_),
    .A2(_01471_),
    .Y(_01472_),
    .B1(_01464_));
 sg13g2_xnor2_1 _06987_ (.Y(_01473_),
    .A(_01443_),
    .B(_01444_));
 sg13g2_o21ai_1 _06988_ (.B1(_01445_),
    .Y(_01474_),
    .A1(_01472_),
    .A2(_01473_));
 sg13g2_nand2_1 _06989_ (.Y(_01475_),
    .A(_01363_),
    .B(_01446_));
 sg13g2_o21ai_1 _06990_ (.B1(_01475_),
    .Y(_01476_),
    .A1(_01363_),
    .A2(_01450_));
 sg13g2_a22oi_1 _06991_ (.Y(_01477_),
    .B1(_01476_),
    .B2(_01361_),
    .A2(_01442_),
    .A1(_01391_));
 sg13g2_xor2_1 _06992_ (.B(_01404_),
    .A(_01402_),
    .X(_01478_));
 sg13g2_nor2_1 _06993_ (.A(_01477_),
    .B(_01478_),
    .Y(_01479_));
 sg13g2_xor2_1 _06994_ (.B(_01478_),
    .A(_01477_),
    .X(_01480_));
 sg13g2_a221oi_1 _06995_ (.B2(_01480_),
    .C1(_01479_),
    .B1(_01474_),
    .A1(_01427_),
    .Y(_01481_),
    .A2(_01429_));
 sg13g2_or2_1 _06996_ (.X(_01482_),
    .B(_01481_),
    .A(_01430_));
 sg13g2_or2_1 _06997_ (.X(_01483_),
    .B(_01441_),
    .A(net1476));
 sg13g2_nand2_1 _06998_ (.Y(_01484_),
    .A(_01362_),
    .B(_01483_));
 sg13g2_xor2_1 _06999_ (.B(_01412_),
    .A(_01394_),
    .X(_01485_));
 sg13g2_nand2b_1 _07000_ (.Y(_01486_),
    .B(_01485_),
    .A_N(_01484_));
 sg13g2_nand2_1 _07001_ (.Y(_01487_),
    .A(_01360_),
    .B(_01447_));
 sg13g2_xnor2_1 _07002_ (.Y(_01488_),
    .A(_01409_),
    .B(_01410_));
 sg13g2_nand3_1 _07003_ (.B(_01487_),
    .C(_01488_),
    .A(_01362_),
    .Y(_01489_));
 sg13g2_and2_1 _07004_ (.A(_01486_),
    .B(_01489_),
    .X(_01490_));
 sg13g2_o21ai_1 _07005_ (.B1(_01490_),
    .Y(_01491_),
    .A1(_01430_),
    .A2(_01481_));
 sg13g2_a21oi_1 _07006_ (.A1(_01362_),
    .A2(_01483_),
    .Y(_01492_),
    .B1(_01485_));
 sg13g2_a21o_1 _07007_ (.A2(_01487_),
    .A1(_01362_),
    .B1(_01488_),
    .X(_01493_));
 sg13g2_inv_1 _07008_ (.Y(_01494_),
    .A(_01493_));
 sg13g2_o21ai_1 _07009_ (.B1(_01486_),
    .Y(_01495_),
    .A1(_01492_),
    .A2(_01494_));
 sg13g2_nand2_1 _07010_ (.Y(_01496_),
    .A(_01491_),
    .B(_01495_));
 sg13g2_nand3b_1 _07011_ (.B(_01491_),
    .C(_01495_),
    .Y(_01497_),
    .A_N(_01415_));
 sg13g2_a21oi_1 _07012_ (.A1(_01414_),
    .A2(_01497_),
    .Y(_01498_),
    .B1(_01358_));
 sg13g2_nand3_1 _07013_ (.B(_01414_),
    .C(_01497_),
    .A(_01358_),
    .Y(_01499_));
 sg13g2_nor2b_1 _07014_ (.A(net1463),
    .B_N(_01499_),
    .Y(_01500_));
 sg13g2_xnor2_1 _07015_ (.Y(_01501_),
    .A(_01484_),
    .B(_01485_));
 sg13g2_and2_1 _07016_ (.A(_01489_),
    .B(_01493_),
    .X(_01502_));
 sg13g2_o21ai_1 _07017_ (.B1(_01489_),
    .Y(_01503_),
    .A1(_01482_),
    .A2(_01494_));
 sg13g2_xnor2_1 _07018_ (.Y(_01504_),
    .A(_01501_),
    .B(_01503_));
 sg13g2_xor2_1 _07019_ (.B(_01502_),
    .A(_01482_),
    .X(_01505_));
 sg13g2_xnor2_1 _07020_ (.Y(_01506_),
    .A(_01427_),
    .B(_01429_));
 sg13g2_a21oi_1 _07021_ (.A1(_01474_),
    .A2(_01480_),
    .Y(_01507_),
    .B1(_01479_));
 sg13g2_xnor2_1 _07022_ (.Y(_01508_),
    .A(_01506_),
    .B(_01507_));
 sg13g2_xnor2_1 _07023_ (.Y(_01509_),
    .A(_01474_),
    .B(_01480_));
 sg13g2_xnor2_1 _07024_ (.Y(_01510_),
    .A(_01472_),
    .B(_01473_));
 sg13g2_xnor2_1 _07025_ (.Y(_01511_),
    .A(_01466_),
    .B(_01471_));
 sg13g2_o21ai_1 _07026_ (.B1(_01397_),
    .Y(_01512_),
    .A1(_01348_),
    .A2(_01470_));
 sg13g2_nor2b_2 _07027_ (.A(_01471_),
    .B_N(_01512_),
    .Y(_01513_));
 sg13g2_nand3_1 _07028_ (.B(_01375_),
    .C(_01437_),
    .A(_01367_),
    .Y(_01514_));
 sg13g2_a22oi_1 _07029_ (.Y(_01515_),
    .B1(_01476_),
    .B2(net1476),
    .A2(_01458_),
    .A1(_01439_));
 sg13g2_a21o_1 _07030_ (.A2(_01515_),
    .A1(_01514_),
    .B1(_01348_),
    .X(_01516_));
 sg13g2_nor2b_1 _07031_ (.A(_01513_),
    .B_N(_01516_),
    .Y(_01517_));
 sg13g2_and4_1 _07032_ (.A(_01509_),
    .B(_01510_),
    .C(_01511_),
    .D(_01517_),
    .X(_01518_));
 sg13g2_nand4_1 _07033_ (.B(_01505_),
    .C(_01508_),
    .A(_01504_),
    .Y(_01519_),
    .D(_01518_));
 sg13g2_xor2_1 _07034_ (.B(_01496_),
    .A(_01415_),
    .X(_01520_));
 sg13g2_inv_1 _07035_ (.Y(_01521_),
    .A(_01520_));
 sg13g2_nor3_1 _07036_ (.A(_01500_),
    .B(_01519_),
    .C(_01520_),
    .Y(_01522_));
 sg13g2_nor2_1 _07037_ (.A(net1669),
    .B(_01522_),
    .Y(_01523_));
 sg13g2_or2_1 _07038_ (.X(_01524_),
    .B(_01522_),
    .A(net1669));
 sg13g2_mux2_2 _07039_ (.A0(_00073_),
    .A1(_01237_),
    .S(net1496),
    .X(_01525_));
 sg13g2_nor2_2 _07040_ (.A(_01357_),
    .B(net1463),
    .Y(_01526_));
 sg13g2_nor2_1 _07041_ (.A(_01437_),
    .B(_01467_),
    .Y(_01527_));
 sg13g2_nor2_1 _07042_ (.A(_01420_),
    .B(_01431_),
    .Y(_01528_));
 sg13g2_a21oi_1 _07043_ (.A1(_01419_),
    .A2(_01528_),
    .Y(_01529_),
    .B1(_01364_));
 sg13g2_nand3b_1 _07044_ (.B(_01454_),
    .C(_01432_),
    .Y(_01530_),
    .A_N(_01435_));
 sg13g2_o21ai_1 _07045_ (.B1(net1476),
    .Y(_01531_),
    .A1(_01529_),
    .A2(_01530_));
 sg13g2_nor2b_1 _07046_ (.A(_01527_),
    .B_N(_01531_),
    .Y(_01532_));
 sg13g2_or2_2 _07047_ (.X(_01533_),
    .B(_01532_),
    .A(_01348_));
 sg13g2_inv_1 _07048_ (.Y(_01534_),
    .A(_01533_));
 sg13g2_nand2_1 _07049_ (.Y(_01535_),
    .A(_01516_),
    .B(_01533_));
 sg13g2_xor2_1 _07050_ (.B(_01535_),
    .A(_01513_),
    .X(_01536_));
 sg13g2_or3_1 _07051_ (.A(_01357_),
    .B(net1463),
    .C(_01536_),
    .X(_01537_));
 sg13g2_mux2_2 _07052_ (.A0(_01513_),
    .A1(_01536_),
    .S(_01526_),
    .X(_01538_));
 sg13g2_o21ai_1 _07053_ (.B1(_01537_),
    .Y(_01539_),
    .A1(_01513_),
    .A2(_01526_));
 sg13g2_o21ai_1 _07054_ (.B1(_01535_),
    .Y(_01540_),
    .A1(_01516_),
    .A2(_01532_));
 sg13g2_mux2_2 _07055_ (.A0(_01516_),
    .A1(_01540_),
    .S(_01526_),
    .X(_01541_));
 sg13g2_inv_1 _07056_ (.Y(_01542_),
    .A(_01541_));
 sg13g2_and2_1 _07057_ (.A(_01539_),
    .B(_01541_),
    .X(_01543_));
 sg13g2_a221oi_1 _07058_ (.B2(_01533_),
    .C1(net1463),
    .B1(_01517_),
    .A1(_01353_),
    .Y(_01544_),
    .A2(_01355_));
 sg13g2_xor2_1 _07059_ (.B(_01544_),
    .A(_01511_),
    .X(_01545_));
 sg13g2_inv_1 _07060_ (.Y(_01546_),
    .A(_01545_));
 sg13g2_and3_1 _07061_ (.X(_01547_),
    .A(_01511_),
    .B(_01517_),
    .C(_01533_));
 sg13g2_nor3_1 _07062_ (.A(_01357_),
    .B(_01498_),
    .C(_01547_),
    .Y(_01548_));
 sg13g2_xor2_1 _07063_ (.B(_01548_),
    .A(_01510_),
    .X(_01549_));
 sg13g2_nand2_1 _07064_ (.Y(_01550_),
    .A(_01545_),
    .B(_01549_));
 sg13g2_nand4_1 _07065_ (.B(_01541_),
    .C(_01545_),
    .A(_01539_),
    .Y(_01551_),
    .D(net1434));
 sg13g2_and2_1 _07066_ (.A(_01510_),
    .B(_01547_),
    .X(_01552_));
 sg13g2_nand2_1 _07067_ (.Y(_01553_),
    .A(_01518_),
    .B(_01533_));
 sg13g2_inv_1 _07068_ (.Y(_01554_),
    .A(_01553_));
 sg13g2_nor2b_1 _07069_ (.A(_01553_),
    .B_N(_01508_),
    .Y(_01555_));
 sg13g2_nor3_2 _07070_ (.A(_01357_),
    .B(net1463),
    .C(_01554_),
    .Y(_01556_));
 sg13g2_nor3_1 _07071_ (.A(_01357_),
    .B(net1463),
    .C(_01555_),
    .Y(_01557_));
 sg13g2_xnor2_1 _07072_ (.Y(_01558_),
    .A(_01505_),
    .B(_01557_));
 sg13g2_a221oi_1 _07073_ (.B2(_01555_),
    .C1(net1463),
    .B1(_01505_),
    .A1(_01353_),
    .Y(_01559_),
    .A2(_01355_));
 sg13g2_xnor2_1 _07074_ (.Y(_01560_),
    .A(_01504_),
    .B(_01559_));
 sg13g2_inv_1 _07075_ (.Y(_01561_),
    .A(net1431));
 sg13g2_nor2_2 _07076_ (.A(net1433),
    .B(net1431),
    .Y(_01562_));
 sg13g2_xnor2_1 _07077_ (.Y(_01563_),
    .A(_01508_),
    .B(_01556_));
 sg13g2_xor2_1 _07078_ (.B(_01556_),
    .A(_01508_),
    .X(_01564_));
 sg13g2_nor3_1 _07079_ (.A(_01357_),
    .B(net1463),
    .C(_01552_),
    .Y(_01565_));
 sg13g2_xor2_1 _07080_ (.B(_01565_),
    .A(_01509_),
    .X(_01566_));
 sg13g2_xnor2_1 _07081_ (.Y(_01567_),
    .A(_01509_),
    .B(_01565_));
 sg13g2_nor2_2 _07082_ (.A(net1430),
    .B(_01567_),
    .Y(_01568_));
 sg13g2_nand3_1 _07083_ (.B(_01562_),
    .C(_01568_),
    .A(_01551_),
    .Y(_01569_));
 sg13g2_nand4_1 _07084_ (.B(_01551_),
    .C(_01562_),
    .A(_01525_),
    .Y(_01570_),
    .D(_01568_));
 sg13g2_nand2_1 _07085_ (.Y(_01571_),
    .A(_01249_),
    .B(net1495));
 sg13g2_nand2_2 _07086_ (.Y(_01572_),
    .A(_01337_),
    .B(_01571_));
 sg13g2_o21ai_1 _07087_ (.B1(_01545_),
    .Y(_01573_),
    .A1(_01538_),
    .A2(_01541_));
 sg13g2_and2_1 _07088_ (.A(net1434),
    .B(_01564_),
    .X(_01574_));
 sg13g2_a21o_1 _07089_ (.A2(_01567_),
    .A1(_01564_),
    .B1(net1432),
    .X(_01575_));
 sg13g2_a21o_1 _07090_ (.A2(_01574_),
    .A1(_01573_),
    .B1(_01575_),
    .X(_01576_));
 sg13g2_and2_1 _07091_ (.A(_01561_),
    .B(_01576_),
    .X(_01577_));
 sg13g2_and3_1 _07092_ (.X(_01578_),
    .A(net1490),
    .B(net1429),
    .C(_01576_));
 sg13g2_a21oi_2 _07093_ (.B1(_01321_),
    .Y(_01579_),
    .A2(net1495),
    .A1(_01232_));
 sg13g2_o21ai_1 _07094_ (.B1(_01568_),
    .Y(_01580_),
    .A1(_01543_),
    .A2(_01550_));
 sg13g2_a21oi_1 _07095_ (.A1(_01562_),
    .A2(_01580_),
    .Y(_01581_),
    .B1(_01579_));
 sg13g2_a21o_1 _07096_ (.A2(_01580_),
    .A1(_01562_),
    .B1(_01579_),
    .X(_01582_));
 sg13g2_o21ai_1 _07097_ (.B1(_01572_),
    .Y(_01583_),
    .A1(_01578_),
    .A2(_01582_));
 sg13g2_nand2b_1 _07098_ (.Y(_01584_),
    .B(_01569_),
    .A_N(_01525_));
 sg13g2_nand2_1 _07099_ (.Y(_01585_),
    .A(_01572_),
    .B(_01584_));
 sg13g2_nand3_1 _07100_ (.B(_01579_),
    .C(_01580_),
    .A(_01562_),
    .Y(_01586_));
 sg13g2_nand4_1 _07101_ (.B(_01578_),
    .C(_01579_),
    .A(_01562_),
    .Y(_01587_),
    .D(_01580_));
 sg13g2_mux2_2 _07102_ (.A0(_00081_),
    .A1(_01248_),
    .S(net1496),
    .X(_01588_));
 sg13g2_a21oi_2 _07103_ (.B1(_01327_),
    .Y(_01589_),
    .A2(net1496),
    .A1(_01240_));
 sg13g2_o21ai_1 _07104_ (.B1(_01526_),
    .Y(_01590_),
    .A1(_01519_),
    .A2(_01534_));
 sg13g2_or2_1 _07105_ (.X(_01591_),
    .B(_01590_),
    .A(_01521_));
 sg13g2_nand2_1 _07106_ (.Y(_01592_),
    .A(_01521_),
    .B(_01590_));
 sg13g2_xnor2_1 _07107_ (.Y(_01593_),
    .A(_01521_),
    .B(_01590_));
 sg13g2_nand2_1 _07108_ (.Y(_01594_),
    .A(_01520_),
    .B(_01526_));
 sg13g2_and2_1 _07109_ (.A(_01590_),
    .B(_01594_),
    .X(_01595_));
 sg13g2_xnor2_1 _07110_ (.Y(_01596_),
    .A(_01500_),
    .B(_01595_));
 sg13g2_inv_2 _07111_ (.Y(_01597_),
    .A(net1425));
 sg13g2_nor2_1 _07112_ (.A(_01252_),
    .B(net1499),
    .Y(_01598_));
 sg13g2_a21oi_2 _07113_ (.B1(_01598_),
    .Y(_01599_),
    .A2(net1499),
    .A1(_00703_));
 sg13g2_nor2_1 _07114_ (.A(_01245_),
    .B(net1499),
    .Y(_01600_));
 sg13g2_a21oi_2 _07115_ (.B1(_01600_),
    .Y(_01601_),
    .A2(net1499),
    .A1(_00704_));
 sg13g2_and4_1 _07116_ (.A(_01588_),
    .B(_01589_),
    .C(net1428),
    .D(_01599_),
    .X(_01602_));
 sg13g2_and2_1 _07117_ (.A(_01601_),
    .B(_01602_),
    .X(_01603_));
 sg13g2_nand2_1 _07118_ (.Y(_01604_),
    .A(_01597_),
    .B(_01603_));
 sg13g2_a221oi_1 _07119_ (.B2(_01587_),
    .C1(_01604_),
    .B1(_01585_),
    .A1(_01570_),
    .Y(_01605_),
    .A2(_01583_));
 sg13g2_xnor2_1 _07120_ (.Y(_01606_),
    .A(_01521_),
    .B(_01590_));
 sg13g2_inv_1 _07121_ (.Y(_01607_),
    .A(_01606_));
 sg13g2_nor2_2 _07122_ (.A(_01524_),
    .B(_01605_),
    .Y(_01608_));
 sg13g2_or2_2 _07123_ (.X(_01609_),
    .B(_01579_),
    .A(_01525_));
 sg13g2_nor3_1 _07124_ (.A(_01572_),
    .B(_01599_),
    .C(_01609_),
    .Y(_01610_));
 sg13g2_or2_1 _07125_ (.X(_01611_),
    .B(_01589_),
    .A(_01588_));
 sg13g2_inv_1 _07126_ (.Y(_01612_),
    .A(_01611_));
 sg13g2_nor2b_1 _07127_ (.A(_01601_),
    .B_N(net1490),
    .Y(_01613_));
 sg13g2_and4_1 _07128_ (.A(net1425),
    .B(_01610_),
    .C(_01612_),
    .D(_01613_),
    .X(_01614_));
 sg13g2_nor3_2 _07129_ (.A(_01524_),
    .B(_01605_),
    .C(_01614_),
    .Y(_01615_));
 sg13g2_and2_1 _07130_ (.A(_01560_),
    .B(net1427),
    .X(_01616_));
 sg13g2_a221oi_1 _07131_ (.B2(_01542_),
    .C1(net1423),
    .B1(_01616_),
    .A1(_01538_),
    .Y(_01617_),
    .A2(_01607_));
 sg13g2_a21oi_1 _07132_ (.A1(_01545_),
    .A2(net1423),
    .Y(_01618_),
    .B1(_01617_));
 sg13g2_a21oi_1 _07133_ (.A1(_01229_),
    .A2(_01254_),
    .Y(_01619_),
    .B1(_01266_));
 sg13g2_a21o_1 _07134_ (.A2(_01254_),
    .A1(_01229_),
    .B1(_01266_),
    .X(_01620_));
 sg13g2_a221oi_1 _07135_ (.B2(_01618_),
    .C1(net1486),
    .B1(_01615_),
    .A1(_01219_),
    .Y(_01621_),
    .A2(net1669));
 sg13g2_o21ai_1 _07136_ (.B1(net1500),
    .Y(_01622_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[0] ),
    .A2(net1487));
 sg13g2_o21ai_1 _07137_ (.B1(_01269_),
    .Y(_01623_),
    .A1(_01621_),
    .A2(_01622_));
 sg13g2_nor4_1 _07138_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][12] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][11] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][14] ),
    .D(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][13] ),
    .Y(_01624_));
 sg13g2_nor4_1 _07139_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][8] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][7] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][10] ),
    .D(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][9] ),
    .Y(_01625_));
 sg13g2_and2_1 _07140_ (.A(_01624_),
    .B(_01625_),
    .X(_01626_));
 sg13g2_nand4_1 _07141_ (.B(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][11] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][14] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][12] ),
    .Y(_01627_),
    .D(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][13] ));
 sg13g2_nand4_1 _07142_ (.B(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][7] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][10] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][8] ),
    .Y(_01628_),
    .D(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][9] ));
 sg13g2_nor2_2 _07143_ (.A(_01627_),
    .B(_01628_),
    .Y(_01629_));
 sg13g2_or4_1 _07144_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][3] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][2] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][5] ),
    .D(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][4] ),
    .X(_01630_));
 sg13g2_nor3_1 _07145_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][1] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][0] ),
    .C(_01630_),
    .Y(_01631_));
 sg13g2_nand2_1 _07146_ (.Y(_01632_),
    .A(_00141_),
    .B(_01631_));
 sg13g2_o21ai_1 _07147_ (.B1(_01632_),
    .Y(_01633_),
    .A1(_01626_),
    .A2(_01629_));
 sg13g2_nor4_1 _07148_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][11] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][12] ),
    .C(net1787),
    .D(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][14] ),
    .Y(_01634_));
 sg13g2_nor3_1 _07149_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][7] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][8] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][9] ),
    .Y(_01635_));
 sg13g2_nand3_1 _07150_ (.B(_01634_),
    .C(_01635_),
    .A(_00769_),
    .Y(_01636_));
 sg13g2_inv_1 _07151_ (.Y(_01637_),
    .A(_01636_));
 sg13g2_nand4_1 _07152_ (.B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][12] ),
    .C(net1787),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][11] ),
    .Y(_01638_),
    .D(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][14] ));
 sg13g2_nand4_1 _07153_ (.B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][8] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][9] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][7] ),
    .Y(_01639_),
    .D(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][10] ));
 sg13g2_o21ai_1 _07154_ (.B1(_01636_),
    .Y(_01640_),
    .A1(_01638_),
    .A2(_01639_));
 sg13g2_nor4_1 _07155_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][1] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][0] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][3] ),
    .D(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][4] ),
    .Y(_01641_));
 sg13g2_nand3_1 _07156_ (.B(_00766_),
    .C(_01641_),
    .A(_00765_),
    .Y(_01642_));
 sg13g2_o21ai_1 _07157_ (.B1(_01640_),
    .Y(_01643_),
    .A1(_00768_),
    .A2(_01642_));
 sg13g2_a22oi_1 _07158_ (.Y(_01644_),
    .B1(_01637_),
    .B2(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][15] ),
    .A2(_01626_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][15] ));
 sg13g2_nand4_1 _07159_ (.B(_01633_),
    .C(_01643_),
    .A(net1531),
    .Y(_01645_),
    .D(_01644_));
 sg13g2_nor2b_1 _07160_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][6] ),
    .B_N(_01631_),
    .Y(_01646_));
 sg13g2_and2_1 _07161_ (.A(_01629_),
    .B(_01646_),
    .X(_01647_));
 sg13g2_nand2_1 _07162_ (.Y(_01648_),
    .A(_01629_),
    .B(_01646_));
 sg13g2_nor4_2 _07163_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][6] ),
    .B(_01638_),
    .C(_01639_),
    .Y(_01649_),
    .D(_01642_));
 sg13g2_a21oi_1 _07164_ (.A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][15] ),
    .A2(_01649_),
    .Y(_01650_),
    .B1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][15] ));
 sg13g2_nand2b_1 _07165_ (.Y(_01651_),
    .B(_01647_),
    .A_N(_01650_));
 sg13g2_nand2b_1 _07166_ (.Y(_01652_),
    .B(_01649_),
    .A_N(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][15] ));
 sg13g2_a21oi_1 _07167_ (.A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][15] ),
    .A2(_01652_),
    .Y(_01653_),
    .B1(_01651_));
 sg13g2_or2_2 _07168_ (.X(_01654_),
    .B(_01653_),
    .A(_01645_));
 sg13g2_nand2b_1 _07169_ (.Y(_01655_),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][12] ),
    .A_N(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][12] ));
 sg13g2_xor2_1 _07170_ (.B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][12] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][12] ),
    .X(_01656_));
 sg13g2_xor2_1 _07171_ (.B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][11] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][11] ),
    .X(_01657_));
 sg13g2_nand2_1 _07172_ (.Y(_01658_),
    .A(_00763_),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][13] ));
 sg13g2_xnor2_1 _07173_ (.Y(_01659_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][13] ),
    .B(net1787));
 sg13g2_xor2_1 _07174_ (.B(net1787),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][13] ),
    .X(_01660_));
 sg13g2_nor3_2 _07175_ (.A(_01656_),
    .B(_01657_),
    .C(_01660_),
    .Y(_01661_));
 sg13g2_nand2b_1 _07176_ (.Y(_01662_),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][10] ),
    .A_N(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][10] ));
 sg13g2_nor2b_1 _07177_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][10] ),
    .B_N(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][10] ),
    .Y(_01663_));
 sg13g2_xnor2_1 _07178_ (.Y(_01664_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][10] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][10] ));
 sg13g2_nor2b_1 _07179_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][9] ),
    .B_N(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][9] ),
    .Y(_01665_));
 sg13g2_xnor2_1 _07180_ (.Y(_01666_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][9] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][9] ));
 sg13g2_xor2_1 _07181_ (.B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][9] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][9] ),
    .X(_01667_));
 sg13g2_nor2b_1 _07182_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][8] ),
    .B_N(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][8] ),
    .Y(_01668_));
 sg13g2_nand2b_1 _07183_ (.Y(_01669_),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][8] ),
    .A_N(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][8] ));
 sg13g2_nor2b_1 _07184_ (.A(_01668_),
    .B_N(_01669_),
    .Y(_01670_));
 sg13g2_nor2_1 _07185_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][14] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][14] ),
    .Y(_01671_));
 sg13g2_xnor2_1 _07186_ (.Y(_01672_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][14] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][14] ));
 sg13g2_and2_1 _07187_ (.A(_01661_),
    .B(_01672_),
    .X(_01673_));
 sg13g2_nand2_1 _07188_ (.Y(_01674_),
    .A(_01664_),
    .B(_01666_));
 sg13g2_nand2b_1 _07189_ (.Y(_01675_),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][7] ),
    .A_N(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][7] ));
 sg13g2_xnor2_1 _07190_ (.Y(_01676_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][7] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][7] ));
 sg13g2_xor2_1 _07191_ (.B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][7] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][7] ),
    .X(_01677_));
 sg13g2_and4_1 _07192_ (.A(_01664_),
    .B(_01666_),
    .C(_01670_),
    .D(_01676_),
    .X(_01678_));
 sg13g2_and2_2 _07193_ (.A(_01673_),
    .B(_01678_),
    .X(_01679_));
 sg13g2_nand2_1 _07194_ (.Y(_01680_),
    .A(_01673_),
    .B(_01678_));
 sg13g2_a21oi_1 _07195_ (.A1(_01669_),
    .A2(_01675_),
    .Y(_01681_),
    .B1(_01668_));
 sg13g2_a21oi_1 _07196_ (.A1(_01662_),
    .A2(_01665_),
    .Y(_01682_),
    .B1(_01663_));
 sg13g2_o21ai_1 _07197_ (.B1(_01682_),
    .Y(_01683_),
    .A1(_01674_),
    .A2(_01681_));
 sg13g2_nor2b_1 _07198_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][14] ),
    .B_N(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][14] ),
    .Y(_01684_));
 sg13g2_a22oi_1 _07199_ (.Y(_01685_),
    .B1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][12] ),
    .B2(_00761_),
    .A2(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][11] ),
    .A1(_00762_));
 sg13g2_o21ai_1 _07200_ (.B1(_01655_),
    .Y(_01686_),
    .A1(_00763_),
    .A2(net1787));
 sg13g2_o21ai_1 _07201_ (.B1(_01658_),
    .Y(_01687_),
    .A1(_01685_),
    .A2(_01686_));
 sg13g2_a221oi_1 _07202_ (.B2(_01672_),
    .C1(_01684_),
    .B1(_01687_),
    .A1(_01673_),
    .Y(_01688_),
    .A2(_01683_));
 sg13g2_nor2_1 _07203_ (.A(_01679_),
    .B(net1667),
    .Y(_01689_));
 sg13g2_nand3b_1 _07204_ (.B(_00145_),
    .C(_01680_),
    .Y(_01690_),
    .A_N(net1667));
 sg13g2_o21ai_1 _07205_ (.B1(_00146_),
    .Y(_01691_),
    .A1(_01679_),
    .A2(net1667));
 sg13g2_nand2_2 _07206_ (.Y(_01692_),
    .A(_01690_),
    .B(_01691_));
 sg13g2_and2_1 _07207_ (.A(_00146_),
    .B(_00145_),
    .X(_01693_));
 sg13g2_a21o_1 _07208_ (.A2(_01691_),
    .A1(_01690_),
    .B1(_01693_),
    .X(_01694_));
 sg13g2_or3_2 _07209_ (.A(_00153_),
    .B(_01679_),
    .C(net1667),
    .X(_01695_));
 sg13g2_o21ai_1 _07210_ (.B1(_00773_),
    .Y(_01696_),
    .A1(_01679_),
    .A2(net1667));
 sg13g2_and2_2 _07211_ (.A(_01695_),
    .B(_01696_),
    .X(_01697_));
 sg13g2_nand2_2 _07212_ (.Y(_01698_),
    .A(_01695_),
    .B(_01696_));
 sg13g2_a22oi_1 _07213_ (.Y(_01699_),
    .B1(_01696_),
    .B2(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][8] ),
    .A2(_01695_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][8] ));
 sg13g2_a22oi_1 _07214_ (.Y(_01700_),
    .B1(_01698_),
    .B2(_01699_),
    .A2(_01694_),
    .A1(_01670_));
 sg13g2_nor2b_1 _07215_ (.A(net1553),
    .B_N(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][9] ),
    .Y(_01701_));
 sg13g2_a21oi_2 _07216_ (.B1(_01701_),
    .Y(_01702_),
    .A2(net1553),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][9] ));
 sg13g2_mux2_1 _07217_ (.A0(_01700_),
    .A1(_01702_),
    .S(_01667_),
    .X(_01703_));
 sg13g2_nand2b_1 _07218_ (.Y(_01704_),
    .B(_01664_),
    .A_N(_01703_));
 sg13g2_nor2b_1 _07219_ (.A(net1549),
    .B_N(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][10] ),
    .Y(_01705_));
 sg13g2_a21o_1 _07220_ (.A2(net1549),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][10] ),
    .B1(_01705_),
    .X(_01706_));
 sg13g2_a21oi_2 _07221_ (.B1(_01705_),
    .Y(_01707_),
    .A2(net1549),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][10] ));
 sg13g2_mux2_1 _07222_ (.A0(_01707_),
    .A1(_01703_),
    .S(_01664_),
    .X(_01708_));
 sg13g2_or2_2 _07223_ (.X(_01709_),
    .B(_01708_),
    .A(_01661_));
 sg13g2_mux2_2 _07224_ (.A0(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][11] ),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][11] ),
    .S(net1549),
    .X(_01710_));
 sg13g2_a21o_1 _07225_ (.A2(_01710_),
    .A1(_01659_),
    .B1(_01656_),
    .X(_01711_));
 sg13g2_mux2_1 _07226_ (.A0(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][12] ),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][12] ),
    .S(net1549),
    .X(_01712_));
 sg13g2_nor2_2 _07227_ (.A(_01710_),
    .B(_01712_),
    .Y(_01713_));
 sg13g2_nand3_1 _07228_ (.B(_01659_),
    .C(_01710_),
    .A(_01656_),
    .Y(_01714_));
 sg13g2_xnor2_1 _07229_ (.Y(_01715_),
    .A(_01660_),
    .B(_01713_));
 sg13g2_nand4_1 _07230_ (.B(_01711_),
    .C(_01714_),
    .A(_01657_),
    .Y(_01716_),
    .D(_01715_));
 sg13g2_nor2_1 _07231_ (.A(_00763_),
    .B(net1549),
    .Y(_01717_));
 sg13g2_a21oi_2 _07232_ (.B1(_01717_),
    .Y(_01718_),
    .A2(net1549),
    .A1(net1787));
 sg13g2_a21oi_1 _07233_ (.A1(_01660_),
    .A2(_01718_),
    .Y(_01719_),
    .B1(_01672_));
 sg13g2_nand2b_1 _07234_ (.Y(_01720_),
    .B(_01703_),
    .A_N(_01664_));
 sg13g2_a221oi_1 _07235_ (.B2(_01704_),
    .C1(_01719_),
    .B1(_01720_),
    .A1(_01708_),
    .Y(_01721_),
    .A2(_01716_));
 sg13g2_and2_2 _07236_ (.A(_01709_),
    .B(_01721_),
    .X(_01722_));
 sg13g2_nand2_1 _07237_ (.Y(_01723_),
    .A(_00772_),
    .B(net1551));
 sg13g2_mux2_2 _07238_ (.A0(_00150_),
    .A1(_00149_),
    .S(net1551),
    .X(_01724_));
 sg13g2_o21ai_1 _07239_ (.B1(_01723_),
    .Y(_01725_),
    .A1(_00150_),
    .A2(net1551));
 sg13g2_nor2_1 _07240_ (.A(_00772_),
    .B(net1551),
    .Y(_01726_));
 sg13g2_a21o_1 _07241_ (.A2(net1551),
    .A1(_00150_),
    .B1(_01726_),
    .X(_01727_));
 sg13g2_a21oi_2 _07242_ (.B1(_01726_),
    .Y(_01728_),
    .A2(net1552),
    .A1(_00150_));
 sg13g2_a21oi_2 _07243_ (.B1(_01728_),
    .Y(_01729_),
    .A2(_01725_),
    .A1(_01722_));
 sg13g2_nand3_1 _07244_ (.B(_00772_),
    .C(_01722_),
    .A(_00771_),
    .Y(_01730_));
 sg13g2_nor2b_2 _07245_ (.A(_01729_),
    .B_N(_01730_),
    .Y(_01731_));
 sg13g2_xnor2_1 _07246_ (.Y(_01732_),
    .A(_01666_),
    .B(_01700_));
 sg13g2_xnor2_1 _07247_ (.Y(_01733_),
    .A(_01667_),
    .B(_01700_));
 sg13g2_and3_2 _07248_ (.X(_01734_),
    .A(_01709_),
    .B(_01721_),
    .C(_01733_));
 sg13g2_a21oi_1 _07249_ (.A1(_01722_),
    .A2(_01725_),
    .Y(_01735_),
    .B1(_01734_));
 sg13g2_xnor2_1 _07250_ (.Y(_01736_),
    .A(_01670_),
    .B(_01694_));
 sg13g2_inv_2 _07251_ (.Y(_01737_),
    .A(net1506));
 sg13g2_nor2_1 _07252_ (.A(_01725_),
    .B(_01736_),
    .Y(_01738_));
 sg13g2_nand3b_1 _07253_ (.B(_00144_),
    .C(_01680_),
    .Y(_01739_),
    .A_N(_01688_));
 sg13g2_o21ai_1 _07254_ (.B1(_00143_),
    .Y(_01740_),
    .A1(_01679_),
    .A2(net1667));
 sg13g2_nand2_2 _07255_ (.Y(_01741_),
    .A(_01739_),
    .B(_01740_));
 sg13g2_nand3b_1 _07256_ (.B(_00152_),
    .C(_01680_),
    .Y(_01742_),
    .A_N(net1667));
 sg13g2_o21ai_1 _07257_ (.B1(_00151_),
    .Y(_01743_),
    .A1(_01679_),
    .A2(net1667));
 sg13g2_nand2_1 _07258_ (.Y(_01744_),
    .A(_01742_),
    .B(_01743_));
 sg13g2_a22oi_1 _07259_ (.Y(_01745_),
    .B1(_01742_),
    .B2(_01743_),
    .A2(_01740_),
    .A1(_01739_));
 sg13g2_mux2_2 _07260_ (.A0(_00147_),
    .A1(_00148_),
    .S(net1551),
    .X(_01746_));
 sg13g2_nor2_1 _07261_ (.A(_01724_),
    .B(_01745_),
    .Y(_01747_));
 sg13g2_xnor2_1 _07262_ (.Y(_01748_),
    .A(_01746_),
    .B(_01747_));
 sg13g2_nand2_1 _07263_ (.Y(_01749_),
    .A(_01745_),
    .B(_01746_));
 sg13g2_mux2_1 _07264_ (.A0(_00157_),
    .A1(_00158_),
    .S(net1552),
    .X(_01750_));
 sg13g2_mux2_1 _07265_ (.A0(_00155_),
    .A1(_00156_),
    .S(net1552),
    .X(_01751_));
 sg13g2_nand4_1 _07266_ (.B(_01746_),
    .C(_01750_),
    .A(_01745_),
    .Y(_01752_),
    .D(_01751_));
 sg13g2_mux2_1 _07267_ (.A0(_00159_),
    .A1(_00160_),
    .S(net1550),
    .X(_01753_));
 sg13g2_inv_1 _07268_ (.Y(_01754_),
    .A(_01753_));
 sg13g2_a21oi_1 _07269_ (.A1(_01745_),
    .A2(_01746_),
    .Y(_01755_),
    .B1(_01724_));
 sg13g2_nor2_1 _07270_ (.A(_01724_),
    .B(_01750_),
    .Y(_01756_));
 sg13g2_nor2_1 _07271_ (.A(_01755_),
    .B(_01756_),
    .Y(_01757_));
 sg13g2_nand2_1 _07272_ (.Y(_01758_),
    .A(_01725_),
    .B(_01752_));
 sg13g2_o21ai_1 _07273_ (.B1(_01725_),
    .Y(_01759_),
    .A1(_01752_),
    .A2(_01754_));
 sg13g2_nand2_1 _07274_ (.Y(_01760_),
    .A(_00141_),
    .B(net1550));
 sg13g2_o21ai_1 _07275_ (.B1(_01760_),
    .Y(_01761_),
    .A1(_00768_),
    .A2(net1549));
 sg13g2_a21o_1 _07276_ (.A2(_01761_),
    .A1(_01759_),
    .B1(_01724_),
    .X(_01762_));
 sg13g2_nor2_1 _07277_ (.A(net1748),
    .B(_01724_),
    .Y(_01763_));
 sg13g2_a21oi_1 _07278_ (.A1(net1749),
    .A2(_01762_),
    .Y(_01764_),
    .B1(_01763_));
 sg13g2_a21oi_1 _07279_ (.A1(_01736_),
    .A2(_01764_),
    .Y(_01765_),
    .B1(_01738_));
 sg13g2_nor2_1 _07280_ (.A(_01732_),
    .B(_01765_),
    .Y(_01766_));
 sg13g2_or2_1 _07281_ (.X(_01767_),
    .B(_01766_),
    .A(_01735_));
 sg13g2_nor2b_1 _07282_ (.A(net1550),
    .B_N(_00141_),
    .Y(_01768_));
 sg13g2_a21oi_2 _07283_ (.B1(_01768_),
    .Y(_01769_),
    .A2(net1550),
    .A1(_00142_));
 sg13g2_mux2_2 _07284_ (.A0(_00144_),
    .A1(_00143_),
    .S(net1553),
    .X(_01770_));
 sg13g2_mux2_1 _07285_ (.A0(_00152_),
    .A1(_00151_),
    .S(net1551),
    .X(_01771_));
 sg13g2_nor2_1 _07286_ (.A(_01727_),
    .B(_01770_),
    .Y(_01772_));
 sg13g2_a21oi_1 _07287_ (.A1(_01770_),
    .A2(_01771_),
    .Y(_01773_),
    .B1(_01727_));
 sg13g2_mux2_1 _07288_ (.A0(_00148_),
    .A1(_00147_),
    .S(net1552),
    .X(_01774_));
 sg13g2_nand2b_1 _07289_ (.Y(_01775_),
    .B(_01774_),
    .A_N(_01773_));
 sg13g2_nand2_1 _07290_ (.Y(_01776_),
    .A(_01728_),
    .B(_01775_));
 sg13g2_nand2b_1 _07291_ (.Y(_01777_),
    .B(net1552),
    .A_N(_00157_));
 sg13g2_o21ai_1 _07292_ (.B1(_01777_),
    .Y(_01778_),
    .A1(_00158_),
    .A2(net1551));
 sg13g2_o21ai_1 _07293_ (.B1(_01728_),
    .Y(_01779_),
    .A1(_01775_),
    .A2(_01778_));
 sg13g2_mux2_1 _07294_ (.A0(_00156_),
    .A1(_00155_),
    .S(net1552),
    .X(_01780_));
 sg13g2_and2_1 _07295_ (.A(_01779_),
    .B(_01780_),
    .X(_01781_));
 sg13g2_nor2_1 _07296_ (.A(_01727_),
    .B(_01781_),
    .Y(_01782_));
 sg13g2_mux2_1 _07297_ (.A0(_00160_),
    .A1(_00159_),
    .S(net1550),
    .X(_01783_));
 sg13g2_nand2_1 _07298_ (.Y(_01784_),
    .A(_01781_),
    .B(_01783_));
 sg13g2_nand2_1 _07299_ (.Y(_01785_),
    .A(_01728_),
    .B(_01784_));
 sg13g2_o21ai_1 _07300_ (.B1(_01728_),
    .Y(_01786_),
    .A1(_01769_),
    .A2(_01784_));
 sg13g2_nand2b_1 _07301_ (.Y(_01787_),
    .B(_01786_),
    .A_N(_01767_));
 sg13g2_xor2_1 _07302_ (.B(_01761_),
    .A(_01759_),
    .X(_01788_));
 sg13g2_mux2_1 _07303_ (.A0(_01762_),
    .A1(_01788_),
    .S(net1748),
    .X(_01789_));
 sg13g2_mux2_1 _07304_ (.A0(_01725_),
    .A1(_01789_),
    .S(net1506),
    .X(_01790_));
 sg13g2_nor2_1 _07305_ (.A(_01732_),
    .B(_01790_),
    .Y(_01791_));
 sg13g2_or2_1 _07306_ (.X(_01792_),
    .B(_01791_),
    .A(_01735_));
 sg13g2_xor2_1 _07307_ (.B(_01785_),
    .A(_01769_),
    .X(_01793_));
 sg13g2_nor2_1 _07308_ (.A(_01792_),
    .B(_01793_),
    .Y(_01794_));
 sg13g2_xnor2_1 _07309_ (.Y(_01795_),
    .A(_01792_),
    .B(_01793_));
 sg13g2_inv_1 _07310_ (.Y(_01796_),
    .A(_01795_));
 sg13g2_xnor2_1 _07311_ (.Y(_01797_),
    .A(_01754_),
    .B(_01758_));
 sg13g2_mux4_1 _07312_ (.S0(net1748),
    .A0(_01725_),
    .A1(_01762_),
    .A2(_01788_),
    .A3(_01797_),
    .S1(net1506),
    .X(_01798_));
 sg13g2_nor2_1 _07313_ (.A(_01732_),
    .B(_01798_),
    .Y(_01799_));
 sg13g2_or2_1 _07314_ (.X(_01800_),
    .B(_01799_),
    .A(_01735_));
 sg13g2_xor2_1 _07315_ (.B(_01783_),
    .A(_01782_),
    .X(_01801_));
 sg13g2_or2_1 _07316_ (.X(_01802_),
    .B(_01801_),
    .A(_01800_));
 sg13g2_xor2_1 _07317_ (.B(_01801_),
    .A(_01800_),
    .X(_01803_));
 sg13g2_inv_1 _07318_ (.Y(_01804_),
    .A(_01803_));
 sg13g2_nand2_1 _07319_ (.Y(_01805_),
    .A(_01677_),
    .B(_01797_));
 sg13g2_xor2_1 _07320_ (.B(_01757_),
    .A(_01751_),
    .X(_01806_));
 sg13g2_mux4_1 _07321_ (.S0(net1748),
    .A0(_01762_),
    .A1(_01788_),
    .A2(_01797_),
    .A3(_01806_),
    .S1(net1506),
    .X(_01807_));
 sg13g2_nor2_1 _07322_ (.A(_01732_),
    .B(_01807_),
    .Y(_01808_));
 sg13g2_or2_1 _07323_ (.X(_01809_),
    .B(_01808_),
    .A(_01735_));
 sg13g2_xnor2_1 _07324_ (.Y(_01810_),
    .A(_01779_),
    .B(_01780_));
 sg13g2_nor2_1 _07325_ (.A(_01809_),
    .B(_01810_),
    .Y(_01811_));
 sg13g2_xor2_1 _07326_ (.B(_01810_),
    .A(_01809_),
    .X(_01812_));
 sg13g2_and3_1 _07327_ (.X(_01813_),
    .A(_01709_),
    .B(_01721_),
    .C(_01732_));
 sg13g2_xnor2_1 _07328_ (.Y(_01814_),
    .A(_01750_),
    .B(_01755_));
 sg13g2_mux4_1 _07329_ (.S0(net1748),
    .A0(_01788_),
    .A1(_01797_),
    .A2(_01806_),
    .A3(_01814_),
    .S1(net1506),
    .X(_01815_));
 sg13g2_a22oi_1 _07330_ (.Y(_01816_),
    .B1(_01815_),
    .B2(_01734_),
    .A2(_01813_),
    .A1(_01765_));
 sg13g2_xnor2_1 _07331_ (.Y(_01817_),
    .A(_01776_),
    .B(_01778_));
 sg13g2_nand2b_1 _07332_ (.Y(_01818_),
    .B(_01817_),
    .A_N(_01816_));
 sg13g2_nand2_1 _07333_ (.Y(_01819_),
    .A(_01677_),
    .B(_01814_));
 sg13g2_mux4_1 _07334_ (.S0(_01737_),
    .A0(_01748_),
    .A1(_01806_),
    .A2(_01814_),
    .A3(_01797_),
    .S1(_01677_),
    .X(_01820_));
 sg13g2_a22oi_1 _07335_ (.Y(_01821_),
    .B1(_01820_),
    .B2(_01734_),
    .A2(_01813_),
    .A1(_01790_));
 sg13g2_xor2_1 _07336_ (.B(_01774_),
    .A(_01773_),
    .X(_01822_));
 sg13g2_nor2_1 _07337_ (.A(_01821_),
    .B(_01822_),
    .Y(_01823_));
 sg13g2_nand4_1 _07338_ (.B(_01721_),
    .C(_01732_),
    .A(_01709_),
    .Y(_01824_),
    .D(_01798_));
 sg13g2_nor2_1 _07339_ (.A(_01724_),
    .B(_01741_),
    .Y(_01825_));
 sg13g2_xnor2_1 _07340_ (.Y(_01826_),
    .A(_01744_),
    .B(_01825_));
 sg13g2_and2_1 _07341_ (.A(net1748),
    .B(_01826_),
    .X(_01827_));
 sg13g2_a21oi_1 _07342_ (.A1(_01677_),
    .A2(_01748_),
    .Y(_01828_),
    .B1(_01827_));
 sg13g2_mux4_1 _07343_ (.S0(_01737_),
    .A0(_01748_),
    .A1(_01806_),
    .A2(_01826_),
    .A3(_01814_),
    .S1(net1748),
    .X(_01829_));
 sg13g2_nand4_1 _07344_ (.B(_01721_),
    .C(_01733_),
    .A(_01709_),
    .Y(_01830_),
    .D(_01829_));
 sg13g2_xnor2_1 _07345_ (.Y(_01831_),
    .A(_01771_),
    .B(_01772_));
 sg13g2_inv_1 _07346_ (.Y(_01832_),
    .A(_01831_));
 sg13g2_a21oi_1 _07347_ (.A1(_01824_),
    .A2(_01830_),
    .Y(_01833_),
    .B1(_01832_));
 sg13g2_nand4_1 _07348_ (.B(_01721_),
    .C(_01732_),
    .A(_01709_),
    .Y(_01834_),
    .D(_01807_));
 sg13g2_a21oi_1 _07349_ (.A1(net1748),
    .A2(_01748_),
    .Y(_01835_),
    .B1(net1506));
 sg13g2_nor2_1 _07350_ (.A(_01677_),
    .B(_01741_),
    .Y(_01836_));
 sg13g2_a21oi_1 _07351_ (.A1(_01677_),
    .A2(_01826_),
    .Y(_01837_),
    .B1(_01836_));
 sg13g2_a22oi_1 _07352_ (.Y(_01838_),
    .B1(_01837_),
    .B2(net1506),
    .A2(_01835_),
    .A1(_01819_));
 sg13g2_nand4_1 _07353_ (.B(_01721_),
    .C(_01733_),
    .A(_01709_),
    .Y(_01839_),
    .D(_01838_));
 sg13g2_a21oi_1 _07354_ (.A1(_01834_),
    .A2(_01839_),
    .Y(_01840_),
    .B1(_01770_));
 sg13g2_nand3_1 _07355_ (.B(_01830_),
    .C(_01832_),
    .A(_01824_),
    .Y(_01841_));
 sg13g2_nor2b_1 _07356_ (.A(_01833_),
    .B_N(_01841_),
    .Y(_01842_));
 sg13g2_a21o_1 _07357_ (.A2(_01841_),
    .A1(_01840_),
    .B1(_01833_),
    .X(_01843_));
 sg13g2_xor2_1 _07358_ (.B(_01822_),
    .A(_01821_),
    .X(_01844_));
 sg13g2_a21oi_1 _07359_ (.A1(_01843_),
    .A2(_01844_),
    .Y(_01845_),
    .B1(_01823_));
 sg13g2_xor2_1 _07360_ (.B(_01817_),
    .A(_01816_),
    .X(_01846_));
 sg13g2_o21ai_1 _07361_ (.B1(_01818_),
    .Y(_01847_),
    .A1(_01845_),
    .A2(_01846_));
 sg13g2_a21oi_1 _07362_ (.A1(_01812_),
    .A2(_01847_),
    .Y(_01848_),
    .B1(_01811_));
 sg13g2_o21ai_1 _07363_ (.B1(_01802_),
    .Y(_01849_),
    .A1(_01804_),
    .A2(_01848_));
 sg13g2_a21oi_1 _07364_ (.A1(_01796_),
    .A2(_01849_),
    .Y(_01850_),
    .B1(_01794_));
 sg13g2_xnor2_1 _07365_ (.Y(_01851_),
    .A(_01767_),
    .B(_01786_));
 sg13g2_inv_1 _07366_ (.Y(_01852_),
    .A(_01851_));
 sg13g2_o21ai_1 _07367_ (.B1(_01787_),
    .Y(_01853_),
    .A1(_01850_),
    .A2(_01852_));
 sg13g2_xor2_1 _07368_ (.B(_01853_),
    .A(_01731_),
    .X(_01854_));
 sg13g2_a21oi_2 _07369_ (.B1(_01729_),
    .Y(_01855_),
    .A2(_01853_),
    .A1(_01730_));
 sg13g2_xnor2_1 _07370_ (.Y(_01856_),
    .A(_01850_),
    .B(_01851_));
 sg13g2_nand2_1 _07371_ (.Y(_01857_),
    .A(_01855_),
    .B(_01856_));
 sg13g2_nor2_1 _07372_ (.A(_01806_),
    .B(_01814_),
    .Y(_01858_));
 sg13g2_a22oi_1 _07373_ (.Y(_01859_),
    .B1(_01858_),
    .B2(_01805_),
    .A2(_01819_),
    .A1(net1506));
 sg13g2_o21ai_1 _07374_ (.B1(_01741_),
    .Y(_01860_),
    .A1(net1749),
    .A2(_01744_));
 sg13g2_a21o_1 _07375_ (.A2(_01860_),
    .A1(_01737_),
    .B1(_01732_),
    .X(_01861_));
 sg13g2_and2_1 _07376_ (.A(_01722_),
    .B(_01861_),
    .X(_01862_));
 sg13g2_o21ai_1 _07377_ (.B1(_01862_),
    .Y(_01863_),
    .A1(_01749_),
    .A2(_01859_));
 sg13g2_inv_1 _07378_ (.Y(_01864_),
    .A(_01863_));
 sg13g2_xnor2_1 _07379_ (.Y(_01865_),
    .A(_01803_),
    .B(_01848_));
 sg13g2_xor2_1 _07380_ (.B(_01847_),
    .A(_01812_),
    .X(_01866_));
 sg13g2_xor2_1 _07381_ (.B(_01846_),
    .A(_01845_),
    .X(_01867_));
 sg13g2_inv_1 _07382_ (.Y(_01868_),
    .A(_01867_));
 sg13g2_xnor2_1 _07383_ (.Y(_01869_),
    .A(_01843_),
    .B(_01844_));
 sg13g2_nand3_1 _07384_ (.B(_01834_),
    .C(_01839_),
    .A(_01770_),
    .Y(_01870_));
 sg13g2_nand2b_2 _07385_ (.Y(_01871_),
    .B(_01870_),
    .A_N(_01840_));
 sg13g2_nor2_1 _07386_ (.A(net1749),
    .B(_01741_),
    .Y(_01872_));
 sg13g2_nor2_1 _07387_ (.A(_01737_),
    .B(_01872_),
    .Y(_01873_));
 sg13g2_a21oi_1 _07388_ (.A1(_01737_),
    .A2(_01828_),
    .Y(_01874_),
    .B1(_01873_));
 sg13g2_a22oi_1 _07389_ (.Y(_01875_),
    .B1(_01874_),
    .B2(_01734_),
    .A2(_01815_),
    .A1(_01813_));
 sg13g2_inv_1 _07390_ (.Y(_01876_),
    .A(_01875_));
 sg13g2_nand2_1 _07391_ (.Y(_01877_),
    .A(_01871_),
    .B(_01875_));
 sg13g2_inv_1 _07392_ (.Y(_01878_),
    .A(_01877_));
 sg13g2_xnor2_1 _07393_ (.Y(_01879_),
    .A(_01840_),
    .B(_01842_));
 sg13g2_nand2_1 _07394_ (.Y(_01880_),
    .A(_01869_),
    .B(_01879_));
 sg13g2_inv_1 _07395_ (.Y(_01881_),
    .A(_01880_));
 sg13g2_or4_1 _07396_ (.A(_01866_),
    .B(_01867_),
    .C(_01877_),
    .D(_01880_),
    .X(_01882_));
 sg13g2_nor2_1 _07397_ (.A(_01865_),
    .B(_01882_),
    .Y(_01883_));
 sg13g2_nand2_1 _07398_ (.Y(_01884_),
    .A(_01863_),
    .B(_01883_));
 sg13g2_nor2_1 _07399_ (.A(_01864_),
    .B(_01877_),
    .Y(_01885_));
 sg13g2_nor2b_1 _07400_ (.A(_01880_),
    .B_N(_01885_),
    .Y(_01886_));
 sg13g2_a221oi_1 _07401_ (.B2(_01875_),
    .C1(_01729_),
    .B1(_01863_),
    .A1(_01731_),
    .Y(_01887_),
    .A2(_01853_));
 sg13g2_a221oi_1 _07402_ (.B2(_01878_),
    .C1(_01729_),
    .B1(_01863_),
    .A1(_01730_),
    .Y(_01888_),
    .A2(_01853_));
 sg13g2_a221oi_1 _07403_ (.B2(_01885_),
    .C1(_01729_),
    .B1(_01881_),
    .A1(_01731_),
    .Y(_01889_),
    .A2(_01853_));
 sg13g2_a221oi_1 _07404_ (.B2(_01886_),
    .C1(_01729_),
    .B1(_01868_),
    .A1(_01731_),
    .Y(_01890_),
    .A2(_01853_));
 sg13g2_o21ai_1 _07405_ (.B1(_01855_),
    .Y(_01891_),
    .A1(_01864_),
    .A2(_01882_));
 sg13g2_nand2_1 _07406_ (.Y(_01892_),
    .A(_01855_),
    .B(_01884_));
 sg13g2_xnor2_1 _07407_ (.Y(_01893_),
    .A(_01796_),
    .B(_01849_));
 sg13g2_inv_1 _07408_ (.Y(_01894_),
    .A(_01893_));
 sg13g2_o21ai_1 _07409_ (.B1(_01855_),
    .Y(_01895_),
    .A1(_01884_),
    .A2(_01894_));
 sg13g2_and2_1 _07410_ (.A(_01857_),
    .B(_01895_),
    .X(_01896_));
 sg13g2_xor2_1 _07411_ (.B(_01896_),
    .A(_01854_),
    .X(_01897_));
 sg13g2_xnor2_1 _07412_ (.Y(_01898_),
    .A(_01854_),
    .B(_01896_));
 sg13g2_nor4_1 _07413_ (.A(_01697_),
    .B(_01702_),
    .C(_01707_),
    .D(_01718_),
    .Y(_01899_));
 sg13g2_nand2_1 _07414_ (.Y(_01900_),
    .A(_01710_),
    .B(_01712_));
 sg13g2_nand3b_1 _07415_ (.B(_01692_),
    .C(_01899_),
    .Y(_01901_),
    .A_N(_01671_));
 sg13g2_nor3_1 _07416_ (.A(net1451),
    .B(_01900_),
    .C(_01901_),
    .Y(_01902_));
 sg13g2_and3_1 _07417_ (.X(_01903_),
    .A(_01855_),
    .B(_01864_),
    .C(_01876_));
 sg13g2_a21oi_2 _07418_ (.B1(_01876_),
    .Y(_01904_),
    .A2(_01864_),
    .A1(_01855_));
 sg13g2_nor2_2 _07419_ (.A(_01903_),
    .B(_01904_),
    .Y(_01905_));
 sg13g2_xor2_1 _07420_ (.B(_01887_),
    .A(_01871_),
    .X(_01906_));
 sg13g2_xnor2_1 _07421_ (.Y(_01907_),
    .A(_01871_),
    .B(_01887_));
 sg13g2_o21ai_1 _07422_ (.B1(_01906_),
    .Y(_01908_),
    .A1(_01903_),
    .A2(_01904_));
 sg13g2_xnor2_1 _07423_ (.Y(_01909_),
    .A(_01879_),
    .B(_01888_));
 sg13g2_xor2_1 _07424_ (.B(_01888_),
    .A(_01879_),
    .X(_01910_));
 sg13g2_a221oi_1 _07425_ (.B2(_01885_),
    .C1(_01729_),
    .B1(_01879_),
    .A1(_01730_),
    .Y(_01911_),
    .A2(_01853_));
 sg13g2_xnor2_1 _07426_ (.Y(_01912_),
    .A(_01869_),
    .B(_01911_));
 sg13g2_inv_1 _07427_ (.Y(_01913_),
    .A(_01912_));
 sg13g2_nor2_1 _07428_ (.A(_01909_),
    .B(_01912_),
    .Y(_01914_));
 sg13g2_nand2b_1 _07429_ (.Y(_01915_),
    .B(_01914_),
    .A_N(_01908_));
 sg13g2_xnor2_1 _07430_ (.Y(_01916_),
    .A(_01865_),
    .B(_01891_));
 sg13g2_xor2_1 _07431_ (.B(_01891_),
    .A(_01865_),
    .X(_01917_));
 sg13g2_xnor2_1 _07432_ (.Y(_01918_),
    .A(_01892_),
    .B(_01894_));
 sg13g2_xnor2_1 _07433_ (.Y(_01919_),
    .A(_01892_),
    .B(_01893_));
 sg13g2_nor2_1 _07434_ (.A(_01916_),
    .B(net1462),
    .Y(_01920_));
 sg13g2_nand2_1 _07435_ (.Y(_01921_),
    .A(_01917_),
    .B(_01919_));
 sg13g2_xnor2_1 _07436_ (.Y(_01922_),
    .A(_01867_),
    .B(_01889_));
 sg13g2_inv_1 _07437_ (.Y(_01923_),
    .A(_01922_));
 sg13g2_xor2_1 _07438_ (.B(_01890_),
    .A(_01866_),
    .X(_01924_));
 sg13g2_xnor2_1 _07439_ (.Y(_01925_),
    .A(_01866_),
    .B(_01890_));
 sg13g2_nand2_1 _07440_ (.Y(_01926_),
    .A(net1469),
    .B(_01925_));
 sg13g2_nor3_1 _07441_ (.A(_01916_),
    .B(net1462),
    .C(_01926_),
    .Y(_01927_));
 sg13g2_nand3_1 _07442_ (.B(_01915_),
    .C(_01927_),
    .A(_01702_),
    .Y(_01928_));
 sg13g2_nor2_2 _07443_ (.A(_01917_),
    .B(net1462),
    .Y(_01929_));
 sg13g2_nor3_1 _07444_ (.A(_01903_),
    .B(_01904_),
    .C(_01912_),
    .Y(_01930_));
 sg13g2_nor2_1 _07445_ (.A(_01923_),
    .B(_01930_),
    .Y(_01931_));
 sg13g2_a21oi_1 _07446_ (.A1(_01907_),
    .A2(net1469),
    .Y(_01932_),
    .B1(_01924_));
 sg13g2_o21ai_1 _07447_ (.B1(_01925_),
    .Y(_01933_),
    .A1(_01906_),
    .A2(_01923_));
 sg13g2_o21ai_1 _07448_ (.B1(_01932_),
    .Y(_01934_),
    .A1(_01923_),
    .A2(_01930_));
 sg13g2_nand2_1 _07449_ (.Y(_01935_),
    .A(_01909_),
    .B(_01925_));
 sg13g2_nand2b_1 _07450_ (.Y(_01936_),
    .B(_01913_),
    .A_N(_01935_));
 sg13g2_nand2_1 _07451_ (.Y(_01937_),
    .A(_01934_),
    .B(_01936_));
 sg13g2_nand3_1 _07452_ (.B(_01934_),
    .C(_01936_),
    .A(_01917_),
    .Y(_01938_));
 sg13g2_and2_1 _07453_ (.A(_01919_),
    .B(_01938_),
    .X(_01939_));
 sg13g2_a21oi_1 _07454_ (.A1(_01908_),
    .A2(_01914_),
    .Y(_01940_),
    .B1(_01926_));
 sg13g2_nor2_1 _07455_ (.A(_01921_),
    .B(_01940_),
    .Y(_01941_));
 sg13g2_nor2_1 _07456_ (.A(_01697_),
    .B(_01941_),
    .Y(_01942_));
 sg13g2_a221oi_1 _07457_ (.B2(_01692_),
    .C1(_01941_),
    .B1(_01939_),
    .A1(_01695_),
    .Y(_01943_),
    .A2(_01696_));
 sg13g2_o21ai_1 _07458_ (.B1(_01928_),
    .Y(_01944_),
    .A1(_01706_),
    .A2(_01943_));
 sg13g2_xor2_1 _07459_ (.B(_01895_),
    .A(_01856_),
    .X(_01945_));
 sg13g2_inv_2 _07460_ (.Y(_01946_),
    .A(net1460));
 sg13g2_nor2_2 _07461_ (.A(net1449),
    .B(_01946_),
    .Y(_01947_));
 sg13g2_nand4_1 _07462_ (.B(_01713_),
    .C(_01718_),
    .A(_01671_),
    .Y(_01948_),
    .D(_01947_));
 sg13g2_a21o_1 _07463_ (.A2(_01927_),
    .A1(_01915_),
    .B1(_01702_),
    .X(_01949_));
 sg13g2_and2_1 _07464_ (.A(_01707_),
    .B(_01949_),
    .X(_01950_));
 sg13g2_inv_1 _07465_ (.Y(_01951_),
    .A(_01950_));
 sg13g2_nand2b_1 _07466_ (.Y(_01952_),
    .B(_01919_),
    .A_N(_01692_));
 sg13g2_nand4_1 _07467_ (.B(_01937_),
    .C(_01941_),
    .A(_01697_),
    .Y(_01953_),
    .D(_01952_));
 sg13g2_a21oi_1 _07468_ (.A1(_01951_),
    .A2(_01953_),
    .Y(_01954_),
    .B1(_01948_));
 sg13g2_nor4_2 _07469_ (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][6] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][15] ),
    .C(_01636_),
    .Y(_01955_),
    .D(_01642_));
 sg13g2_nand2_1 _07470_ (.Y(_01956_),
    .A(_01883_),
    .B(_01893_));
 sg13g2_nor3_1 _07471_ (.A(_01854_),
    .B(_01856_),
    .C(_01956_),
    .Y(_01957_));
 sg13g2_or2_1 _07472_ (.X(_01958_),
    .B(_01957_),
    .A(net1723));
 sg13g2_nand2b_1 _07473_ (.Y(_01959_),
    .B(_01698_),
    .A_N(_01692_));
 sg13g2_a21o_2 _07474_ (.A2(_01954_),
    .A1(_01944_),
    .B1(_01958_),
    .X(_01960_));
 sg13g2_inv_1 _07475_ (.Y(_01961_),
    .A(_01960_));
 sg13g2_nor2_2 _07476_ (.A(_01902_),
    .B(_01960_),
    .Y(_01962_));
 sg13g2_nor2_1 _07477_ (.A(_01919_),
    .B(_01946_),
    .Y(_01963_));
 sg13g2_a221oi_1 _07478_ (.B2(_01905_),
    .C1(net1450),
    .B1(_01963_),
    .A1(_01907_),
    .Y(_01964_),
    .A2(_01946_));
 sg13g2_a21oi_1 _07479_ (.A1(net1449),
    .A2(_01910_),
    .Y(_01965_),
    .B1(_01964_));
 sg13g2_nand3b_1 _07480_ (.B(_01626_),
    .C(_01646_),
    .Y(_01966_),
    .A_N(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][15] ));
 sg13g2_nor2b_1 _07481_ (.A(_01649_),
    .B_N(_01966_),
    .Y(_01967_));
 sg13g2_nand2b_1 _07482_ (.Y(_01968_),
    .B(_01966_),
    .A_N(_01649_));
 sg13g2_a221oi_1 _07483_ (.B2(_01965_),
    .C1(net1547),
    .B1(_01962_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][0] ),
    .Y(_01969_),
    .A2(net1723));
 sg13g2_o21ai_1 _07484_ (.B1(net1668),
    .Y(_01970_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][0] ),
    .A2(net1548));
 sg13g2_nor2_1 _07485_ (.A(_01969_),
    .B(_01970_),
    .Y(_01971_));
 sg13g2_nor2_1 _07486_ (.A(_01654_),
    .B(_01971_),
    .Y(_01972_));
 sg13g2_nor2_1 _07487_ (.A(net1675),
    .B(_01972_),
    .Y(_01973_));
 sg13g2_o21ai_1 _07488_ (.B1(_01973_),
    .Y(_01974_),
    .A1(net1530),
    .A2(_01623_));
 sg13g2_nor4_1 _07489_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][11] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][12] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][13] ),
    .D(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][14] ),
    .Y(_01975_));
 sg13g2_nor4_1 _07490_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][7] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][8] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][9] ),
    .D(net1786),
    .Y(_01976_));
 sg13g2_nand2_1 _07491_ (.Y(_01977_),
    .A(_01975_),
    .B(_01976_));
 sg13g2_inv_1 _07492_ (.Y(_01978_),
    .A(_01977_));
 sg13g2_nand4_1 _07493_ (.B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][12] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][13] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][11] ),
    .Y(_01979_),
    .D(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][14] ));
 sg13g2_nand4_1 _07494_ (.B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][8] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][9] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][7] ),
    .Y(_01980_),
    .D(net1786));
 sg13g2_o21ai_1 _07495_ (.B1(_01977_),
    .Y(_01981_),
    .A1(_01979_),
    .A2(_01980_));
 sg13g2_nor2_1 _07496_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][1] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][0] ),
    .Y(_01982_));
 sg13g2_nor4_1 _07497_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][3] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][2] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][5] ),
    .D(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][4] ),
    .Y(_01983_));
 sg13g2_nand2_2 _07498_ (.Y(_01984_),
    .A(_01982_),
    .B(_01983_));
 sg13g2_o21ai_1 _07499_ (.B1(_01981_),
    .Y(_01985_),
    .A1(_00675_),
    .A2(_01984_));
 sg13g2_nor3_1 _07500_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][12] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][11] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][14] ),
    .Y(_01986_));
 sg13g2_nor4_1 _07501_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][8] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][7] ),
    .C(net1785),
    .D(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][9] ),
    .Y(_01987_));
 sg13g2_nand3_1 _07502_ (.B(_01986_),
    .C(_01987_),
    .A(_00674_),
    .Y(_01988_));
 sg13g2_inv_1 _07503_ (.Y(_01989_),
    .A(_01988_));
 sg13g2_nand4_1 _07504_ (.B(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][11] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][14] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][12] ),
    .Y(_01990_),
    .D(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][13] ));
 sg13g2_nand4_1 _07505_ (.B(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][7] ),
    .C(net1785),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][8] ),
    .Y(_01991_),
    .D(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][9] ));
 sg13g2_or2_1 _07506_ (.X(_01992_),
    .B(_01991_),
    .A(_01990_));
 sg13g2_nor2_1 _07507_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][1] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][0] ),
    .Y(_01993_));
 sg13g2_nor4_1 _07508_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][3] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][2] ),
    .C(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][5] ),
    .D(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][4] ),
    .Y(_01994_));
 sg13g2_nand2_2 _07509_ (.Y(_01995_),
    .A(_01993_),
    .B(_01994_));
 sg13g2_inv_1 _07510_ (.Y(_01996_),
    .A(_01995_));
 sg13g2_a22oi_1 _07511_ (.Y(_01997_),
    .B1(_01996_),
    .B2(_00018_),
    .A2(_01992_),
    .A1(_01988_));
 sg13g2_a221oi_1 _07512_ (.B2(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][15] ),
    .C1(_01997_),
    .B1(_01989_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][15] ),
    .Y(_01998_),
    .A2(_01978_));
 sg13g2_nand2_1 _07513_ (.Y(_01999_),
    .A(_01985_),
    .B(_01998_));
 sg13g2_nor4_2 _07514_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][6] ),
    .B(_01979_),
    .C(_01980_),
    .Y(_02000_),
    .D(_01984_));
 sg13g2_a21o_1 _07515_ (.A2(_02000_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][15] ),
    .B1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][15] ),
    .X(_02001_));
 sg13g2_nor3_2 _07516_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][6] ),
    .B(_01992_),
    .C(_01995_),
    .Y(_02002_));
 sg13g2_or3_2 _07517_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][6] ),
    .B(_01992_),
    .C(_01995_),
    .X(_02003_));
 sg13g2_a21oi_1 _07518_ (.A1(_02001_),
    .A2(_02002_),
    .Y(_02004_),
    .B1(_01999_));
 sg13g2_xor2_1 _07519_ (.B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][15] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][15] ),
    .X(_02005_));
 sg13g2_nand3_1 _07520_ (.B(_02002_),
    .C(_02005_),
    .A(_02000_),
    .Y(_02006_));
 sg13g2_nand3_1 _07521_ (.B(_01998_),
    .C(_02006_),
    .A(_01985_),
    .Y(_02007_));
 sg13g2_nand2b_1 _07522_ (.Y(_02008_),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][11] ),
    .A_N(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][11] ));
 sg13g2_xor2_1 _07523_ (.B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][11] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][11] ),
    .X(_02009_));
 sg13g2_nand2b_1 _07524_ (.Y(_02010_),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][12] ),
    .A_N(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][12] ));
 sg13g2_nor2b_1 _07525_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][12] ),
    .B_N(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][12] ),
    .Y(_02011_));
 sg13g2_xor2_1 _07526_ (.B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][12] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][12] ),
    .X(_02012_));
 sg13g2_xor2_1 _07527_ (.B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][13] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][13] ),
    .X(_02013_));
 sg13g2_inv_1 _07528_ (.Y(_02014_),
    .A(_02013_));
 sg13g2_nor3_2 _07529_ (.A(_02009_),
    .B(_02012_),
    .C(_02013_),
    .Y(_02015_));
 sg13g2_nand2b_1 _07530_ (.Y(_02016_),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][10] ),
    .A_N(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][10] ));
 sg13g2_nor2b_1 _07531_ (.A(net1786),
    .B_N(net1785),
    .Y(_02017_));
 sg13g2_xnor2_1 _07532_ (.Y(_02018_),
    .A(net1785),
    .B(net1786));
 sg13g2_xor2_1 _07533_ (.B(net1786),
    .A(net1785),
    .X(_02019_));
 sg13g2_nand2b_1 _07534_ (.Y(_02020_),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][9] ),
    .A_N(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][9] ));
 sg13g2_xnor2_1 _07535_ (.Y(_02021_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][9] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][9] ));
 sg13g2_nand2b_1 _07536_ (.Y(_02022_),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][8] ),
    .A_N(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][8] ));
 sg13g2_nor2b_1 _07537_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][8] ),
    .B_N(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][8] ),
    .Y(_02023_));
 sg13g2_xnor2_1 _07538_ (.Y(_02024_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][8] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][8] ));
 sg13g2_nor2b_1 _07539_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][14] ),
    .B_N(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][14] ),
    .Y(_02025_));
 sg13g2_nor2_2 _07540_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][14] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][14] ),
    .Y(_02026_));
 sg13g2_xor2_1 _07541_ (.B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][14] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][14] ),
    .X(_02027_));
 sg13g2_nor2b_1 _07542_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][7] ),
    .B_N(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][7] ),
    .Y(_02028_));
 sg13g2_o21ai_1 _07543_ (.B1(_02022_),
    .Y(_02029_),
    .A1(_02023_),
    .A2(_02028_));
 sg13g2_nand4_1 _07544_ (.B(_02018_),
    .C(_02021_),
    .A(_02015_),
    .Y(_02030_),
    .D(_02029_));
 sg13g2_o21ai_1 _07545_ (.B1(_02016_),
    .Y(_02031_),
    .A1(_02017_),
    .A2(_02020_));
 sg13g2_a221oi_1 _07546_ (.B2(_02010_),
    .C1(_02011_),
    .B1(_02008_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][13] ),
    .Y(_02032_),
    .A2(_00678_));
 sg13g2_a221oi_1 _07547_ (.B2(_02031_),
    .C1(_02032_),
    .B1(_02015_),
    .A1(_00674_),
    .Y(_02033_),
    .A2(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][13] ));
 sg13g2_a21oi_1 _07548_ (.A1(_02030_),
    .A2(_02033_),
    .Y(_02034_),
    .B1(_02027_));
 sg13g2_nor2_1 _07549_ (.A(_02025_),
    .B(_02034_),
    .Y(_02035_));
 sg13g2_xnor2_1 _07550_ (.Y(_02036_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][7] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][7] ));
 sg13g2_xor2_1 _07551_ (.B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][7] ),
    .A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][7] ),
    .X(_02037_));
 sg13g2_and4_1 _07552_ (.A(_02015_),
    .B(_02018_),
    .C(_02021_),
    .D(_02036_),
    .X(_02038_));
 sg13g2_nand3b_1 _07553_ (.B(_02038_),
    .C(_02024_),
    .Y(_02039_),
    .A_N(_02027_));
 sg13g2_o21ai_1 _07554_ (.B1(_02039_),
    .Y(_02040_),
    .A1(_02025_),
    .A2(_02034_));
 sg13g2_nand2b_1 _07555_ (.Y(_02041_),
    .B(net1543),
    .A_N(_00023_));
 sg13g2_mux2_2 _07556_ (.A0(_00022_),
    .A1(_00023_),
    .S(net1543),
    .X(_02042_));
 sg13g2_o21ai_1 _07557_ (.B1(_02041_),
    .Y(_02043_),
    .A1(_00022_),
    .A2(net1544));
 sg13g2_nand2_1 _07558_ (.Y(_02044_),
    .A(_00023_),
    .B(_00022_));
 sg13g2_nand2_1 _07559_ (.Y(_02045_),
    .A(_02042_),
    .B(_02044_));
 sg13g2_nand3_1 _07560_ (.B(_02042_),
    .C(_02044_),
    .A(_02024_),
    .Y(_02046_));
 sg13g2_mux2_1 _07561_ (.A0(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][8] ),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][8] ),
    .S(_02035_),
    .X(_02047_));
 sg13g2_inv_1 _07562_ (.Y(_02048_),
    .A(_02047_));
 sg13g2_or2_1 _07563_ (.X(_02049_),
    .B(net1527),
    .A(_02024_));
 sg13g2_and3_1 _07564_ (.X(_02050_),
    .A(_02021_),
    .B(_02046_),
    .C(_02049_));
 sg13g2_mux2_1 _07565_ (.A0(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][9] ),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][9] ),
    .S(_02035_),
    .X(_02051_));
 sg13g2_inv_2 _07566_ (.Y(_02052_),
    .A(_02051_));
 sg13g2_nor2_1 _07567_ (.A(_02021_),
    .B(_02052_),
    .Y(_02053_));
 sg13g2_nor3_1 _07568_ (.A(_02019_),
    .B(_02050_),
    .C(_02053_),
    .Y(_02054_));
 sg13g2_or3_1 _07569_ (.A(_02019_),
    .B(_02050_),
    .C(_02053_),
    .X(_02055_));
 sg13g2_mux2_2 _07570_ (.A0(net1786),
    .A1(net1785),
    .S(net1544),
    .X(_02056_));
 sg13g2_inv_1 _07571_ (.Y(_02057_),
    .A(_02056_));
 sg13g2_nor2_1 _07572_ (.A(_02018_),
    .B(_02056_),
    .Y(_02058_));
 sg13g2_nand2_1 _07573_ (.Y(_02059_),
    .A(_02019_),
    .B(_02057_));
 sg13g2_nor3_2 _07574_ (.A(_02015_),
    .B(_02054_),
    .C(_02058_),
    .Y(_02060_));
 sg13g2_nand2b_1 _07575_ (.Y(_02061_),
    .B(net1543),
    .A_N(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][11] ));
 sg13g2_mux2_2 _07576_ (.A0(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][11] ),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][11] ),
    .S(net1543),
    .X(_02062_));
 sg13g2_o21ai_1 _07577_ (.B1(_02061_),
    .Y(_02063_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][11] ),
    .A2(net1543));
 sg13g2_mux2_2 _07578_ (.A0(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][12] ),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][12] ),
    .S(net1543),
    .X(_02064_));
 sg13g2_nor2_2 _07579_ (.A(_02062_),
    .B(_02064_),
    .Y(_02065_));
 sg13g2_a21oi_1 _07580_ (.A1(_02014_),
    .A2(_02062_),
    .Y(_02066_),
    .B1(_02012_));
 sg13g2_a21oi_1 _07581_ (.A1(_02014_),
    .A2(_02065_),
    .Y(_02067_),
    .B1(_02066_));
 sg13g2_a22oi_1 _07582_ (.Y(_02068_),
    .B1(_02064_),
    .B2(_02013_),
    .A2(_02062_),
    .A1(_02012_));
 sg13g2_and2_1 _07583_ (.A(_02067_),
    .B(_02068_),
    .X(_02069_));
 sg13g2_a22oi_1 _07584_ (.Y(_02070_),
    .B1(_02069_),
    .B2(_02009_),
    .A2(_02059_),
    .A1(_02055_));
 sg13g2_o21ai_1 _07585_ (.B1(_02019_),
    .Y(_02071_),
    .A1(_02050_),
    .A2(_02053_));
 sg13g2_nor2_1 _07586_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][13] ),
    .B(net1543),
    .Y(_02072_));
 sg13g2_a21oi_2 _07587_ (.B1(_02072_),
    .Y(_02073_),
    .A2(net1543),
    .A1(_00674_));
 sg13g2_o21ai_1 _07588_ (.B1(_02027_),
    .Y(_02074_),
    .A1(_02014_),
    .A2(_02073_));
 sg13g2_nand3_1 _07589_ (.B(_02071_),
    .C(_02074_),
    .A(_02055_),
    .Y(_02075_));
 sg13g2_nor3_2 _07590_ (.A(_02060_),
    .B(_02070_),
    .C(_02075_),
    .Y(_02076_));
 sg13g2_nand2b_1 _07591_ (.Y(_02077_),
    .B(net1541),
    .A_N(_00021_));
 sg13g2_mux2_1 _07592_ (.A0(_00020_),
    .A1(_00021_),
    .S(net1541),
    .X(_02078_));
 sg13g2_o21ai_1 _07593_ (.B1(_02077_),
    .Y(_02079_),
    .A1(_00020_),
    .A2(net1541));
 sg13g2_nand2_2 _07594_ (.Y(_02080_),
    .A(_02076_),
    .B(_02079_));
 sg13g2_mux2_1 _07595_ (.A0(_00021_),
    .A1(_00020_),
    .S(net1541),
    .X(_02081_));
 sg13g2_and2_2 _07596_ (.A(_02080_),
    .B(net1526),
    .X(_02082_));
 sg13g2_xor2_1 _07597_ (.B(net1526),
    .A(_02080_),
    .X(_02083_));
 sg13g2_a21oi_1 _07598_ (.A1(_02046_),
    .A2(_02049_),
    .Y(_02084_),
    .B1(_02021_));
 sg13g2_nor2_2 _07599_ (.A(_02050_),
    .B(_02084_),
    .Y(_02085_));
 sg13g2_inv_1 _07600_ (.Y(_02086_),
    .A(_02085_));
 sg13g2_nor4_2 _07601_ (.A(_02060_),
    .B(_02070_),
    .C(_02075_),
    .Y(_02087_),
    .D(_02085_));
 sg13g2_nand2_1 _07602_ (.Y(_02088_),
    .A(_02076_),
    .B(_02086_));
 sg13g2_nand2_2 _07603_ (.Y(_02089_),
    .A(_02080_),
    .B(_02088_));
 sg13g2_xnor2_1 _07604_ (.Y(_02090_),
    .A(_02024_),
    .B(_02045_));
 sg13g2_xor2_1 _07605_ (.B(_02045_),
    .A(_02024_),
    .X(_02091_));
 sg13g2_nor2_1 _07606_ (.A(_02079_),
    .B(net1502),
    .Y(_02092_));
 sg13g2_mux2_2 _07607_ (.A0(_00035_),
    .A1(_00034_),
    .S(net1542),
    .X(_02093_));
 sg13g2_mux2_2 _07608_ (.A0(_00033_),
    .A1(_00032_),
    .S(net1540),
    .X(_02094_));
 sg13g2_mux2_1 _07609_ (.A0(_00031_),
    .A1(_00030_),
    .S(net1542),
    .X(_02095_));
 sg13g2_nand3_1 _07610_ (.B(_02094_),
    .C(_02095_),
    .A(_02093_),
    .Y(_02096_));
 sg13g2_mux2_1 _07611_ (.A0(_00029_),
    .A1(_00028_),
    .S(net1540),
    .X(_02097_));
 sg13g2_nand4_1 _07612_ (.B(_02094_),
    .C(_02095_),
    .A(_02093_),
    .Y(_02098_),
    .D(_02097_));
 sg13g2_nand2b_1 _07613_ (.Y(_02099_),
    .B(net1540),
    .A_N(_00026_));
 sg13g2_o21ai_1 _07614_ (.B1(_02099_),
    .Y(_02100_),
    .A1(_00027_),
    .A2(net1541));
 sg13g2_mux2_1 _07615_ (.A0(_00025_),
    .A1(_00024_),
    .S(net1540),
    .X(_02101_));
 sg13g2_nand2_1 _07616_ (.Y(_02102_),
    .A(_02079_),
    .B(_02096_));
 sg13g2_nand2_1 _07617_ (.Y(_02103_),
    .A(_02079_),
    .B(_02098_));
 sg13g2_o21ai_1 _07618_ (.B1(_02079_),
    .Y(_02104_),
    .A1(_02098_),
    .A2(_02100_));
 sg13g2_or2_1 _07619_ (.X(_02105_),
    .B(_02101_),
    .A(_02078_));
 sg13g2_nor2_1 _07620_ (.A(_00018_),
    .B(net1541),
    .Y(_02106_));
 sg13g2_a21oi_1 _07621_ (.A1(_00675_),
    .A2(net1541),
    .Y(_02107_),
    .B1(_02106_));
 sg13g2_nand3_1 _07622_ (.B(_02105_),
    .C(_02107_),
    .A(_02104_),
    .Y(_02108_));
 sg13g2_nand2_1 _07623_ (.Y(_02109_),
    .A(_02079_),
    .B(_02108_));
 sg13g2_nor2_1 _07624_ (.A(net1746),
    .B(_02078_),
    .Y(_02110_));
 sg13g2_a21oi_1 _07625_ (.A1(net1746),
    .A2(_02109_),
    .Y(_02111_),
    .B1(_02110_));
 sg13g2_a21oi_1 _07626_ (.A1(net1502),
    .A2(_02111_),
    .Y(_02112_),
    .B1(_02092_));
 sg13g2_o21ai_1 _07627_ (.B1(_02089_),
    .Y(_02113_),
    .A1(_02085_),
    .A2(_02112_));
 sg13g2_mux2_2 _07628_ (.A0(_00034_),
    .A1(_00035_),
    .S(net1542),
    .X(_02114_));
 sg13g2_mux2_1 _07629_ (.A0(_00032_),
    .A1(_00033_),
    .S(net1540),
    .X(_02115_));
 sg13g2_nor2_1 _07630_ (.A(net1526),
    .B(_02114_),
    .Y(_02116_));
 sg13g2_a21oi_1 _07631_ (.A1(_02114_),
    .A2(_02115_),
    .Y(_02117_),
    .B1(net1526));
 sg13g2_mux2_1 _07632_ (.A0(_00030_),
    .A1(_00031_),
    .S(net1542),
    .X(_02118_));
 sg13g2_nor2b_1 _07633_ (.A(_02117_),
    .B_N(_02118_),
    .Y(_02119_));
 sg13g2_mux2_1 _07634_ (.A0(_00028_),
    .A1(_00029_),
    .S(net1540),
    .X(_02120_));
 sg13g2_mux2_1 _07635_ (.A0(_00026_),
    .A1(_00027_),
    .S(net1540),
    .X(_02121_));
 sg13g2_mux2_1 _07636_ (.A0(_00024_),
    .A1(_00025_),
    .S(net1540),
    .X(_02122_));
 sg13g2_nand2_1 _07637_ (.Y(_02123_),
    .A(_00018_),
    .B(net1542));
 sg13g2_o21ai_1 _07638_ (.B1(_02123_),
    .Y(_02124_),
    .A1(_00675_),
    .A2(net1542));
 sg13g2_nor2_1 _07639_ (.A(_02081_),
    .B(_02119_),
    .Y(_02125_));
 sg13g2_a21o_1 _07640_ (.A2(_02120_),
    .A1(_02119_),
    .B1(net1526),
    .X(_02126_));
 sg13g2_o21ai_1 _07641_ (.B1(_02126_),
    .Y(_02127_),
    .A1(net1526),
    .A2(_02121_));
 sg13g2_nor2_1 _07642_ (.A(net1526),
    .B(_02122_),
    .Y(_02128_));
 sg13g2_nor2_1 _07643_ (.A(_02127_),
    .B(_02128_),
    .Y(_02129_));
 sg13g2_o21ai_1 _07644_ (.B1(_02129_),
    .Y(_02130_),
    .A1(net1526),
    .A2(_02124_));
 sg13g2_or2_1 _07645_ (.X(_02131_),
    .B(_02130_),
    .A(_02113_));
 sg13g2_a21o_1 _07646_ (.A2(_02105_),
    .A1(_02104_),
    .B1(_02107_),
    .X(_02132_));
 sg13g2_and2_1 _07647_ (.A(_02108_),
    .B(_02132_),
    .X(_02133_));
 sg13g2_mux2_1 _07648_ (.A0(_02109_),
    .A1(_02133_),
    .S(net1746),
    .X(_02134_));
 sg13g2_mux2_1 _07649_ (.A0(_02079_),
    .A1(_02134_),
    .S(net1502),
    .X(_02135_));
 sg13g2_o21ai_1 _07650_ (.B1(_02089_),
    .Y(_02136_),
    .A1(_02085_),
    .A2(_02135_));
 sg13g2_xor2_1 _07651_ (.B(_02129_),
    .A(_02124_),
    .X(_02137_));
 sg13g2_nor2b_1 _07652_ (.A(_02136_),
    .B_N(_02137_),
    .Y(_02138_));
 sg13g2_xor2_1 _07653_ (.B(_02104_),
    .A(_02101_),
    .X(_02139_));
 sg13g2_and2_1 _07654_ (.A(net1746),
    .B(_02139_),
    .X(_02140_));
 sg13g2_a21oi_1 _07655_ (.A1(_02037_),
    .A2(_02133_),
    .Y(_02141_),
    .B1(_02140_));
 sg13g2_mux4_1 _07656_ (.S0(net1746),
    .A0(_02079_),
    .A1(_02109_),
    .A2(_02133_),
    .A3(_02139_),
    .S1(net1502),
    .X(_02142_));
 sg13g2_o21ai_1 _07657_ (.B1(_02089_),
    .Y(_02143_),
    .A1(_02085_),
    .A2(_02142_));
 sg13g2_xnor2_1 _07658_ (.Y(_02144_),
    .A(_02122_),
    .B(_02127_));
 sg13g2_nand2b_1 _07659_ (.Y(_02145_),
    .B(_02144_),
    .A_N(_02143_));
 sg13g2_xor2_1 _07660_ (.B(_02144_),
    .A(_02143_),
    .X(_02146_));
 sg13g2_nand2_1 _07661_ (.Y(_02147_),
    .A(_02037_),
    .B(_02139_));
 sg13g2_xnor2_1 _07662_ (.Y(_02148_),
    .A(_02100_),
    .B(_02103_));
 sg13g2_nand2_1 _07663_ (.Y(_02149_),
    .A(net1746),
    .B(_02148_));
 sg13g2_mux4_1 _07664_ (.S0(net1746),
    .A0(_02109_),
    .A1(_02133_),
    .A2(_02139_),
    .A3(_02148_),
    .S1(net1502),
    .X(_02150_));
 sg13g2_o21ai_1 _07665_ (.B1(_02089_),
    .Y(_02151_),
    .A1(_02085_),
    .A2(_02150_));
 sg13g2_xor2_1 _07666_ (.B(_02126_),
    .A(_02121_),
    .X(_02152_));
 sg13g2_nor2b_1 _07667_ (.A(_02151_),
    .B_N(_02152_),
    .Y(_02153_));
 sg13g2_xor2_1 _07668_ (.B(_02152_),
    .A(_02151_),
    .X(_02154_));
 sg13g2_inv_1 _07669_ (.Y(_02155_),
    .A(_02154_));
 sg13g2_nor4_2 _07670_ (.A(_02060_),
    .B(_02070_),
    .C(_02075_),
    .Y(_02156_),
    .D(_02086_));
 sg13g2_xor2_1 _07671_ (.B(_02102_),
    .A(_02097_),
    .X(_02157_));
 sg13g2_mux2_1 _07672_ (.A0(_02148_),
    .A1(_02157_),
    .S(net1746),
    .X(_02158_));
 sg13g2_nor2_1 _07673_ (.A(_02091_),
    .B(_02158_),
    .Y(_02159_));
 sg13g2_a21oi_1 _07674_ (.A1(_02091_),
    .A2(_02141_),
    .Y(_02160_),
    .B1(_02159_));
 sg13g2_a22oi_1 _07675_ (.Y(_02161_),
    .B1(_02160_),
    .B2(_02087_),
    .A2(_02156_),
    .A1(_02112_));
 sg13g2_xnor2_1 _07676_ (.Y(_02162_),
    .A(_02120_),
    .B(_02125_));
 sg13g2_nand2b_1 _07677_ (.Y(_02163_),
    .B(_02162_),
    .A_N(_02161_));
 sg13g2_xor2_1 _07678_ (.B(_02162_),
    .A(_02161_),
    .X(_02164_));
 sg13g2_nand3_1 _07679_ (.B(_02147_),
    .C(_02149_),
    .A(_02091_),
    .Y(_02165_));
 sg13g2_a21oi_1 _07680_ (.A1(_02093_),
    .A2(_02094_),
    .Y(_02166_),
    .B1(_02078_));
 sg13g2_xor2_1 _07681_ (.B(_02166_),
    .A(_02095_),
    .X(_02167_));
 sg13g2_nor2_1 _07682_ (.A(_02037_),
    .B(_02167_),
    .Y(_02168_));
 sg13g2_a21oi_1 _07683_ (.A1(_02037_),
    .A2(_02157_),
    .Y(_02169_),
    .B1(_02091_));
 sg13g2_a21oi_1 _07684_ (.A1(_02037_),
    .A2(_02157_),
    .Y(_02170_),
    .B1(_02168_));
 sg13g2_nand2_1 _07685_ (.Y(_02171_),
    .A(net1502),
    .B(_02170_));
 sg13g2_and2_1 _07686_ (.A(_02087_),
    .B(_02171_),
    .X(_02172_));
 sg13g2_a22oi_1 _07687_ (.Y(_02173_),
    .B1(_02165_),
    .B2(_02172_),
    .A2(_02156_),
    .A1(_02135_));
 sg13g2_xor2_1 _07688_ (.B(_02118_),
    .A(_02117_),
    .X(_02174_));
 sg13g2_nor2_1 _07689_ (.A(_02173_),
    .B(_02174_),
    .Y(_02175_));
 sg13g2_nor2_1 _07690_ (.A(_02078_),
    .B(_02093_),
    .Y(_02176_));
 sg13g2_xnor2_1 _07691_ (.Y(_02177_),
    .A(_02094_),
    .B(_02176_));
 sg13g2_nand2_1 _07692_ (.Y(_02178_),
    .A(net1747),
    .B(_02177_));
 sg13g2_o21ai_1 _07693_ (.B1(_02178_),
    .Y(_02179_),
    .A1(net1747),
    .A2(_02167_));
 sg13g2_mux2_1 _07694_ (.A0(_02158_),
    .A1(_02179_),
    .S(net1502),
    .X(_02180_));
 sg13g2_a22oi_1 _07695_ (.Y(_02181_),
    .B1(_02180_),
    .B2(_02087_),
    .A2(_02156_),
    .A1(_02142_));
 sg13g2_xnor2_1 _07696_ (.Y(_02182_),
    .A(_02115_),
    .B(_02116_));
 sg13g2_nor2b_1 _07697_ (.A(_02181_),
    .B_N(_02182_),
    .Y(_02183_));
 sg13g2_o21ai_1 _07698_ (.B1(_02090_),
    .Y(_02184_),
    .A1(_02037_),
    .A2(_02093_));
 sg13g2_a21oi_1 _07699_ (.A1(_02037_),
    .A2(_02177_),
    .Y(_02185_),
    .B1(_02184_));
 sg13g2_a21oi_1 _07700_ (.A1(_02091_),
    .A2(_02170_),
    .Y(_02186_),
    .B1(_02185_));
 sg13g2_a22oi_1 _07701_ (.Y(_02187_),
    .B1(_02186_),
    .B2(_02087_),
    .A2(_02156_),
    .A1(_02150_));
 sg13g2_nor2_1 _07702_ (.A(_02114_),
    .B(_02187_),
    .Y(_02188_));
 sg13g2_xnor2_1 _07703_ (.Y(_02189_),
    .A(_02181_),
    .B(_02182_));
 sg13g2_a21o_1 _07704_ (.A2(_02189_),
    .A1(_02188_),
    .B1(_02183_),
    .X(_02190_));
 sg13g2_xor2_1 _07705_ (.B(_02174_),
    .A(_02173_),
    .X(_02191_));
 sg13g2_a21oi_1 _07706_ (.A1(_02190_),
    .A2(_02191_),
    .Y(_02192_),
    .B1(_02175_));
 sg13g2_o21ai_1 _07707_ (.B1(_02163_),
    .Y(_02193_),
    .A1(_02164_),
    .A2(_02192_));
 sg13g2_a21oi_1 _07708_ (.A1(_02155_),
    .A2(_02193_),
    .Y(_02194_),
    .B1(_02153_));
 sg13g2_o21ai_1 _07709_ (.B1(_02145_),
    .Y(_02195_),
    .A1(_02146_),
    .A2(_02194_));
 sg13g2_xnor2_1 _07710_ (.Y(_02196_),
    .A(_02136_),
    .B(_02137_));
 sg13g2_a21oi_1 _07711_ (.A1(_02195_),
    .A2(_02196_),
    .Y(_02197_),
    .B1(_02138_));
 sg13g2_xor2_1 _07712_ (.B(_02130_),
    .A(_02113_),
    .X(_02198_));
 sg13g2_inv_1 _07713_ (.Y(_02199_),
    .A(_02198_));
 sg13g2_o21ai_1 _07714_ (.B1(_02131_),
    .Y(_02200_),
    .A1(_02197_),
    .A2(_02199_));
 sg13g2_a21oi_2 _07715_ (.B1(_02082_),
    .Y(_02201_),
    .A2(_02200_),
    .A1(_02083_));
 sg13g2_nor2_1 _07716_ (.A(_02148_),
    .B(_02157_),
    .Y(_02202_));
 sg13g2_a21oi_1 _07717_ (.A1(_02147_),
    .A2(_02202_),
    .Y(_02203_),
    .B1(_02169_));
 sg13g2_o21ai_1 _07718_ (.B1(_02093_),
    .Y(_02204_),
    .A1(net1747),
    .A2(_02094_));
 sg13g2_a21oi_1 _07719_ (.A1(_02091_),
    .A2(_02204_),
    .Y(_02205_),
    .B1(_02085_));
 sg13g2_nor2b_1 _07720_ (.A(_02205_),
    .B_N(_02076_),
    .Y(_02206_));
 sg13g2_o21ai_1 _07721_ (.B1(_02206_),
    .Y(_02207_),
    .A1(_02096_),
    .A2(_02203_));
 sg13g2_inv_1 _07722_ (.Y(_02208_),
    .A(_02207_));
 sg13g2_xnor2_1 _07723_ (.Y(_02209_),
    .A(_02114_),
    .B(_02187_));
 sg13g2_o21ai_1 _07724_ (.B1(_02090_),
    .Y(_02210_),
    .A1(net1747),
    .A2(_02093_));
 sg13g2_nor2_1 _07725_ (.A(net1502),
    .B(_02179_),
    .Y(_02211_));
 sg13g2_nor2_1 _07726_ (.A(_02088_),
    .B(_02211_),
    .Y(_02212_));
 sg13g2_a22oi_1 _07727_ (.Y(_02213_),
    .B1(_02210_),
    .B2(_02212_),
    .A2(_02160_),
    .A1(_02156_));
 sg13g2_inv_1 _07728_ (.Y(_02214_),
    .A(_02213_));
 sg13g2_nand2_1 _07729_ (.Y(_02215_),
    .A(_02209_),
    .B(_02213_));
 sg13g2_inv_1 _07730_ (.Y(_02216_),
    .A(_02215_));
 sg13g2_xor2_1 _07731_ (.B(_02189_),
    .A(_02188_),
    .X(_02217_));
 sg13g2_nor2_1 _07732_ (.A(_02215_),
    .B(_02217_),
    .Y(_02218_));
 sg13g2_xnor2_1 _07733_ (.Y(_02219_),
    .A(_02190_),
    .B(_02191_));
 sg13g2_and2_1 _07734_ (.A(_02218_),
    .B(_02219_),
    .X(_02220_));
 sg13g2_xnor2_1 _07735_ (.Y(_02221_),
    .A(_02164_),
    .B(_02192_));
 sg13g2_and2_1 _07736_ (.A(_02220_),
    .B(_02221_),
    .X(_02222_));
 sg13g2_xnor2_1 _07737_ (.Y(_02223_),
    .A(_02155_),
    .B(_02193_));
 sg13g2_and2_1 _07738_ (.A(_02222_),
    .B(_02223_),
    .X(_02224_));
 sg13g2_xnor2_1 _07739_ (.Y(_02225_),
    .A(_02146_),
    .B(_02194_));
 sg13g2_and2_1 _07740_ (.A(_02224_),
    .B(_02225_),
    .X(_02226_));
 sg13g2_xnor2_1 _07741_ (.Y(_02227_),
    .A(_02195_),
    .B(_02196_));
 sg13g2_nand2_1 _07742_ (.Y(_02228_),
    .A(_02226_),
    .B(_02227_));
 sg13g2_xnor2_1 _07743_ (.Y(_02229_),
    .A(_02197_),
    .B(_02199_));
 sg13g2_nand3_1 _07744_ (.B(_02227_),
    .C(_02229_),
    .A(_02226_),
    .Y(_02230_));
 sg13g2_o21ai_1 _07745_ (.B1(_02201_),
    .Y(_02231_),
    .A1(_02208_),
    .A2(_02230_));
 sg13g2_xnor2_1 _07746_ (.Y(_02232_),
    .A(net1475),
    .B(net1470));
 sg13g2_xor2_1 _07747_ (.B(_02232_),
    .A(_02231_),
    .X(_02233_));
 sg13g2_nand3b_1 _07748_ (.B(_02042_),
    .C(net1527),
    .Y(_02234_),
    .A_N(_02026_));
 sg13g2_nand2_1 _07749_ (.Y(_02235_),
    .A(_02064_),
    .B(_02073_));
 sg13g2_nand2_1 _07750_ (.Y(_02236_),
    .A(_02051_),
    .B(_02056_));
 sg13g2_nor4_1 _07751_ (.A(_02063_),
    .B(_02234_),
    .C(_02235_),
    .D(_02236_),
    .Y(_02237_));
 sg13g2_nand2_1 _07752_ (.Y(_02238_),
    .A(net1445),
    .B(_02237_));
 sg13g2_nor4_1 _07753_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][6] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][15] ),
    .C(_01977_),
    .D(_01984_),
    .Y(_02239_));
 sg13g2_nand2b_1 _07754_ (.Y(_02240_),
    .B(_02232_),
    .A_N(_02230_));
 sg13g2_nand2b_1 _07755_ (.Y(_02241_),
    .B(_02240_),
    .A_N(net1721));
 sg13g2_a221oi_1 _07756_ (.B2(_02226_),
    .C1(_02082_),
    .B1(_02207_),
    .A1(net1475),
    .Y(_02242_),
    .A2(net1470));
 sg13g2_xnor2_1 _07757_ (.Y(_02243_),
    .A(_02227_),
    .B(_02242_));
 sg13g2_a221oi_1 _07758_ (.B2(_02224_),
    .C1(_02082_),
    .B1(_02207_),
    .A1(net1475),
    .Y(_02244_),
    .A2(net1470));
 sg13g2_xor2_1 _07759_ (.B(_02244_),
    .A(_02225_),
    .X(_02245_));
 sg13g2_nor2_2 _07760_ (.A(net1458),
    .B(net1457),
    .Y(_02246_));
 sg13g2_a221oi_1 _07761_ (.B2(_02222_),
    .C1(_02082_),
    .B1(_02207_),
    .A1(net1475),
    .Y(_02247_),
    .A2(net1470));
 sg13g2_xor2_1 _07762_ (.B(_02247_),
    .A(_02223_),
    .X(_02248_));
 sg13g2_a221oi_1 _07763_ (.B2(_02213_),
    .C1(_02082_),
    .B1(_02207_),
    .A1(net1475),
    .Y(_02249_),
    .A2(net1470));
 sg13g2_xnor2_1 _07764_ (.Y(_02250_),
    .A(_02209_),
    .B(_02249_));
 sg13g2_xor2_1 _07765_ (.B(_02249_),
    .A(_02209_),
    .X(_02251_));
 sg13g2_and2_1 _07766_ (.A(net1456),
    .B(_02251_),
    .X(_02252_));
 sg13g2_a221oi_1 _07767_ (.B2(_02218_),
    .C1(_02082_),
    .B1(_02207_),
    .A1(net1475),
    .Y(_02253_),
    .A2(net1470));
 sg13g2_xor2_1 _07768_ (.B(_02253_),
    .A(_02219_),
    .X(_02254_));
 sg13g2_xnor2_1 _07769_ (.Y(_02255_),
    .A(_02219_),
    .B(_02253_));
 sg13g2_a21oi_2 _07770_ (.B1(_02214_),
    .Y(_02256_),
    .A2(_02208_),
    .A1(_02201_));
 sg13g2_and3_1 _07771_ (.X(_02257_),
    .A(_02201_),
    .B(_02208_),
    .C(_02214_));
 sg13g2_nor2_2 _07772_ (.A(_02256_),
    .B(_02257_),
    .Y(_02258_));
 sg13g2_nor3_1 _07773_ (.A(_02255_),
    .B(_02256_),
    .C(_02257_),
    .Y(_02259_));
 sg13g2_nand2_1 _07774_ (.Y(_02260_),
    .A(_02254_),
    .B(_02258_));
 sg13g2_a221oi_1 _07775_ (.B2(_02220_),
    .C1(_02082_),
    .B1(_02207_),
    .A1(net1475),
    .Y(_02261_),
    .A2(net1470));
 sg13g2_xor2_1 _07776_ (.B(_02261_),
    .A(_02221_),
    .X(_02262_));
 sg13g2_nor2b_2 _07777_ (.A(_02262_),
    .B_N(net1456),
    .Y(_02263_));
 sg13g2_a221oi_1 _07778_ (.B2(_02216_),
    .C1(_02082_),
    .B1(_02207_),
    .A1(net1475),
    .Y(_02264_),
    .A2(net1470));
 sg13g2_xnor2_1 _07779_ (.Y(_02265_),
    .A(_02217_),
    .B(_02264_));
 sg13g2_nor2b_1 _07780_ (.A(_02265_),
    .B_N(net1455),
    .Y(_02266_));
 sg13g2_inv_1 _07781_ (.Y(_02267_),
    .A(_02266_));
 sg13g2_a221oi_1 _07782_ (.B2(_02254_),
    .C1(_02263_),
    .B1(_02266_),
    .A1(_02252_),
    .Y(_02268_),
    .A2(_02259_));
 sg13g2_a21oi_2 _07783_ (.B1(net1459),
    .Y(_02269_),
    .A2(_02268_),
    .A1(net1457));
 sg13g2_o21ai_1 _07784_ (.B1(_02251_),
    .Y(_02270_),
    .A1(_02256_),
    .A2(_02257_));
 sg13g2_and2_1 _07785_ (.A(_02254_),
    .B(_02265_),
    .X(_02271_));
 sg13g2_nand2b_1 _07786_ (.Y(_02272_),
    .B(_02271_),
    .A_N(_02270_));
 sg13g2_nand2_1 _07787_ (.Y(_02273_),
    .A(net1455),
    .B(_02262_));
 sg13g2_nor2b_1 _07788_ (.A(net1458),
    .B_N(net1457),
    .Y(_02274_));
 sg13g2_nand2b_2 _07789_ (.Y(_02275_),
    .B(net1457),
    .A_N(net1458));
 sg13g2_nor2_1 _07790_ (.A(_02273_),
    .B(_02275_),
    .Y(_02276_));
 sg13g2_and3_1 _07791_ (.X(_02277_),
    .A(_02052_),
    .B(_02272_),
    .C(_02276_));
 sg13g2_nand3_1 _07792_ (.B(_02272_),
    .C(_02276_),
    .A(_02052_),
    .Y(_02278_));
 sg13g2_a21oi_1 _07793_ (.A1(_02270_),
    .A2(_02271_),
    .Y(_02279_),
    .B1(_02273_));
 sg13g2_a21o_1 _07794_ (.A2(_02271_),
    .A1(_02270_),
    .B1(_02273_),
    .X(_02280_));
 sg13g2_nor3_1 _07795_ (.A(net1527),
    .B(_02275_),
    .C(_02279_),
    .Y(_02281_));
 sg13g2_or4_1 _07796_ (.A(net1527),
    .B(_02268_),
    .C(_02275_),
    .D(_02279_),
    .X(_02282_));
 sg13g2_a221oi_1 _07797_ (.B2(_02056_),
    .C1(_02282_),
    .B1(_02278_),
    .A1(_02043_),
    .Y(_02283_),
    .A2(_02269_));
 sg13g2_nand2_1 _07798_ (.Y(_02284_),
    .A(_02043_),
    .B(net1527));
 sg13g2_a221oi_1 _07799_ (.B2(_02268_),
    .C1(net1458),
    .B1(net1457),
    .A1(_02043_),
    .Y(_02285_),
    .A2(net1527));
 sg13g2_a21oi_2 _07800_ (.B1(_02048_),
    .Y(_02286_),
    .A2(_02280_),
    .A1(_02274_));
 sg13g2_o21ai_1 _07801_ (.B1(net1527),
    .Y(_02287_),
    .A1(_02275_),
    .A2(_02279_));
 sg13g2_or3_1 _07802_ (.A(_02277_),
    .B(_02285_),
    .C(_02287_),
    .X(_02288_));
 sg13g2_a21o_1 _07803_ (.A2(_02276_),
    .A1(_02272_),
    .B1(_02052_),
    .X(_02289_));
 sg13g2_and2_1 _07804_ (.A(_02057_),
    .B(_02289_),
    .X(_02290_));
 sg13g2_a21o_1 _07805_ (.A2(_02290_),
    .A1(_02288_),
    .B1(_02283_),
    .X(_02291_));
 sg13g2_o21ai_1 _07806_ (.B1(_02201_),
    .Y(_02292_),
    .A1(_02208_),
    .A2(_02228_));
 sg13g2_xnor2_1 _07807_ (.Y(_02293_),
    .A(_02229_),
    .B(_02292_));
 sg13g2_inv_2 _07808_ (.Y(_02294_),
    .A(net1444));
 sg13g2_nor4_1 _07809_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][14] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][14] ),
    .C(_02073_),
    .D(net1446),
    .Y(_02295_));
 sg13g2_and3_1 _07810_ (.X(_02296_),
    .A(_02065_),
    .B(net1444),
    .C(_02295_));
 sg13g2_nand2_1 _07811_ (.Y(_02297_),
    .A(_02291_),
    .B(_02296_));
 sg13g2_a21o_1 _07812_ (.A2(_02296_),
    .A1(_02291_),
    .B1(_02241_),
    .X(_02298_));
 sg13g2_nor2b_2 _07813_ (.A(net1422),
    .B_N(_02238_),
    .Y(_02299_));
 sg13g2_and2_1 _07814_ (.A(net1458),
    .B(net1443),
    .X(_02300_));
 sg13g2_nand2_1 _07815_ (.Y(_02301_),
    .A(_02258_),
    .B(_02300_));
 sg13g2_a21oi_1 _07816_ (.A1(_02250_),
    .A2(_02294_),
    .Y(_02302_),
    .B1(net1448));
 sg13g2_a22oi_1 _07817_ (.Y(_02303_),
    .B1(_02301_),
    .B2(_02302_),
    .A2(_02265_),
    .A1(net1448));
 sg13g2_nor4_1 _07818_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][6] ),
    .B(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][15] ),
    .C(_01988_),
    .D(_01995_),
    .Y(_02304_));
 sg13g2_nor2_1 _07819_ (.A(_02000_),
    .B(_02304_),
    .Y(_02305_));
 sg13g2_or2_2 _07820_ (.X(_02306_),
    .B(_02304_),
    .A(_02000_));
 sg13g2_a22oi_1 _07821_ (.Y(_02307_),
    .B1(_02299_),
    .B2(_02303_),
    .A2(net1719),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][0] ));
 sg13g2_o21ai_1 _07822_ (.B1(_02003_),
    .Y(_02308_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][0] ),
    .A2(net1665));
 sg13g2_a21oi_1 _07823_ (.A1(net1666),
    .A2(_02307_),
    .Y(_02309_),
    .B1(_02308_));
 sg13g2_nor2_2 _07824_ (.A(_02007_),
    .B(_02309_),
    .Y(_02310_));
 sg13g2_nor2b_1 _07825_ (.A(_00166_),
    .B_N(\u_tiny_nn_top.state_q[10] ),
    .Y(_02311_));
 sg13g2_a21oi_1 _07826_ (.A1(_00786_),
    .A2(_02311_),
    .Y(_02312_),
    .B1(\u_tiny_nn_top.state_q[6] ));
 sg13g2_a21oi_2 _07827_ (.B1(_00774_),
    .Y(_02313_),
    .A2(_02312_),
    .A1(net1768));
 sg13g2_nor2_1 _07828_ (.A(_01187_),
    .B(_02313_),
    .Y(_02314_));
 sg13g2_a21o_1 _07829_ (.A2(_02297_),
    .A1(_02201_),
    .B1(net1721),
    .X(_02315_));
 sg13g2_a21oi_1 _07830_ (.A1(_00673_),
    .A2(net1719),
    .Y(_02316_),
    .B1(_02306_));
 sg13g2_a22oi_1 _07831_ (.Y(_02317_),
    .B1(_02315_),
    .B2(_02316_),
    .A2(_02306_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][15] ));
 sg13g2_o21ai_1 _07832_ (.B1(_02004_),
    .Y(_02318_),
    .A1(_02002_),
    .A2(_02317_));
 sg13g2_a21o_2 _07833_ (.A2(_02318_),
    .A1(_02313_),
    .B1(_01187_),
    .X(_02319_));
 sg13g2_a21oi_1 _07834_ (.A1(_02313_),
    .A2(_02318_),
    .Y(_02320_),
    .B1(_01187_));
 sg13g2_nor2_1 _07835_ (.A(_02310_),
    .B(_02319_),
    .Y(_02321_));
 sg13g2_nor2_1 _07836_ (.A(net1507),
    .B(_02321_),
    .Y(_02322_));
 sg13g2_a22oi_1 _07837_ (.Y(_00215_),
    .B1(_01974_),
    .B2(_02322_),
    .A2(net1507),
    .A1(_00705_));
 sg13g2_a21oi_1 _07838_ (.A1(_01546_),
    .A2(_01607_),
    .Y(_02323_),
    .B1(net1423));
 sg13g2_nand2_1 _07839_ (.Y(_02324_),
    .A(_01538_),
    .B(net1431));
 sg13g2_o21ai_1 _07840_ (.B1(_02324_),
    .Y(_02325_),
    .A1(_01541_),
    .A2(net1431));
 sg13g2_nand3b_1 _07841_ (.B(net1427),
    .C(_02325_),
    .Y(_02326_),
    .A_N(_01562_));
 sg13g2_a22oi_1 _07842_ (.Y(_02327_),
    .B1(_02323_),
    .B2(_02326_),
    .A2(net1424),
    .A1(net1434));
 sg13g2_a221oi_1 _07843_ (.B2(_02327_),
    .C1(net1486),
    .B1(_01615_),
    .A1(_01220_),
    .Y(_02328_),
    .A2(net1669));
 sg13g2_o21ai_1 _07844_ (.B1(net1500),
    .Y(_02329_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[1] ),
    .A2(net1487));
 sg13g2_o21ai_1 _07845_ (.B1(_01269_),
    .Y(_02330_),
    .A1(_02328_),
    .A2(_02329_));
 sg13g2_nand2_1 _07846_ (.Y(_02331_),
    .A(_01909_),
    .B(_01946_));
 sg13g2_nand2_1 _07847_ (.Y(_02332_),
    .A(_01905_),
    .B(_01929_));
 sg13g2_o21ai_1 _07848_ (.B1(_02332_),
    .Y(_02333_),
    .A1(_01906_),
    .A2(_01919_));
 sg13g2_a21oi_1 _07849_ (.A1(net1460),
    .A2(_02333_),
    .Y(_02334_),
    .B1(net1449));
 sg13g2_a22oi_1 _07850_ (.Y(_02335_),
    .B1(_02331_),
    .B2(_02334_),
    .A2(_01913_),
    .A1(net1450));
 sg13g2_a221oi_1 _07851_ (.B2(_02335_),
    .C1(net1545),
    .B1(_01962_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][1] ),
    .Y(_02336_),
    .A2(net1723));
 sg13g2_o21ai_1 _07852_ (.B1(net1668),
    .Y(_02337_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][1] ),
    .A2(net1548));
 sg13g2_nor2_1 _07853_ (.A(_02336_),
    .B(_02337_),
    .Y(_02338_));
 sg13g2_nor2_1 _07854_ (.A(_01654_),
    .B(_02338_),
    .Y(_02339_));
 sg13g2_nor2_1 _07855_ (.A(net1674),
    .B(_02339_),
    .Y(_02340_));
 sg13g2_o21ai_1 _07856_ (.B1(_02340_),
    .Y(_02341_),
    .A1(net1530),
    .A2(_02330_));
 sg13g2_nor2_1 _07857_ (.A(net1459),
    .B(_02294_),
    .Y(_02342_));
 sg13g2_nand3_1 _07858_ (.B(_02258_),
    .C(net1443),
    .A(_02246_),
    .Y(_02343_));
 sg13g2_nor2_1 _07859_ (.A(_02265_),
    .B(net1443),
    .Y(_02344_));
 sg13g2_a21oi_1 _07860_ (.A1(_02250_),
    .A2(_02300_),
    .Y(_02345_),
    .B1(_02344_));
 sg13g2_nor2b_1 _07861_ (.A(net1447),
    .B_N(_02345_),
    .Y(_02346_));
 sg13g2_a22oi_1 _07862_ (.Y(_02347_),
    .B1(_02343_),
    .B2(_02346_),
    .A2(_02254_),
    .A1(net1448));
 sg13g2_a22oi_1 _07863_ (.Y(_02348_),
    .B1(_02299_),
    .B2(_02347_),
    .A2(net1719),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][1] ));
 sg13g2_o21ai_1 _07864_ (.B1(_02003_),
    .Y(_02349_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][1] ),
    .A2(net1664));
 sg13g2_a21oi_1 _07865_ (.A1(net1664),
    .A2(_02348_),
    .Y(_02350_),
    .B1(_02349_));
 sg13g2_nor2_2 _07866_ (.A(net1528),
    .B(_02350_),
    .Y(_02351_));
 sg13g2_nor2_1 _07867_ (.A(_02319_),
    .B(_02351_),
    .Y(_02352_));
 sg13g2_nor2_1 _07868_ (.A(net1507),
    .B(_02352_),
    .Y(_02353_));
 sg13g2_a22oi_1 _07869_ (.Y(_00216_),
    .B1(_02341_),
    .B2(_02353_),
    .A2(net1509),
    .A1(_00707_));
 sg13g2_a21oi_1 _07870_ (.A1(_01542_),
    .A2(net1430),
    .Y(_02354_),
    .B1(net1432));
 sg13g2_a21oi_1 _07871_ (.A1(_01539_),
    .A2(net1432),
    .Y(_02355_),
    .B1(_02354_));
 sg13g2_o21ai_1 _07872_ (.B1(net1427),
    .Y(_02356_),
    .A1(_01545_),
    .A2(net1429));
 sg13g2_a21oi_1 _07873_ (.A1(net1429),
    .A2(_02355_),
    .Y(_02357_),
    .B1(_02356_));
 sg13g2_a21o_1 _07874_ (.A2(_01607_),
    .A1(_01549_),
    .B1(_02357_),
    .X(_02358_));
 sg13g2_nand2_1 _07875_ (.Y(_02359_),
    .A(_01567_),
    .B(net1423));
 sg13g2_o21ai_1 _07876_ (.B1(_02359_),
    .Y(_02360_),
    .A1(_01596_),
    .A2(_02358_));
 sg13g2_a221oi_1 _07877_ (.B2(_02360_),
    .C1(net1486),
    .B1(_01615_),
    .A1(_01223_),
    .Y(_02361_),
    .A2(net1669));
 sg13g2_o21ai_1 _07878_ (.B1(net1500),
    .Y(_02362_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[2] ),
    .A2(net1487));
 sg13g2_o21ai_1 _07879_ (.B1(_01269_),
    .Y(_02363_),
    .A1(_02361_),
    .A2(_02362_));
 sg13g2_nand2_1 _07880_ (.Y(_02364_),
    .A(_01907_),
    .B(_01929_));
 sg13g2_nand2_1 _07881_ (.Y(_02365_),
    .A(_01909_),
    .B(net1462));
 sg13g2_nand3_1 _07882_ (.B(_01920_),
    .C(_01924_),
    .A(_01905_),
    .Y(_02366_));
 sg13g2_nand4_1 _07883_ (.B(_02364_),
    .C(_02365_),
    .A(net1460),
    .Y(_02367_),
    .D(_02366_));
 sg13g2_nand2_1 _07884_ (.Y(_02368_),
    .A(_01913_),
    .B(_01946_));
 sg13g2_nand3_1 _07885_ (.B(_02367_),
    .C(_02368_),
    .A(net1452),
    .Y(_02369_));
 sg13g2_o21ai_1 _07886_ (.B1(_02369_),
    .Y(_02370_),
    .A1(net1452),
    .A2(net1469));
 sg13g2_a221oi_1 _07887_ (.B2(_02370_),
    .C1(net1547),
    .B1(_01962_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][2] ),
    .Y(_02371_),
    .A2(net1723));
 sg13g2_a21oi_1 _07888_ (.A1(_00765_),
    .A2(_01968_),
    .Y(_02372_),
    .B1(_02371_));
 sg13g2_a21oi_1 _07889_ (.A1(_01648_),
    .A2(_02372_),
    .Y(_02373_),
    .B1(_01654_));
 sg13g2_nor2_1 _07890_ (.A(net1674),
    .B(_02373_),
    .Y(_02374_));
 sg13g2_o21ai_1 _07891_ (.B1(_02374_),
    .Y(_02375_),
    .A1(net1531),
    .A2(_02363_));
 sg13g2_nor3_1 _07892_ (.A(net1455),
    .B(_02256_),
    .C(_02257_),
    .Y(_02376_));
 sg13g2_a221oi_1 _07893_ (.B2(net1458),
    .C1(_02294_),
    .B1(_02265_),
    .A1(_02246_),
    .Y(_02377_),
    .A2(_02251_));
 sg13g2_o21ai_1 _07894_ (.B1(_02377_),
    .Y(_02378_),
    .A1(_02275_),
    .A2(_02376_));
 sg13g2_a21oi_1 _07895_ (.A1(_02255_),
    .A2(_02294_),
    .Y(_02379_),
    .B1(net1447));
 sg13g2_a22oi_1 _07896_ (.Y(_02380_),
    .B1(_02378_),
    .B2(_02379_),
    .A2(_02262_),
    .A1(net1447));
 sg13g2_a221oi_1 _07897_ (.B2(_02380_),
    .C1(_02306_),
    .B1(_02299_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][2] ),
    .Y(_02381_),
    .A2(net1719));
 sg13g2_o21ai_1 _07898_ (.B1(_02003_),
    .Y(_02382_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][2] ),
    .A2(net1664));
 sg13g2_nor2_1 _07899_ (.A(_02381_),
    .B(_02382_),
    .Y(_02383_));
 sg13g2_nor2_2 _07900_ (.A(net1528),
    .B(_02383_),
    .Y(_02384_));
 sg13g2_inv_1 _07901_ (.Y(_02385_),
    .A(_02384_));
 sg13g2_a21oi_1 _07902_ (.A1(net1418),
    .A2(_02385_),
    .Y(_02386_),
    .B1(net1510));
 sg13g2_a22oi_1 _07903_ (.Y(_00217_),
    .B1(_02375_),
    .B2(_02386_),
    .A2(net1510),
    .A1(_00710_));
 sg13g2_nor2_1 _07904_ (.A(net1433),
    .B(_01568_),
    .Y(_02387_));
 sg13g2_nand2_1 _07905_ (.Y(_02388_),
    .A(_01538_),
    .B(net1430));
 sg13g2_o21ai_1 _07906_ (.B1(_02388_),
    .Y(_02389_),
    .A1(_01541_),
    .A2(net1430));
 sg13g2_nand2_1 _07907_ (.Y(_02390_),
    .A(_02387_),
    .B(_02389_));
 sg13g2_nand2_1 _07908_ (.Y(_02391_),
    .A(_01546_),
    .B(net1432));
 sg13g2_nand4_1 _07909_ (.B(net1427),
    .C(_02390_),
    .A(net1429),
    .Y(_02392_),
    .D(_02391_));
 sg13g2_a221oi_1 _07910_ (.B2(net1434),
    .C1(net1424),
    .B1(_01616_),
    .A1(_01566_),
    .Y(_02393_),
    .A2(_01607_));
 sg13g2_a22oi_1 _07911_ (.Y(_02394_),
    .B1(_02392_),
    .B2(_02393_),
    .A2(net1424),
    .A1(_01563_));
 sg13g2_nor2b_1 _07912_ (.A(_02394_),
    .B_N(_01615_),
    .Y(_02395_));
 sg13g2_o21ai_1 _07913_ (.B1(net1487),
    .Y(_02396_),
    .A1(_01217_),
    .A2(_01271_));
 sg13g2_nor2_1 _07914_ (.A(_02395_),
    .B(_02396_),
    .Y(_02397_));
 sg13g2_o21ai_1 _07915_ (.B1(net1500),
    .Y(_02398_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[3] ),
    .A2(net1487));
 sg13g2_o21ai_1 _07916_ (.B1(_01269_),
    .Y(_02399_),
    .A1(_02397_),
    .A2(_02398_));
 sg13g2_nand3_1 _07917_ (.B(_01920_),
    .C(_01925_),
    .A(_01905_),
    .Y(_02400_));
 sg13g2_a22oi_1 _07918_ (.Y(_02401_),
    .B1(_01947_),
    .B2(_02400_),
    .A2(net1469),
    .A1(net1452));
 sg13g2_nand2_1 _07919_ (.Y(_02402_),
    .A(_01907_),
    .B(_01924_));
 sg13g2_o21ai_1 _07920_ (.B1(net1460),
    .Y(_02403_),
    .A1(_01912_),
    .A2(_01919_));
 sg13g2_a221oi_1 _07921_ (.B2(_01920_),
    .C1(_02403_),
    .B1(_02402_),
    .A1(_01910_),
    .Y(_02404_),
    .A2(_01929_));
 sg13g2_nor2_1 _07922_ (.A(_02401_),
    .B(_02404_),
    .Y(_02405_));
 sg13g2_a21oi_1 _07923_ (.A1(net1449),
    .A2(_01925_),
    .Y(_02406_),
    .B1(_02405_));
 sg13g2_a221oi_1 _07924_ (.B2(_02406_),
    .C1(net1547),
    .B1(_01962_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][3] ),
    .Y(_02407_),
    .A2(net1723));
 sg13g2_a21oi_1 _07925_ (.A1(_00764_),
    .A2(net1545),
    .Y(_02408_),
    .B1(_02407_));
 sg13g2_a21oi_1 _07926_ (.A1(net1668),
    .A2(_02408_),
    .Y(_02409_),
    .B1(_01654_));
 sg13g2_nor2_1 _07927_ (.A(net1674),
    .B(_02409_),
    .Y(_02410_));
 sg13g2_o21ai_1 _07928_ (.B1(_02410_),
    .Y(_02411_),
    .A1(net1530),
    .A2(_02399_));
 sg13g2_nor2_1 _07929_ (.A(_02262_),
    .B(net1443),
    .Y(_02412_));
 sg13g2_nor2_1 _07930_ (.A(net1447),
    .B(_02412_),
    .Y(_02413_));
 sg13g2_a21oi_1 _07931_ (.A1(_02258_),
    .A2(_02263_),
    .Y(_02414_),
    .B1(_02275_));
 sg13g2_o21ai_1 _07932_ (.B1(_02414_),
    .Y(_02415_),
    .A1(net1455),
    .A2(_02251_));
 sg13g2_a22oi_1 _07933_ (.Y(_02416_),
    .B1(_02265_),
    .B2(_02246_),
    .A2(_02254_),
    .A1(net1458));
 sg13g2_nand3_1 _07934_ (.B(_02415_),
    .C(_02416_),
    .A(net1443),
    .Y(_02417_));
 sg13g2_a22oi_1 _07935_ (.Y(_02418_),
    .B1(_02413_),
    .B2(_02417_),
    .A2(net1455),
    .A1(net1447));
 sg13g2_a22oi_1 _07936_ (.Y(_02419_),
    .B1(_02299_),
    .B2(_02418_),
    .A2(net1720),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][3] ));
 sg13g2_o21ai_1 _07937_ (.B1(_02003_),
    .Y(_02420_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][3] ),
    .A2(net1664));
 sg13g2_a21oi_1 _07938_ (.A1(net1664),
    .A2(_02419_),
    .Y(_02421_),
    .B1(_02420_));
 sg13g2_nor2_2 _07939_ (.A(net1528),
    .B(_02421_),
    .Y(_02422_));
 sg13g2_nor2_1 _07940_ (.A(_02319_),
    .B(_02422_),
    .Y(_02423_));
 sg13g2_nor2_1 _07941_ (.A(net1508),
    .B(_02423_),
    .Y(_02424_));
 sg13g2_a22oi_1 _07942_ (.Y(_00218_),
    .B1(_02411_),
    .B2(_02424_),
    .A2(net1508),
    .A1(_00712_));
 sg13g2_nand2_1 _07943_ (.Y(_02425_),
    .A(net1433),
    .B(net1423));
 sg13g2_nor2_1 _07944_ (.A(_01542_),
    .B(net1432),
    .Y(_02426_));
 sg13g2_nor3_1 _07945_ (.A(net1434),
    .B(_02387_),
    .C(_02426_),
    .Y(_02427_));
 sg13g2_o21ai_1 _07946_ (.B1(_02387_),
    .Y(_02428_),
    .A1(_01538_),
    .A2(net1430));
 sg13g2_a21oi_1 _07947_ (.A1(_01545_),
    .A2(net1430),
    .Y(_02429_),
    .B1(_02428_));
 sg13g2_o21ai_1 _07948_ (.B1(_01597_),
    .Y(_02430_),
    .A1(_01563_),
    .A2(net1427));
 sg13g2_or2_1 _07949_ (.X(_02431_),
    .B(_02429_),
    .A(_02427_));
 sg13g2_o21ai_1 _07950_ (.B1(net1427),
    .Y(_02432_),
    .A1(net1429),
    .A2(_01566_));
 sg13g2_a21oi_1 _07951_ (.A1(net1429),
    .A2(_02431_),
    .Y(_02433_),
    .B1(_02432_));
 sg13g2_o21ai_1 _07952_ (.B1(_02425_),
    .Y(_02434_),
    .A1(_02430_),
    .A2(_02433_));
 sg13g2_o21ai_1 _07953_ (.B1(net1487),
    .Y(_02435_),
    .A1(_01214_),
    .A2(_01271_));
 sg13g2_a21oi_1 _07954_ (.A1(_01615_),
    .A2(_02434_),
    .Y(_02436_),
    .B1(_02435_));
 sg13g2_o21ai_1 _07955_ (.B1(net1500),
    .Y(_02437_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[4] ),
    .A2(net1487));
 sg13g2_o21ai_1 _07956_ (.B1(_01269_),
    .Y(_02438_),
    .A1(_02436_),
    .A2(_02437_));
 sg13g2_nor3_1 _07957_ (.A(_01906_),
    .B(_01916_),
    .C(_01924_),
    .Y(_02439_));
 sg13g2_nor2_1 _07958_ (.A(_01918_),
    .B(_02439_),
    .Y(_02440_));
 sg13g2_nor2b_1 _07959_ (.A(_01926_),
    .B_N(_01905_),
    .Y(_02441_));
 sg13g2_nor2_1 _07960_ (.A(_01913_),
    .B(_01918_),
    .Y(_02442_));
 sg13g2_o21ai_1 _07961_ (.B1(_02442_),
    .Y(_02443_),
    .A1(_01916_),
    .A2(_02441_));
 sg13g2_o21ai_1 _07962_ (.B1(_02443_),
    .Y(_02444_),
    .A1(net1469),
    .A2(_02440_));
 sg13g2_o21ai_1 _07963_ (.B1(net1461),
    .Y(_02445_),
    .A1(_01910_),
    .A2(_01921_));
 sg13g2_a221oi_1 _07964_ (.B2(_01924_),
    .C1(net1449),
    .B1(_02445_),
    .A1(net1460),
    .Y(_02446_),
    .A2(_02444_));
 sg13g2_a21oi_1 _07965_ (.A1(net1449),
    .A2(_01917_),
    .Y(_02447_),
    .B1(_02446_));
 sg13g2_a221oi_1 _07966_ (.B2(_02447_),
    .C1(net1545),
    .B1(_01962_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][4] ),
    .Y(_02448_),
    .A2(_01955_));
 sg13g2_a21oi_1 _07967_ (.A1(_00767_),
    .A2(net1545),
    .Y(_02449_),
    .B1(_02448_));
 sg13g2_a21oi_1 _07968_ (.A1(net1668),
    .A2(_02449_),
    .Y(_02450_),
    .B1(_01654_));
 sg13g2_nor2_1 _07969_ (.A(net1674),
    .B(_02450_),
    .Y(_02451_));
 sg13g2_o21ai_1 _07970_ (.B1(_02451_),
    .Y(_02452_),
    .A1(_01182_),
    .A2(_02438_));
 sg13g2_nand2b_1 _07971_ (.Y(_02453_),
    .B(_02258_),
    .A_N(_02273_));
 sg13g2_a21oi_1 _07972_ (.A1(_02245_),
    .A2(_02453_),
    .Y(_02454_),
    .B1(_02254_));
 sg13g2_nor2_1 _07973_ (.A(net1455),
    .B(_02265_),
    .Y(_02455_));
 sg13g2_o21ai_1 _07974_ (.B1(net1457),
    .Y(_02456_),
    .A1(_02263_),
    .A2(_02455_));
 sg13g2_nor2_1 _07975_ (.A(_02252_),
    .B(_02456_),
    .Y(_02457_));
 sg13g2_o21ai_1 _07976_ (.B1(_02342_),
    .Y(_02458_),
    .A1(_02454_),
    .A2(_02457_));
 sg13g2_nor2b_1 _07977_ (.A(_02262_),
    .B_N(_02300_),
    .Y(_02459_));
 sg13g2_nor2_1 _07978_ (.A(net1456),
    .B(net1444),
    .Y(_02460_));
 sg13g2_nor3_1 _07979_ (.A(net1447),
    .B(_02459_),
    .C(_02460_),
    .Y(_02461_));
 sg13g2_a22oi_1 _07980_ (.Y(_02462_),
    .B1(_02458_),
    .B2(_02461_),
    .A2(_02245_),
    .A1(net1447));
 sg13g2_a22oi_1 _07981_ (.Y(_02463_),
    .B1(_02299_),
    .B2(_02462_),
    .A2(net1720),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][4] ));
 sg13g2_o21ai_1 _07982_ (.B1(_02003_),
    .Y(_02464_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][4] ),
    .A2(net1664));
 sg13g2_a21oi_1 _07983_ (.A1(net1665),
    .A2(_02463_),
    .Y(_02465_),
    .B1(_02464_));
 sg13g2_nor2_2 _07984_ (.A(net1528),
    .B(_02465_),
    .Y(_02466_));
 sg13g2_inv_1 _07985_ (.Y(_02467_),
    .A(_02466_));
 sg13g2_a21oi_1 _07986_ (.A1(_02320_),
    .A2(_02467_),
    .Y(_02468_),
    .B1(net1509));
 sg13g2_a22oi_1 _07987_ (.Y(_00219_),
    .B1(_02452_),
    .B2(_02468_),
    .A2(net1512),
    .A1(_00714_));
 sg13g2_nor2_1 _07988_ (.A(net1433),
    .B(net1427),
    .Y(_02469_));
 sg13g2_nor2_1 _07989_ (.A(net1423),
    .B(_02469_),
    .Y(_02470_));
 sg13g2_a21oi_1 _07990_ (.A1(_01538_),
    .A2(_01566_),
    .Y(_02471_),
    .B1(net1430));
 sg13g2_nor2_1 _07991_ (.A(net1434),
    .B(_02471_),
    .Y(_02472_));
 sg13g2_nand3_1 _07992_ (.B(net1434),
    .C(_01564_),
    .A(_01542_),
    .Y(_02473_));
 sg13g2_nor2_1 _07993_ (.A(_01545_),
    .B(_02473_),
    .Y(_02474_));
 sg13g2_o21ai_1 _07994_ (.B1(_01562_),
    .Y(_02475_),
    .A1(_02472_),
    .A2(_02474_));
 sg13g2_a21oi_1 _07995_ (.A1(_01546_),
    .A2(_01564_),
    .Y(_02476_),
    .B1(net1432));
 sg13g2_nor3_1 _07996_ (.A(net1431),
    .B(_01566_),
    .C(_02476_),
    .Y(_02477_));
 sg13g2_a21oi_1 _07997_ (.A1(net1431),
    .A2(net1430),
    .Y(_02478_),
    .B1(_02477_));
 sg13g2_nand3_1 _07998_ (.B(_02475_),
    .C(_02478_),
    .A(_01606_),
    .Y(_02479_));
 sg13g2_a22oi_1 _07999_ (.Y(_02480_),
    .B1(_02470_),
    .B2(_02479_),
    .A2(net1423),
    .A1(net1431));
 sg13g2_inv_1 _08000_ (.Y(_02481_),
    .A(_02480_));
 sg13g2_a221oi_1 _08001_ (.B2(_02481_),
    .C1(net1486),
    .B1(_01615_),
    .A1(_01212_),
    .Y(_02482_),
    .A2(net1669));
 sg13g2_o21ai_1 _08002_ (.B1(net1500),
    .Y(_02483_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[5] ),
    .A2(net1487));
 sg13g2_o21ai_1 _08003_ (.B1(_01269_),
    .Y(_02484_),
    .A1(_02482_),
    .A2(_02483_));
 sg13g2_a22oi_1 _08004_ (.Y(_02485_),
    .B1(_01929_),
    .B2(net1469),
    .A2(_01925_),
    .A1(net1462));
 sg13g2_o21ai_1 _08005_ (.B1(net1452),
    .Y(_02486_),
    .A1(_01917_),
    .A2(net1460));
 sg13g2_a21oi_1 _08006_ (.A1(net1460),
    .A2(_02485_),
    .Y(_02487_),
    .B1(_02486_));
 sg13g2_nor2_1 _08007_ (.A(_01931_),
    .B(_01935_),
    .Y(_02488_));
 sg13g2_a21oi_1 _08008_ (.A1(_01912_),
    .A2(_01933_),
    .Y(_02489_),
    .B1(_02488_));
 sg13g2_a221oi_1 _08009_ (.B2(_02489_),
    .C1(_02487_),
    .B1(_01920_),
    .A1(net1449),
    .Y(_02490_),
    .A2(_01919_));
 sg13g2_a221oi_1 _08010_ (.B2(_02490_),
    .C1(net1545),
    .B1(_01962_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][5] ),
    .Y(_02491_),
    .A2(net1723));
 sg13g2_a21oi_1 _08011_ (.A1(_00766_),
    .A2(net1545),
    .Y(_02492_),
    .B1(_02491_));
 sg13g2_a21oi_1 _08012_ (.A1(net1668),
    .A2(_02492_),
    .Y(_02493_),
    .B1(_01654_));
 sg13g2_nor2_1 _08013_ (.A(net1674),
    .B(_02493_),
    .Y(_02494_));
 sg13g2_o21ai_1 _08014_ (.B1(_02494_),
    .Y(_02495_),
    .A1(net1531),
    .A2(_02484_));
 sg13g2_nand2_1 _08015_ (.Y(_02496_),
    .A(net1455),
    .B(_02259_));
 sg13g2_a21oi_1 _08016_ (.A1(_02260_),
    .A2(_02262_),
    .Y(_02497_),
    .B1(_02267_));
 sg13g2_nor3_1 _08017_ (.A(_02252_),
    .B(_02254_),
    .C(_02263_),
    .Y(_02498_));
 sg13g2_nor3_1 _08018_ (.A(net1459),
    .B(_02497_),
    .C(_02498_),
    .Y(_02499_));
 sg13g2_o21ai_1 _08019_ (.B1(net1457),
    .Y(_02500_),
    .A1(_02294_),
    .A2(_02499_));
 sg13g2_nand3_1 _08020_ (.B(_02262_),
    .C(net1443),
    .A(_02246_),
    .Y(_02501_));
 sg13g2_a21oi_1 _08021_ (.A1(net1455),
    .A2(_02300_),
    .Y(_02502_),
    .B1(net1447));
 sg13g2_nand3_1 _08022_ (.B(_02501_),
    .C(_02502_),
    .A(_02500_),
    .Y(_02503_));
 sg13g2_nand2_1 _08023_ (.Y(_02504_),
    .A(net1448),
    .B(net1458));
 sg13g2_nand2_1 _08024_ (.Y(_02505_),
    .A(_02503_),
    .B(_02504_));
 sg13g2_a22oi_1 _08025_ (.Y(_02506_),
    .B1(_02299_),
    .B2(_02505_),
    .A2(net1720),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][5] ));
 sg13g2_o21ai_1 _08026_ (.B1(_02003_),
    .Y(_02507_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][5] ),
    .A2(net1664));
 sg13g2_a21oi_1 _08027_ (.A1(net1664),
    .A2(_02506_),
    .Y(_02508_),
    .B1(_02507_));
 sg13g2_nor2_2 _08028_ (.A(net1528),
    .B(_02508_),
    .Y(_02509_));
 sg13g2_inv_1 _08029_ (.Y(_02510_),
    .A(_02509_));
 sg13g2_a21oi_1 _08030_ (.A1(_02320_),
    .A2(_02510_),
    .Y(_02511_),
    .B1(net1510));
 sg13g2_a22oi_1 _08031_ (.Y(_00220_),
    .B1(_02495_),
    .B2(_02511_),
    .A2(net1510),
    .A1(_00716_));
 sg13g2_nor2_1 _08032_ (.A(net1431),
    .B(net1423),
    .Y(_02512_));
 sg13g2_nand2_1 _08033_ (.Y(_02513_),
    .A(net1434),
    .B(_02471_));
 sg13g2_nand3_1 _08034_ (.B(_02473_),
    .C(_02476_),
    .A(_01566_),
    .Y(_02514_));
 sg13g2_nand2_1 _08035_ (.Y(_02515_),
    .A(net1432),
    .B(_01564_));
 sg13g2_nand4_1 _08036_ (.B(_02513_),
    .C(_02514_),
    .A(net1427),
    .Y(_02516_),
    .D(_02515_));
 sg13g2_o21ai_1 _08037_ (.B1(_01597_),
    .Y(_02517_),
    .A1(net1432),
    .A2(net1429));
 sg13g2_a22oi_1 _08038_ (.Y(_02518_),
    .B1(_02517_),
    .B2(net1428),
    .A2(_02516_),
    .A1(_02512_));
 sg13g2_a221oi_1 _08039_ (.B2(_02518_),
    .C1(net1486),
    .B1(_01615_),
    .A1(_01209_),
    .Y(_02519_),
    .A2(net1669));
 sg13g2_o21ai_1 _08040_ (.B1(net1500),
    .Y(_02520_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[6] ),
    .A2(net1489));
 sg13g2_o21ai_1 _08041_ (.B1(_01269_),
    .Y(_02521_),
    .A1(_02519_),
    .A2(_02520_));
 sg13g2_nor2_1 _08042_ (.A(net1449),
    .B(net1462),
    .Y(_02522_));
 sg13g2_a221oi_1 _08043_ (.B2(_01910_),
    .C1(net1462),
    .B1(_01931_),
    .A1(net1469),
    .Y(_02523_),
    .A2(_01924_));
 sg13g2_or2_1 _08044_ (.X(_02524_),
    .B(_02523_),
    .A(_01916_));
 sg13g2_a21oi_1 _08045_ (.A1(_01907_),
    .A2(net1469),
    .Y(_02525_),
    .B1(_01912_));
 sg13g2_nor2_1 _08046_ (.A(net1462),
    .B(_01924_),
    .Y(_02526_));
 sg13g2_o21ai_1 _08047_ (.B1(_02526_),
    .Y(_02527_),
    .A1(_01916_),
    .A2(_02525_));
 sg13g2_nand3_1 _08048_ (.B(_02524_),
    .C(_02527_),
    .A(_01947_),
    .Y(_02528_));
 sg13g2_o21ai_1 _08049_ (.B1(_02528_),
    .Y(_02529_),
    .A1(net1460),
    .A2(_02522_));
 sg13g2_a221oi_1 _08050_ (.B2(_02529_),
    .C1(net1545),
    .B1(_01962_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][6] ),
    .Y(_02530_),
    .A2(_01955_));
 sg13g2_o21ai_1 _08051_ (.B1(net1668),
    .Y(_02531_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][6] ),
    .A2(net1548));
 sg13g2_nor2_1 _08052_ (.A(_02530_),
    .B(_02531_),
    .Y(_02532_));
 sg13g2_nor2_1 _08053_ (.A(_01654_),
    .B(_02532_),
    .Y(_02533_));
 sg13g2_nor2_1 _08054_ (.A(net1674),
    .B(_02533_),
    .Y(_02534_));
 sg13g2_o21ai_1 _08055_ (.B1(_02534_),
    .Y(_02535_),
    .A1(net1530),
    .A2(_02521_));
 sg13g2_nor2_1 _08056_ (.A(net1448),
    .B(net1459),
    .Y(_02536_));
 sg13g2_o21ai_1 _08057_ (.B1(_02254_),
    .Y(_02537_),
    .A1(_02252_),
    .A2(_02263_));
 sg13g2_nand2b_1 _08058_ (.Y(_02538_),
    .B(net1456),
    .A_N(net1457));
 sg13g2_nand3_1 _08059_ (.B(_02537_),
    .C(_02538_),
    .A(net1443),
    .Y(_02539_));
 sg13g2_nand3_1 _08060_ (.B(_02267_),
    .C(_02496_),
    .A(_02262_),
    .Y(_02540_));
 sg13g2_nor2_1 _08061_ (.A(net1448),
    .B(_02245_),
    .Y(_02541_));
 sg13g2_a21oi_1 _08062_ (.A1(_02536_),
    .A2(_02540_),
    .Y(_02542_),
    .B1(_02541_));
 sg13g2_a22oi_1 _08063_ (.Y(_02543_),
    .B1(_02542_),
    .B2(net1443),
    .A2(_02539_),
    .A1(_02536_));
 sg13g2_a22oi_1 _08064_ (.Y(_02544_),
    .B1(_02299_),
    .B2(_02543_),
    .A2(net1719),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][6] ));
 sg13g2_o21ai_1 _08065_ (.B1(_02003_),
    .Y(_02545_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][6] ),
    .A2(net1665));
 sg13g2_a21oi_1 _08066_ (.A1(net1666),
    .A2(_02544_),
    .Y(_02546_),
    .B1(_02545_));
 sg13g2_nor2_2 _08067_ (.A(net1528),
    .B(_02546_),
    .Y(_02547_));
 sg13g2_nor2_1 _08068_ (.A(_02319_),
    .B(_02547_),
    .Y(_02548_));
 sg13g2_nor2_1 _08069_ (.A(net1508),
    .B(_02548_),
    .Y(_02549_));
 sg13g2_a22oi_1 _08070_ (.Y(_00221_),
    .B1(_02535_),
    .B2(_02549_),
    .A2(net1510),
    .A1(_00718_));
 sg13g2_o21ai_1 _08071_ (.B1(_01597_),
    .Y(_02550_),
    .A1(_01577_),
    .A2(_01607_));
 sg13g2_xnor2_1 _08072_ (.Y(_02551_),
    .A(net1490),
    .B(_02550_));
 sg13g2_a221oi_1 _08073_ (.B2(_02551_),
    .C1(_01620_),
    .B1(_01608_),
    .A1(_01236_),
    .Y(_02552_),
    .A2(net1670));
 sg13g2_o21ai_1 _08074_ (.B1(net1501),
    .Y(_02553_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[7] ),
    .A2(net1488));
 sg13g2_o21ai_1 _08075_ (.B1(_01261_),
    .Y(_02554_),
    .A1(_02552_),
    .A2(_02553_));
 sg13g2_o21ai_1 _08076_ (.B1(net1452),
    .Y(_02555_),
    .A1(_01939_),
    .A2(_01946_));
 sg13g2_xor2_1 _08077_ (.B(_02555_),
    .A(_01692_),
    .X(_02556_));
 sg13g2_a21oi_1 _08078_ (.A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][7] ),
    .A2(net1722),
    .Y(_02557_),
    .B1(net1546));
 sg13g2_o21ai_1 _08079_ (.B1(_02557_),
    .Y(_02558_),
    .A1(_01960_),
    .A2(_02556_));
 sg13g2_o21ai_1 _08080_ (.B1(_02558_),
    .Y(_02559_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][7] ),
    .A2(net1548));
 sg13g2_nor2_2 _08081_ (.A(_01645_),
    .B(_01647_),
    .Y(_02560_));
 sg13g2_nand2b_1 _08082_ (.Y(_02561_),
    .B(net1668),
    .A_N(_01645_));
 sg13g2_a21oi_1 _08083_ (.A1(_02559_),
    .A2(_02560_),
    .Y(_02562_),
    .B1(net1675));
 sg13g2_o21ai_1 _08084_ (.B1(_02562_),
    .Y(_02563_),
    .A1(net1530),
    .A2(_02554_));
 sg13g2_nor2_2 _08085_ (.A(_02002_),
    .B(net1528),
    .Y(_02564_));
 sg13g2_or2_2 _08086_ (.X(_02565_),
    .B(net1528),
    .A(_02002_));
 sg13g2_nand2_1 _08087_ (.Y(_02566_),
    .A(_00676_),
    .B(_02306_));
 sg13g2_nor2_1 _08088_ (.A(_02269_),
    .B(_02294_),
    .Y(_02567_));
 sg13g2_nor2_1 _08089_ (.A(net1446),
    .B(_02567_),
    .Y(_02568_));
 sg13g2_xnor2_1 _08090_ (.Y(_02569_),
    .A(_02042_),
    .B(_02568_));
 sg13g2_a21oi_1 _08091_ (.A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][7] ),
    .A2(net1719),
    .Y(_02570_),
    .B1(_02306_));
 sg13g2_o21ai_1 _08092_ (.B1(_02570_),
    .Y(_02571_),
    .A1(net1422),
    .A2(_02569_));
 sg13g2_a21oi_2 _08093_ (.B1(_02565_),
    .Y(_02572_),
    .A2(_02571_),
    .A1(_02566_));
 sg13g2_inv_1 _08094_ (.Y(_02573_),
    .A(_02572_));
 sg13g2_a21oi_1 _08095_ (.A1(net1418),
    .A2(_02573_),
    .Y(_02574_),
    .B1(net1511));
 sg13g2_a22oi_1 _08096_ (.Y(_00222_),
    .B1(_02563_),
    .B2(_02574_),
    .A2(net1511),
    .A1(_00720_));
 sg13g2_xor2_1 _08097_ (.B(_01579_),
    .A(_01318_),
    .X(_02575_));
 sg13g2_a21oi_1 _08098_ (.A1(net1429),
    .A2(_01576_),
    .Y(_02576_),
    .B1(net1490));
 sg13g2_nand2_1 _08099_ (.Y(_02577_),
    .A(_01582_),
    .B(_01586_));
 sg13g2_xor2_1 _08100_ (.B(_02577_),
    .A(_02576_),
    .X(_02578_));
 sg13g2_mux2_1 _08101_ (.A0(_01579_),
    .A1(_02578_),
    .S(net1428),
    .X(_02579_));
 sg13g2_nand2_1 _08102_ (.Y(_02580_),
    .A(net1426),
    .B(_02575_));
 sg13g2_o21ai_1 _08103_ (.B1(_02580_),
    .Y(_02581_),
    .A1(net1426),
    .A2(_02579_));
 sg13g2_a21oi_1 _08104_ (.A1(_01523_),
    .A2(_01614_),
    .Y(_02582_),
    .B1(_01620_));
 sg13g2_o21ai_1 _08105_ (.B1(_02582_),
    .Y(_02583_),
    .A1(_01233_),
    .A2(_01271_));
 sg13g2_a21oi_1 _08106_ (.A1(_01608_),
    .A2(_02581_),
    .Y(_02584_),
    .B1(_02583_));
 sg13g2_nor2_1 _08107_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[8] ),
    .B(net1488),
    .Y(_02585_));
 sg13g2_o21ai_1 _08108_ (.B1(_01261_),
    .Y(_02586_),
    .A1(_02584_),
    .A2(_02585_));
 sg13g2_nor2_1 _08109_ (.A(_01692_),
    .B(_01939_),
    .Y(_02587_));
 sg13g2_o21ai_1 _08110_ (.B1(_01697_),
    .Y(_02588_),
    .A1(_01921_),
    .A2(_01940_));
 sg13g2_or3_1 _08111_ (.A(_01697_),
    .B(_01921_),
    .C(_01940_),
    .X(_02589_));
 sg13g2_and2_1 _08112_ (.A(_02588_),
    .B(_02589_),
    .X(_02590_));
 sg13g2_a221oi_1 _08113_ (.B2(_02589_),
    .C1(_01692_),
    .B1(_02588_),
    .A1(_01919_),
    .Y(_02591_),
    .A2(_01938_));
 sg13g2_xnor2_1 _08114_ (.Y(_02592_),
    .A(_02587_),
    .B(_02590_));
 sg13g2_xnor2_1 _08115_ (.Y(_02593_),
    .A(_01692_),
    .B(_01698_));
 sg13g2_o21ai_1 _08116_ (.B1(net1451),
    .Y(_02594_),
    .A1(_01697_),
    .A2(net1461));
 sg13g2_a21o_1 _08117_ (.A2(_02592_),
    .A1(net1461),
    .B1(_02594_),
    .X(_02595_));
 sg13g2_o21ai_1 _08118_ (.B1(_02595_),
    .Y(_02596_),
    .A1(net1452),
    .A2(_02593_));
 sg13g2_a21oi_1 _08119_ (.A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][8] ),
    .A2(net1722),
    .Y(_02597_),
    .B1(net1546));
 sg13g2_o21ai_1 _08120_ (.B1(_02597_),
    .Y(_02598_),
    .A1(_01960_),
    .A2(_02596_));
 sg13g2_o21ai_1 _08121_ (.B1(_02598_),
    .Y(_02599_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][8] ),
    .A2(net1548));
 sg13g2_a21oi_1 _08122_ (.A1(_02560_),
    .A2(_02599_),
    .Y(_02600_),
    .B1(net1675));
 sg13g2_o21ai_1 _08123_ (.B1(_02600_),
    .Y(_02601_),
    .A1(net1530),
    .A2(_02586_));
 sg13g2_nand2b_1 _08124_ (.Y(_02602_),
    .B(_02306_),
    .A_N(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][8] ));
 sg13g2_xor2_1 _08125_ (.B(_02047_),
    .A(_02042_),
    .X(_02603_));
 sg13g2_nand2b_1 _08126_ (.Y(_02604_),
    .B(_02043_),
    .A_N(_02269_));
 sg13g2_nor4_2 _08127_ (.A(_02042_),
    .B(_02269_),
    .C(_02281_),
    .Y(_02605_),
    .D(_02286_));
 sg13g2_o21ai_1 _08128_ (.B1(_02604_),
    .Y(_02606_),
    .A1(_02281_),
    .A2(_02286_));
 sg13g2_nand3b_1 _08129_ (.B(_02606_),
    .C(net1444),
    .Y(_02607_),
    .A_N(_02605_));
 sg13g2_a21oi_1 _08130_ (.A1(net1527),
    .A2(_02294_),
    .Y(_02608_),
    .B1(net1448));
 sg13g2_a221oi_1 _08131_ (.B2(_02608_),
    .C1(_02298_),
    .B1(_02607_),
    .A1(net1446),
    .Y(_02609_),
    .A2(_02603_));
 sg13g2_nand2_2 _08132_ (.Y(_02610_),
    .A(_02238_),
    .B(net1666));
 sg13g2_a21oi_1 _08133_ (.A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][8] ),
    .A2(net1720),
    .Y(_02611_),
    .B1(_02610_));
 sg13g2_nand2b_1 _08134_ (.Y(_02612_),
    .B(_02611_),
    .A_N(_02609_));
 sg13g2_a21oi_2 _08135_ (.B1(_02565_),
    .Y(_02613_),
    .A2(_02612_),
    .A1(_02602_));
 sg13g2_inv_1 _08136_ (.Y(_02614_),
    .A(_02613_));
 sg13g2_a21oi_1 _08137_ (.A1(net1418),
    .A2(_02614_),
    .Y(_02615_),
    .B1(net1507));
 sg13g2_a22oi_1 _08138_ (.Y(_00223_),
    .B1(_02601_),
    .B2(_02615_),
    .A2(net1509),
    .A1(_00706_));
 sg13g2_and2_1 _08139_ (.A(_02278_),
    .B(_02289_),
    .X(_02616_));
 sg13g2_o21ai_1 _08140_ (.B1(_02616_),
    .Y(_02617_),
    .A1(_02286_),
    .A2(_02605_));
 sg13g2_nand2_1 _08141_ (.Y(_02618_),
    .A(net1444),
    .B(_02617_));
 sg13g2_nor3_1 _08142_ (.A(_02286_),
    .B(_02605_),
    .C(_02616_),
    .Y(_02619_));
 sg13g2_a21oi_1 _08143_ (.A1(_02051_),
    .A2(_02294_),
    .Y(_02620_),
    .B1(net1446));
 sg13g2_o21ai_1 _08144_ (.B1(_02620_),
    .Y(_02621_),
    .A1(_02618_),
    .A2(_02619_));
 sg13g2_xnor2_1 _08145_ (.Y(_02622_),
    .A(_02052_),
    .B(_02284_));
 sg13g2_a21oi_1 _08146_ (.A1(net1446),
    .A2(_02622_),
    .Y(_02623_),
    .B1(net1422));
 sg13g2_a221oi_1 _08147_ (.B2(_02623_),
    .C1(_02610_),
    .B1(_02621_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][9] ),
    .Y(_02624_),
    .A2(net1721));
 sg13g2_a21oi_1 _08148_ (.A1(_00677_),
    .A2(_02306_),
    .Y(_02625_),
    .B1(_02624_));
 sg13g2_nor2_2 _08149_ (.A(_02565_),
    .B(_02625_),
    .Y(_02626_));
 sg13g2_or2_1 _08150_ (.X(_02627_),
    .B(_02626_),
    .A(_02319_));
 sg13g2_nor2_1 _08151_ (.A(_01525_),
    .B(net1428),
    .Y(_02628_));
 sg13g2_nor2_1 _08152_ (.A(net1426),
    .B(_02628_),
    .Y(_02629_));
 sg13g2_and2_1 _08153_ (.A(_01570_),
    .B(_01584_),
    .X(_02630_));
 sg13g2_a21o_1 _08154_ (.A2(_02576_),
    .A1(_01586_),
    .B1(_01581_),
    .X(_02631_));
 sg13g2_a22oi_1 _08155_ (.Y(_02632_),
    .B1(_02630_),
    .B2(_02631_),
    .A2(_01592_),
    .A1(_01591_));
 sg13g2_o21ai_1 _08156_ (.B1(_02632_),
    .Y(_02633_),
    .A1(_02630_),
    .A2(_02631_));
 sg13g2_o21ai_1 _08157_ (.B1(_01525_),
    .Y(_02634_),
    .A1(net1490),
    .A2(_01579_));
 sg13g2_o21ai_1 _08158_ (.B1(_02634_),
    .Y(_02635_),
    .A1(net1490),
    .A2(_01609_));
 sg13g2_a22oi_1 _08159_ (.Y(_02636_),
    .B1(_02635_),
    .B2(net1426),
    .A2(_02633_),
    .A1(_02629_));
 sg13g2_o21ai_1 _08160_ (.B1(_02582_),
    .Y(_02637_),
    .A1(_01237_),
    .A2(_01271_));
 sg13g2_a21oi_1 _08161_ (.A1(_01608_),
    .A2(_02636_),
    .Y(_02638_),
    .B1(_02637_));
 sg13g2_nor2_1 _08162_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[9] ),
    .B(net1489),
    .Y(_02639_));
 sg13g2_o21ai_1 _08163_ (.B1(_01261_),
    .Y(_02640_),
    .A1(_02638_),
    .A2(_02639_));
 sg13g2_and2_1 _08164_ (.A(_01928_),
    .B(_01949_),
    .X(_02641_));
 sg13g2_or3_1 _08165_ (.A(_01942_),
    .B(_02591_),
    .C(_02641_),
    .X(_02642_));
 sg13g2_o21ai_1 _08166_ (.B1(_02641_),
    .Y(_02643_),
    .A1(_01942_),
    .A2(_02591_));
 sg13g2_nand3_1 _08167_ (.B(_02642_),
    .C(_02643_),
    .A(net1461),
    .Y(_02644_));
 sg13g2_o21ai_1 _08168_ (.B1(net1451),
    .Y(_02645_),
    .A1(_01702_),
    .A2(net1461));
 sg13g2_nor2b_1 _08169_ (.A(_02645_),
    .B_N(_02644_),
    .Y(_02646_));
 sg13g2_nor2_1 _08170_ (.A(_01702_),
    .B(_01959_),
    .Y(_02647_));
 sg13g2_xor2_1 _08171_ (.B(_01959_),
    .A(_01702_),
    .X(_02648_));
 sg13g2_nor2_1 _08172_ (.A(net1451),
    .B(_02648_),
    .Y(_02649_));
 sg13g2_nor2_1 _08173_ (.A(_02646_),
    .B(_02649_),
    .Y(_02650_));
 sg13g2_nand2_1 _08174_ (.Y(_02651_),
    .A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][9] ),
    .B(net1546));
 sg13g2_a22oi_1 _08175_ (.Y(_02652_),
    .B1(_01961_),
    .B2(_02650_),
    .A2(net1722),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][9] ));
 sg13g2_o21ai_1 _08176_ (.B1(_02651_),
    .Y(_02653_),
    .A1(net1547),
    .A2(_02652_));
 sg13g2_o21ai_1 _08177_ (.B1(_01187_),
    .Y(_02654_),
    .A1(_02561_),
    .A2(_02653_));
 sg13g2_nand2b_1 _08178_ (.Y(_02655_),
    .B(_02654_),
    .A_N(net1507));
 sg13g2_o21ai_1 _08179_ (.B1(_02655_),
    .Y(_02656_),
    .A1(net1530),
    .A2(_02640_));
 sg13g2_a22oi_1 _08180_ (.Y(_00224_),
    .B1(_02627_),
    .B2(_02656_),
    .A2(net1509),
    .A1(_00708_));
 sg13g2_a21o_1 _08181_ (.A2(_02632_),
    .A1(_01584_),
    .B1(_01572_),
    .X(_02657_));
 sg13g2_a221oi_1 _08182_ (.B2(_02631_),
    .C1(_01585_),
    .B1(_02630_),
    .A1(_01591_),
    .Y(_02658_),
    .A2(_01592_));
 sg13g2_a21oi_2 _08183_ (.B1(_01585_),
    .Y(_02659_),
    .A2(_02631_),
    .A1(_02630_));
 sg13g2_nor2_1 _08184_ (.A(net1425),
    .B(_02658_),
    .Y(_02660_));
 sg13g2_nor3_2 _08185_ (.A(net1490),
    .B(_01572_),
    .C(_01609_),
    .Y(_02661_));
 sg13g2_o21ai_1 _08186_ (.B1(_01572_),
    .Y(_02662_),
    .A1(net1490),
    .A2(_01609_));
 sg13g2_nand2b_1 _08187_ (.Y(_02663_),
    .B(_02662_),
    .A_N(_02661_));
 sg13g2_a22oi_1 _08188_ (.Y(_02664_),
    .B1(_02663_),
    .B2(net1426),
    .A2(_02660_),
    .A1(_02657_));
 sg13g2_o21ai_1 _08189_ (.B1(net1488),
    .Y(_02665_),
    .A1(_01249_),
    .A2(_01271_));
 sg13g2_a21oi_1 _08190_ (.A1(_01608_),
    .A2(_02664_),
    .Y(_02666_),
    .B1(_02665_));
 sg13g2_o21ai_1 _08191_ (.B1(net1501),
    .Y(_02667_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[10] ),
    .A2(net1488));
 sg13g2_o21ai_1 _08192_ (.B1(_01261_),
    .Y(_02668_),
    .A1(_02666_),
    .A2(_02667_));
 sg13g2_nand2_1 _08193_ (.Y(_02669_),
    .A(net1450),
    .B(_02647_));
 sg13g2_nand3_1 _08194_ (.B(_01949_),
    .C(_02643_),
    .A(_01947_),
    .Y(_02670_));
 sg13g2_nand2_1 _08195_ (.Y(_02671_),
    .A(_02669_),
    .B(_02670_));
 sg13g2_xnor2_1 _08196_ (.Y(_02672_),
    .A(_01707_),
    .B(_02671_));
 sg13g2_a221oi_1 _08197_ (.B2(_02672_),
    .C1(net1547),
    .B1(_01961_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][10] ),
    .Y(_02673_),
    .A2(net1722));
 sg13g2_a21oi_1 _08198_ (.A1(_00769_),
    .A2(net1547),
    .Y(_02674_),
    .B1(_02673_));
 sg13g2_nor2_1 _08199_ (.A(_02561_),
    .B(_02674_),
    .Y(_02675_));
 sg13g2_nor2_1 _08200_ (.A(net1674),
    .B(_02675_),
    .Y(_02676_));
 sg13g2_o21ai_1 _08201_ (.B1(_02676_),
    .Y(_02677_),
    .A1(net1531),
    .A2(_02668_));
 sg13g2_nor2_1 _08202_ (.A(net1786),
    .B(net1666),
    .Y(_02678_));
 sg13g2_nor2b_1 _08203_ (.A(_02618_),
    .B_N(_02289_),
    .Y(_02679_));
 sg13g2_nand3_1 _08204_ (.B(net1444),
    .C(_02617_),
    .A(_02290_),
    .Y(_02680_));
 sg13g2_nor2b_1 _08205_ (.A(net1446),
    .B_N(_02680_),
    .Y(_02681_));
 sg13g2_o21ai_1 _08206_ (.B1(_02681_),
    .Y(_02682_),
    .A1(_02057_),
    .A2(_02679_));
 sg13g2_or2_1 _08207_ (.X(_02683_),
    .B(_02284_),
    .A(_02236_));
 sg13g2_o21ai_1 _08208_ (.B1(_02057_),
    .Y(_02684_),
    .A1(_02052_),
    .A2(_02284_));
 sg13g2_nand2_1 _08209_ (.Y(_02685_),
    .A(_02683_),
    .B(_02684_));
 sg13g2_a21oi_1 _08210_ (.A1(net1445),
    .A2(_02685_),
    .Y(_02686_),
    .B1(net1422));
 sg13g2_a221oi_1 _08211_ (.B2(_02686_),
    .C1(_02610_),
    .B1(_02682_),
    .A1(net1785),
    .Y(_02687_),
    .A2(net1721));
 sg13g2_o21ai_1 _08212_ (.B1(_02564_),
    .Y(_02688_),
    .A1(_02678_),
    .A2(_02687_));
 sg13g2_a21oi_1 _08213_ (.A1(net1418),
    .A2(_02688_),
    .Y(_02689_),
    .B1(net1511));
 sg13g2_a22oi_1 _08214_ (.Y(_00225_),
    .B1(_02677_),
    .B2(_02689_),
    .A2(net1510),
    .A1(_00711_));
 sg13g2_mux2_1 _08215_ (.A0(_02658_),
    .A1(_02661_),
    .S(net1425),
    .X(_02690_));
 sg13g2_xnor2_1 _08216_ (.Y(_02691_),
    .A(_01589_),
    .B(_02690_));
 sg13g2_a221oi_1 _08217_ (.B2(_02691_),
    .C1(net1486),
    .B1(_01608_),
    .A1(_01240_),
    .Y(_02692_),
    .A2(net1669));
 sg13g2_nor2_1 _08218_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[11] ),
    .B(net1489),
    .Y(_02693_));
 sg13g2_o21ai_1 _08219_ (.B1(_01261_),
    .Y(_02694_),
    .A1(_02692_),
    .A2(_02693_));
 sg13g2_nand3_1 _08220_ (.B(_01950_),
    .C(_02643_),
    .A(net1461),
    .Y(_02695_));
 sg13g2_nand2_1 _08221_ (.Y(_02696_),
    .A(_01706_),
    .B(_02647_));
 sg13g2_and2_1 _08222_ (.A(net1450),
    .B(_02696_),
    .X(_02697_));
 sg13g2_a21oi_1 _08223_ (.A1(net1451),
    .A2(_02695_),
    .Y(_02698_),
    .B1(_02697_));
 sg13g2_xnor2_1 _08224_ (.Y(_02699_),
    .A(_01710_),
    .B(_02698_));
 sg13g2_a21oi_1 _08225_ (.A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][11] ),
    .A2(net1722),
    .Y(_02700_),
    .B1(net1546));
 sg13g2_o21ai_1 _08226_ (.B1(_02700_),
    .Y(_02701_),
    .A1(_01960_),
    .A2(_02699_));
 sg13g2_o21ai_1 _08227_ (.B1(_02701_),
    .Y(_02702_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][11] ),
    .A2(_01967_));
 sg13g2_a21oi_1 _08228_ (.A1(_02560_),
    .A2(_02702_),
    .Y(_02703_),
    .B1(net1675));
 sg13g2_o21ai_1 _08229_ (.B1(_02703_),
    .Y(_02704_),
    .A1(net1530),
    .A2(_02694_));
 sg13g2_mux2_1 _08230_ (.A0(_02680_),
    .A1(_02683_),
    .S(net1445),
    .X(_02705_));
 sg13g2_xnor2_1 _08231_ (.Y(_02706_),
    .A(_02063_),
    .B(_02705_));
 sg13g2_a21oi_1 _08232_ (.A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][11] ),
    .A2(net1720),
    .Y(_02707_),
    .B1(_02610_));
 sg13g2_o21ai_1 _08233_ (.B1(_02707_),
    .Y(_02708_),
    .A1(net1422),
    .A2(_02706_));
 sg13g2_o21ai_1 _08234_ (.B1(_02708_),
    .Y(_02709_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][11] ),
    .A2(net1666));
 sg13g2_nand2_2 _08235_ (.Y(_02710_),
    .A(_02564_),
    .B(_02709_));
 sg13g2_a21oi_1 _08236_ (.A1(net1418),
    .A2(_02710_),
    .Y(_02711_),
    .B1(net1507));
 sg13g2_a22oi_1 _08237_ (.Y(_00226_),
    .B1(_02704_),
    .B2(_02711_),
    .A2(net1508),
    .A1(_00713_));
 sg13g2_nor2_1 _08238_ (.A(_01588_),
    .B(_02658_),
    .Y(_02712_));
 sg13g2_and4_1 _08239_ (.A(_01588_),
    .B(_01589_),
    .C(_01606_),
    .D(_02659_),
    .X(_02713_));
 sg13g2_nor4_1 _08240_ (.A(net1426),
    .B(_01612_),
    .C(_02712_),
    .D(_02713_),
    .Y(_02714_));
 sg13g2_nor2b_1 _08241_ (.A(_01589_),
    .B_N(_02661_),
    .Y(_02715_));
 sg13g2_nand2_1 _08242_ (.Y(_02716_),
    .A(_01612_),
    .B(_02661_));
 sg13g2_xnor2_1 _08243_ (.Y(_02717_),
    .A(_01588_),
    .B(_02715_));
 sg13g2_o21ai_1 _08244_ (.B1(_01608_),
    .Y(_02718_),
    .A1(_01597_),
    .A2(_02717_));
 sg13g2_o21ai_1 _08245_ (.B1(net1670),
    .Y(_02719_),
    .A1(_01246_),
    .A2(_01247_));
 sg13g2_o21ai_1 _08246_ (.B1(_02719_),
    .Y(_02720_),
    .A1(_02714_),
    .A2(_02718_));
 sg13g2_o21ai_1 _08247_ (.B1(_01261_),
    .Y(_02721_),
    .A1(_00699_),
    .A2(net1488));
 sg13g2_a21oi_1 _08248_ (.A1(net1488),
    .A2(_02720_),
    .Y(_02722_),
    .B1(_02721_));
 sg13g2_nand2b_1 _08249_ (.Y(_02723_),
    .B(_01900_),
    .A_N(_01713_));
 sg13g2_mux2_1 _08250_ (.A0(_02723_),
    .A1(_01712_),
    .S(_02695_),
    .X(_02724_));
 sg13g2_o21ai_1 _08251_ (.B1(net1450),
    .Y(_02725_),
    .A1(_02696_),
    .A2(_02723_));
 sg13g2_a21oi_1 _08252_ (.A1(_01712_),
    .A2(_02696_),
    .Y(_02726_),
    .B1(_02725_));
 sg13g2_nor2_1 _08253_ (.A(_01960_),
    .B(_02726_),
    .Y(_02727_));
 sg13g2_o21ai_1 _08254_ (.B1(_02727_),
    .Y(_02728_),
    .A1(net1450),
    .A2(_02724_));
 sg13g2_a21oi_1 _08255_ (.A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][12] ),
    .A2(net1722),
    .Y(_02729_),
    .B1(net1546));
 sg13g2_a22oi_1 _08256_ (.Y(_02730_),
    .B1(_02728_),
    .B2(_02729_),
    .A2(net1545),
    .A1(_00770_));
 sg13g2_o21ai_1 _08257_ (.B1(_01187_),
    .Y(_02731_),
    .A1(_02561_),
    .A2(_02730_));
 sg13g2_a21o_1 _08258_ (.A2(_02722_),
    .A1(_01183_),
    .B1(_02731_),
    .X(_02732_));
 sg13g2_o21ai_1 _08259_ (.B1(_02064_),
    .Y(_02733_),
    .A1(_02062_),
    .A2(_02680_));
 sg13g2_nand4_1 _08260_ (.B(_02290_),
    .C(net1444),
    .A(_02065_),
    .Y(_02734_),
    .D(_02617_));
 sg13g2_nor2b_1 _08261_ (.A(net1445),
    .B_N(_02733_),
    .Y(_02735_));
 sg13g2_nor2_1 _08262_ (.A(_02063_),
    .B(_02683_),
    .Y(_02736_));
 sg13g2_nand2_1 _08263_ (.Y(_02737_),
    .A(_02064_),
    .B(_02736_));
 sg13g2_xnor2_1 _08264_ (.Y(_02738_),
    .A(_02064_),
    .B(_02736_));
 sg13g2_nand2_1 _08265_ (.Y(_02739_),
    .A(net1445),
    .B(_02738_));
 sg13g2_a21oi_1 _08266_ (.A1(_02734_),
    .A2(_02735_),
    .Y(_02740_),
    .B1(net1422));
 sg13g2_a221oi_1 _08267_ (.B2(_02740_),
    .C1(_02610_),
    .B1(_02739_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][12] ),
    .Y(_02741_),
    .A2(net1719));
 sg13g2_nor2_1 _08268_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][12] ),
    .B(net1666),
    .Y(_02742_));
 sg13g2_o21ai_1 _08269_ (.B1(_02564_),
    .Y(_02743_),
    .A1(_02741_),
    .A2(_02742_));
 sg13g2_a21oi_2 _08270_ (.B1(net1507),
    .Y(_02744_),
    .A2(_02743_),
    .A1(net1418));
 sg13g2_a22oi_1 _08271_ (.Y(_00227_),
    .B1(_02732_),
    .B2(_02744_),
    .A2(net1512),
    .A1(_00715_));
 sg13g2_a21oi_1 _08272_ (.A1(_01602_),
    .A2(_02659_),
    .Y(_02745_),
    .B1(net1425));
 sg13g2_o21ai_1 _08273_ (.B1(_02745_),
    .Y(_02746_),
    .A1(_01599_),
    .A2(_02713_));
 sg13g2_nor2_1 _08274_ (.A(_01599_),
    .B(_02716_),
    .Y(_02747_));
 sg13g2_and2_1 _08275_ (.A(_01599_),
    .B(_02716_),
    .X(_02748_));
 sg13g2_o21ai_1 _08276_ (.B1(net1425),
    .Y(_02749_),
    .A1(_02747_),
    .A2(_02748_));
 sg13g2_and2_1 _08277_ (.A(_01608_),
    .B(_02749_),
    .X(_02750_));
 sg13g2_o21ai_1 _08278_ (.B1(net1488),
    .Y(_02751_),
    .A1(_01252_),
    .A2(_01271_));
 sg13g2_a21o_1 _08279_ (.A2(_02750_),
    .A1(_02746_),
    .B1(_02751_),
    .X(_02752_));
 sg13g2_o21ai_1 _08280_ (.B1(net1501),
    .Y(_02753_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[13] ),
    .A2(net1488));
 sg13g2_inv_1 _08281_ (.Y(_02754_),
    .A(_02753_));
 sg13g2_a21oi_1 _08282_ (.A1(_02752_),
    .A2(_02754_),
    .Y(_02755_),
    .B1(_01262_));
 sg13g2_nor2_1 _08283_ (.A(_01900_),
    .B(_02696_),
    .Y(_02756_));
 sg13g2_nor2_1 _08284_ (.A(net1451),
    .B(_02756_),
    .Y(_02757_));
 sg13g2_nand4_1 _08285_ (.B(net1461),
    .C(_01950_),
    .A(_01713_),
    .Y(_02758_),
    .D(_02643_));
 sg13g2_a21oi_1 _08286_ (.A1(net1451),
    .A2(_02758_),
    .Y(_02759_),
    .B1(_02757_));
 sg13g2_xor2_1 _08287_ (.B(_02759_),
    .A(_01718_),
    .X(_02760_));
 sg13g2_a21oi_1 _08288_ (.A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][13] ),
    .A2(net1722),
    .Y(_02761_),
    .B1(net1546));
 sg13g2_o21ai_1 _08289_ (.B1(_02761_),
    .Y(_02762_),
    .A1(_01960_),
    .A2(_02760_));
 sg13g2_o21ai_1 _08290_ (.B1(_02762_),
    .Y(_02763_),
    .A1(net1787),
    .A2(net1548));
 sg13g2_a21o_1 _08291_ (.A2(_02763_),
    .A1(_02560_),
    .B1(net1675),
    .X(_02764_));
 sg13g2_a21o_1 _08292_ (.A2(_02755_),
    .A1(_01183_),
    .B1(_02764_),
    .X(_02765_));
 sg13g2_nand2_1 _08293_ (.Y(_02766_),
    .A(_00678_),
    .B(_02306_));
 sg13g2_mux2_1 _08294_ (.A0(_02734_),
    .A1(_02737_),
    .S(net1445),
    .X(_02767_));
 sg13g2_nor3_1 _08295_ (.A(_02063_),
    .B(_02235_),
    .C(_02683_),
    .Y(_02768_));
 sg13g2_nor2_1 _08296_ (.A(_02073_),
    .B(_02734_),
    .Y(_02769_));
 sg13g2_xor2_1 _08297_ (.B(_02767_),
    .A(_02073_),
    .X(_02770_));
 sg13g2_a21oi_1 _08298_ (.A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][13] ),
    .A2(net1719),
    .Y(_02771_),
    .B1(_02610_));
 sg13g2_o21ai_1 _08299_ (.B1(_02771_),
    .Y(_02772_),
    .A1(net1422),
    .A2(_02770_));
 sg13g2_a21oi_2 _08300_ (.B1(_02565_),
    .Y(_02773_),
    .A2(_02772_),
    .A1(_02766_));
 sg13g2_inv_1 _08301_ (.Y(_02774_),
    .A(_02773_));
 sg13g2_a21oi_1 _08302_ (.A1(net1418),
    .A2(_02774_),
    .Y(_02775_),
    .B1(net1508));
 sg13g2_a22oi_1 _08303_ (.Y(_00228_),
    .B1(_02765_),
    .B2(_02775_),
    .A2(net1512),
    .A1(_00717_));
 sg13g2_xnor2_1 _08304_ (.Y(_02776_),
    .A(_01718_),
    .B(net1451));
 sg13g2_nand2_1 _08305_ (.Y(_02777_),
    .A(_02759_),
    .B(_02776_));
 sg13g2_xnor2_1 _08306_ (.Y(_02778_),
    .A(_01671_),
    .B(_02777_));
 sg13g2_a21oi_1 _08307_ (.A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][14] ),
    .A2(net1723),
    .Y(_02779_),
    .B1(net1546));
 sg13g2_o21ai_1 _08308_ (.B1(_02779_),
    .Y(_02780_),
    .A1(_01960_),
    .A2(_02778_));
 sg13g2_o21ai_1 _08309_ (.B1(_02780_),
    .Y(_02781_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][14] ),
    .A2(net1548));
 sg13g2_a21oi_1 _08310_ (.A1(_01602_),
    .A2(_02659_),
    .Y(_02782_),
    .B1(_01601_));
 sg13g2_a21oi_1 _08311_ (.A1(_01603_),
    .A2(_02659_),
    .Y(_02783_),
    .B1(net1425));
 sg13g2_nand2b_1 _08312_ (.Y(_02784_),
    .B(_02783_),
    .A_N(_02782_));
 sg13g2_o21ai_1 _08313_ (.B1(net1425),
    .Y(_02785_),
    .A1(_01601_),
    .A2(_02747_));
 sg13g2_a21oi_1 _08314_ (.A1(_01601_),
    .A2(_02747_),
    .Y(_02786_),
    .B1(_02785_));
 sg13g2_nor3_1 _08315_ (.A(_01524_),
    .B(_01605_),
    .C(_02786_),
    .Y(_02787_));
 sg13g2_o21ai_1 _08316_ (.B1(_02582_),
    .Y(_02788_),
    .A1(_01245_),
    .A2(_01271_));
 sg13g2_a21o_1 _08317_ (.A2(_02787_),
    .A1(_02784_),
    .B1(_02788_),
    .X(_02789_));
 sg13g2_nand2_1 _08318_ (.Y(_02790_),
    .A(_00701_),
    .B(net1486));
 sg13g2_a21oi_1 _08319_ (.A1(_02789_),
    .A2(_02790_),
    .Y(_02791_),
    .B1(_01262_));
 sg13g2_a21o_1 _08320_ (.A2(_02781_),
    .A1(_02560_),
    .B1(net1675),
    .X(_02792_));
 sg13g2_a21o_1 _08321_ (.A2(_02791_),
    .A1(_01183_),
    .B1(_02792_),
    .X(_02793_));
 sg13g2_xor2_1 _08322_ (.B(_02768_),
    .A(_02026_),
    .X(_02794_));
 sg13g2_a21oi_1 _08323_ (.A1(net1445),
    .A2(_02794_),
    .Y(_02795_),
    .B1(net1422));
 sg13g2_xor2_1 _08324_ (.B(_02769_),
    .A(_02026_),
    .X(_02796_));
 sg13g2_nand2b_1 _08325_ (.Y(_02797_),
    .B(_02796_),
    .A_N(net1445));
 sg13g2_a221oi_1 _08326_ (.B2(_02797_),
    .C1(_02610_),
    .B1(_02795_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][14] ),
    .Y(_02798_),
    .A2(net1721));
 sg13g2_nor2_1 _08327_ (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][14] ),
    .B(net1666),
    .Y(_02799_));
 sg13g2_o21ai_1 _08328_ (.B1(_02564_),
    .Y(_02800_),
    .A1(_02798_),
    .A2(_02799_));
 sg13g2_a21oi_1 _08329_ (.A1(net1418),
    .A2(_02800_),
    .Y(_02801_),
    .B1(net1507));
 sg13g2_a22oi_1 _08330_ (.Y(_00229_),
    .B1(_02793_),
    .B2(_02801_),
    .A2(net1512),
    .A1(_00719_));
 sg13g2_nand2_1 _08331_ (.Y(_02802_),
    .A(_01271_),
    .B(_01526_));
 sg13g2_a21oi_1 _08332_ (.A1(_01228_),
    .A2(net1670),
    .Y(_02803_),
    .B1(net1486));
 sg13g2_o21ai_1 _08333_ (.B1(_02803_),
    .Y(_02804_),
    .A1(_01605_),
    .A2(_02802_));
 sg13g2_o21ai_1 _08334_ (.B1(net1501),
    .Y(_02805_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[15] ),
    .A2(net1489));
 sg13g2_inv_1 _08335_ (.Y(_02806_),
    .A(_02805_));
 sg13g2_a21oi_1 _08336_ (.A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[15] ),
    .A2(_01266_),
    .Y(_02807_),
    .B1(_01228_));
 sg13g2_o21ai_1 _08337_ (.B1(_01263_),
    .Y(_02808_),
    .A1(net1500),
    .A2(_02807_));
 sg13g2_a21oi_2 _08338_ (.B1(_02808_),
    .Y(_02809_),
    .A2(_02806_),
    .A1(_02804_));
 sg13g2_a221oi_1 _08339_ (.B2(_01855_),
    .C1(net1546),
    .B1(_01961_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][15] ),
    .Y(_02810_),
    .A2(net1722));
 sg13g2_o21ai_1 _08340_ (.B1(net1668),
    .Y(_02811_),
    .A1(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][15] ),
    .A2(net1548));
 sg13g2_o21ai_1 _08341_ (.B1(_01651_),
    .Y(_02812_),
    .A1(_02810_),
    .A2(_02811_));
 sg13g2_a21oi_1 _08342_ (.A1(_01183_),
    .A2(_02809_),
    .Y(_02813_),
    .B1(net1674));
 sg13g2_o21ai_1 _08343_ (.B1(_02813_),
    .Y(_02814_),
    .A1(_01645_),
    .A2(_02812_));
 sg13g2_a21oi_1 _08344_ (.A1(_02314_),
    .A2(_02318_),
    .Y(_02815_),
    .B1(net1510));
 sg13g2_a22oi_1 _08345_ (.Y(_00230_),
    .B1(_02814_),
    .B2(_02815_),
    .A2(net1510),
    .A1(_00721_));
 sg13g2_a22oi_1 _08346_ (.Y(_00231_),
    .B1(_01049_),
    .B2(_00651_),
    .A2(_00800_),
    .A1(net674));
 sg13g2_a21oi_1 _08347_ (.A1(_00652_),
    .A2(_00660_),
    .Y(_02816_),
    .B1(_00799_));
 sg13g2_nand3_1 _08348_ (.B(_01048_),
    .C(net1717),
    .A(net1822),
    .Y(_02817_));
 sg13g2_o21ai_1 _08349_ (.B1(_02817_),
    .Y(_00232_),
    .A1(_00650_),
    .A2(net1717));
 sg13g2_nand3_1 _08350_ (.B(_01048_),
    .C(net1717),
    .A(net1817),
    .Y(_02818_));
 sg13g2_o21ai_1 _08351_ (.B1(_02818_),
    .Y(_00233_),
    .A1(_00649_),
    .A2(net1717));
 sg13g2_nand3_1 _08352_ (.B(_01048_),
    .C(net1717),
    .A(net1813),
    .Y(_02819_));
 sg13g2_o21ai_1 _08353_ (.B1(_02819_),
    .Y(_00234_),
    .A1(_00648_),
    .A2(net1717));
 sg13g2_nand3_1 _08354_ (.B(_01048_),
    .C(net1717),
    .A(net1809),
    .Y(_02820_));
 sg13g2_o21ai_1 _08355_ (.B1(_02820_),
    .Y(_00235_),
    .A1(_00647_),
    .A2(net1718));
 sg13g2_nand3_1 _08356_ (.B(_01048_),
    .C(net1718),
    .A(net1802),
    .Y(_02821_));
 sg13g2_o21ai_1 _08357_ (.B1(_02821_),
    .Y(_00236_),
    .A1(_00723_),
    .A2(net1718));
 sg13g2_nand3_1 _08358_ (.B(_01048_),
    .C(net1718),
    .A(net1865),
    .Y(_02822_));
 sg13g2_o21ai_1 _08359_ (.B1(_02822_),
    .Y(_00237_),
    .A1(_00656_),
    .A2(net1717));
 sg13g2_o21ai_1 _08360_ (.B1(_01039_),
    .Y(_02823_),
    .A1(_00655_),
    .A2(net1793));
 sg13g2_o21ai_1 _08361_ (.B1(_02823_),
    .Y(_02824_),
    .A1(net1727),
    .A2(_01018_));
 sg13g2_nand2b_1 _08362_ (.Y(_02825_),
    .B(net1477),
    .A_N(net1727));
 sg13g2_and2_1 _08363_ (.A(_02823_),
    .B(_02825_),
    .X(_02826_));
 sg13g2_o21ai_1 _08364_ (.B1(_02824_),
    .Y(_02827_),
    .A1(net1033),
    .A2(net1472));
 sg13g2_inv_1 _08365_ (.Y(_00238_),
    .A(_02827_));
 sg13g2_o21ai_1 _08366_ (.B1(_02823_),
    .Y(_02828_),
    .A1(net1727),
    .A2(_01004_));
 sg13g2_o21ai_1 _08367_ (.B1(_02828_),
    .Y(_02829_),
    .A1(net1015),
    .A2(net1472));
 sg13g2_inv_1 _08368_ (.Y(_00239_),
    .A(_02829_));
 sg13g2_o21ai_1 _08369_ (.B1(_02823_),
    .Y(_02830_),
    .A1(net1727),
    .A2(_00990_));
 sg13g2_o21ai_1 _08370_ (.B1(_02830_),
    .Y(_02831_),
    .A1(net999),
    .A2(net1471));
 sg13g2_inv_1 _08371_ (.Y(_00240_),
    .A(_02831_));
 sg13g2_o21ai_1 _08372_ (.B1(_02823_),
    .Y(_02832_),
    .A1(net1727),
    .A2(_00978_));
 sg13g2_o21ai_1 _08373_ (.B1(_02832_),
    .Y(_02833_),
    .A1(net971),
    .A2(net1471));
 sg13g2_inv_1 _08374_ (.Y(_00241_),
    .A(_02833_));
 sg13g2_o21ai_1 _08375_ (.B1(_02823_),
    .Y(_02834_),
    .A1(net1727),
    .A2(_00968_));
 sg13g2_o21ai_1 _08376_ (.B1(_02834_),
    .Y(_02835_),
    .A1(net1001),
    .A2(net1472));
 sg13g2_inv_1 _08377_ (.Y(_00242_),
    .A(_02835_));
 sg13g2_o21ai_1 _08378_ (.B1(_02823_),
    .Y(_02836_),
    .A1(net1727),
    .A2(_00953_));
 sg13g2_o21ai_1 _08379_ (.B1(_02836_),
    .Y(_02837_),
    .A1(net980),
    .A2(net1471));
 sg13g2_inv_1 _08380_ (.Y(_00243_),
    .A(_02837_));
 sg13g2_o21ai_1 _08381_ (.B1(_02823_),
    .Y(_02838_),
    .A1(net1727),
    .A2(_00942_));
 sg13g2_o21ai_1 _08382_ (.B1(_02838_),
    .Y(_02839_),
    .A1(net1020),
    .A2(net1474));
 sg13g2_inv_1 _08383_ (.Y(_00244_),
    .A(_02839_));
 sg13g2_nor2_1 _08384_ (.A(net1002),
    .B(net1471),
    .Y(_02840_));
 sg13g2_nor2_1 _08385_ (.A(net1833),
    .B(net1728),
    .Y(_02841_));
 sg13g2_a21oi_1 _08386_ (.A1(net1471),
    .A2(_02841_),
    .Y(_00245_),
    .B1(_02840_));
 sg13g2_nor2_1 _08387_ (.A(net946),
    .B(net1471),
    .Y(_02842_));
 sg13g2_nor2_1 _08388_ (.A(net1830),
    .B(net1728),
    .Y(_02843_));
 sg13g2_a21oi_1 _08389_ (.A1(net1471),
    .A2(_02843_),
    .Y(_00246_),
    .B1(_02842_));
 sg13g2_nor2_1 _08390_ (.A(net954),
    .B(net1473),
    .Y(_02844_));
 sg13g2_nor2_1 _08391_ (.A(\u_tiny_nn_top.data_i_q[9] ),
    .B(net1729),
    .Y(_02845_));
 sg13g2_a21oi_1 _08392_ (.A1(net1473),
    .A2(_02845_),
    .Y(_00247_),
    .B1(_02844_));
 sg13g2_nor2_1 _08393_ (.A(net981),
    .B(net1473),
    .Y(_02846_));
 sg13g2_nor2_1 _08394_ (.A(\u_tiny_nn_top.data_i_q[10] ),
    .B(net1728),
    .Y(_02847_));
 sg13g2_a21oi_1 _08395_ (.A1(net1471),
    .A2(_02847_),
    .Y(_00248_),
    .B1(_02846_));
 sg13g2_nor2_1 _08396_ (.A(net995),
    .B(net1473),
    .Y(_02848_));
 sg13g2_nor2_1 _08397_ (.A(\u_tiny_nn_top.data_i_q[11] ),
    .B(net1729),
    .Y(_02849_));
 sg13g2_a21oi_1 _08398_ (.A1(net1473),
    .A2(_02849_),
    .Y(_00249_),
    .B1(_02848_));
 sg13g2_nor2_1 _08399_ (.A(net960),
    .B(net1473),
    .Y(_02850_));
 sg13g2_nor2_1 _08400_ (.A(net1828),
    .B(net1729),
    .Y(_02851_));
 sg13g2_a21oi_1 _08401_ (.A1(net1473),
    .A2(_02851_),
    .Y(_00250_),
    .B1(_02850_));
 sg13g2_nor2_1 _08402_ (.A(net973),
    .B(net1473),
    .Y(_02852_));
 sg13g2_nor2_1 _08403_ (.A(\u_tiny_nn_top.data_i_q[13] ),
    .B(net1729),
    .Y(_02853_));
 sg13g2_a21oi_1 _08404_ (.A1(net1474),
    .A2(_02853_),
    .Y(_00251_),
    .B1(_02852_));
 sg13g2_nor2_1 _08405_ (.A(net970),
    .B(net1474),
    .Y(_02854_));
 sg13g2_nor2_1 _08406_ (.A(net1827),
    .B(net1729),
    .Y(_02855_));
 sg13g2_a21oi_1 _08407_ (.A1(net1474),
    .A2(_02855_),
    .Y(_00252_),
    .B1(_02854_));
 sg13g2_nor2_1 _08408_ (.A(net987),
    .B(net1474),
    .Y(_02856_));
 sg13g2_nor2_1 _08409_ (.A(net1823),
    .B(net1728),
    .Y(_02857_));
 sg13g2_a21oi_1 _08410_ (.A1(net1472),
    .A2(_02857_),
    .Y(_00253_),
    .B1(_02856_));
 sg13g2_nor2_1 _08411_ (.A(net1819),
    .B(net530),
    .Y(_02858_));
 sg13g2_a21oi_1 _08412_ (.A1(net1770),
    .A2(net1819),
    .Y(_00254_),
    .B1(_02858_));
 sg13g2_mux2_1 _08413_ (.A0(net532),
    .A1(net1851),
    .S(net1819),
    .X(_00255_));
 sg13g2_nor2_1 _08414_ (.A(net1819),
    .B(net514),
    .Y(_02859_));
 sg13g2_a21oi_1 _08415_ (.A1(net1772),
    .A2(net1819),
    .Y(_00256_),
    .B1(_02859_));
 sg13g2_mux2_1 _08416_ (.A0(net664),
    .A1(net1848),
    .S(net1819),
    .X(_00257_));
 sg13g2_mux2_1 _08417_ (.A0(net517),
    .A1(net1845),
    .S(net1820),
    .X(_00258_));
 sg13g2_mux2_1 _08418_ (.A0(net620),
    .A1(net1842),
    .S(net1819),
    .X(_00259_));
 sg13g2_mux2_1 _08419_ (.A0(net594),
    .A1(net1839),
    .S(net1819),
    .X(_00260_));
 sg13g2_mux2_1 _08420_ (.A0(net766),
    .A1(net1836),
    .S(net1820),
    .X(_00261_));
 sg13g2_nor2_1 _08421_ (.A(net1822),
    .B(net655),
    .Y(_02860_));
 sg13g2_a21oi_1 _08422_ (.A1(_00644_),
    .A2(net1822),
    .Y(_00262_),
    .B1(net656));
 sg13g2_nor2_1 _08423_ (.A(net1821),
    .B(net604),
    .Y(_02861_));
 sg13g2_a21oi_1 _08424_ (.A1(net1773),
    .A2(net1821),
    .Y(_00263_),
    .B1(_02861_));
 sg13g2_nor2_1 _08425_ (.A(net1821),
    .B(net617),
    .Y(_02862_));
 sg13g2_a21oi_1 _08426_ (.A1(net1775),
    .A2(net1821),
    .Y(_00264_),
    .B1(_02862_));
 sg13g2_nor2_1 _08427_ (.A(net1820),
    .B(net611),
    .Y(_02863_));
 sg13g2_a21oi_1 _08428_ (.A1(net1778),
    .A2(net1820),
    .Y(_00265_),
    .B1(_02863_));
 sg13g2_nor2_1 _08429_ (.A(net1820),
    .B(net518),
    .Y(_02864_));
 sg13g2_a21oi_1 _08430_ (.A1(net1780),
    .A2(net1820),
    .Y(_00266_),
    .B1(_02864_));
 sg13g2_nor2_1 _08431_ (.A(net1821),
    .B(net500),
    .Y(_02865_));
 sg13g2_a21oi_1 _08432_ (.A1(net1781),
    .A2(net1821),
    .Y(_00267_),
    .B1(_02865_));
 sg13g2_nor2_1 _08433_ (.A(net1822),
    .B(net599),
    .Y(_02866_));
 sg13g2_a21oi_1 _08434_ (.A1(net1784),
    .A2(net1822),
    .Y(_00268_),
    .B1(net600));
 sg13g2_mux2_1 _08435_ (.A0(net639),
    .A1(net1826),
    .S(net1822),
    .X(_00269_));
 sg13g2_nor2_1 _08436_ (.A(\u_tiny_nn_top.state_q[15] ),
    .B(net1792),
    .Y(_02867_));
 sg13g2_nand2_1 _08437_ (.Y(_02868_),
    .A(net1761),
    .B(_02867_));
 sg13g2_nand2b_2 _08438_ (.Y(_02869_),
    .B(_01180_),
    .A_N(_02868_));
 sg13g2_nand2_1 _08439_ (.Y(_02870_),
    .A(net1764),
    .B(_02869_));
 sg13g2_nand2_1 _08440_ (.Y(_02871_),
    .A(net688),
    .B(net1660));
 sg13g2_o21ai_1 _08441_ (.B1(_02871_),
    .Y(_00270_),
    .A1(_02310_),
    .A2(net1661));
 sg13g2_nand2_1 _08442_ (.Y(_02872_),
    .A(net719),
    .B(net1659));
 sg13g2_o21ai_1 _08443_ (.B1(_02872_),
    .Y(_00271_),
    .A1(_02351_),
    .A2(net1659));
 sg13g2_nand2_1 _08444_ (.Y(_02873_),
    .A(net531),
    .B(net1659));
 sg13g2_o21ai_1 _08445_ (.B1(_02873_),
    .Y(_00272_),
    .A1(_02384_),
    .A2(net1659));
 sg13g2_nand2_1 _08446_ (.Y(_02874_),
    .A(net610),
    .B(net1659));
 sg13g2_o21ai_1 _08447_ (.B1(_02874_),
    .Y(_00273_),
    .A1(_02422_),
    .A2(net1659));
 sg13g2_nand2_1 _08448_ (.Y(_02875_),
    .A(net696),
    .B(net1659));
 sg13g2_o21ai_1 _08449_ (.B1(_02875_),
    .Y(_00274_),
    .A1(_02466_),
    .A2(net1659));
 sg13g2_nand2_1 _08450_ (.Y(_02876_),
    .A(net515),
    .B(net1660));
 sg13g2_o21ai_1 _08451_ (.B1(_02876_),
    .Y(_00275_),
    .A1(_02509_),
    .A2(net1660));
 sg13g2_nand2_1 _08452_ (.Y(_02877_),
    .A(net957),
    .B(net1661));
 sg13g2_o21ai_1 _08453_ (.B1(_02877_),
    .Y(_00276_),
    .A1(_02547_),
    .A2(net1661));
 sg13g2_nand2_1 _08454_ (.Y(_02878_),
    .A(net1050),
    .B(net1662));
 sg13g2_o21ai_1 _08455_ (.B1(_02878_),
    .Y(_00277_),
    .A1(_02572_),
    .A2(net1662));
 sg13g2_nand2_1 _08456_ (.Y(_02879_),
    .A(net991),
    .B(net1662));
 sg13g2_o21ai_1 _08457_ (.B1(_02879_),
    .Y(_00278_),
    .A1(_02613_),
    .A2(net1663));
 sg13g2_nand2_1 _08458_ (.Y(_02880_),
    .A(net1076),
    .B(net1662));
 sg13g2_o21ai_1 _08459_ (.B1(_02880_),
    .Y(_00279_),
    .A1(_02626_),
    .A2(net1662));
 sg13g2_nor2_1 _08460_ (.A(_02688_),
    .B(net1662),
    .Y(_02881_));
 sg13g2_a21oi_1 _08461_ (.A1(_00769_),
    .A2(net1662),
    .Y(_00280_),
    .B1(_02881_));
 sg13g2_mux2_1 _08462_ (.A0(_02710_),
    .A1(net1078),
    .S(net1661),
    .X(_00281_));
 sg13g2_nor2_1 _08463_ (.A(_02743_),
    .B(net1661),
    .Y(_02882_));
 sg13g2_a21oi_1 _08464_ (.A1(_00770_),
    .A2(net1661),
    .Y(_00282_),
    .B1(_02882_));
 sg13g2_nand2_1 _08465_ (.Y(_02883_),
    .A(net1787),
    .B(net1661));
 sg13g2_o21ai_1 _08466_ (.B1(_02883_),
    .Y(_00283_),
    .A1(_02773_),
    .A2(net1661));
 sg13g2_mux2_1 _08467_ (.A0(_02800_),
    .A1(net1074),
    .S(net1662),
    .X(_00284_));
 sg13g2_mux2_1 _08468_ (.A0(_02318_),
    .A1(net1046),
    .S(net1660),
    .X(_00285_));
 sg13g2_nor2_1 _08469_ (.A(net1766),
    .B(_02869_),
    .Y(_02884_));
 sg13g2_nor2_1 _08470_ (.A(net972),
    .B(net1654),
    .Y(_02885_));
 sg13g2_a21oi_1 _08471_ (.A1(_02310_),
    .A2(net1654),
    .Y(_00286_),
    .B1(_02885_));
 sg13g2_nor2_1 _08472_ (.A(net876),
    .B(net1655),
    .Y(_02886_));
 sg13g2_a21oi_1 _08473_ (.A1(_02351_),
    .A2(net1655),
    .Y(_00287_),
    .B1(_02886_));
 sg13g2_nor2_1 _08474_ (.A(net855),
    .B(net1656),
    .Y(_02887_));
 sg13g2_a21oi_1 _08475_ (.A1(_02384_),
    .A2(net1655),
    .Y(_00288_),
    .B1(_02887_));
 sg13g2_nor2_1 _08476_ (.A(net802),
    .B(net1656),
    .Y(_02888_));
 sg13g2_a21oi_1 _08477_ (.A1(_02422_),
    .A2(net1656),
    .Y(_00289_),
    .B1(_02888_));
 sg13g2_nor2_1 _08478_ (.A(net805),
    .B(net1655),
    .Y(_02889_));
 sg13g2_a21oi_1 _08479_ (.A1(_02466_),
    .A2(net1655),
    .Y(_00290_),
    .B1(_02889_));
 sg13g2_nor2_1 _08480_ (.A(net768),
    .B(net1655),
    .Y(_02890_));
 sg13g2_a21oi_1 _08481_ (.A1(_02509_),
    .A2(net1655),
    .Y(_00291_),
    .B1(_02890_));
 sg13g2_nor2_1 _08482_ (.A(net763),
    .B(net1656),
    .Y(_02891_));
 sg13g2_a21oi_1 _08483_ (.A1(_02547_),
    .A2(net1655),
    .Y(_00292_),
    .B1(_02891_));
 sg13g2_nor2_1 _08484_ (.A(net1068),
    .B(net1658),
    .Y(_02892_));
 sg13g2_a21oi_1 _08485_ (.A1(_02572_),
    .A2(net1658),
    .Y(_00293_),
    .B1(_02892_));
 sg13g2_nor2_1 _08486_ (.A(net1038),
    .B(net1658),
    .Y(_02893_));
 sg13g2_a21oi_1 _08487_ (.A1(_02613_),
    .A2(net1658),
    .Y(_00294_),
    .B1(_02893_));
 sg13g2_nor2_1 _08488_ (.A(net1082),
    .B(net1658),
    .Y(_02894_));
 sg13g2_a21oi_1 _08489_ (.A1(_02626_),
    .A2(net1658),
    .Y(_00295_),
    .B1(_02894_));
 sg13g2_mux2_1 _08490_ (.A0(net1090),
    .A1(_02688_),
    .S(net1658),
    .X(_00296_));
 sg13g2_nand2_1 _08491_ (.Y(_02895_),
    .A(_02710_),
    .B(net1654));
 sg13g2_o21ai_1 _08492_ (.B1(_02895_),
    .Y(_00297_),
    .A1(_00762_),
    .A2(net1654));
 sg13g2_nand2_1 _08493_ (.Y(_02896_),
    .A(_02743_),
    .B(net1654));
 sg13g2_o21ai_1 _08494_ (.B1(_02896_),
    .Y(_00298_),
    .A1(_00761_),
    .A2(net1654));
 sg13g2_nor2_1 _08495_ (.A(net1036),
    .B(net1654),
    .Y(_02897_));
 sg13g2_a21oi_1 _08496_ (.A1(_02773_),
    .A2(net1654),
    .Y(_00299_),
    .B1(_02897_));
 sg13g2_mux2_1 _08497_ (.A0(net1037),
    .A1(_02800_),
    .S(net1657),
    .X(_00300_));
 sg13g2_mux2_1 _08498_ (.A0(net998),
    .A1(_02318_),
    .S(net1657),
    .X(_00301_));
 sg13g2_a21oi_1 _08499_ (.A1(net1854),
    .A2(net1792),
    .Y(_02898_),
    .B1(net1789));
 sg13g2_a22oi_1 _08500_ (.Y(_02899_),
    .B1(_02898_),
    .B2(_01045_),
    .A2(_01205_),
    .A1(_00161_));
 sg13g2_nor3_1 _08501_ (.A(\u_tiny_nn_top.state_q[15] ),
    .B(net1764),
    .C(_02899_),
    .Y(_02900_));
 sg13g2_mux2_1 _08502_ (.A0(_01623_),
    .A1(net1018),
    .S(net1651),
    .X(_00302_));
 sg13g2_mux2_1 _08503_ (.A0(_02330_),
    .A1(net1007),
    .S(net1651),
    .X(_00303_));
 sg13g2_mux2_1 _08504_ (.A0(_02363_),
    .A1(net1014),
    .S(net1651),
    .X(_00304_));
 sg13g2_mux2_1 _08505_ (.A0(_02399_),
    .A1(net1019),
    .S(net1651),
    .X(_00305_));
 sg13g2_mux2_1 _08506_ (.A0(_02438_),
    .A1(net1042),
    .S(net1651),
    .X(_00306_));
 sg13g2_mux2_1 _08507_ (.A0(_02484_),
    .A1(net1070),
    .S(net1651),
    .X(_00307_));
 sg13g2_mux2_1 _08508_ (.A0(_02521_),
    .A1(net1057),
    .S(net1652),
    .X(_00308_));
 sg13g2_nor2_1 _08509_ (.A(_02554_),
    .B(net1652),
    .Y(_02901_));
 sg13g2_a21oi_1 _08510_ (.A1(_00676_),
    .A2(net1652),
    .Y(_00309_),
    .B1(_02901_));
 sg13g2_mux2_1 _08511_ (.A0(_02586_),
    .A1(net1105),
    .S(net1653),
    .X(_00310_));
 sg13g2_nor2_1 _08512_ (.A(_02640_),
    .B(net1652),
    .Y(_02902_));
 sg13g2_a21oi_1 _08513_ (.A1(_00677_),
    .A2(net1652),
    .Y(_00311_),
    .B1(_02902_));
 sg13g2_mux2_1 _08514_ (.A0(_02668_),
    .A1(net1786),
    .S(net1652),
    .X(_00312_));
 sg13g2_mux2_1 _08515_ (.A0(_02694_),
    .A1(net1072),
    .S(net1652),
    .X(_00313_));
 sg13g2_nand2_1 _08516_ (.Y(_02903_),
    .A(net1043),
    .B(net1653));
 sg13g2_o21ai_1 _08517_ (.B1(_02903_),
    .Y(_00314_),
    .A1(_02722_),
    .A2(net1653));
 sg13g2_nand2_1 _08518_ (.Y(_02904_),
    .A(net1029),
    .B(net1653));
 sg13g2_o21ai_1 _08519_ (.B1(_02904_),
    .Y(_00315_),
    .A1(_02755_),
    .A2(net1653));
 sg13g2_nand2_1 _08520_ (.Y(_02905_),
    .A(net1077),
    .B(net1653));
 sg13g2_o21ai_1 _08521_ (.B1(_02905_),
    .Y(_00316_),
    .A1(_02791_),
    .A2(net1653));
 sg13g2_nand2_1 _08522_ (.Y(_02906_),
    .A(net1087),
    .B(net1651));
 sg13g2_o21ai_1 _08523_ (.B1(_02906_),
    .Y(_00317_),
    .A1(_02809_),
    .A2(net1651));
 sg13g2_a21oi_2 _08524_ (.B1(\u_tiny_nn_top.state_q[16] ),
    .Y(_02907_),
    .A2(_01032_),
    .A1(_00826_));
 sg13g2_nand2_1 _08525_ (.Y(_02908_),
    .A(_00163_),
    .B(net1765));
 sg13g2_a21oi_2 _08526_ (.B1(_02908_),
    .Y(_02909_),
    .A2(_01057_),
    .A1(_00957_));
 sg13g2_and2_1 _08527_ (.A(_02907_),
    .B(net1650),
    .X(_02910_));
 sg13g2_nor2b_2 _08528_ (.A(net1650),
    .B_N(_02907_),
    .Y(_02911_));
 sg13g2_nand2b_1 _08529_ (.Y(_02912_),
    .B(_02907_),
    .A_N(net1650));
 sg13g2_nand3_1 _08530_ (.B(net1765),
    .C(_02867_),
    .A(_00036_),
    .Y(_02913_));
 sg13g2_o21ai_1 _08531_ (.B1(_02913_),
    .Y(_02914_),
    .A1(_01179_),
    .A2(_02868_));
 sg13g2_nand2b_1 _08532_ (.Y(_02915_),
    .B(net1689),
    .A_N(\u_tiny_nn_top.u_core.mul_val_op_q[5][2] ));
 sg13g2_mux2_1 _08533_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][2] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][2] ),
    .S(net1690),
    .X(_02916_));
 sg13g2_o21ai_1 _08534_ (.B1(_02915_),
    .Y(_02917_),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[4][2] ),
    .A2(net1690));
 sg13g2_mux2_1 _08535_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][6] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][6] ),
    .S(net1695),
    .X(_02918_));
 sg13g2_mux2_1 _08536_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][1] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][1] ),
    .S(net1689),
    .X(_02919_));
 sg13g2_nor3_1 _08537_ (.A(net1643),
    .B(net1641),
    .C(net1639),
    .Y(_02920_));
 sg13g2_mux2_1 _08538_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][3] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][3] ),
    .S(net1694),
    .X(_02921_));
 sg13g2_mux2_1 _08539_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][4] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][4] ),
    .S(net1694),
    .X(_02922_));
 sg13g2_mux2_1 _08540_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][5] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][5] ),
    .S(net1689),
    .X(_02923_));
 sg13g2_nand2b_1 _08541_ (.Y(_02924_),
    .B(net1689),
    .A_N(\u_tiny_nn_top.u_core.mul_val_op_q[5][0] ));
 sg13g2_mux2_1 _08542_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][0] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][0] ),
    .S(net1689),
    .X(_02925_));
 sg13g2_o21ai_1 _08543_ (.B1(_02924_),
    .Y(_02926_),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[4][0] ),
    .A2(net1689));
 sg13g2_nor4_1 _08544_ (.A(net1636),
    .B(net1633),
    .C(net1631),
    .D(net1630),
    .Y(_02927_));
 sg13g2_nand2_2 _08545_ (.Y(_02928_),
    .A(_02920_),
    .B(_02927_));
 sg13g2_inv_1 _08546_ (.Y(_02929_),
    .A(_02928_));
 sg13g2_mux2_2 _08547_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][15] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][15] ),
    .S(net1715),
    .X(_02930_));
 sg13g2_nor2_1 _08548_ (.A(_02928_),
    .B(_02930_),
    .Y(_02931_));
 sg13g2_mux2_2 _08549_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][12] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][12] ),
    .S(net1696),
    .X(_02932_));
 sg13g2_mux2_2 _08550_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][11] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][11] ),
    .S(net1696),
    .X(_02933_));
 sg13g2_mux2_1 _08551_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][9] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][9] ),
    .S(net1696),
    .X(_02934_));
 sg13g2_mux2_2 _08552_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][7] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][7] ),
    .S(net1696),
    .X(_02935_));
 sg13g2_mux2_2 _08553_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][10] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][10] ),
    .S(net1698),
    .X(_02936_));
 sg13g2_mux2_2 _08554_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][13] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][13] ),
    .S(net1703),
    .X(_02937_));
 sg13g2_mux2_2 _08555_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][8] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][8] ),
    .S(net1703),
    .X(_02938_));
 sg13g2_mux2_2 _08556_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][14] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][14] ),
    .S(net1703),
    .X(_02939_));
 sg13g2_nor4_1 _08557_ (.A(_02932_),
    .B(_02933_),
    .C(_02936_),
    .D(_02937_),
    .Y(_02940_));
 sg13g2_nor4_1 _08558_ (.A(_02934_),
    .B(_02935_),
    .C(_02938_),
    .D(_02939_),
    .Y(_02941_));
 sg13g2_nand2_1 _08559_ (.Y(_02942_),
    .A(_00053_),
    .B(net1693));
 sg13g2_mux2_1 _08560_ (.A0(_00691_),
    .A1(_00692_),
    .S(net1693),
    .X(_02943_));
 sg13g2_o21ai_1 _08561_ (.B1(_02942_),
    .Y(_02944_),
    .A1(_00691_),
    .A2(net1693));
 sg13g2_nand2b_1 _08562_ (.Y(_02945_),
    .B(net1693),
    .A_N(_00051_));
 sg13g2_o21ai_1 _08563_ (.B1(_02945_),
    .Y(_02946_),
    .A1(_00052_),
    .A2(net1692));
 sg13g2_mux2_1 _08564_ (.A0(_00052_),
    .A1(_00051_),
    .S(net1692),
    .X(_02947_));
 sg13g2_mux2_1 _08565_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[4][6] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[5][6] ),
    .S(net1692),
    .X(_02948_));
 sg13g2_nand2b_1 _08566_ (.Y(_02949_),
    .B(net1692),
    .A_N(\u_tiny_nn_top.u_core.param_val_op_q[5][2] ));
 sg13g2_mux2_1 _08567_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[4][2] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[5][2] ),
    .S(net1692),
    .X(_02950_));
 sg13g2_o21ai_1 _08568_ (.B1(_02949_),
    .Y(_02951_),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[4][2] ),
    .A2(net1692));
 sg13g2_mux2_1 _08569_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[4][0] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[5][0] ),
    .S(net1692),
    .X(_02952_));
 sg13g2_nor2_1 _08570_ (.A(net1624),
    .B(net1622),
    .Y(_02953_));
 sg13g2_mux2_1 _08571_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[4][1] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[5][1] ),
    .S(net1691),
    .X(_02954_));
 sg13g2_mux2_1 _08572_ (.A0(_00693_),
    .A1(_00694_),
    .S(net1692),
    .X(_02955_));
 sg13g2_nor3_1 _08573_ (.A(net1625),
    .B(net1621),
    .C(net1620),
    .Y(_02956_));
 sg13g2_nand4_1 _08574_ (.B(_02947_),
    .C(_02953_),
    .A(_02944_),
    .Y(_02957_),
    .D(_02956_));
 sg13g2_inv_1 _08575_ (.Y(_02958_),
    .A(_02957_));
 sg13g2_mux2_2 _08576_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[4][15] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[5][15] ),
    .S(net1702),
    .X(_02959_));
 sg13g2_nor2_1 _08577_ (.A(_02957_),
    .B(_02959_),
    .Y(_02960_));
 sg13g2_mux2_2 _08578_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[4][12] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[5][12] ),
    .S(net1702),
    .X(_02961_));
 sg13g2_mux2_2 _08579_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[4][9] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[5][9] ),
    .S(net1702),
    .X(_02962_));
 sg13g2_mux2_2 _08580_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[4][11] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[5][11] ),
    .S(net1702),
    .X(_02963_));
 sg13g2_mux2_2 _08581_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[4][14] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[5][14] ),
    .S(net1702),
    .X(_02964_));
 sg13g2_mux2_2 _08582_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[4][13] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[5][13] ),
    .S(net1702),
    .X(_02965_));
 sg13g2_mux2_2 _08583_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[4][8] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[5][8] ),
    .S(net1702),
    .X(_02966_));
 sg13g2_mux2_2 _08584_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[4][10] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[5][10] ),
    .S(net1702),
    .X(_02967_));
 sg13g2_nand2b_1 _08585_ (.Y(_02968_),
    .B(net1697),
    .A_N(\u_tiny_nn_top.u_core.param_val_op_q[5][7] ));
 sg13g2_mux2_1 _08586_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[4][7] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[5][7] ),
    .S(net1697),
    .X(_02969_));
 sg13g2_o21ai_1 _08587_ (.B1(_02968_),
    .Y(_02970_),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[4][7] ),
    .A2(net1697));
 sg13g2_nor4_1 _08588_ (.A(_02961_),
    .B(_02963_),
    .C(_02964_),
    .D(_02967_),
    .Y(_02971_));
 sg13g2_nor4_1 _08589_ (.A(_02962_),
    .B(_02965_),
    .C(_02966_),
    .D(_02969_),
    .Y(_02972_));
 sg13g2_nand4_1 _08590_ (.B(_02963_),
    .C(_02964_),
    .A(_02962_),
    .Y(_02973_),
    .D(_02965_));
 sg13g2_nand4_1 _08591_ (.B(_02966_),
    .C(_02967_),
    .A(_02961_),
    .Y(_02974_),
    .D(_02969_));
 sg13g2_nor2_1 _08592_ (.A(_02973_),
    .B(_02974_),
    .Y(_02975_));
 sg13g2_nand4_1 _08593_ (.B(_02933_),
    .C(_02936_),
    .A(_02932_),
    .Y(_02976_),
    .D(_02937_));
 sg13g2_nand4_1 _08594_ (.B(_02935_),
    .C(_02938_),
    .A(_02934_),
    .Y(_02977_),
    .D(_02939_));
 sg13g2_nor2_1 _08595_ (.A(_02976_),
    .B(_02977_),
    .Y(_02978_));
 sg13g2_a22oi_1 _08596_ (.Y(_02979_),
    .B1(_02975_),
    .B2(_02957_),
    .A2(_02972_),
    .A1(_02971_));
 sg13g2_nor2_1 _08597_ (.A(_02960_),
    .B(_02979_),
    .Y(_02980_));
 sg13g2_a22oi_1 _08598_ (.Y(_02981_),
    .B1(_02978_),
    .B2(_02928_),
    .A2(_02941_),
    .A1(_02940_));
 sg13g2_nor2_1 _08599_ (.A(_02931_),
    .B(_02981_),
    .Y(_02982_));
 sg13g2_nor2_1 _08600_ (.A(_02980_),
    .B(_02982_),
    .Y(_02983_));
 sg13g2_nand2_1 _08601_ (.Y(_02984_),
    .A(_02937_),
    .B(_02965_));
 sg13g2_xnor2_1 _08602_ (.Y(_02985_),
    .A(_02937_),
    .B(_02965_));
 sg13g2_or2_1 _08603_ (.X(_02986_),
    .B(_02961_),
    .A(_02932_));
 sg13g2_nand2_1 _08604_ (.Y(_02987_),
    .A(_02932_),
    .B(_02961_));
 sg13g2_and2_1 _08605_ (.A(_02933_),
    .B(_02963_),
    .X(_02988_));
 sg13g2_xnor2_1 _08606_ (.Y(_02989_),
    .A(_02933_),
    .B(_02963_));
 sg13g2_nor2_1 _08607_ (.A(_02936_),
    .B(_02967_),
    .Y(_02990_));
 sg13g2_and2_1 _08608_ (.A(_02934_),
    .B(_02962_),
    .X(_02991_));
 sg13g2_nand2_1 _08609_ (.Y(_02992_),
    .A(_02938_),
    .B(_02966_));
 sg13g2_nand2_1 _08610_ (.Y(_02993_),
    .A(net1641),
    .B(net1626));
 sg13g2_xor2_1 _08611_ (.B(_02993_),
    .A(net1632),
    .X(_02994_));
 sg13g2_xnor2_1 _08612_ (.Y(_02995_),
    .A(_02944_),
    .B(_02994_));
 sg13g2_nand2_1 _08613_ (.Y(_02996_),
    .A(net1632),
    .B(net1626));
 sg13g2_nand3_1 _08614_ (.B(net1632),
    .C(net1626),
    .A(net1634),
    .Y(_02997_));
 sg13g2_nand2_1 _08615_ (.Y(_02998_),
    .A(net1640),
    .B(net1628));
 sg13g2_xor2_1 _08616_ (.B(_02996_),
    .A(net1634),
    .X(_02999_));
 sg13g2_o21ai_1 _08617_ (.B1(_02997_),
    .Y(_03000_),
    .A1(_02998_),
    .A2(_02999_));
 sg13g2_nand2b_1 _08618_ (.Y(_03001_),
    .B(_03000_),
    .A_N(_02995_));
 sg13g2_xor2_1 _08619_ (.B(net1626),
    .A(net1640),
    .X(_03002_));
 sg13g2_nand2_1 _08620_ (.Y(_03003_),
    .A(net1632),
    .B(net1628));
 sg13g2_nand3_1 _08621_ (.B(net1628),
    .C(_03002_),
    .A(net1632),
    .Y(_03004_));
 sg13g2_nand3_1 _08622_ (.B(_03001_),
    .C(_03004_),
    .A(_02993_),
    .Y(_03005_));
 sg13g2_o21ai_1 _08623_ (.B1(_02996_),
    .Y(_03006_),
    .A1(_02944_),
    .A2(_02994_));
 sg13g2_o21ai_1 _08624_ (.B1(_03004_),
    .Y(_03007_),
    .A1(_03002_),
    .A2(_03006_));
 sg13g2_nand2b_1 _08625_ (.Y(_03008_),
    .B(_03001_),
    .A_N(_03007_));
 sg13g2_xnor2_1 _08626_ (.Y(_03009_),
    .A(_02995_),
    .B(_03000_));
 sg13g2_nand3_1 _08627_ (.B(net1634),
    .C(net1626),
    .A(net1636),
    .Y(_03010_));
 sg13g2_a21o_1 _08628_ (.A2(net1626),
    .A1(net1634),
    .B1(net1635),
    .X(_03011_));
 sg13g2_nand2_1 _08629_ (.Y(_03012_),
    .A(_03010_),
    .B(_03011_));
 sg13g2_o21ai_1 _08630_ (.B1(_03010_),
    .Y(_03013_),
    .A1(_03003_),
    .A2(_03012_));
 sg13g2_xor2_1 _08631_ (.B(_02999_),
    .A(_02998_),
    .X(_03014_));
 sg13g2_and2_1 _08632_ (.A(_03013_),
    .B(_03014_),
    .X(_03015_));
 sg13g2_or2_1 _08633_ (.X(_03016_),
    .B(_03014_),
    .A(_03013_));
 sg13g2_nand2b_1 _08634_ (.Y(_03017_),
    .B(_03016_),
    .A_N(_03015_));
 sg13g2_a21o_1 _08635_ (.A2(_03016_),
    .A1(net1620),
    .B1(_03015_),
    .X(_03018_));
 sg13g2_nand2_1 _08636_ (.Y(_03019_),
    .A(_03009_),
    .B(_03018_));
 sg13g2_or2_1 _08637_ (.X(_03020_),
    .B(_03019_),
    .A(_03008_));
 sg13g2_nand4_1 _08638_ (.B(net1631),
    .C(net1628),
    .A(net1640),
    .Y(_03021_),
    .D(net1626));
 sg13g2_nand2_1 _08639_ (.Y(_03022_),
    .A(_03005_),
    .B(_03021_));
 sg13g2_nor2b_1 _08640_ (.A(_03005_),
    .B_N(_03020_),
    .Y(_03023_));
 sg13g2_xnor2_1 _08641_ (.Y(_03024_),
    .A(net1620),
    .B(_03017_));
 sg13g2_nand3_1 _08642_ (.B(net1635),
    .C(net1625),
    .A(net1642),
    .Y(_03025_));
 sg13g2_nand2_1 _08643_ (.Y(_03026_),
    .A(net1633),
    .B(net1627));
 sg13g2_a21o_1 _08644_ (.A2(net1625),
    .A1(net1635),
    .B1(net1642),
    .X(_03027_));
 sg13g2_nand2_1 _08645_ (.Y(_03028_),
    .A(_03025_),
    .B(_03027_));
 sg13g2_o21ai_1 _08646_ (.B1(_03025_),
    .Y(_03029_),
    .A1(_03026_),
    .A2(_03028_));
 sg13g2_xor2_1 _08647_ (.B(_03012_),
    .A(_03003_),
    .X(_03030_));
 sg13g2_nand2_1 _08648_ (.Y(_03031_),
    .A(_03029_),
    .B(_03030_));
 sg13g2_nand2_1 _08649_ (.Y(_03032_),
    .A(net1640),
    .B(net1620));
 sg13g2_xnor2_1 _08650_ (.Y(_03033_),
    .A(_03029_),
    .B(_03030_));
 sg13g2_o21ai_1 _08651_ (.B1(_03031_),
    .Y(_03034_),
    .A1(_03032_),
    .A2(_03033_));
 sg13g2_nand2_1 _08652_ (.Y(_03035_),
    .A(_03024_),
    .B(_03034_));
 sg13g2_xor2_1 _08653_ (.B(_03018_),
    .A(_03009_),
    .X(_03036_));
 sg13g2_nand2b_1 _08654_ (.Y(_03037_),
    .B(_03036_),
    .A_N(_03035_));
 sg13g2_nor2_1 _08655_ (.A(_03008_),
    .B(_03037_),
    .Y(_03038_));
 sg13g2_xor2_1 _08656_ (.B(_03034_),
    .A(_03024_),
    .X(_03039_));
 sg13g2_nand3_1 _08657_ (.B(net1638),
    .C(net1625),
    .A(net1643),
    .Y(_03040_));
 sg13g2_nand2_1 _08658_ (.Y(_03041_),
    .A(net1635),
    .B(net1627));
 sg13g2_a21o_1 _08659_ (.A2(net1625),
    .A1(net1643),
    .B1(net1638),
    .X(_03042_));
 sg13g2_nand2_1 _08660_ (.Y(_03043_),
    .A(_03040_),
    .B(_03042_));
 sg13g2_o21ai_1 _08661_ (.B1(_03040_),
    .Y(_03044_),
    .A1(_03041_),
    .A2(_03043_));
 sg13g2_xor2_1 _08662_ (.B(_03028_),
    .A(_03026_),
    .X(_03045_));
 sg13g2_nand2_1 _08663_ (.Y(_03046_),
    .A(_03044_),
    .B(_03045_));
 sg13g2_nand2_1 _08664_ (.Y(_03047_),
    .A(net1631),
    .B(net1620));
 sg13g2_xnor2_1 _08665_ (.Y(_03048_),
    .A(_03044_),
    .B(_03045_));
 sg13g2_o21ai_1 _08666_ (.B1(_03046_),
    .Y(_03049_),
    .A1(_03047_),
    .A2(_03048_));
 sg13g2_xor2_1 _08667_ (.B(_03033_),
    .A(_03032_),
    .X(_03050_));
 sg13g2_nand2_1 _08668_ (.Y(_03051_),
    .A(_03049_),
    .B(_03050_));
 sg13g2_xnor2_1 _08669_ (.Y(_03052_),
    .A(_03049_),
    .B(_03050_));
 sg13g2_o21ai_1 _08670_ (.B1(_03051_),
    .Y(_03053_),
    .A1(_02947_),
    .A2(_03052_));
 sg13g2_nand2_1 _08671_ (.Y(_03054_),
    .A(_03039_),
    .B(_03053_));
 sg13g2_nand3_1 _08672_ (.B(_03039_),
    .C(_03053_),
    .A(_03036_),
    .Y(_03055_));
 sg13g2_xor2_1 _08673_ (.B(_03053_),
    .A(_03039_),
    .X(_03056_));
 sg13g2_and2_1 _08674_ (.A(net1629),
    .B(net1625),
    .X(_03057_));
 sg13g2_nand3_1 _08675_ (.B(net1629),
    .C(net1625),
    .A(net1637),
    .Y(_03058_));
 sg13g2_a21o_1 _08676_ (.A2(net1625),
    .A1(net1637),
    .B1(net1629),
    .X(_03059_));
 sg13g2_and4_1 _08677_ (.A(net1643),
    .B(net1627),
    .C(_03058_),
    .D(_03059_),
    .X(_03060_));
 sg13g2_a21o_1 _08678_ (.A2(_03057_),
    .A1(net1638),
    .B1(_03060_),
    .X(_03061_));
 sg13g2_xor2_1 _08679_ (.B(_03043_),
    .A(_03041_),
    .X(_03062_));
 sg13g2_nand2_1 _08680_ (.Y(_03063_),
    .A(_03061_),
    .B(_03062_));
 sg13g2_xnor2_1 _08681_ (.Y(_03064_),
    .A(_03061_),
    .B(_03062_));
 sg13g2_nand2_1 _08682_ (.Y(_03065_),
    .A(net1633),
    .B(net1621));
 sg13g2_nand3_1 _08683_ (.B(_02954_),
    .C(net1619),
    .A(net1634),
    .Y(_03066_));
 sg13g2_a21o_1 _08684_ (.A2(net1619),
    .A1(net1634),
    .B1(net1621),
    .X(_03067_));
 sg13g2_nand2_1 _08685_ (.Y(_03068_),
    .A(_03066_),
    .B(_03067_));
 sg13g2_o21ai_1 _08686_ (.B1(_03063_),
    .Y(_03069_),
    .A1(_03064_),
    .A2(_03068_));
 sg13g2_xor2_1 _08687_ (.B(_03048_),
    .A(_03047_),
    .X(_03070_));
 sg13g2_nand2_1 _08688_ (.Y(_03071_),
    .A(_03069_),
    .B(_03070_));
 sg13g2_or2_1 _08689_ (.X(_03072_),
    .B(_03066_),
    .A(_02951_));
 sg13g2_xnor2_1 _08690_ (.Y(_03073_),
    .A(_02951_),
    .B(_03066_));
 sg13g2_nand2_1 _08691_ (.Y(_03074_),
    .A(net1641),
    .B(_02946_));
 sg13g2_xnor2_1 _08692_ (.Y(_03075_),
    .A(_03073_),
    .B(_03074_));
 sg13g2_xnor2_1 _08693_ (.Y(_03076_),
    .A(_03069_),
    .B(_03070_));
 sg13g2_o21ai_1 _08694_ (.B1(_03071_),
    .Y(_03077_),
    .A1(_03075_),
    .A2(_03076_));
 sg13g2_xnor2_1 _08695_ (.Y(_03078_),
    .A(_02946_),
    .B(_03052_));
 sg13g2_o21ai_1 _08696_ (.B1(_03072_),
    .Y(_03079_),
    .A1(_03073_),
    .A2(_03074_));
 sg13g2_xnor2_1 _08697_ (.Y(_03080_),
    .A(_03077_),
    .B(_03078_));
 sg13g2_nor2b_1 _08698_ (.A(_03080_),
    .B_N(_03079_),
    .Y(_03081_));
 sg13g2_a21o_1 _08699_ (.A2(_03078_),
    .A1(_03077_),
    .B1(_03081_),
    .X(_03082_));
 sg13g2_and2_1 _08700_ (.A(_03056_),
    .B(_03082_),
    .X(_03083_));
 sg13g2_nand2_1 _08701_ (.Y(_03084_),
    .A(net1630),
    .B(net1627));
 sg13g2_and3_1 _08702_ (.X(_03085_),
    .A(net1629),
    .B(net1627),
    .C(_02948_));
 sg13g2_nand2_1 _08703_ (.Y(_03086_),
    .A(net1638),
    .B(_03085_));
 sg13g2_a22oi_1 _08704_ (.Y(_03087_),
    .B1(_03058_),
    .B2(_03059_),
    .A2(net1627),
    .A1(net1642));
 sg13g2_or3_1 _08705_ (.A(_03060_),
    .B(_03086_),
    .C(_03087_),
    .X(_03088_));
 sg13g2_o21ai_1 _08706_ (.B1(_03086_),
    .Y(_03089_),
    .A1(_03060_),
    .A2(_03087_));
 sg13g2_nand2_1 _08707_ (.Y(_03090_),
    .A(net1640),
    .B(net1621));
 sg13g2_and2_1 _08708_ (.A(net1635),
    .B(net1622),
    .X(_03091_));
 sg13g2_nand2_1 _08709_ (.Y(_03092_),
    .A(net1618),
    .B(_03091_));
 sg13g2_a21oi_1 _08710_ (.A1(net1635),
    .A2(net1618),
    .Y(_03093_),
    .B1(net1622));
 sg13g2_a21o_1 _08711_ (.A2(_03091_),
    .A1(net1618),
    .B1(_03093_),
    .X(_03094_));
 sg13g2_xor2_1 _08712_ (.B(_03094_),
    .A(_03090_),
    .X(_03095_));
 sg13g2_nand3_1 _08713_ (.B(_03089_),
    .C(_03095_),
    .A(_03088_),
    .Y(_03096_));
 sg13g2_and2_1 _08714_ (.A(_03088_),
    .B(_03096_),
    .X(_03097_));
 sg13g2_xor2_1 _08715_ (.B(_03068_),
    .A(_03064_),
    .X(_03098_));
 sg13g2_nor2b_1 _08716_ (.A(_03097_),
    .B_N(_03098_),
    .Y(_03099_));
 sg13g2_xnor2_1 _08717_ (.Y(_03100_),
    .A(_03097_),
    .B(_03098_));
 sg13g2_nand2_1 _08718_ (.Y(_03101_),
    .A(net1632),
    .B(_02946_));
 sg13g2_o21ai_1 _08719_ (.B1(_03092_),
    .Y(_03102_),
    .A1(_03090_),
    .A2(_03094_));
 sg13g2_nand2_1 _08720_ (.Y(_03103_),
    .A(net1640),
    .B(_02950_));
 sg13g2_nand2b_1 _08721_ (.Y(_03104_),
    .B(_03102_),
    .A_N(_03103_));
 sg13g2_xor2_1 _08722_ (.B(_03103_),
    .A(_03102_),
    .X(_03105_));
 sg13g2_xor2_1 _08723_ (.B(_03105_),
    .A(_03101_),
    .X(_03106_));
 sg13g2_a21o_1 _08724_ (.A2(_03106_),
    .A1(_03100_),
    .B1(_03099_),
    .X(_03107_));
 sg13g2_xnor2_1 _08725_ (.Y(_03108_),
    .A(_03075_),
    .B(_03076_));
 sg13g2_nand2b_1 _08726_ (.Y(_03109_),
    .B(_03107_),
    .A_N(_03108_));
 sg13g2_o21ai_1 _08727_ (.B1(_03104_),
    .Y(_03110_),
    .A1(_03101_),
    .A2(_03105_));
 sg13g2_inv_1 _08728_ (.Y(_03111_),
    .A(_03110_));
 sg13g2_xor2_1 _08729_ (.B(_03108_),
    .A(_03107_),
    .X(_03112_));
 sg13g2_o21ai_1 _08730_ (.B1(_03109_),
    .Y(_03113_),
    .A1(_03111_),
    .A2(_03112_));
 sg13g2_xor2_1 _08731_ (.B(_03080_),
    .A(_03079_),
    .X(_03114_));
 sg13g2_nand2b_1 _08732_ (.Y(_03115_),
    .B(_03113_),
    .A_N(_03114_));
 sg13g2_nand2_1 _08733_ (.Y(_03116_),
    .A(net1631),
    .B(net1621));
 sg13g2_nand2_1 _08734_ (.Y(_03117_),
    .A(net1642),
    .B(net1622));
 sg13g2_and4_1 _08735_ (.A(net1642),
    .B(net1640),
    .C(net1623),
    .D(net1618),
    .X(_03118_));
 sg13g2_a22oi_1 _08736_ (.Y(_03119_),
    .B1(net1618),
    .B2(net1643),
    .A2(net1623),
    .A1(net1640));
 sg13g2_o21ai_1 _08737_ (.B1(_03116_),
    .Y(_03120_),
    .A1(_03118_),
    .A2(_03119_));
 sg13g2_or3_1 _08738_ (.A(_03116_),
    .B(_03118_),
    .C(_03119_),
    .X(_03121_));
 sg13g2_a22oi_1 _08739_ (.Y(_03122_),
    .B1(_02948_),
    .B2(net1630),
    .A2(net1627),
    .A1(net1638));
 sg13g2_a21oi_1 _08740_ (.A1(net1637),
    .A2(_03085_),
    .Y(_03123_),
    .B1(_03122_));
 sg13g2_and3_1 _08741_ (.X(_03124_),
    .A(_03120_),
    .B(_03121_),
    .C(_03123_));
 sg13g2_a21o_1 _08742_ (.A2(_03089_),
    .A1(_03088_),
    .B1(_03095_),
    .X(_03125_));
 sg13g2_nand3_1 _08743_ (.B(_03124_),
    .C(_03125_),
    .A(_03096_),
    .Y(_03126_));
 sg13g2_a21o_1 _08744_ (.A2(_03125_),
    .A1(_03096_),
    .B1(_03124_),
    .X(_03127_));
 sg13g2_and2_1 _08745_ (.A(net1633),
    .B(_02946_),
    .X(_03128_));
 sg13g2_nor2b_1 _08746_ (.A(_03118_),
    .B_N(_03121_),
    .Y(_03129_));
 sg13g2_nand2_1 _08747_ (.Y(_03130_),
    .A(net1631),
    .B(net1624));
 sg13g2_xor2_1 _08748_ (.B(_03130_),
    .A(_03129_),
    .X(_03131_));
 sg13g2_nand2_1 _08749_ (.Y(_03132_),
    .A(_03128_),
    .B(_03131_));
 sg13g2_xor2_1 _08750_ (.B(_03131_),
    .A(_03128_),
    .X(_03133_));
 sg13g2_and3_1 _08751_ (.X(_03134_),
    .A(_03126_),
    .B(_03127_),
    .C(_03133_));
 sg13g2_nand3_1 _08752_ (.B(_03127_),
    .C(_03133_),
    .A(_03126_),
    .Y(_03135_));
 sg13g2_and2_1 _08753_ (.A(_03126_),
    .B(_03135_),
    .X(_03136_));
 sg13g2_xnor2_1 _08754_ (.Y(_03137_),
    .A(_03100_),
    .B(_03106_));
 sg13g2_nor2_1 _08755_ (.A(_03136_),
    .B(_03137_),
    .Y(_03138_));
 sg13g2_o21ai_1 _08756_ (.B1(_03132_),
    .Y(_03139_),
    .A1(_03129_),
    .A2(_03130_));
 sg13g2_xor2_1 _08757_ (.B(_03137_),
    .A(_03136_),
    .X(_03140_));
 sg13g2_a21oi_1 _08758_ (.A1(_03139_),
    .A2(_03140_),
    .Y(_03141_),
    .B1(_03138_));
 sg13g2_xnor2_1 _08759_ (.Y(_03142_),
    .A(_03111_),
    .B(_03112_));
 sg13g2_nor2_1 _08760_ (.A(_03141_),
    .B(_03142_),
    .Y(_03143_));
 sg13g2_a21oi_1 _08761_ (.A1(_03120_),
    .A2(_03121_),
    .Y(_03144_),
    .B1(_03123_));
 sg13g2_and4_1 _08762_ (.A(net1637),
    .B(net1631),
    .C(net1623),
    .D(net1619),
    .X(_03145_));
 sg13g2_nand4_1 _08763_ (.B(net1631),
    .C(net1623),
    .A(net1639),
    .Y(_03146_),
    .D(net1619));
 sg13g2_a22oi_1 _08764_ (.Y(_03147_),
    .B1(net1619),
    .B2(net1637),
    .A2(net1623),
    .A1(net1631));
 sg13g2_o21ai_1 _08765_ (.B1(_03065_),
    .Y(_03148_),
    .A1(_03145_),
    .A2(_03147_));
 sg13g2_or3_1 _08766_ (.A(_03065_),
    .B(_03145_),
    .C(_03147_),
    .X(_03149_));
 sg13g2_and2_1 _08767_ (.A(_03148_),
    .B(_03149_),
    .X(_03150_));
 sg13g2_nand4_1 _08768_ (.B(net1627),
    .C(_03148_),
    .A(net1630),
    .Y(_03151_),
    .D(_03149_));
 sg13g2_or3_1 _08769_ (.A(_03124_),
    .B(_03144_),
    .C(_03151_),
    .X(_03152_));
 sg13g2_o21ai_1 _08770_ (.B1(_03151_),
    .Y(_03153_),
    .A1(_03124_),
    .A2(_03144_));
 sg13g2_and2_1 _08771_ (.A(net1636),
    .B(_02946_),
    .X(_03154_));
 sg13g2_o21ai_1 _08772_ (.B1(_03146_),
    .Y(_03155_),
    .A1(_03065_),
    .A2(_03147_));
 sg13g2_nand2_1 _08773_ (.Y(_03156_),
    .A(net1633),
    .B(net1624));
 sg13g2_nand2b_1 _08774_ (.Y(_03157_),
    .B(_03155_),
    .A_N(_03156_));
 sg13g2_xnor2_1 _08775_ (.Y(_03158_),
    .A(_03155_),
    .B(_03156_));
 sg13g2_nand2_1 _08776_ (.Y(_03159_),
    .A(_03154_),
    .B(_03158_));
 sg13g2_xor2_1 _08777_ (.B(_03158_),
    .A(_03154_),
    .X(_03160_));
 sg13g2_nand3_1 _08778_ (.B(_03153_),
    .C(_03160_),
    .A(_03152_),
    .Y(_03161_));
 sg13g2_and2_1 _08779_ (.A(_03152_),
    .B(_03161_),
    .X(_03162_));
 sg13g2_a21oi_1 _08780_ (.A1(_03126_),
    .A2(_03127_),
    .Y(_03163_),
    .B1(_03133_));
 sg13g2_nor3_1 _08781_ (.A(_03134_),
    .B(_03162_),
    .C(_03163_),
    .Y(_03164_));
 sg13g2_or3_1 _08782_ (.A(_03134_),
    .B(_03162_),
    .C(_03163_),
    .X(_03165_));
 sg13g2_nand2_1 _08783_ (.Y(_03166_),
    .A(_03157_),
    .B(_03159_));
 sg13g2_o21ai_1 _08784_ (.B1(_03162_),
    .Y(_03167_),
    .A1(_03134_),
    .A2(_03163_));
 sg13g2_and3_1 _08785_ (.X(_03168_),
    .A(_03165_),
    .B(_03166_),
    .C(_03167_));
 sg13g2_nor2_1 _08786_ (.A(_03164_),
    .B(_03168_),
    .Y(_03169_));
 sg13g2_xnor2_1 _08787_ (.Y(_03170_),
    .A(_03139_),
    .B(_03140_));
 sg13g2_or2_1 _08788_ (.X(_03171_),
    .B(_03170_),
    .A(_03169_));
 sg13g2_nand2_1 _08789_ (.Y(_03172_),
    .A(net1642),
    .B(_02946_));
 sg13g2_and4_1 _08790_ (.A(net1633),
    .B(net1629),
    .C(net1622),
    .D(net1618),
    .X(_03173_));
 sg13g2_nand4_1 _08791_ (.B(net1629),
    .C(net1622),
    .A(net1633),
    .Y(_03174_),
    .D(net1618));
 sg13g2_nand2_1 _08792_ (.Y(_03175_),
    .A(net1635),
    .B(net1621));
 sg13g2_a22oi_1 _08793_ (.Y(_03176_),
    .B1(net1618),
    .B2(net1629),
    .A2(net1622),
    .A1(net1633));
 sg13g2_or2_1 _08794_ (.X(_03177_),
    .B(_03176_),
    .A(_03173_));
 sg13g2_o21ai_1 _08795_ (.B1(_03174_),
    .Y(_03178_),
    .A1(_03175_),
    .A2(_03176_));
 sg13g2_nand2_1 _08796_ (.Y(_03179_),
    .A(net1635),
    .B(net1624));
 sg13g2_nand2b_1 _08797_ (.Y(_03180_),
    .B(_03178_),
    .A_N(_03179_));
 sg13g2_xnor2_1 _08798_ (.Y(_03181_),
    .A(_03178_),
    .B(_03179_));
 sg13g2_nand2b_1 _08799_ (.Y(_03182_),
    .B(_03181_),
    .A_N(_03172_));
 sg13g2_xor2_1 _08800_ (.B(_03181_),
    .A(_03172_),
    .X(_03183_));
 sg13g2_xnor2_1 _08801_ (.Y(_03184_),
    .A(_03084_),
    .B(_03150_));
 sg13g2_nor2b_1 _08802_ (.A(_03183_),
    .B_N(_03184_),
    .Y(_03185_));
 sg13g2_a21o_1 _08803_ (.A2(_03153_),
    .A1(_03152_),
    .B1(_03160_),
    .X(_03186_));
 sg13g2_nand3_1 _08804_ (.B(_03185_),
    .C(_03186_),
    .A(_03161_),
    .Y(_03187_));
 sg13g2_nand2_1 _08805_ (.Y(_03188_),
    .A(_03180_),
    .B(_03182_));
 sg13g2_a21o_1 _08806_ (.A2(_03186_),
    .A1(_03161_),
    .B1(_03185_),
    .X(_03189_));
 sg13g2_nand3_1 _08807_ (.B(_03188_),
    .C(_03189_),
    .A(_03187_),
    .Y(_03190_));
 sg13g2_and2_1 _08808_ (.A(_03187_),
    .B(_03190_),
    .X(_03191_));
 sg13g2_a21oi_1 _08809_ (.A1(_03165_),
    .A2(_03167_),
    .Y(_03192_),
    .B1(_03166_));
 sg13g2_nor3_1 _08810_ (.A(_03168_),
    .B(_03191_),
    .C(_03192_),
    .Y(_03193_));
 sg13g2_o21ai_1 _08811_ (.B1(_03191_),
    .Y(_03194_),
    .A1(_03168_),
    .A2(_03192_));
 sg13g2_nor2b_1 _08812_ (.A(_03193_),
    .B_N(_03194_),
    .Y(_03195_));
 sg13g2_a21o_1 _08813_ (.A2(_03189_),
    .A1(_03187_),
    .B1(_03188_),
    .X(_03196_));
 sg13g2_or2_1 _08814_ (.X(_03197_),
    .B(_03175_),
    .A(_03117_));
 sg13g2_nor2_1 _08815_ (.A(_02951_),
    .B(_03197_),
    .Y(_03198_));
 sg13g2_nand2_1 _08816_ (.Y(_03199_),
    .A(net1642),
    .B(net1624));
 sg13g2_mux2_1 _08817_ (.A0(net1624),
    .A1(_03199_),
    .S(_03197_),
    .X(_03200_));
 sg13g2_nand2_1 _08818_ (.Y(_03201_),
    .A(net1637),
    .B(_02946_));
 sg13g2_nor2_1 _08819_ (.A(_03200_),
    .B(_03201_),
    .Y(_03202_));
 sg13g2_nor2_1 _08820_ (.A(_03198_),
    .B(_03202_),
    .Y(_03203_));
 sg13g2_xnor2_1 _08821_ (.Y(_03204_),
    .A(_03183_),
    .B(_03184_));
 sg13g2_xor2_1 _08822_ (.B(_03201_),
    .A(_03200_),
    .X(_03205_));
 sg13g2_xor2_1 _08823_ (.B(_03177_),
    .A(_03175_),
    .X(_03206_));
 sg13g2_nand2_1 _08824_ (.Y(_03207_),
    .A(_03205_),
    .B(_03206_));
 sg13g2_nand3_1 _08825_ (.B(_03205_),
    .C(_03206_),
    .A(_03204_),
    .Y(_03208_));
 sg13g2_inv_1 _08826_ (.Y(_03209_),
    .A(_03208_));
 sg13g2_xor2_1 _08827_ (.B(_03207_),
    .A(_03204_),
    .X(_03210_));
 sg13g2_nand2_1 _08828_ (.Y(_03211_),
    .A(net1637),
    .B(net1621));
 sg13g2_or3_1 _08829_ (.A(_02951_),
    .B(_03117_),
    .C(_03211_),
    .X(_03212_));
 sg13g2_nand2_1 _08830_ (.Y(_03213_),
    .A(net1637),
    .B(net1624));
 sg13g2_o21ai_1 _08831_ (.B1(_03213_),
    .Y(_03214_),
    .A1(_03117_),
    .A2(_03211_));
 sg13g2_nand2_1 _08832_ (.Y(_03215_),
    .A(_03212_),
    .B(_03214_));
 sg13g2_nand2_1 _08833_ (.Y(_03216_),
    .A(net1629),
    .B(_02946_));
 sg13g2_o21ai_1 _08834_ (.B1(_03212_),
    .Y(_03217_),
    .A1(_03215_),
    .A2(_03216_));
 sg13g2_xor2_1 _08835_ (.B(_03206_),
    .A(_03205_),
    .X(_03218_));
 sg13g2_nand2_1 _08836_ (.Y(_03219_),
    .A(_03117_),
    .B(_03211_));
 sg13g2_a21oi_1 _08837_ (.A1(_02917_),
    .A2(net1622),
    .Y(_03220_),
    .B1(net1624));
 sg13g2_nor2_1 _08838_ (.A(_02926_),
    .B(_03220_),
    .Y(_03221_));
 sg13g2_a21o_1 _08839_ (.A2(net1621),
    .A1(net1642),
    .B1(_03091_),
    .X(_03222_));
 sg13g2_xnor2_1 _08840_ (.Y(_03223_),
    .A(_03215_),
    .B(_03216_));
 sg13g2_a22oi_1 _08841_ (.Y(_03224_),
    .B1(_03222_),
    .B2(_03197_),
    .A2(_03221_),
    .A1(_03219_));
 sg13g2_nand4_1 _08842_ (.B(_03219_),
    .C(_03221_),
    .A(_03197_),
    .Y(_03225_),
    .D(_03222_));
 sg13g2_o21ai_1 _08843_ (.B1(_03225_),
    .Y(_03226_),
    .A1(_03223_),
    .A2(_03224_));
 sg13g2_a21oi_1 _08844_ (.A1(_03218_),
    .A2(_03226_),
    .Y(_03227_),
    .B1(_03217_));
 sg13g2_nor2_1 _08845_ (.A(_03218_),
    .B(_03226_),
    .Y(_03228_));
 sg13g2_a21oi_1 _08846_ (.A1(_03190_),
    .A2(_03196_),
    .Y(_03229_),
    .B1(_03209_));
 sg13g2_o21ai_1 _08847_ (.B1(_03208_),
    .Y(_03230_),
    .A1(_03203_),
    .A2(_03210_));
 sg13g2_nand3_1 _08848_ (.B(_03196_),
    .C(_03230_),
    .A(_03190_),
    .Y(_03231_));
 sg13g2_xnor2_1 _08849_ (.Y(_03232_),
    .A(_03203_),
    .B(_03210_));
 sg13g2_or3_1 _08850_ (.A(_03227_),
    .B(_03228_),
    .C(_03232_),
    .X(_03233_));
 sg13g2_o21ai_1 _08851_ (.B1(_03231_),
    .Y(_03234_),
    .A1(_03229_),
    .A2(_03233_));
 sg13g2_a21oi_2 _08852_ (.B1(_03193_),
    .Y(_03235_),
    .A2(_03234_),
    .A1(_03194_));
 sg13g2_and2_1 _08853_ (.A(_03169_),
    .B(_03170_),
    .X(_03236_));
 sg13g2_xor2_1 _08854_ (.B(_03170_),
    .A(_03169_),
    .X(_03237_));
 sg13g2_o21ai_1 _08855_ (.B1(_03171_),
    .Y(_03238_),
    .A1(_03235_),
    .A2(_03236_));
 sg13g2_xor2_1 _08856_ (.B(_03142_),
    .A(_03141_),
    .X(_03239_));
 sg13g2_a21oi_1 _08857_ (.A1(_03238_),
    .A2(_03239_),
    .Y(_03240_),
    .B1(_03143_));
 sg13g2_xor2_1 _08858_ (.B(_03114_),
    .A(_03113_),
    .X(_03241_));
 sg13g2_o21ai_1 _08859_ (.B1(_03115_),
    .Y(_03242_),
    .A1(_03240_),
    .A2(_03241_));
 sg13g2_xor2_1 _08860_ (.B(_03082_),
    .A(_03056_),
    .X(_03243_));
 sg13g2_a21oi_1 _08861_ (.A1(_03242_),
    .A2(_03243_),
    .Y(_03244_),
    .B1(_03083_));
 sg13g2_nand2_1 _08862_ (.Y(_03245_),
    .A(_03035_),
    .B(_03054_));
 sg13g2_xor2_1 _08863_ (.B(_03245_),
    .A(_03036_),
    .X(_03246_));
 sg13g2_inv_1 _08864_ (.Y(_03247_),
    .A(_03246_));
 sg13g2_o21ai_1 _08865_ (.B1(_03055_),
    .Y(_03248_),
    .A1(_03244_),
    .A2(_03247_));
 sg13g2_nand2_1 _08866_ (.Y(_03249_),
    .A(_03019_),
    .B(_03037_));
 sg13g2_xnor2_1 _08867_ (.Y(_03250_),
    .A(_03008_),
    .B(_03249_));
 sg13g2_a21oi_2 _08868_ (.B1(_03038_),
    .Y(_03251_),
    .A2(_03250_),
    .A1(_03248_));
 sg13g2_xnor2_1 _08869_ (.Y(_03252_),
    .A(_03020_),
    .B(_03022_));
 sg13g2_and2_1 _08870_ (.A(_03023_),
    .B(_03251_),
    .X(_03253_));
 sg13g2_a21oi_1 _08871_ (.A1(_03023_),
    .A2(_03251_),
    .Y(_03254_),
    .B1(_02970_));
 sg13g2_nand3_1 _08872_ (.B(_03023_),
    .C(_03251_),
    .A(_02970_),
    .Y(_03255_));
 sg13g2_nor2b_1 _08873_ (.A(_03254_),
    .B_N(_03255_),
    .Y(_03256_));
 sg13g2_a21oi_1 _08874_ (.A1(_02935_),
    .A2(_03255_),
    .Y(_03257_),
    .B1(_03254_));
 sg13g2_nor2_1 _08875_ (.A(_02938_),
    .B(_02966_),
    .Y(_03258_));
 sg13g2_xor2_1 _08876_ (.B(_02966_),
    .A(_02938_),
    .X(_03259_));
 sg13g2_o21ai_1 _08877_ (.B1(_02992_),
    .Y(_03260_),
    .A1(_03257_),
    .A2(_03258_));
 sg13g2_xor2_1 _08878_ (.B(_02962_),
    .A(_02934_),
    .X(_03261_));
 sg13g2_a21oi_1 _08879_ (.A1(_03260_),
    .A2(_03261_),
    .Y(_03262_),
    .B1(_02991_));
 sg13g2_a221oi_1 _08880_ (.B2(_03261_),
    .C1(_02991_),
    .B1(_03260_),
    .A1(_02936_),
    .Y(_03263_),
    .A2(_02967_));
 sg13g2_nor3_1 _08881_ (.A(_02989_),
    .B(_02990_),
    .C(_03263_),
    .Y(_03264_));
 sg13g2_nor2_1 _08882_ (.A(_02988_),
    .B(_03264_),
    .Y(_03265_));
 sg13g2_o21ai_1 _08883_ (.B1(_02986_),
    .Y(_03266_),
    .A1(_02988_),
    .A2(_03264_));
 sg13g2_a21o_2 _08884_ (.A2(_03266_),
    .A1(_02987_),
    .B1(_02985_),
    .X(_03267_));
 sg13g2_and2_1 _08885_ (.A(_02984_),
    .B(_03267_),
    .X(_03268_));
 sg13g2_nor2_1 _08886_ (.A(_02939_),
    .B(_02964_),
    .Y(_03269_));
 sg13g2_nand3_1 _08887_ (.B(_03267_),
    .C(_03269_),
    .A(_02984_),
    .Y(_03270_));
 sg13g2_nand2_1 _08888_ (.Y(_03271_),
    .A(_02939_),
    .B(_02964_));
 sg13g2_o21ai_1 _08889_ (.B1(_03271_),
    .Y(_03272_),
    .A1(_03268_),
    .A2(_03269_));
 sg13g2_nand2b_1 _08890_ (.Y(_03273_),
    .B(_03271_),
    .A_N(_03269_));
 sg13g2_a21o_1 _08891_ (.A2(_03267_),
    .A1(_02984_),
    .B1(_03273_),
    .X(_03274_));
 sg13g2_nand3_1 _08892_ (.B(_03267_),
    .C(_03273_),
    .A(_02984_),
    .Y(_03275_));
 sg13g2_and2_1 _08893_ (.A(_03274_),
    .B(_03275_),
    .X(_03276_));
 sg13g2_nand3_1 _08894_ (.B(_02987_),
    .C(_03266_),
    .A(_02985_),
    .Y(_03277_));
 sg13g2_nand2_1 _08895_ (.Y(_03278_),
    .A(_02986_),
    .B(_02987_));
 sg13g2_xor2_1 _08896_ (.B(_03278_),
    .A(_03265_),
    .X(_03279_));
 sg13g2_o21ai_1 _08897_ (.B1(_02989_),
    .Y(_03280_),
    .A1(_02990_),
    .A2(_03263_));
 sg13g2_nand2b_1 _08898_ (.Y(_03281_),
    .B(_03280_),
    .A_N(_03264_));
 sg13g2_xor2_1 _08899_ (.B(_02967_),
    .A(_02936_),
    .X(_03282_));
 sg13g2_xnor2_1 _08900_ (.Y(_03283_),
    .A(_03262_),
    .B(_03282_));
 sg13g2_xnor2_1 _08901_ (.Y(_03284_),
    .A(_03260_),
    .B(_03261_));
 sg13g2_xnor2_1 _08902_ (.Y(_03285_),
    .A(_03257_),
    .B(_03259_));
 sg13g2_xor2_1 _08903_ (.B(_03256_),
    .A(_02935_),
    .X(_03286_));
 sg13g2_xnor2_1 _08904_ (.Y(_03287_),
    .A(_02935_),
    .B(_03256_));
 sg13g2_nand2_1 _08905_ (.Y(_03288_),
    .A(_03285_),
    .B(_03286_));
 sg13g2_nor2_1 _08906_ (.A(_03284_),
    .B(_03288_),
    .Y(_03289_));
 sg13g2_nand2_1 _08907_ (.Y(_03290_),
    .A(_03283_),
    .B(_03289_));
 sg13g2_nor2_1 _08908_ (.A(_03281_),
    .B(_03290_),
    .Y(_03291_));
 sg13g2_and4_1 _08909_ (.A(_03267_),
    .B(_03277_),
    .C(_03279_),
    .D(_03291_),
    .X(_03292_));
 sg13g2_a22oi_1 _08910_ (.Y(_03293_),
    .B1(_03279_),
    .B2(_03291_),
    .A2(_03277_),
    .A1(_03267_));
 sg13g2_or2_1 _08911_ (.X(_03294_),
    .B(_03293_),
    .A(_03292_));
 sg13g2_xnor2_1 _08912_ (.Y(_03295_),
    .A(_03281_),
    .B(_03290_));
 sg13g2_nor2_1 _08913_ (.A(_03284_),
    .B(_03286_),
    .Y(_03296_));
 sg13g2_nand4_1 _08914_ (.B(_03283_),
    .C(_03285_),
    .A(_03279_),
    .Y(_03297_),
    .D(_03296_));
 sg13g2_nor4_1 _08915_ (.A(_03276_),
    .B(_03294_),
    .C(_03295_),
    .D(_03297_),
    .Y(_03298_));
 sg13g2_a21o_1 _08916_ (.A2(_03275_),
    .A1(_03274_),
    .B1(_03292_),
    .X(_03299_));
 sg13g2_nor2_1 _08917_ (.A(_03270_),
    .B(_03292_),
    .Y(_03300_));
 sg13g2_a21oi_1 _08918_ (.A1(_03272_),
    .A2(_03299_),
    .Y(_03301_),
    .B1(_03300_));
 sg13g2_nand2b_2 _08919_ (.Y(_03302_),
    .B(_03301_),
    .A_N(_03298_));
 sg13g2_nand3_1 _08920_ (.B(_02940_),
    .C(_02941_),
    .A(_02931_),
    .Y(_03303_));
 sg13g2_nand3_1 _08921_ (.B(_02971_),
    .C(_02972_),
    .A(_02960_),
    .Y(_03304_));
 sg13g2_and2_1 _08922_ (.A(_03303_),
    .B(_03304_),
    .X(_03305_));
 sg13g2_a22oi_1 _08923_ (.Y(_03306_),
    .B1(_02978_),
    .B2(_02929_),
    .A2(_02975_),
    .A1(_02958_));
 sg13g2_and2_1 _08924_ (.A(_03305_),
    .B(_03306_),
    .X(_03307_));
 sg13g2_nor2b_1 _08925_ (.A(_03302_),
    .B_N(_03307_),
    .Y(_03308_));
 sg13g2_xnor2_1 _08926_ (.Y(_03309_),
    .A(_03235_),
    .B(_03237_));
 sg13g2_xnor2_1 _08927_ (.Y(_03310_),
    .A(_03195_),
    .B(_03234_));
 sg13g2_nor2_1 _08928_ (.A(net1467),
    .B(_03309_),
    .Y(_03311_));
 sg13g2_a21oi_1 _08929_ (.A1(net1467),
    .A2(_03310_),
    .Y(_03312_),
    .B1(_03311_));
 sg13g2_nand3_1 _08930_ (.B(_03308_),
    .C(_03312_),
    .A(net1421),
    .Y(_03313_));
 sg13g2_a21oi_1 _08931_ (.A1(net1493),
    .A2(_03313_),
    .Y(_03314_),
    .B1(net1522));
 sg13g2_a21o_1 _08932_ (.A2(net1525),
    .A1(net1011),
    .B1(_03314_),
    .X(_00318_));
 sg13g2_nand2b_1 _08933_ (.Y(_03315_),
    .B(net1467),
    .A_N(_03309_));
 sg13g2_xnor2_1 _08934_ (.Y(_03316_),
    .A(_03238_),
    .B(_03239_));
 sg13g2_nand2b_1 _08935_ (.Y(_03317_),
    .B(_03316_),
    .A_N(net1468));
 sg13g2_nand4_1 _08936_ (.B(_03307_),
    .C(_03315_),
    .A(net1421),
    .Y(_03318_),
    .D(_03317_));
 sg13g2_o21ai_1 _08937_ (.B1(net1493),
    .Y(_03319_),
    .A1(_03302_),
    .A2(_03318_));
 sg13g2_a22oi_1 _08938_ (.Y(_03320_),
    .B1(_02911_),
    .B2(_03319_),
    .A2(net1524),
    .A1(net905));
 sg13g2_inv_1 _08939_ (.Y(_00319_),
    .A(net906));
 sg13g2_xnor2_1 _08940_ (.Y(_03321_),
    .A(_03240_),
    .B(_03241_));
 sg13g2_nand2b_1 _08941_ (.Y(_03322_),
    .B(_03321_),
    .A_N(net1467));
 sg13g2_nand2_1 _08942_ (.Y(_03323_),
    .A(net1467),
    .B(_03316_));
 sg13g2_nand4_1 _08943_ (.B(_03307_),
    .C(_03322_),
    .A(net1421),
    .Y(_03324_),
    .D(_03323_));
 sg13g2_o21ai_1 _08944_ (.B1(net1493),
    .Y(_03325_),
    .A1(_03302_),
    .A2(_03324_));
 sg13g2_a22oi_1 _08945_ (.Y(_03326_),
    .B1(_02911_),
    .B2(_03325_),
    .A2(net1525),
    .A1(net890));
 sg13g2_inv_1 _08946_ (.Y(_00320_),
    .A(net891));
 sg13g2_xnor2_1 _08947_ (.Y(_03327_),
    .A(_03242_),
    .B(_03243_));
 sg13g2_nand2b_1 _08948_ (.Y(_03328_),
    .B(_03327_),
    .A_N(net1467));
 sg13g2_nand2_1 _08949_ (.Y(_03329_),
    .A(net1467),
    .B(_03321_));
 sg13g2_nand4_1 _08950_ (.B(_03307_),
    .C(_03328_),
    .A(net1421),
    .Y(_03330_),
    .D(_03329_));
 sg13g2_o21ai_1 _08951_ (.B1(net1493),
    .Y(_03331_),
    .A1(_03302_),
    .A2(_03330_));
 sg13g2_a22oi_1 _08952_ (.Y(_03332_),
    .B1(_02911_),
    .B2(_03331_),
    .A2(_02910_),
    .A1(net868));
 sg13g2_inv_1 _08953_ (.Y(_00321_),
    .A(net869));
 sg13g2_xnor2_1 _08954_ (.Y(_03333_),
    .A(_03244_),
    .B(_03246_));
 sg13g2_o21ai_1 _08955_ (.B1(_03307_),
    .Y(_03334_),
    .A1(net1468),
    .A2(_03333_));
 sg13g2_a21oi_1 _08956_ (.A1(net1467),
    .A2(_03327_),
    .Y(_03335_),
    .B1(_03334_));
 sg13g2_nand2_1 _08957_ (.Y(_03336_),
    .A(net1421),
    .B(_03335_));
 sg13g2_o21ai_1 _08958_ (.B1(net1493),
    .Y(_03337_),
    .A1(_03302_),
    .A2(_03336_));
 sg13g2_a22oi_1 _08959_ (.Y(_03338_),
    .B1(_02911_),
    .B2(_03337_),
    .A2(net1524),
    .A1(net874));
 sg13g2_inv_1 _08960_ (.Y(_00322_),
    .A(net875));
 sg13g2_xor2_1 _08961_ (.B(_03250_),
    .A(_03248_),
    .X(_03339_));
 sg13g2_mux2_1 _08962_ (.A0(_03339_),
    .A1(_03333_),
    .S(net1468),
    .X(_03340_));
 sg13g2_nand3_1 _08963_ (.B(_03308_),
    .C(_03340_),
    .A(net1421),
    .Y(_03341_));
 sg13g2_a21oi_1 _08964_ (.A1(net1493),
    .A2(_03341_),
    .Y(_03342_),
    .B1(net1522));
 sg13g2_a21o_1 _08965_ (.A2(net1525),
    .A1(net1021),
    .B1(_03342_),
    .X(_00323_));
 sg13g2_nand2b_1 _08966_ (.Y(_03343_),
    .B(net1468),
    .A_N(_03339_));
 sg13g2_xnor2_1 _08967_ (.Y(_03344_),
    .A(_03251_),
    .B(_03252_));
 sg13g2_nand4_1 _08968_ (.B(_03308_),
    .C(_03343_),
    .A(net1421),
    .Y(_03345_),
    .D(_03344_));
 sg13g2_a21oi_1 _08969_ (.A1(net1493),
    .A2(_03345_),
    .Y(_03346_),
    .B1(net1522));
 sg13g2_a21o_1 _08970_ (.A2(net1525),
    .A1(net1016),
    .B1(_03346_),
    .X(_00324_));
 sg13g2_and2_2 _08971_ (.A(net1421),
    .B(_03305_),
    .X(_03347_));
 sg13g2_inv_1 _08972_ (.Y(_03348_),
    .A(_03347_));
 sg13g2_and2_1 _08973_ (.A(_03301_),
    .B(_03306_),
    .X(_03349_));
 sg13g2_nand2b_2 _08974_ (.Y(_03350_),
    .B(_03306_),
    .A_N(_03302_));
 sg13g2_o21ai_1 _08975_ (.B1(_03347_),
    .Y(_03351_),
    .A1(_03287_),
    .A2(_03350_));
 sg13g2_a21oi_1 _08976_ (.A1(net1494),
    .A2(_03351_),
    .Y(_03352_),
    .B1(net1522));
 sg13g2_a21o_1 _08977_ (.A2(net1524),
    .A1(net1000),
    .B1(_03352_),
    .X(_00325_));
 sg13g2_xnor2_1 _08978_ (.Y(_03353_),
    .A(_03285_),
    .B(_03287_));
 sg13g2_o21ai_1 _08979_ (.B1(_03347_),
    .Y(_03354_),
    .A1(_03350_),
    .A2(_03353_));
 sg13g2_a21oi_1 _08980_ (.A1(net1494),
    .A2(_03354_),
    .Y(_03355_),
    .B1(net1523));
 sg13g2_a21o_1 _08981_ (.A2(net1524),
    .A1(net613),
    .B1(_03355_),
    .X(_00326_));
 sg13g2_xor2_1 _08982_ (.B(_03288_),
    .A(_03284_),
    .X(_03356_));
 sg13g2_o21ai_1 _08983_ (.B1(_03347_),
    .Y(_03357_),
    .A1(_03350_),
    .A2(_03356_));
 sg13g2_a21oi_1 _08984_ (.A1(net1494),
    .A2(_03357_),
    .Y(_03358_),
    .B1(net1522));
 sg13g2_a21o_1 _08985_ (.A2(net1524),
    .A1(net578),
    .B1(_03358_),
    .X(_00327_));
 sg13g2_xor2_1 _08986_ (.B(_03289_),
    .A(_03283_),
    .X(_03359_));
 sg13g2_o21ai_1 _08987_ (.B1(_03347_),
    .Y(_03360_),
    .A1(_03350_),
    .A2(_03359_));
 sg13g2_a21oi_1 _08988_ (.A1(net1494),
    .A2(_03360_),
    .Y(_03361_),
    .B1(net1522));
 sg13g2_a21o_1 _08989_ (.A2(net1524),
    .A1(net650),
    .B1(_03361_),
    .X(_00328_));
 sg13g2_a21o_1 _08990_ (.A2(_03349_),
    .A1(_03295_),
    .B1(_03348_),
    .X(_03362_));
 sg13g2_a21oi_1 _08991_ (.A1(net1494),
    .A2(_03362_),
    .Y(_03363_),
    .B1(net1523));
 sg13g2_a21o_1 _08992_ (.A2(net1525),
    .A1(net641),
    .B1(_03363_),
    .X(_00329_));
 sg13g2_xor2_1 _08993_ (.B(_03291_),
    .A(_03279_),
    .X(_03364_));
 sg13g2_o21ai_1 _08994_ (.B1(_03347_),
    .Y(_03365_),
    .A1(_03350_),
    .A2(_03364_));
 sg13g2_a21oi_1 _08995_ (.A1(net1494),
    .A2(_03365_),
    .Y(_03366_),
    .B1(net1523));
 sg13g2_a21o_1 _08996_ (.A2(net1524),
    .A1(net603),
    .B1(_03366_),
    .X(_00330_));
 sg13g2_a21o_1 _08997_ (.A2(_03349_),
    .A1(_03294_),
    .B1(_03348_),
    .X(_03367_));
 sg13g2_a21oi_1 _08998_ (.A1(net1493),
    .A2(_03367_),
    .Y(_03368_),
    .B1(net1522));
 sg13g2_a21o_1 _08999_ (.A2(net1525),
    .A1(net647),
    .B1(_03368_),
    .X(_00331_));
 sg13g2_xnor2_1 _09000_ (.Y(_03369_),
    .A(_03276_),
    .B(_03292_));
 sg13g2_o21ai_1 _09001_ (.B1(_03347_),
    .Y(_03370_),
    .A1(_03350_),
    .A2(_03369_));
 sg13g2_a21oi_1 _09002_ (.A1(net1494),
    .A2(_03370_),
    .Y(_03371_),
    .B1(net1523));
 sg13g2_a21o_1 _09003_ (.A2(net1525),
    .A1(net602),
    .B1(_03371_),
    .X(_00332_));
 sg13g2_xor2_1 _09004_ (.B(_02959_),
    .A(_02930_),
    .X(_03372_));
 sg13g2_nand2_1 _09005_ (.Y(_03373_),
    .A(_03347_),
    .B(_03372_));
 sg13g2_a21oi_1 _09006_ (.A1(net1494),
    .A2(_03373_),
    .Y(_03374_),
    .B1(net1522));
 sg13g2_a21o_1 _09007_ (.A2(net1524),
    .A1(net978),
    .B1(_03374_),
    .X(_00333_));
 sg13g2_and2_1 _09008_ (.A(net1767),
    .B(net1650),
    .X(_03375_));
 sg13g2_nand2_1 _09009_ (.Y(_03376_),
    .A(net1767),
    .B(net1650));
 sg13g2_nand2_1 _09010_ (.Y(_03377_),
    .A(net969),
    .B(net1538));
 sg13g2_mux2_1 _09011_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[6][14] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[7][14] ),
    .S(net1704),
    .X(_03378_));
 sg13g2_mux2_2 _09012_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[6][13] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[7][13] ),
    .S(net1701),
    .X(_03379_));
 sg13g2_mux2_1 _09013_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[6][8] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[7][8] ),
    .S(net1704),
    .X(_03380_));
 sg13g2_mux2_2 _09014_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[6][11] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[7][11] ),
    .S(net1701),
    .X(_03381_));
 sg13g2_mux2_2 _09015_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[6][9] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[7][9] ),
    .S(net1701),
    .X(_03382_));
 sg13g2_mux2_2 _09016_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[6][12] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[7][12] ),
    .S(net1700),
    .X(_03383_));
 sg13g2_mux2_2 _09017_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[6][10] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[7][10] ),
    .S(net1700),
    .X(_03384_));
 sg13g2_mux2_2 _09018_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[6][7] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[7][7] ),
    .S(net1704),
    .X(_03385_));
 sg13g2_nor4_1 _09019_ (.A(_03378_),
    .B(_03379_),
    .C(_03381_),
    .D(_03383_),
    .Y(_03386_));
 sg13g2_nor4_1 _09020_ (.A(_03380_),
    .B(_03382_),
    .C(_03384_),
    .D(_03385_),
    .Y(_03387_));
 sg13g2_nand2_1 _09021_ (.Y(_03388_),
    .A(_03386_),
    .B(_03387_));
 sg13g2_inv_1 _09022_ (.Y(_03389_),
    .A(_03388_));
 sg13g2_mux2_1 _09023_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[6][0] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[7][0] ),
    .S(net1700),
    .X(_03390_));
 sg13g2_mux2_1 _09024_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[6][6] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[7][6] ),
    .S(net1700),
    .X(_03391_));
 sg13g2_nand2_1 _09025_ (.Y(_03392_),
    .A(_00137_),
    .B(net1701));
 sg13g2_mux2_2 _09026_ (.A0(_00757_),
    .A1(_00758_),
    .S(net1701),
    .X(_03393_));
 sg13g2_o21ai_1 _09027_ (.B1(_03392_),
    .Y(_03394_),
    .A1(_00757_),
    .A2(net1701));
 sg13g2_nor3_1 _09028_ (.A(net1617),
    .B(net1614),
    .C(net1613),
    .Y(_03395_));
 sg13g2_mux2_2 _09029_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[6][2] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[7][2] ),
    .S(net1700),
    .X(_03396_));
 sg13g2_inv_1 _09030_ (.Y(_03397_),
    .A(_03396_));
 sg13g2_mux2_1 _09031_ (.A0(_00136_),
    .A1(_00135_),
    .S(net1700),
    .X(_03398_));
 sg13g2_mux2_1 _09032_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[6][1] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[7][1] ),
    .S(net1700),
    .X(_03399_));
 sg13g2_mux2_1 _09033_ (.A0(_00759_),
    .A1(_00760_),
    .S(net1700),
    .X(_03400_));
 sg13g2_nor2_1 _09034_ (.A(_03399_),
    .B(net1607),
    .Y(_03401_));
 sg13g2_and4_1 _09035_ (.A(_03395_),
    .B(_03397_),
    .C(net1611),
    .D(_03401_),
    .X(_03402_));
 sg13g2_nand4_1 _09036_ (.B(_03397_),
    .C(net1610),
    .A(_03395_),
    .Y(_03403_),
    .D(_03401_));
 sg13g2_mux2_2 _09037_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[6][15] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[7][15] ),
    .S(net1704),
    .X(_03404_));
 sg13g2_nor2_1 _09038_ (.A(_03403_),
    .B(_03404_),
    .Y(_03405_));
 sg13g2_nand2b_1 _09039_ (.Y(_03406_),
    .B(_03389_),
    .A_N(_03405_));
 sg13g2_mux2_2 _09040_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][12] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][12] ),
    .S(net1696),
    .X(_03407_));
 sg13g2_mux2_1 _09041_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][8] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][8] ),
    .S(net1703),
    .X(_03408_));
 sg13g2_mux2_2 _09042_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][10] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][10] ),
    .S(net1696),
    .X(_03409_));
 sg13g2_mux2_2 _09043_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][14] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][14] ),
    .S(net1703),
    .X(_03410_));
 sg13g2_mux2_2 _09044_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][7] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][7] ),
    .S(net1696),
    .X(_03411_));
 sg13g2_inv_1 _09045_ (.Y(_03412_),
    .A(_03411_));
 sg13g2_mux2_2 _09046_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][11] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][11] ),
    .S(net1696),
    .X(_03413_));
 sg13g2_mux2_2 _09047_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][13] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][13] ),
    .S(net1703),
    .X(_03414_));
 sg13g2_mux2_2 _09048_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][9] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][9] ),
    .S(net1703),
    .X(_03415_));
 sg13g2_nor4_1 _09049_ (.A(_03407_),
    .B(_03409_),
    .C(_03410_),
    .D(_03414_),
    .Y(_03416_));
 sg13g2_nor4_1 _09050_ (.A(_03408_),
    .B(_03411_),
    .C(_03413_),
    .D(_03415_),
    .Y(_03417_));
 sg13g2_and2_1 _09051_ (.A(_03416_),
    .B(_03417_),
    .X(_03418_));
 sg13g2_mux2_2 _09052_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][3] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][3] ),
    .S(net1690),
    .X(_03419_));
 sg13g2_mux2_2 _09053_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][6] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][6] ),
    .S(net1694),
    .X(_03420_));
 sg13g2_mux2_2 _09054_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][1] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][1] ),
    .S(net1689),
    .X(_03421_));
 sg13g2_mux2_2 _09055_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][2] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][2] ),
    .S(net1690),
    .X(_03422_));
 sg13g2_mux2_2 _09056_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][0] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][0] ),
    .S(net1691),
    .X(_03423_));
 sg13g2_mux2_2 _09057_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][5] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][5] ),
    .S(net1689),
    .X(_03424_));
 sg13g2_inv_2 _09058_ (.Y(_03425_),
    .A(net1596));
 sg13g2_mux2_2 _09059_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][4] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][4] ),
    .S(net1694),
    .X(_03426_));
 sg13g2_nor3_1 _09060_ (.A(net1603),
    .B(net1601),
    .C(net1595),
    .Y(_03427_));
 sg13g2_nor3_1 _09061_ (.A(net1605),
    .B(net1600),
    .C(net1597),
    .Y(_03428_));
 sg13g2_nand3_1 _09062_ (.B(_03427_),
    .C(_03428_),
    .A(_03425_),
    .Y(_03429_));
 sg13g2_mux2_2 _09063_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[6][15] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[7][15] ),
    .S(net1703),
    .X(_03430_));
 sg13g2_nor2_1 _09064_ (.A(_03429_),
    .B(_03430_),
    .Y(_03431_));
 sg13g2_o21ai_1 _09065_ (.B1(_03418_),
    .Y(_03432_),
    .A1(_03429_),
    .A2(_03430_));
 sg13g2_nand4_1 _09066_ (.B(_03380_),
    .C(_03382_),
    .A(_03378_),
    .Y(_03433_),
    .D(_03383_));
 sg13g2_nand4_1 _09067_ (.B(_03381_),
    .C(_03384_),
    .A(_03379_),
    .Y(_03434_),
    .D(_03385_));
 sg13g2_nor2_1 _09068_ (.A(_03433_),
    .B(_03434_),
    .Y(_03435_));
 sg13g2_nand4_1 _09069_ (.B(_03409_),
    .C(_03410_),
    .A(_03407_),
    .Y(_03436_),
    .D(_03414_));
 sg13g2_nand3_1 _09070_ (.B(_03413_),
    .C(_03415_),
    .A(_03408_),
    .Y(_03437_));
 sg13g2_nor3_1 _09071_ (.A(_03412_),
    .B(_03436_),
    .C(_03437_),
    .Y(_03438_));
 sg13g2_a22oi_1 _09072_ (.Y(_03439_),
    .B1(_03438_),
    .B2(_03429_),
    .A2(_03435_),
    .A1(_03403_));
 sg13g2_nand4_1 _09073_ (.B(_03406_),
    .C(_03432_),
    .A(net1768),
    .Y(_03440_),
    .D(_03439_));
 sg13g2_or2_1 _09074_ (.X(_03441_),
    .B(_03410_),
    .A(_03378_));
 sg13g2_nand2_1 _09075_ (.Y(_03442_),
    .A(_03379_),
    .B(_03414_));
 sg13g2_xnor2_1 _09076_ (.Y(_03443_),
    .A(_03379_),
    .B(_03414_));
 sg13g2_or2_1 _09077_ (.X(_03444_),
    .B(_03407_),
    .A(_03383_));
 sg13g2_nand2_1 _09078_ (.Y(_03445_),
    .A(_03383_),
    .B(_03407_));
 sg13g2_and2_1 _09079_ (.A(_03381_),
    .B(_03413_),
    .X(_03446_));
 sg13g2_xnor2_1 _09080_ (.Y(_03447_),
    .A(_03381_),
    .B(_03413_));
 sg13g2_nor2_1 _09081_ (.A(_03384_),
    .B(_03409_),
    .Y(_03448_));
 sg13g2_and2_1 _09082_ (.A(_03382_),
    .B(_03415_),
    .X(_03449_));
 sg13g2_and2_1 _09083_ (.A(_03380_),
    .B(_03408_),
    .X(_03450_));
 sg13g2_nand2_1 _09084_ (.Y(_03451_),
    .A(net1615),
    .B(net1603));
 sg13g2_xnor2_1 _09085_ (.Y(_03452_),
    .A(_03425_),
    .B(_03451_));
 sg13g2_xnor2_1 _09086_ (.Y(_03453_),
    .A(_03394_),
    .B(_03452_));
 sg13g2_nand2_1 _09087_ (.Y(_03454_),
    .A(net1615),
    .B(net1596));
 sg13g2_nand3_1 _09088_ (.B(net1596),
    .C(net1595),
    .A(net1615),
    .Y(_03455_));
 sg13g2_nand2_1 _09089_ (.Y(_03456_),
    .A(_03393_),
    .B(_03420_));
 sg13g2_xor2_1 _09090_ (.B(_03454_),
    .A(net1595),
    .X(_03457_));
 sg13g2_o21ai_1 _09091_ (.B1(_03455_),
    .Y(_03458_),
    .A1(_03456_),
    .A2(_03457_));
 sg13g2_nand2b_1 _09092_ (.Y(_03459_),
    .B(_03458_),
    .A_N(_03453_));
 sg13g2_xor2_1 _09093_ (.B(net1603),
    .A(net1615),
    .X(_03460_));
 sg13g2_nor2_2 _09094_ (.A(_03394_),
    .B(_03425_),
    .Y(_03461_));
 sg13g2_inv_1 _09095_ (.Y(_03462_),
    .A(_03461_));
 sg13g2_nand2_1 _09096_ (.Y(_03463_),
    .A(_03460_),
    .B(_03461_));
 sg13g2_o21ai_1 _09097_ (.B1(_03454_),
    .Y(_03464_),
    .A1(_03394_),
    .A2(_03452_));
 sg13g2_o21ai_1 _09098_ (.B1(_03463_),
    .Y(_03465_),
    .A1(_03460_),
    .A2(_03464_));
 sg13g2_nand2b_1 _09099_ (.Y(_03466_),
    .B(_03459_),
    .A_N(_03465_));
 sg13g2_xnor2_1 _09100_ (.Y(_03467_),
    .A(_03453_),
    .B(_03458_));
 sg13g2_nand3_1 _09101_ (.B(net1605),
    .C(net1595),
    .A(net1615),
    .Y(_03468_));
 sg13g2_a21o_1 _09102_ (.A2(net1594),
    .A1(net1615),
    .B1(net1605),
    .X(_03469_));
 sg13g2_nand2_1 _09103_ (.Y(_03470_),
    .A(_03468_),
    .B(_03469_));
 sg13g2_o21ai_1 _09104_ (.B1(_03468_),
    .Y(_03471_),
    .A1(_03462_),
    .A2(_03470_));
 sg13g2_xor2_1 _09105_ (.B(_03457_),
    .A(_03456_),
    .X(_03472_));
 sg13g2_and2_1 _09106_ (.A(_03471_),
    .B(_03472_),
    .X(_03473_));
 sg13g2_or2_1 _09107_ (.X(_03474_),
    .B(_03472_),
    .A(_03471_));
 sg13g2_nand2b_1 _09108_ (.Y(_03475_),
    .B(_03474_),
    .A_N(_03473_));
 sg13g2_a21o_1 _09109_ (.A2(_03474_),
    .A1(net1608),
    .B1(_03473_),
    .X(_03476_));
 sg13g2_nand2_1 _09110_ (.Y(_03477_),
    .A(_03467_),
    .B(_03476_));
 sg13g2_xor2_1 _09111_ (.B(_03476_),
    .A(_03467_),
    .X(_03478_));
 sg13g2_xnor2_1 _09112_ (.Y(_03479_),
    .A(net1608),
    .B(_03475_));
 sg13g2_nand3_1 _09113_ (.B(net1605),
    .C(net1600),
    .A(net1615),
    .Y(_03480_));
 sg13g2_nand2_1 _09114_ (.Y(_03481_),
    .A(_03393_),
    .B(net1595));
 sg13g2_a21o_1 _09115_ (.A2(net1604),
    .A1(net1615),
    .B1(net1600),
    .X(_03482_));
 sg13g2_nand2_1 _09116_ (.Y(_03483_),
    .A(_03480_),
    .B(_03482_));
 sg13g2_o21ai_1 _09117_ (.B1(_03480_),
    .Y(_03484_),
    .A1(_03481_),
    .A2(_03483_));
 sg13g2_xor2_1 _09118_ (.B(_03470_),
    .A(_03461_),
    .X(_03485_));
 sg13g2_nand2b_1 _09119_ (.Y(_03486_),
    .B(_03484_),
    .A_N(_03485_));
 sg13g2_nand2_1 _09120_ (.Y(_03487_),
    .A(net1608),
    .B(_03420_));
 sg13g2_xor2_1 _09121_ (.B(_03485_),
    .A(_03484_),
    .X(_03488_));
 sg13g2_o21ai_1 _09122_ (.B1(_03486_),
    .Y(_03489_),
    .A1(_03487_),
    .A2(_03488_));
 sg13g2_and2_1 _09123_ (.A(_03479_),
    .B(_03489_),
    .X(_03490_));
 sg13g2_nand2_1 _09124_ (.Y(_03491_),
    .A(_03478_),
    .B(_03490_));
 sg13g2_or2_1 _09125_ (.X(_03492_),
    .B(_03491_),
    .A(_03466_));
 sg13g2_inv_1 _09126_ (.Y(_03493_),
    .A(_03492_));
 sg13g2_xor2_1 _09127_ (.B(_03489_),
    .A(_03479_),
    .X(_03494_));
 sg13g2_inv_1 _09128_ (.Y(_03495_),
    .A(_03494_));
 sg13g2_nand3_1 _09129_ (.B(net1602),
    .C(net1600),
    .A(net1614),
    .Y(_03496_));
 sg13g2_nand2_1 _09130_ (.Y(_03497_),
    .A(_03393_),
    .B(net1605));
 sg13g2_a21o_1 _09131_ (.A2(net1600),
    .A1(net1614),
    .B1(net1601),
    .X(_03498_));
 sg13g2_nand2_1 _09132_ (.Y(_03499_),
    .A(_03496_),
    .B(_03498_));
 sg13g2_o21ai_1 _09133_ (.B1(_03496_),
    .Y(_03500_),
    .A1(_03497_),
    .A2(_03499_));
 sg13g2_xor2_1 _09134_ (.B(_03483_),
    .A(_03481_),
    .X(_03501_));
 sg13g2_nand2_1 _09135_ (.Y(_03502_),
    .A(_03500_),
    .B(_03501_));
 sg13g2_nand2_1 _09136_ (.Y(_03503_),
    .A(net1608),
    .B(_03424_));
 sg13g2_xnor2_1 _09137_ (.Y(_03504_),
    .A(_03500_),
    .B(_03501_));
 sg13g2_o21ai_1 _09138_ (.B1(_03502_),
    .Y(_03505_),
    .A1(_03503_),
    .A2(_03504_));
 sg13g2_xor2_1 _09139_ (.B(_03488_),
    .A(_03487_),
    .X(_03506_));
 sg13g2_nand2_1 _09140_ (.Y(_03507_),
    .A(_03505_),
    .B(_03506_));
 sg13g2_xnor2_1 _09141_ (.Y(_03508_),
    .A(_03505_),
    .B(_03506_));
 sg13g2_or2_1 _09142_ (.X(_03509_),
    .B(_03508_),
    .A(net1610));
 sg13g2_a21oi_1 _09143_ (.A1(_03507_),
    .A2(_03509_),
    .Y(_03510_),
    .B1(_03495_));
 sg13g2_nand2_1 _09144_ (.Y(_03511_),
    .A(_03478_),
    .B(_03510_));
 sg13g2_nand3_1 _09145_ (.B(_03507_),
    .C(_03509_),
    .A(_03495_),
    .Y(_03512_));
 sg13g2_nor2b_1 _09146_ (.A(_03510_),
    .B_N(_03512_),
    .Y(_03513_));
 sg13g2_and3_1 _09147_ (.X(_03514_),
    .A(net1614),
    .B(net1602),
    .C(net1598));
 sg13g2_nand3_1 _09148_ (.B(net1602),
    .C(net1598),
    .A(net1614),
    .Y(_03515_));
 sg13g2_nand2_1 _09149_ (.Y(_03516_),
    .A(net1613),
    .B(net1600));
 sg13g2_a21oi_1 _09150_ (.A1(net1614),
    .A2(net1602),
    .Y(_03517_),
    .B1(net1598));
 sg13g2_a21o_1 _09151_ (.A2(net1602),
    .A1(net1614),
    .B1(net1598),
    .X(_03518_));
 sg13g2_nor3_1 _09152_ (.A(_03514_),
    .B(_03516_),
    .C(_03517_),
    .Y(_03519_));
 sg13g2_o21ai_1 _09153_ (.B1(_03515_),
    .Y(_03520_),
    .A1(_03516_),
    .A2(_03517_));
 sg13g2_xor2_1 _09154_ (.B(_03499_),
    .A(_03497_),
    .X(_03521_));
 sg13g2_nand2_1 _09155_ (.Y(_03522_),
    .A(_03520_),
    .B(_03521_));
 sg13g2_xnor2_1 _09156_ (.Y(_03523_),
    .A(_03520_),
    .B(_03521_));
 sg13g2_nand2_1 _09157_ (.Y(_03524_),
    .A(net1609),
    .B(net1594));
 sg13g2_nand3_1 _09158_ (.B(net1607),
    .C(net1594),
    .A(net1609),
    .Y(_03525_));
 sg13g2_a21o_1 _09159_ (.A2(net1595),
    .A1(net1607),
    .B1(net1609),
    .X(_03526_));
 sg13g2_nand2_1 _09160_ (.Y(_03527_),
    .A(_03525_),
    .B(_03526_));
 sg13g2_o21ai_1 _09161_ (.B1(_03522_),
    .Y(_03528_),
    .A1(_03523_),
    .A2(_03527_));
 sg13g2_xor2_1 _09162_ (.B(_03504_),
    .A(_03503_),
    .X(_03529_));
 sg13g2_nand2_1 _09163_ (.Y(_03530_),
    .A(_03528_),
    .B(_03529_));
 sg13g2_xnor2_1 _09164_ (.Y(_03531_),
    .A(_03397_),
    .B(_03525_));
 sg13g2_nand2b_1 _09165_ (.Y(_03532_),
    .B(net1603),
    .A_N(net1611));
 sg13g2_or2_1 _09166_ (.X(_03533_),
    .B(_03532_),
    .A(_03531_));
 sg13g2_xnor2_1 _09167_ (.Y(_03534_),
    .A(_03531_),
    .B(_03532_));
 sg13g2_xnor2_1 _09168_ (.Y(_03535_),
    .A(_03528_),
    .B(_03529_));
 sg13g2_o21ai_1 _09169_ (.B1(_03530_),
    .Y(_03536_),
    .A1(_03534_),
    .A2(_03535_));
 sg13g2_xor2_1 _09170_ (.B(_03508_),
    .A(net1610),
    .X(_03537_));
 sg13g2_nand2_1 _09171_ (.Y(_03538_),
    .A(_03536_),
    .B(_03537_));
 sg13g2_o21ai_1 _09172_ (.B1(_03533_),
    .Y(_03539_),
    .A1(_03397_),
    .A2(_03525_));
 sg13g2_inv_1 _09173_ (.Y(_03540_),
    .A(_03539_));
 sg13g2_xnor2_1 _09174_ (.Y(_03541_),
    .A(_03536_),
    .B(_03537_));
 sg13g2_o21ai_1 _09175_ (.B1(_03538_),
    .Y(_03542_),
    .A1(_03540_),
    .A2(_03541_));
 sg13g2_and2_1 _09176_ (.A(_03513_),
    .B(_03542_),
    .X(_03543_));
 sg13g2_nand2_1 _09177_ (.Y(_03544_),
    .A(net1613),
    .B(_03514_));
 sg13g2_a22oi_1 _09178_ (.Y(_03545_),
    .B1(_03515_),
    .B2(_03518_),
    .A2(net1600),
    .A1(net1613));
 sg13g2_nand3_1 _09179_ (.B(net1599),
    .C(_03514_),
    .A(net1613),
    .Y(_03546_));
 sg13g2_o21ai_1 _09180_ (.B1(_03544_),
    .Y(_03547_),
    .A1(_03519_),
    .A2(_03545_));
 sg13g2_nand2_1 _09181_ (.Y(_03548_),
    .A(_03399_),
    .B(net1603));
 sg13g2_nand3_1 _09182_ (.B(net1606),
    .C(net1604),
    .A(net1617),
    .Y(_03549_));
 sg13g2_a21o_1 _09183_ (.A2(net1604),
    .A1(net1607),
    .B1(net1617),
    .X(_03550_));
 sg13g2_nand2_1 _09184_ (.Y(_03551_),
    .A(_03549_),
    .B(_03550_));
 sg13g2_xor2_1 _09185_ (.B(_03551_),
    .A(_03548_),
    .X(_03552_));
 sg13g2_nand3_1 _09186_ (.B(_03547_),
    .C(_03552_),
    .A(_03546_),
    .Y(_03553_));
 sg13g2_nand2_1 _09187_ (.Y(_03554_),
    .A(_03546_),
    .B(_03553_));
 sg13g2_xor2_1 _09188_ (.B(_03527_),
    .A(_03523_),
    .X(_03555_));
 sg13g2_nand2_1 _09189_ (.Y(_03556_),
    .A(_03554_),
    .B(_03555_));
 sg13g2_xnor2_1 _09190_ (.Y(_03557_),
    .A(_03554_),
    .B(_03555_));
 sg13g2_o21ai_1 _09191_ (.B1(_03549_),
    .Y(_03558_),
    .A1(_03548_),
    .A2(_03551_));
 sg13g2_nand2_1 _09192_ (.Y(_03559_),
    .A(_03396_),
    .B(net1603));
 sg13g2_inv_1 _09193_ (.Y(_03560_),
    .A(_03559_));
 sg13g2_xnor2_1 _09194_ (.Y(_03561_),
    .A(_03558_),
    .B(_03560_));
 sg13g2_nor3_1 _09195_ (.A(net1611),
    .B(_03425_),
    .C(_03561_),
    .Y(_03562_));
 sg13g2_o21ai_1 _09196_ (.B1(_03561_),
    .Y(_03563_),
    .A1(net1611),
    .A2(_03425_));
 sg13g2_nand2b_1 _09197_ (.Y(_03564_),
    .B(_03563_),
    .A_N(_03562_));
 sg13g2_o21ai_1 _09198_ (.B1(_03556_),
    .Y(_03565_),
    .A1(_03557_),
    .A2(_03564_));
 sg13g2_xor2_1 _09199_ (.B(_03535_),
    .A(_03534_),
    .X(_03566_));
 sg13g2_nand2_1 _09200_ (.Y(_03567_),
    .A(_03565_),
    .B(_03566_));
 sg13g2_a21oi_1 _09201_ (.A1(_03558_),
    .A2(_03560_),
    .Y(_03568_),
    .B1(_03562_));
 sg13g2_xnor2_1 _09202_ (.Y(_03569_),
    .A(_03565_),
    .B(_03566_));
 sg13g2_o21ai_1 _09203_ (.B1(_03567_),
    .Y(_03570_),
    .A1(_03568_),
    .A2(_03569_));
 sg13g2_xnor2_1 _09204_ (.Y(_03571_),
    .A(_03539_),
    .B(_03541_));
 sg13g2_nand2_1 _09205_ (.Y(_03572_),
    .A(_03570_),
    .B(_03571_));
 sg13g2_nand2_1 _09206_ (.Y(_03573_),
    .A(net1609),
    .B(net1596));
 sg13g2_and2_1 _09207_ (.A(net1616),
    .B(net1599),
    .X(_03574_));
 sg13g2_and4_1 _09208_ (.A(net1617),
    .B(net1607),
    .C(net1603),
    .D(net1599),
    .X(_03575_));
 sg13g2_a22oi_1 _09209_ (.Y(_03576_),
    .B1(net1599),
    .B2(net1606),
    .A2(net1603),
    .A1(net1617));
 sg13g2_o21ai_1 _09210_ (.B1(_03573_),
    .Y(_03577_),
    .A1(_03575_),
    .A2(_03576_));
 sg13g2_or3_1 _09211_ (.A(_03573_),
    .B(_03575_),
    .C(_03576_),
    .X(_03578_));
 sg13g2_a22oi_1 _09212_ (.Y(_03579_),
    .B1(net1597),
    .B2(net1614),
    .A2(net1602),
    .A1(net1613));
 sg13g2_a21oi_1 _09213_ (.A1(net1613),
    .A2(_03514_),
    .Y(_03580_),
    .B1(_03579_));
 sg13g2_and3_1 _09214_ (.X(_03581_),
    .A(_03577_),
    .B(_03578_),
    .C(_03580_));
 sg13g2_a21o_1 _09215_ (.A2(_03547_),
    .A1(_03546_),
    .B1(_03552_),
    .X(_03582_));
 sg13g2_and3_1 _09216_ (.X(_03583_),
    .A(_03553_),
    .B(_03581_),
    .C(_03582_));
 sg13g2_nand3_1 _09217_ (.B(_03581_),
    .C(_03582_),
    .A(_03553_),
    .Y(_03584_));
 sg13g2_a21o_1 _09218_ (.A2(_03582_),
    .A1(_03553_),
    .B1(_03581_),
    .X(_03585_));
 sg13g2_nor2b_1 _09219_ (.A(net1610),
    .B_N(net1594),
    .Y(_03586_));
 sg13g2_nor2b_1 _09220_ (.A(_03575_),
    .B_N(_03578_),
    .Y(_03587_));
 sg13g2_nand2_1 _09221_ (.Y(_03588_),
    .A(_03396_),
    .B(net1596));
 sg13g2_xor2_1 _09222_ (.B(_03588_),
    .A(_03587_),
    .X(_03589_));
 sg13g2_nand2_1 _09223_ (.Y(_03590_),
    .A(_03586_),
    .B(_03589_));
 sg13g2_or2_1 _09224_ (.X(_03591_),
    .B(_03589_),
    .A(_03586_));
 sg13g2_and4_1 _09225_ (.A(_03584_),
    .B(_03585_),
    .C(_03590_),
    .D(_03591_),
    .X(_03592_));
 sg13g2_nor2_1 _09226_ (.A(_03583_),
    .B(_03592_),
    .Y(_03593_));
 sg13g2_xnor2_1 _09227_ (.Y(_03594_),
    .A(_03557_),
    .B(_03564_));
 sg13g2_nor2_1 _09228_ (.A(_03593_),
    .B(_03594_),
    .Y(_03595_));
 sg13g2_o21ai_1 _09229_ (.B1(_03590_),
    .Y(_03596_),
    .A1(_03587_),
    .A2(_03588_));
 sg13g2_xor2_1 _09230_ (.B(_03594_),
    .A(_03593_),
    .X(_03597_));
 sg13g2_a21oi_2 _09231_ (.B1(_03595_),
    .Y(_03598_),
    .A2(_03597_),
    .A1(_03596_));
 sg13g2_xnor2_1 _09232_ (.Y(_03599_),
    .A(_03568_),
    .B(_03569_));
 sg13g2_nor2_1 _09233_ (.A(_03598_),
    .B(_03599_),
    .Y(_03600_));
 sg13g2_a21oi_1 _09234_ (.A1(_03577_),
    .A2(_03578_),
    .Y(_03601_),
    .B1(_03580_));
 sg13g2_and2_1 _09235_ (.A(net1613),
    .B(net1597),
    .X(_03602_));
 sg13g2_and4_1 _09236_ (.A(net1617),
    .B(net1606),
    .C(net1601),
    .D(net1596),
    .X(_03603_));
 sg13g2_nand4_1 _09237_ (.B(net1606),
    .C(net1601),
    .A(net1616),
    .Y(_03604_),
    .D(net1596));
 sg13g2_a22oi_1 _09238_ (.Y(_03605_),
    .B1(net1596),
    .B2(net1616),
    .A2(net1601),
    .A1(net1606));
 sg13g2_o21ai_1 _09239_ (.B1(_03524_),
    .Y(_03606_),
    .A1(_03603_),
    .A2(_03605_));
 sg13g2_or3_1 _09240_ (.A(_03524_),
    .B(_03603_),
    .C(_03605_),
    .X(_03607_));
 sg13g2_nand3_1 _09241_ (.B(_03606_),
    .C(_03607_),
    .A(_03602_),
    .Y(_03608_));
 sg13g2_or3_1 _09242_ (.A(_03581_),
    .B(_03601_),
    .C(_03608_),
    .X(_03609_));
 sg13g2_o21ai_1 _09243_ (.B1(_03608_),
    .Y(_03610_),
    .A1(_03581_),
    .A2(_03601_));
 sg13g2_nor2b_1 _09244_ (.A(net1610),
    .B_N(net1604),
    .Y(_03611_));
 sg13g2_o21ai_1 _09245_ (.B1(_03604_),
    .Y(_03612_),
    .A1(_03524_),
    .A2(_03605_));
 sg13g2_nand2_1 _09246_ (.Y(_03613_),
    .A(net1612),
    .B(net1594));
 sg13g2_nand2b_1 _09247_ (.Y(_03614_),
    .B(_03612_),
    .A_N(_03613_));
 sg13g2_xnor2_1 _09248_ (.Y(_03615_),
    .A(_03612_),
    .B(_03613_));
 sg13g2_nand2_1 _09249_ (.Y(_03616_),
    .A(_03611_),
    .B(_03615_));
 sg13g2_xor2_1 _09250_ (.B(_03615_),
    .A(_03611_),
    .X(_03617_));
 sg13g2_nand3_1 _09251_ (.B(_03610_),
    .C(_03617_),
    .A(_03609_),
    .Y(_03618_));
 sg13g2_and2_1 _09252_ (.A(_03609_),
    .B(_03618_),
    .X(_03619_));
 sg13g2_a22oi_1 _09253_ (.Y(_03620_),
    .B1(_03590_),
    .B2(_03591_),
    .A2(_03585_),
    .A1(_03584_));
 sg13g2_nor3_1 _09254_ (.A(_03592_),
    .B(_03619_),
    .C(_03620_),
    .Y(_03621_));
 sg13g2_or3_1 _09255_ (.A(_03592_),
    .B(_03619_),
    .C(_03620_),
    .X(_03622_));
 sg13g2_nand2_1 _09256_ (.Y(_03623_),
    .A(_03614_),
    .B(_03616_));
 sg13g2_o21ai_1 _09257_ (.B1(_03619_),
    .Y(_03624_),
    .A1(_03592_),
    .A2(_03620_));
 sg13g2_and3_1 _09258_ (.X(_03625_),
    .A(_03622_),
    .B(_03623_),
    .C(_03624_));
 sg13g2_nor2_1 _09259_ (.A(_03621_),
    .B(_03625_),
    .Y(_03626_));
 sg13g2_xnor2_1 _09260_ (.Y(_03627_),
    .A(_03596_),
    .B(_03597_));
 sg13g2_or2_1 _09261_ (.X(_03628_),
    .B(_03627_),
    .A(_03626_));
 sg13g2_nor2b_1 _09262_ (.A(net1610),
    .B_N(net1599),
    .Y(_03629_));
 sg13g2_and4_1 _09263_ (.A(net1616),
    .B(net1606),
    .C(net1597),
    .D(net1594),
    .X(_03630_));
 sg13g2_nand4_1 _09264_ (.B(net1606),
    .C(net1597),
    .A(net1616),
    .Y(_03631_),
    .D(net1594));
 sg13g2_nand2_1 _09265_ (.Y(_03632_),
    .A(net1609),
    .B(net1604));
 sg13g2_a22oi_1 _09266_ (.Y(_03633_),
    .B1(net1594),
    .B2(net1616),
    .A2(net1597),
    .A1(net1606));
 sg13g2_nor2_1 _09267_ (.A(_03630_),
    .B(_03633_),
    .Y(_03634_));
 sg13g2_o21ai_1 _09268_ (.B1(_03631_),
    .Y(_03635_),
    .A1(_03632_),
    .A2(_03633_));
 sg13g2_nand2_1 _09269_ (.Y(_03636_),
    .A(net1612),
    .B(net1604));
 sg13g2_nand2b_1 _09270_ (.Y(_03637_),
    .B(_03635_),
    .A_N(_03636_));
 sg13g2_xnor2_1 _09271_ (.Y(_03638_),
    .A(_03635_),
    .B(_03636_));
 sg13g2_nand2_1 _09272_ (.Y(_03639_),
    .A(_03629_),
    .B(_03638_));
 sg13g2_xnor2_1 _09273_ (.Y(_03640_),
    .A(_03629_),
    .B(_03638_));
 sg13g2_a21o_1 _09274_ (.A2(_03607_),
    .A1(_03606_),
    .B1(_03602_),
    .X(_03641_));
 sg13g2_and2_1 _09275_ (.A(_03608_),
    .B(_03641_),
    .X(_03642_));
 sg13g2_nor2b_1 _09276_ (.A(_03640_),
    .B_N(_03642_),
    .Y(_03643_));
 sg13g2_a21o_1 _09277_ (.A2(_03610_),
    .A1(_03609_),
    .B1(_03617_),
    .X(_03644_));
 sg13g2_nand3_1 _09278_ (.B(_03643_),
    .C(_03644_),
    .A(_03618_),
    .Y(_03645_));
 sg13g2_nand2_1 _09279_ (.Y(_03646_),
    .A(_03637_),
    .B(_03639_));
 sg13g2_a21o_1 _09280_ (.A2(_03644_),
    .A1(_03618_),
    .B1(_03643_),
    .X(_03647_));
 sg13g2_nand3_1 _09281_ (.B(_03646_),
    .C(_03647_),
    .A(_03645_),
    .Y(_03648_));
 sg13g2_and2_1 _09282_ (.A(_03645_),
    .B(_03648_),
    .X(_03649_));
 sg13g2_a21oi_1 _09283_ (.A1(_03622_),
    .A2(_03624_),
    .Y(_03650_),
    .B1(_03623_));
 sg13g2_nor3_1 _09284_ (.A(_03625_),
    .B(_03649_),
    .C(_03650_),
    .Y(_03651_));
 sg13g2_o21ai_1 _09285_ (.B1(_03649_),
    .Y(_03652_),
    .A1(_03625_),
    .A2(_03650_));
 sg13g2_nor2b_1 _09286_ (.A(_03651_),
    .B_N(_03652_),
    .Y(_03653_));
 sg13g2_a21o_1 _09287_ (.A2(_03647_),
    .A1(_03645_),
    .B1(_03646_),
    .X(_03654_));
 sg13g2_xnor2_1 _09288_ (.Y(_03655_),
    .A(_03640_),
    .B(_03642_));
 sg13g2_and3_1 _09289_ (.X(_03656_),
    .A(net1609),
    .B(net1604),
    .C(_03574_));
 sg13g2_nand2_1 _09290_ (.Y(_03657_),
    .A(net1612),
    .B(net1599));
 sg13g2_mux2_1 _09291_ (.A0(_03657_),
    .A1(net1612),
    .S(_03656_),
    .X(_03658_));
 sg13g2_nor2b_1 _09292_ (.A(net1610),
    .B_N(net1601),
    .Y(_03659_));
 sg13g2_nor2b_1 _09293_ (.A(_03658_),
    .B_N(_03659_),
    .Y(_03660_));
 sg13g2_xnor2_1 _09294_ (.Y(_03661_),
    .A(_03658_),
    .B(_03659_));
 sg13g2_xnor2_1 _09295_ (.Y(_03662_),
    .A(_03632_),
    .B(_03634_));
 sg13g2_nand2_1 _09296_ (.Y(_03663_),
    .A(_03661_),
    .B(_03662_));
 sg13g2_nand3_1 _09297_ (.B(_03661_),
    .C(_03662_),
    .A(_03655_),
    .Y(_03664_));
 sg13g2_inv_1 _09298_ (.Y(_03665_),
    .A(_03664_));
 sg13g2_a21oi_1 _09299_ (.A1(net1612),
    .A2(_03656_),
    .Y(_03666_),
    .B1(_03660_));
 sg13g2_xor2_1 _09300_ (.B(_03663_),
    .A(_03655_),
    .X(_03667_));
 sg13g2_or2_1 _09301_ (.X(_03668_),
    .B(_03667_),
    .A(_03666_));
 sg13g2_o21ai_1 _09302_ (.B1(_03664_),
    .Y(_03669_),
    .A1(_03666_),
    .A2(_03667_));
 sg13g2_nand3_1 _09303_ (.B(_03654_),
    .C(_03669_),
    .A(_03648_),
    .Y(_03670_));
 sg13g2_a21oi_1 _09304_ (.A1(_03648_),
    .A2(_03654_),
    .Y(_03671_),
    .B1(_03665_));
 sg13g2_nand2_1 _09305_ (.Y(_03672_),
    .A(_03666_),
    .B(_03667_));
 sg13g2_xnor2_1 _09306_ (.Y(_03673_),
    .A(_03661_),
    .B(_03662_));
 sg13g2_a22oi_1 _09307_ (.Y(_03674_),
    .B1(net1599),
    .B2(net1609),
    .A2(net1604),
    .A1(net1616));
 sg13g2_nor2_1 _09308_ (.A(_03656_),
    .B(_03674_),
    .Y(_03675_));
 sg13g2_nor2b_1 _09309_ (.A(net1599),
    .B_N(net1616),
    .Y(_03676_));
 sg13g2_and2_1 _09310_ (.A(net1609),
    .B(net1601),
    .X(_03677_));
 sg13g2_nor2_1 _09311_ (.A(_03574_),
    .B(_03677_),
    .Y(_03678_));
 sg13g2_o21ai_1 _09312_ (.B1(net1597),
    .Y(_03679_),
    .A1(net1612),
    .A2(_03676_));
 sg13g2_nor2_1 _09313_ (.A(_03678_),
    .B(_03679_),
    .Y(_03680_));
 sg13g2_nand2_1 _09314_ (.Y(_03681_),
    .A(_03675_),
    .B(_03680_));
 sg13g2_and3_1 _09315_ (.X(_03682_),
    .A(net1612),
    .B(_03574_),
    .C(_03677_));
 sg13g2_a22oi_1 _09316_ (.Y(_03683_),
    .B1(_03574_),
    .B2(_03677_),
    .A2(net1601),
    .A1(net1612));
 sg13g2_or2_1 _09317_ (.X(_03684_),
    .B(_03683_),
    .A(_03682_));
 sg13g2_nand2b_1 _09318_ (.Y(_03685_),
    .B(net1597),
    .A_N(net1610));
 sg13g2_nor2_1 _09319_ (.A(_03684_),
    .B(_03685_),
    .Y(_03686_));
 sg13g2_and2_1 _09320_ (.A(_03684_),
    .B(_03685_),
    .X(_03687_));
 sg13g2_o21ai_1 _09321_ (.B1(_03681_),
    .Y(_03688_),
    .A1(_03686_),
    .A2(_03687_));
 sg13g2_o21ai_1 _09322_ (.B1(_03688_),
    .Y(_03689_),
    .A1(_03675_),
    .A2(_03680_));
 sg13g2_nand2_1 _09323_ (.Y(_03690_),
    .A(_03673_),
    .B(_03689_));
 sg13g2_nor2_1 _09324_ (.A(_03682_),
    .B(_03686_),
    .Y(_03691_));
 sg13g2_o21ai_1 _09325_ (.B1(_03691_),
    .Y(_03692_),
    .A1(_03673_),
    .A2(_03689_));
 sg13g2_nand4_1 _09326_ (.B(_03672_),
    .C(_03690_),
    .A(_03668_),
    .Y(_03693_),
    .D(_03692_));
 sg13g2_o21ai_1 _09327_ (.B1(_03670_),
    .Y(_03694_),
    .A1(_03671_),
    .A2(_03693_));
 sg13g2_a21oi_2 _09328_ (.B1(_03651_),
    .Y(_03695_),
    .A2(_03694_),
    .A1(_03652_));
 sg13g2_xnor2_1 _09329_ (.Y(_03696_),
    .A(_03626_),
    .B(_03627_));
 sg13g2_o21ai_1 _09330_ (.B1(_03628_),
    .Y(_03697_),
    .A1(_03695_),
    .A2(_03696_));
 sg13g2_xor2_1 _09331_ (.B(_03599_),
    .A(_03598_),
    .X(_03698_));
 sg13g2_a21oi_1 _09332_ (.A1(_03697_),
    .A2(_03698_),
    .Y(_03699_),
    .B1(_03600_));
 sg13g2_xnor2_1 _09333_ (.Y(_03700_),
    .A(_03570_),
    .B(_03571_));
 sg13g2_o21ai_1 _09334_ (.B1(_03572_),
    .Y(_03701_),
    .A1(_03699_),
    .A2(_03700_));
 sg13g2_xor2_1 _09335_ (.B(_03542_),
    .A(_03513_),
    .X(_03702_));
 sg13g2_a21oi_1 _09336_ (.A1(_03701_),
    .A2(_03702_),
    .Y(_03703_),
    .B1(_03543_));
 sg13g2_or2_1 _09337_ (.X(_03704_),
    .B(_03490_),
    .A(_03478_));
 sg13g2_o21ai_1 _09338_ (.B1(_03491_),
    .Y(_03705_),
    .A1(_03510_),
    .A2(_03704_));
 sg13g2_nor2b_1 _09339_ (.A(_03705_),
    .B_N(_03511_),
    .Y(_03706_));
 sg13g2_o21ai_1 _09340_ (.B1(_03511_),
    .Y(_03707_),
    .A1(_03703_),
    .A2(_03705_));
 sg13g2_nand2_1 _09341_ (.Y(_03708_),
    .A(_03477_),
    .B(_03491_));
 sg13g2_xnor2_1 _09342_ (.Y(_03709_),
    .A(_03466_),
    .B(_03708_));
 sg13g2_a21oi_1 _09343_ (.A1(_03707_),
    .A2(_03709_),
    .Y(_03710_),
    .B1(_03493_));
 sg13g2_or2_1 _09344_ (.X(_03711_),
    .B(_03477_),
    .A(_03466_));
 sg13g2_and2_1 _09345_ (.A(_03451_),
    .B(_03463_),
    .X(_03712_));
 sg13g2_xnor2_1 _09346_ (.Y(_03713_),
    .A(_03459_),
    .B(_03712_));
 sg13g2_xor2_1 _09347_ (.B(_03713_),
    .A(_03711_),
    .X(_03714_));
 sg13g2_nand4_1 _09348_ (.B(_03710_),
    .C(_03711_),
    .A(_03459_),
    .Y(_03715_),
    .D(_03712_));
 sg13g2_nand2_1 _09349_ (.Y(_03716_),
    .A(_03385_),
    .B(net1466));
 sg13g2_xnor2_1 _09350_ (.Y(_03717_),
    .A(_03385_),
    .B(net1466));
 sg13g2_o21ai_1 _09351_ (.B1(_03716_),
    .Y(_03718_),
    .A1(_03412_),
    .A2(_03717_));
 sg13g2_or2_1 _09352_ (.X(_03719_),
    .B(_03408_),
    .A(_03380_));
 sg13g2_nor2b_1 _09353_ (.A(_03450_),
    .B_N(_03719_),
    .Y(_03720_));
 sg13g2_a21o_1 _09354_ (.A2(_03719_),
    .A1(_03718_),
    .B1(_03450_),
    .X(_03721_));
 sg13g2_xnor2_1 _09355_ (.Y(_03722_),
    .A(_03382_),
    .B(_03415_));
 sg13g2_inv_1 _09356_ (.Y(_03723_),
    .A(_03722_));
 sg13g2_a21o_1 _09357_ (.A2(_03723_),
    .A1(_03721_),
    .B1(_03449_),
    .X(_03724_));
 sg13g2_a221oi_1 _09358_ (.B2(_03723_),
    .C1(_03449_),
    .B1(_03721_),
    .A1(_03384_),
    .Y(_03725_),
    .A2(_03409_));
 sg13g2_nor3_1 _09359_ (.A(_03447_),
    .B(_03448_),
    .C(_03725_),
    .Y(_03726_));
 sg13g2_nor2_1 _09360_ (.A(_03446_),
    .B(_03726_),
    .Y(_03727_));
 sg13g2_o21ai_1 _09361_ (.B1(_03444_),
    .Y(_03728_),
    .A1(_03446_),
    .A2(_03726_));
 sg13g2_a21o_2 _09362_ (.A2(_03728_),
    .A1(_03445_),
    .B1(_03443_),
    .X(_03729_));
 sg13g2_nand2_1 _09363_ (.Y(_03730_),
    .A(_03442_),
    .B(_03729_));
 sg13g2_nand2_1 _09364_ (.Y(_03731_),
    .A(_03378_),
    .B(_03410_));
 sg13g2_nand3_1 _09365_ (.B(_03729_),
    .C(_03731_),
    .A(_03442_),
    .Y(_03732_));
 sg13g2_and2_1 _09366_ (.A(_03441_),
    .B(_03732_),
    .X(_03733_));
 sg13g2_o21ai_1 _09367_ (.B1(_03447_),
    .Y(_03734_),
    .A1(_03448_),
    .A2(_03725_));
 sg13g2_nand2b_1 _09368_ (.Y(_03735_),
    .B(_03734_),
    .A_N(_03726_));
 sg13g2_xnor2_1 _09369_ (.Y(_03736_),
    .A(_03718_),
    .B(_03720_));
 sg13g2_xnor2_1 _09370_ (.Y(_03737_),
    .A(_03412_),
    .B(_03717_));
 sg13g2_nor2_1 _09371_ (.A(_03736_),
    .B(_03737_),
    .Y(_03738_));
 sg13g2_xnor2_1 _09372_ (.Y(_03739_),
    .A(_03721_),
    .B(_03722_));
 sg13g2_nand2_1 _09373_ (.Y(_03740_),
    .A(_03738_),
    .B(_03739_));
 sg13g2_xor2_1 _09374_ (.B(_03409_),
    .A(_03384_),
    .X(_03741_));
 sg13g2_xnor2_1 _09375_ (.Y(_03742_),
    .A(_03724_),
    .B(_03741_));
 sg13g2_nor2_1 _09376_ (.A(_03740_),
    .B(_03742_),
    .Y(_03743_));
 sg13g2_nor2b_1 _09377_ (.A(_03735_),
    .B_N(_03743_),
    .Y(_03744_));
 sg13g2_nand2_1 _09378_ (.Y(_03745_),
    .A(_03444_),
    .B(_03445_));
 sg13g2_xor2_1 _09379_ (.B(_03745_),
    .A(_03727_),
    .X(_03746_));
 sg13g2_nand3_1 _09380_ (.B(_03445_),
    .C(_03728_),
    .A(_03443_),
    .Y(_03747_));
 sg13g2_and2_1 _09381_ (.A(_03729_),
    .B(_03747_),
    .X(_03748_));
 sg13g2_nand4_1 _09382_ (.B(_03744_),
    .C(_03746_),
    .A(_03729_),
    .Y(_03749_),
    .D(_03747_));
 sg13g2_nor2_1 _09383_ (.A(_03441_),
    .B(_03730_),
    .Y(_03750_));
 sg13g2_and2_1 _09384_ (.A(_03441_),
    .B(_03731_),
    .X(_03751_));
 sg13g2_nand3_1 _09385_ (.B(_03729_),
    .C(_03751_),
    .A(_03442_),
    .Y(_03752_));
 sg13g2_a21o_1 _09386_ (.A2(_03729_),
    .A1(_03442_),
    .B1(_03751_),
    .X(_03753_));
 sg13g2_and3_1 _09387_ (.X(_03754_),
    .A(_03749_),
    .B(_03752_),
    .C(_03753_));
 sg13g2_nand3_1 _09388_ (.B(_03752_),
    .C(_03753_),
    .A(_03749_),
    .Y(_03755_));
 sg13g2_a22oi_1 _09389_ (.Y(_03756_),
    .B1(_03755_),
    .B2(_03733_),
    .A2(_03750_),
    .A1(_03749_));
 sg13g2_a21oi_1 _09390_ (.A1(_03752_),
    .A2(_03753_),
    .Y(_03757_),
    .B1(_03749_));
 sg13g2_nor2_1 _09391_ (.A(_03754_),
    .B(_03757_),
    .Y(_03758_));
 sg13g2_xor2_1 _09392_ (.B(_03746_),
    .A(_03744_),
    .X(_03759_));
 sg13g2_xor2_1 _09393_ (.B(_03743_),
    .A(_03735_),
    .X(_03760_));
 sg13g2_nand2_1 _09394_ (.Y(_03761_),
    .A(_03737_),
    .B(_03739_));
 sg13g2_nor4_1 _09395_ (.A(_03736_),
    .B(_03742_),
    .C(_03760_),
    .D(_03761_),
    .Y(_03762_));
 sg13g2_and3_1 _09396_ (.X(_03763_),
    .A(_03748_),
    .B(_03759_),
    .C(_03762_));
 sg13g2_o21ai_1 _09397_ (.B1(_03763_),
    .Y(_03764_),
    .A1(_03754_),
    .A2(_03757_));
 sg13g2_a21o_1 _09398_ (.A2(_03746_),
    .A1(_03744_),
    .B1(_03748_),
    .X(_03765_));
 sg13g2_nand2_1 _09399_ (.Y(_03766_),
    .A(_03749_),
    .B(_03765_));
 sg13g2_and2_2 _09400_ (.A(_03756_),
    .B(_03764_),
    .X(_03767_));
 sg13g2_xnor2_1 _09401_ (.Y(_03768_),
    .A(_03695_),
    .B(_03696_));
 sg13g2_xor2_1 _09402_ (.B(_03694_),
    .A(_03653_),
    .X(_03769_));
 sg13g2_nand2_1 _09403_ (.Y(_03770_),
    .A(net1465),
    .B(_03768_));
 sg13g2_o21ai_1 _09404_ (.B1(_03770_),
    .Y(_03771_),
    .A1(net1465),
    .A2(_03769_));
 sg13g2_a22oi_1 _09405_ (.Y(_03772_),
    .B1(_03418_),
    .B2(_03431_),
    .A2(_03405_),
    .A1(_03389_));
 sg13g2_nor2b_1 _09406_ (.A(_03429_),
    .B_N(_03438_),
    .Y(_03773_));
 sg13g2_a21o_1 _09407_ (.A2(_03435_),
    .A1(_03402_),
    .B1(_03773_),
    .X(_03774_));
 sg13g2_a221oi_1 _09408_ (.B2(_03431_),
    .C1(_03774_),
    .B1(_03418_),
    .A1(_03389_),
    .Y(_03775_),
    .A2(_03405_));
 sg13g2_inv_2 _09409_ (.Y(_03776_),
    .A(_03775_));
 sg13g2_nor3_1 _09410_ (.A(net1420),
    .B(_03771_),
    .C(_03776_),
    .Y(_03777_));
 sg13g2_a21oi_1 _09411_ (.A1(_03767_),
    .A2(_03777_),
    .Y(_03778_),
    .B1(net1492));
 sg13g2_o21ai_1 _09412_ (.B1(net1537),
    .Y(_03779_),
    .A1(\u_tiny_nn_top.data_i_q[0] ),
    .A2(net1768));
 sg13g2_o21ai_1 _09413_ (.B1(_03377_),
    .Y(_00334_),
    .A1(_03778_),
    .A2(_03779_));
 sg13g2_nand2_1 _09414_ (.Y(_03780_),
    .A(net968),
    .B(net1538));
 sg13g2_xnor2_1 _09415_ (.Y(_03781_),
    .A(_03697_),
    .B(_03698_));
 sg13g2_mux2_1 _09416_ (.A0(_03768_),
    .A1(_03781_),
    .S(net1465),
    .X(_03782_));
 sg13g2_nor3_1 _09417_ (.A(net1420),
    .B(_03776_),
    .C(_03782_),
    .Y(_03783_));
 sg13g2_a21oi_1 _09418_ (.A1(_03767_),
    .A2(_03783_),
    .Y(_03784_),
    .B1(net1492));
 sg13g2_o21ai_1 _09419_ (.B1(net1537),
    .Y(_03785_),
    .A1(net1850),
    .A2(net1768));
 sg13g2_o21ai_1 _09420_ (.B1(_03780_),
    .Y(_00335_),
    .A1(_03784_),
    .A2(_03785_));
 sg13g2_nand2_1 _09421_ (.Y(_03786_),
    .A(net992),
    .B(net1538));
 sg13g2_xnor2_1 _09422_ (.Y(_03787_),
    .A(_03699_),
    .B(_03700_));
 sg13g2_mux2_1 _09423_ (.A0(_03781_),
    .A1(_03787_),
    .S(net1465),
    .X(_03788_));
 sg13g2_nor3_1 _09424_ (.A(net1420),
    .B(_03776_),
    .C(_03788_),
    .Y(_03789_));
 sg13g2_a21oi_1 _09425_ (.A1(_03767_),
    .A2(_03789_),
    .Y(_03790_),
    .B1(net1492));
 sg13g2_o21ai_1 _09426_ (.B1(net1537),
    .Y(_03791_),
    .A1(\u_tiny_nn_top.data_i_q[2] ),
    .A2(net1768));
 sg13g2_o21ai_1 _09427_ (.B1(_03786_),
    .Y(_00336_),
    .A1(_03790_),
    .A2(_03791_));
 sg13g2_nand2_1 _09428_ (.Y(_03792_),
    .A(net986),
    .B(net1538));
 sg13g2_xnor2_1 _09429_ (.Y(_03793_),
    .A(_03701_),
    .B(_03702_));
 sg13g2_mux2_1 _09430_ (.A0(_03787_),
    .A1(_03793_),
    .S(net1466),
    .X(_03794_));
 sg13g2_nor3_1 _09431_ (.A(net1420),
    .B(_03776_),
    .C(_03794_),
    .Y(_03795_));
 sg13g2_a21oi_1 _09432_ (.A1(_03767_),
    .A2(_03795_),
    .Y(_03796_),
    .B1(net1492));
 sg13g2_o21ai_1 _09433_ (.B1(net1537),
    .Y(_03797_),
    .A1(net1846),
    .A2(net1768));
 sg13g2_o21ai_1 _09434_ (.B1(_03792_),
    .Y(_00337_),
    .A1(_03796_),
    .A2(_03797_));
 sg13g2_nand2_1 _09435_ (.Y(_03798_),
    .A(net963),
    .B(net1539));
 sg13g2_xnor2_1 _09436_ (.Y(_03799_),
    .A(_03703_),
    .B(_03706_));
 sg13g2_inv_1 _09437_ (.Y(_03800_),
    .A(_03799_));
 sg13g2_mux2_1 _09438_ (.A0(_03793_),
    .A1(_03800_),
    .S(net1465),
    .X(_03801_));
 sg13g2_nor3_1 _09439_ (.A(net1420),
    .B(_03776_),
    .C(_03801_),
    .Y(_03802_));
 sg13g2_a21oi_1 _09440_ (.A1(_03767_),
    .A2(_03802_),
    .Y(_03803_),
    .B1(net1492));
 sg13g2_o21ai_1 _09441_ (.B1(net1536),
    .Y(_03804_),
    .A1(net1844),
    .A2(net1767));
 sg13g2_o21ai_1 _09442_ (.B1(_03798_),
    .Y(_00338_),
    .A1(_03803_),
    .A2(_03804_));
 sg13g2_nand2_1 _09443_ (.Y(_03805_),
    .A(net939),
    .B(_03375_));
 sg13g2_xnor2_1 _09444_ (.Y(_03806_),
    .A(_03707_),
    .B(_03709_));
 sg13g2_nand2_1 _09445_ (.Y(_03807_),
    .A(net1465),
    .B(_03806_));
 sg13g2_o21ai_1 _09446_ (.B1(_03807_),
    .Y(_03808_),
    .A1(net1465),
    .A2(_03799_));
 sg13g2_nor3_1 _09447_ (.A(net1420),
    .B(_03776_),
    .C(_03808_),
    .Y(_03809_));
 sg13g2_a21oi_1 _09448_ (.A1(_03767_),
    .A2(_03809_),
    .Y(_03810_),
    .B1(net1492));
 sg13g2_o21ai_1 _09449_ (.B1(net1536),
    .Y(_03811_),
    .A1(net1841),
    .A2(net1767));
 sg13g2_o21ai_1 _09450_ (.B1(_03805_),
    .Y(_00339_),
    .A1(_03810_),
    .A2(_03811_));
 sg13g2_nand2_1 _09451_ (.Y(_03812_),
    .A(net935),
    .B(net1539));
 sg13g2_nor2b_1 _09452_ (.A(net1465),
    .B_N(_03806_),
    .Y(_03813_));
 sg13g2_xnor2_1 _09453_ (.Y(_03814_),
    .A(_03710_),
    .B(_03714_));
 sg13g2_nor4_1 _09454_ (.A(net1420),
    .B(_03776_),
    .C(_03813_),
    .D(_03814_),
    .Y(_03815_));
 sg13g2_a21oi_1 _09455_ (.A1(_03767_),
    .A2(_03815_),
    .Y(_03816_),
    .B1(net1492));
 sg13g2_o21ai_1 _09456_ (.B1(net1536),
    .Y(_03817_),
    .A1(net1837),
    .A2(net1767));
 sg13g2_o21ai_1 _09457_ (.B1(_03812_),
    .Y(_00340_),
    .A1(_03816_),
    .A2(_03817_));
 sg13g2_o21ai_1 _09458_ (.B1(_03772_),
    .Y(_03818_),
    .A1(_03441_),
    .A2(_03730_));
 sg13g2_inv_1 _09459_ (.Y(_03819_),
    .A(_03818_));
 sg13g2_a221oi_1 _09460_ (.B2(_03733_),
    .C1(_03774_),
    .B1(_03755_),
    .A1(_03749_),
    .Y(_03820_),
    .A2(net1420));
 sg13g2_and2_1 _09461_ (.A(_03764_),
    .B(_03820_),
    .X(_03821_));
 sg13g2_nand2b_1 _09462_ (.Y(_03822_),
    .B(_03821_),
    .A_N(_03737_));
 sg13g2_a21oi_1 _09463_ (.A1(_03819_),
    .A2(_03822_),
    .Y(_03823_),
    .B1(_03440_));
 sg13g2_o21ai_1 _09464_ (.B1(net1537),
    .Y(_03824_),
    .A1(net1834),
    .A2(net1767));
 sg13g2_nand2_1 _09465_ (.Y(_03825_),
    .A(net1055),
    .B(net1539));
 sg13g2_o21ai_1 _09466_ (.B1(_03825_),
    .Y(_00341_),
    .A1(_03823_),
    .A2(_03824_));
 sg13g2_xnor2_1 _09467_ (.Y(_03826_),
    .A(_03736_),
    .B(_03737_));
 sg13g2_a21oi_1 _09468_ (.A1(_03821_),
    .A2(_03826_),
    .Y(_03827_),
    .B1(_03818_));
 sg13g2_a21oi_1 _09469_ (.A1(_00644_),
    .A2(net1789),
    .Y(_03828_),
    .B1(net1539));
 sg13g2_o21ai_1 _09470_ (.B1(_03828_),
    .Y(_03829_),
    .A1(net1491),
    .A2(_03827_));
 sg13g2_o21ai_1 _09471_ (.B1(_03829_),
    .Y(_00342_),
    .A1(_00696_),
    .A2(_03376_));
 sg13g2_xnor2_1 _09472_ (.Y(_03830_),
    .A(_03738_),
    .B(_03739_));
 sg13g2_a21oi_1 _09473_ (.A1(_03821_),
    .A2(_03830_),
    .Y(_03831_),
    .B1(_03818_));
 sg13g2_a21oi_1 _09474_ (.A1(net1774),
    .A2(net1789),
    .Y(_03832_),
    .B1(net1539));
 sg13g2_o21ai_1 _09475_ (.B1(_03832_),
    .Y(_03833_),
    .A1(net1491),
    .A2(_03831_));
 sg13g2_o21ai_1 _09476_ (.B1(_03833_),
    .Y(_00343_),
    .A1(_00698_),
    .A2(net1537));
 sg13g2_xnor2_1 _09477_ (.Y(_03834_),
    .A(_03740_),
    .B(_03742_));
 sg13g2_a21oi_1 _09478_ (.A1(_03821_),
    .A2(_03834_),
    .Y(_03835_),
    .B1(_03818_));
 sg13g2_a21oi_1 _09479_ (.A1(net1776),
    .A2(net1789),
    .Y(_03836_),
    .B1(net1538));
 sg13g2_o21ai_1 _09480_ (.B1(_03836_),
    .Y(_03837_),
    .A1(net1491),
    .A2(_03835_));
 sg13g2_o21ai_1 _09481_ (.B1(_03837_),
    .Y(_00344_),
    .A1(_00697_),
    .A2(net1536));
 sg13g2_a21oi_1 _09482_ (.A1(_03760_),
    .A2(_03820_),
    .Y(_03838_),
    .B1(_03818_));
 sg13g2_a21oi_1 _09483_ (.A1(net1778),
    .A2(net1789),
    .Y(_03839_),
    .B1(net1538));
 sg13g2_o21ai_1 _09484_ (.B1(_03839_),
    .Y(_03840_),
    .A1(net1491),
    .A2(_03838_));
 sg13g2_o21ai_1 _09485_ (.B1(_03840_),
    .Y(_00345_),
    .A1(_00700_),
    .A2(net1536));
 sg13g2_nand2_1 _09486_ (.Y(_03841_),
    .A(net947),
    .B(net1539));
 sg13g2_nand2b_1 _09487_ (.Y(_03842_),
    .B(_03820_),
    .A_N(_03759_));
 sg13g2_a21oi_1 _09488_ (.A1(_03819_),
    .A2(_03842_),
    .Y(_03843_),
    .B1(net1491));
 sg13g2_o21ai_1 _09489_ (.B1(net1537),
    .Y(_03844_),
    .A1(net1828),
    .A2(net1767));
 sg13g2_o21ai_1 _09490_ (.B1(_03841_),
    .Y(_00346_),
    .A1(_03843_),
    .A2(_03844_));
 sg13g2_a21oi_1 _09491_ (.A1(_03766_),
    .A2(_03820_),
    .Y(_03845_),
    .B1(_03818_));
 sg13g2_a21oi_1 _09492_ (.A1(net1782),
    .A2(net1789),
    .Y(_03846_),
    .B1(net1538));
 sg13g2_o21ai_1 _09493_ (.B1(_03846_),
    .Y(_03847_),
    .A1(net1491),
    .A2(_03845_));
 sg13g2_o21ai_1 _09494_ (.B1(_03847_),
    .Y(_00347_),
    .A1(_00702_),
    .A2(net1536));
 sg13g2_a21oi_1 _09495_ (.A1(_03758_),
    .A2(_03820_),
    .Y(_03848_),
    .B1(_03818_));
 sg13g2_a21oi_1 _09496_ (.A1(net1784),
    .A2(net1789),
    .Y(_03849_),
    .B1(net1538));
 sg13g2_o21ai_1 _09497_ (.B1(_03849_),
    .Y(_03850_),
    .A1(net1491),
    .A2(_03848_));
 sg13g2_o21ai_1 _09498_ (.B1(_03850_),
    .Y(_00348_),
    .A1(_00701_),
    .A2(net1536));
 sg13g2_nand2_1 _09499_ (.Y(_03851_),
    .A(net1030),
    .B(net1539));
 sg13g2_xor2_1 _09500_ (.B(_03430_),
    .A(_03404_),
    .X(_03852_));
 sg13g2_a21oi_1 _09501_ (.A1(_03819_),
    .A2(_03852_),
    .Y(_03853_),
    .B1(net1491));
 sg13g2_o21ai_1 _09502_ (.B1(net1536),
    .Y(_03854_),
    .A1(net1825),
    .A2(net1767));
 sg13g2_o21ai_1 _09503_ (.B1(_03851_),
    .Y(_00349_),
    .A1(_03853_),
    .A2(_03854_));
 sg13g2_mux2_2 _09504_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[2][8] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[3][8] ),
    .S(net1715),
    .X(_03855_));
 sg13g2_mux2_2 _09505_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[2][10] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[3][10] ),
    .S(net1710),
    .X(_03856_));
 sg13g2_mux2_2 _09506_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[2][14] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[3][14] ),
    .S(net1715),
    .X(_03857_));
 sg13g2_mux2_2 _09507_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[2][7] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[3][7] ),
    .S(net1713),
    .X(_03858_));
 sg13g2_mux2_1 _09508_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[2][11] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[3][11] ),
    .S(net1713),
    .X(_03859_));
 sg13g2_mux2_1 _09509_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[2][12] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[3][12] ),
    .S(net1713),
    .X(_03860_));
 sg13g2_mux2_2 _09510_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[2][13] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[3][13] ),
    .S(net1710),
    .X(_03861_));
 sg13g2_mux2_2 _09511_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[2][9] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[3][9] ),
    .S(net1710),
    .X(_03862_));
 sg13g2_nor4_1 _09512_ (.A(_03855_),
    .B(_03856_),
    .C(_03859_),
    .D(_03860_),
    .Y(_03863_));
 sg13g2_nor4_1 _09513_ (.A(_03857_),
    .B(_03858_),
    .C(_03861_),
    .D(_03862_),
    .Y(_03864_));
 sg13g2_nand2_1 _09514_ (.Y(_03865_),
    .A(_03863_),
    .B(_03864_));
 sg13g2_mux2_1 _09515_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[2][3] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[3][3] ),
    .S(net1708),
    .X(_03866_));
 sg13g2_mux2_1 _09516_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[2][6] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[3][6] ),
    .S(net1708),
    .X(_03867_));
 sg13g2_mux2_1 _09517_ (.A0(_00687_),
    .A1(_00688_),
    .S(net1708),
    .X(_03868_));
 sg13g2_nor3_1 _09518_ (.A(net1592),
    .B(net1590),
    .C(net1588),
    .Y(_03869_));
 sg13g2_mux2_2 _09519_ (.A0(_00685_),
    .A1(_00686_),
    .S(net1707),
    .X(_03870_));
 sg13g2_mux2_2 _09520_ (.A0(_00046_),
    .A1(_00045_),
    .S(net1707),
    .X(_03871_));
 sg13g2_mux2_1 _09521_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[2][0] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[3][0] ),
    .S(net1706),
    .X(_03872_));
 sg13g2_nor2_1 _09522_ (.A(_03870_),
    .B(net1587),
    .Y(_03873_));
 sg13g2_nand2_1 _09523_ (.Y(_03874_),
    .A(_00049_),
    .B(net1707));
 sg13g2_mux2_2 _09524_ (.A0(_00689_),
    .A1(_00690_),
    .S(net1707),
    .X(_03875_));
 sg13g2_o21ai_1 _09525_ (.B1(_03874_),
    .Y(_03876_),
    .A1(_00689_),
    .A2(net1707));
 sg13g2_nand2b_1 _09526_ (.Y(_03877_),
    .B(net1707),
    .A_N(_00043_));
 sg13g2_o21ai_1 _09527_ (.B1(_03877_),
    .Y(_03878_),
    .A1(_00044_),
    .A2(net1707));
 sg13g2_mux2_2 _09528_ (.A0(_00044_),
    .A1(_00043_),
    .S(net1707),
    .X(_03879_));
 sg13g2_nand4_1 _09529_ (.B(_03873_),
    .C(_03876_),
    .A(_03869_),
    .Y(_03880_),
    .D(_03879_));
 sg13g2_mux2_1 _09530_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[2][15] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[3][15] ),
    .S(net1715),
    .X(_03881_));
 sg13g2_nor2_1 _09531_ (.A(_03880_),
    .B(_03881_),
    .Y(_03882_));
 sg13g2_mux2_2 _09532_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][8] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][8] ),
    .S(net1710),
    .X(_03883_));
 sg13g2_mux2_2 _09533_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][12] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][12] ),
    .S(net1697),
    .X(_03884_));
 sg13g2_mux2_2 _09534_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][11] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][11] ),
    .S(net1709),
    .X(_03885_));
 sg13g2_mux2_2 _09535_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][14] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][14] ),
    .S(net1715),
    .X(_03886_));
 sg13g2_mux2_2 _09536_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][7] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][7] ),
    .S(net1709),
    .X(_03887_));
 sg13g2_mux2_2 _09537_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][9] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][9] ),
    .S(net1697),
    .X(_03888_));
 sg13g2_mux2_2 _09538_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][13] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][13] ),
    .S(net1709),
    .X(_03889_));
 sg13g2_mux2_2 _09539_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][10] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][10] ),
    .S(net1709),
    .X(_03890_));
 sg13g2_nor4_1 _09540_ (.A(_03883_),
    .B(_03884_),
    .C(_03885_),
    .D(_03889_),
    .Y(_03891_));
 sg13g2_nor4_1 _09541_ (.A(_03886_),
    .B(_03887_),
    .C(_03888_),
    .D(_03890_),
    .Y(_03892_));
 sg13g2_nand2_1 _09542_ (.Y(_03893_),
    .A(_03891_),
    .B(_03892_));
 sg13g2_mux2_1 _09543_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][3] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][3] ),
    .S(net1695),
    .X(_03894_));
 sg13g2_mux2_1 _09544_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][6] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][6] ),
    .S(net1708),
    .X(_03895_));
 sg13g2_mux2_1 _09545_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][1] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][1] ),
    .S(net1706),
    .X(_03896_));
 sg13g2_nor3_1 _09546_ (.A(net1585),
    .B(net1584),
    .C(net1582),
    .Y(_03897_));
 sg13g2_mux2_1 _09547_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][2] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][2] ),
    .S(net1694),
    .X(_03898_));
 sg13g2_mux2_1 _09548_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][0] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][0] ),
    .S(net1706),
    .X(_03899_));
 sg13g2_mux2_1 _09549_ (.A0(_00683_),
    .A1(_00684_),
    .S(net1706),
    .X(_03900_));
 sg13g2_mux2_2 _09550_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][5] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][5] ),
    .S(net1694),
    .X(_03901_));
 sg13g2_mux2_2 _09551_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][4] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][4] ),
    .S(net1695),
    .X(_03902_));
 sg13g2_nor4_1 _09552_ (.A(net1580),
    .B(net1577),
    .C(net1576),
    .D(_03902_),
    .Y(_03903_));
 sg13g2_nand2_2 _09553_ (.Y(_03904_),
    .A(_03897_),
    .B(_03903_));
 sg13g2_mux2_1 _09554_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][15] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][15] ),
    .S(net1709),
    .X(_03905_));
 sg13g2_or2_1 _09555_ (.X(_03906_),
    .B(_03905_),
    .A(_03904_));
 sg13g2_nand2b_1 _09556_ (.Y(_03907_),
    .B(_03906_),
    .A_N(_03893_));
 sg13g2_o21ai_1 _09557_ (.B1(_03907_),
    .Y(_03908_),
    .A1(_03865_),
    .A2(_03882_));
 sg13g2_nand4_1 _09558_ (.B(_03884_),
    .C(_03885_),
    .A(_03883_),
    .Y(_03909_),
    .D(_03889_));
 sg13g2_nand4_1 _09559_ (.B(_03887_),
    .C(_03888_),
    .A(_03886_),
    .Y(_03910_),
    .D(_03890_));
 sg13g2_nor2_1 _09560_ (.A(_03909_),
    .B(_03910_),
    .Y(_03911_));
 sg13g2_nand4_1 _09561_ (.B(_03856_),
    .C(_03859_),
    .A(_03855_),
    .Y(_03912_),
    .D(_03860_));
 sg13g2_nand4_1 _09562_ (.B(_03858_),
    .C(_03861_),
    .A(_03857_),
    .Y(_03913_),
    .D(_03862_));
 sg13g2_nor2_1 _09563_ (.A(_03912_),
    .B(_03913_),
    .Y(_03914_));
 sg13g2_inv_1 _09564_ (.Y(_03915_),
    .A(_03914_));
 sg13g2_a221oi_1 _09565_ (.B2(_03880_),
    .C1(net1650),
    .B1(_03914_),
    .A1(_03904_),
    .Y(_03916_),
    .A2(_03911_));
 sg13g2_nor2b_2 _09566_ (.A(_03908_),
    .B_N(_03916_),
    .Y(_03917_));
 sg13g2_nor2_2 _09567_ (.A(_03857_),
    .B(_03886_),
    .Y(_03918_));
 sg13g2_nand2_1 _09568_ (.Y(_03919_),
    .A(_03857_),
    .B(_03886_));
 sg13g2_xnor2_1 _09569_ (.Y(_03920_),
    .A(_03861_),
    .B(_03889_));
 sg13g2_or2_1 _09570_ (.X(_03921_),
    .B(_03884_),
    .A(_03860_));
 sg13g2_nand2_1 _09571_ (.Y(_03922_),
    .A(_03860_),
    .B(_03884_));
 sg13g2_and2_1 _09572_ (.A(_03859_),
    .B(_03885_),
    .X(_03923_));
 sg13g2_xnor2_1 _09573_ (.Y(_03924_),
    .A(_03859_),
    .B(_03885_));
 sg13g2_nor2_1 _09574_ (.A(_03856_),
    .B(_03890_),
    .Y(_03925_));
 sg13g2_and2_1 _09575_ (.A(_03862_),
    .B(_03888_),
    .X(_03926_));
 sg13g2_nand2_1 _09576_ (.Y(_03927_),
    .A(_03855_),
    .B(_03883_));
 sg13g2_nand2_2 _09577_ (.Y(_03928_),
    .A(net1591),
    .B(net1584));
 sg13g2_xor2_1 _09578_ (.B(_03928_),
    .A(net1576),
    .X(_03929_));
 sg13g2_xnor2_1 _09579_ (.Y(_03930_),
    .A(_03876_),
    .B(_03929_));
 sg13g2_nand3_1 _09580_ (.B(net1576),
    .C(net1575),
    .A(_03867_),
    .Y(_03931_));
 sg13g2_nand2_1 _09581_ (.Y(_03932_),
    .A(_03875_),
    .B(net1584));
 sg13g2_a21o_1 _09582_ (.A2(net1576),
    .A1(net1591),
    .B1(net1575),
    .X(_03933_));
 sg13g2_nand2_1 _09583_ (.Y(_03934_),
    .A(_03931_),
    .B(_03933_));
 sg13g2_o21ai_1 _09584_ (.B1(_03931_),
    .Y(_03935_),
    .A1(_03932_),
    .A2(_03934_));
 sg13g2_nand2b_1 _09585_ (.Y(_03936_),
    .B(_03935_),
    .A_N(_03930_));
 sg13g2_xnor2_1 _09586_ (.Y(_03937_),
    .A(_03930_),
    .B(_03935_));
 sg13g2_nand3_1 _09587_ (.B(net1585),
    .C(net1575),
    .A(net1591),
    .Y(_03938_));
 sg13g2_and2_1 _09588_ (.A(_03875_),
    .B(_03901_),
    .X(_03939_));
 sg13g2_inv_1 _09589_ (.Y(_03940_),
    .A(_03939_));
 sg13g2_a21o_1 _09590_ (.A2(net1575),
    .A1(net1591),
    .B1(net1585),
    .X(_03941_));
 sg13g2_nand2_1 _09591_ (.Y(_03942_),
    .A(_03938_),
    .B(_03941_));
 sg13g2_o21ai_1 _09592_ (.B1(_03938_),
    .Y(_03943_),
    .A1(_03940_),
    .A2(_03942_));
 sg13g2_xor2_1 _09593_ (.B(_03934_),
    .A(_03932_),
    .X(_03944_));
 sg13g2_and2_1 _09594_ (.A(_03943_),
    .B(_03944_),
    .X(_03945_));
 sg13g2_or2_1 _09595_ (.X(_03946_),
    .B(_03944_),
    .A(_03943_));
 sg13g2_nand2b_1 _09596_ (.Y(_03947_),
    .B(_03946_),
    .A_N(_03945_));
 sg13g2_a21o_1 _09597_ (.A2(_03946_),
    .A1(_03868_),
    .B1(_03945_),
    .X(_03948_));
 sg13g2_nand2_1 _09598_ (.Y(_03949_),
    .A(_03937_),
    .B(_03948_));
 sg13g2_xor2_1 _09599_ (.B(_03948_),
    .A(_03937_),
    .X(_03950_));
 sg13g2_nand3_1 _09600_ (.B(net1586),
    .C(net1580),
    .A(net1590),
    .Y(_03951_));
 sg13g2_nand2_1 _09601_ (.Y(_03952_),
    .A(_03875_),
    .B(net1575));
 sg13g2_a21o_1 _09602_ (.A2(net1586),
    .A1(net1590),
    .B1(net1580),
    .X(_03953_));
 sg13g2_nand2_1 _09603_ (.Y(_03954_),
    .A(_03951_),
    .B(_03953_));
 sg13g2_o21ai_1 _09604_ (.B1(_03951_),
    .Y(_03955_),
    .A1(_03952_),
    .A2(_03954_));
 sg13g2_xnor2_1 _09605_ (.Y(_03956_),
    .A(_03939_),
    .B(_03942_));
 sg13g2_nand2_1 _09606_ (.Y(_03957_),
    .A(_03955_),
    .B(_03956_));
 sg13g2_nand3_1 _09607_ (.B(net1589),
    .C(net1584),
    .A(net1593),
    .Y(_03958_));
 sg13g2_a21o_1 _09608_ (.A2(net1584),
    .A1(net1589),
    .B1(net1593),
    .X(_03959_));
 sg13g2_nand2_1 _09609_ (.Y(_03960_),
    .A(_03958_),
    .B(_03959_));
 sg13g2_xnor2_1 _09610_ (.Y(_03961_),
    .A(_03955_),
    .B(_03956_));
 sg13g2_o21ai_1 _09611_ (.B1(_03957_),
    .Y(_03962_),
    .A1(_03960_),
    .A2(_03961_));
 sg13g2_xnor2_1 _09612_ (.Y(_03963_),
    .A(net1589),
    .B(_03947_));
 sg13g2_nand2_1 _09613_ (.Y(_03964_),
    .A(_03962_),
    .B(_03963_));
 sg13g2_xnor2_1 _09614_ (.Y(_03965_),
    .A(_03962_),
    .B(_03963_));
 sg13g2_o21ai_1 _09615_ (.B1(_03964_),
    .Y(_03966_),
    .A1(_03958_),
    .A2(_03965_));
 sg13g2_nand2_1 _09616_ (.Y(_03967_),
    .A(_03950_),
    .B(_03966_));
 sg13g2_or2_1 _09617_ (.X(_03968_),
    .B(net1584),
    .A(net1591));
 sg13g2_nand3_1 _09618_ (.B(_03939_),
    .C(_03968_),
    .A(_03928_),
    .Y(_03969_));
 sg13g2_o21ai_1 _09619_ (.B1(_03968_),
    .Y(_03970_),
    .A1(_03901_),
    .A2(_03928_));
 sg13g2_o21ai_1 _09620_ (.B1(_03970_),
    .Y(_03971_),
    .A1(_03876_),
    .A2(_03929_));
 sg13g2_nand3_1 _09621_ (.B(_03969_),
    .C(_03971_),
    .A(_03936_),
    .Y(_03972_));
 sg13g2_or2_1 _09622_ (.X(_03973_),
    .B(_03972_),
    .A(_03949_));
 sg13g2_xor2_1 _09623_ (.B(_03972_),
    .A(_03949_),
    .X(_03974_));
 sg13g2_nand3_1 _09624_ (.B(_03966_),
    .C(_03974_),
    .A(_03950_),
    .Y(_03975_));
 sg13g2_xor2_1 _09625_ (.B(_03965_),
    .A(_03958_),
    .X(_03976_));
 sg13g2_nand3_1 _09626_ (.B(net1582),
    .C(net1580),
    .A(net1591),
    .Y(_03977_));
 sg13g2_nand2_1 _09627_ (.Y(_03978_),
    .A(_03875_),
    .B(net1586));
 sg13g2_a21o_1 _09628_ (.A2(net1580),
    .A1(net1590),
    .B1(net1582),
    .X(_03979_));
 sg13g2_nand2_1 _09629_ (.Y(_03980_),
    .A(_03977_),
    .B(_03979_));
 sg13g2_o21ai_1 _09630_ (.B1(_03977_),
    .Y(_03981_),
    .A1(_03978_),
    .A2(_03980_));
 sg13g2_xor2_1 _09631_ (.B(_03954_),
    .A(_03952_),
    .X(_03982_));
 sg13g2_nand2_1 _09632_ (.Y(_03983_),
    .A(_03981_),
    .B(_03982_));
 sg13g2_nand2_1 _09633_ (.Y(_03984_),
    .A(net1593),
    .B(_03895_));
 sg13g2_nand2_1 _09634_ (.Y(_03985_),
    .A(net1589),
    .B(net1576));
 sg13g2_nor2_1 _09635_ (.A(_03984_),
    .B(_03985_),
    .Y(_03986_));
 sg13g2_xor2_1 _09636_ (.B(_03985_),
    .A(_03984_),
    .X(_03987_));
 sg13g2_xnor2_1 _09637_ (.Y(_03988_),
    .A(_03871_),
    .B(_03987_));
 sg13g2_inv_1 _09638_ (.Y(_03989_),
    .A(_03988_));
 sg13g2_xnor2_1 _09639_ (.Y(_03990_),
    .A(_03981_),
    .B(_03982_));
 sg13g2_o21ai_1 _09640_ (.B1(_03983_),
    .Y(_03991_),
    .A1(_03989_),
    .A2(_03990_));
 sg13g2_xor2_1 _09641_ (.B(_03961_),
    .A(_03960_),
    .X(_03992_));
 sg13g2_nand2_1 _09642_ (.Y(_03993_),
    .A(_03991_),
    .B(_03992_));
 sg13g2_a21oi_1 _09643_ (.A1(_03870_),
    .A2(_03987_),
    .Y(_03994_),
    .B1(_03986_));
 sg13g2_xnor2_1 _09644_ (.Y(_03995_),
    .A(_03991_),
    .B(_03992_));
 sg13g2_o21ai_1 _09645_ (.B1(_03993_),
    .Y(_03996_),
    .A1(_03994_),
    .A2(_03995_));
 sg13g2_nand2_1 _09646_ (.Y(_03997_),
    .A(_03976_),
    .B(_03996_));
 sg13g2_xor2_1 _09647_ (.B(_03966_),
    .A(_03950_),
    .X(_03998_));
 sg13g2_nand2b_1 _09648_ (.Y(_03999_),
    .B(_03998_),
    .A_N(_03997_));
 sg13g2_xor2_1 _09649_ (.B(_03996_),
    .A(_03976_),
    .X(_04000_));
 sg13g2_inv_1 _09650_ (.Y(_04001_),
    .A(_04000_));
 sg13g2_xor2_1 _09651_ (.B(_03995_),
    .A(_03994_),
    .X(_04002_));
 sg13g2_and2_1 _09652_ (.A(net1591),
    .B(net1577),
    .X(_04003_));
 sg13g2_nand3_1 _09653_ (.B(net1582),
    .C(net1578),
    .A(net1590),
    .Y(_04004_));
 sg13g2_a21o_1 _09654_ (.A2(net1583),
    .A1(net1590),
    .B1(net1578),
    .X(_04005_));
 sg13g2_and4_1 _09655_ (.A(_03875_),
    .B(net1580),
    .C(_04004_),
    .D(_04005_),
    .X(_04006_));
 sg13g2_a21o_1 _09656_ (.A2(_04003_),
    .A1(net1582),
    .B1(_04006_),
    .X(_04007_));
 sg13g2_xor2_1 _09657_ (.B(_03980_),
    .A(_03978_),
    .X(_04008_));
 sg13g2_xnor2_1 _09658_ (.Y(_04009_),
    .A(_04007_),
    .B(_04008_));
 sg13g2_nand2_1 _09659_ (.Y(_04010_),
    .A(_03870_),
    .B(_03895_));
 sg13g2_nand2_1 _09660_ (.Y(_04011_),
    .A(net1593),
    .B(_03902_));
 sg13g2_nor2_1 _09661_ (.A(_03985_),
    .B(_04011_),
    .Y(_04012_));
 sg13g2_a22oi_1 _09662_ (.Y(_04013_),
    .B1(_03902_),
    .B2(net1589),
    .A2(_03901_),
    .A1(net1593));
 sg13g2_nor2_1 _09663_ (.A(_04012_),
    .B(_04013_),
    .Y(_04014_));
 sg13g2_nor2b_1 _09664_ (.A(_04010_),
    .B_N(_04014_),
    .Y(_04015_));
 sg13g2_xnor2_1 _09665_ (.Y(_04016_),
    .A(_04010_),
    .B(_04014_));
 sg13g2_nor2b_1 _09666_ (.A(_04009_),
    .B_N(_04016_),
    .Y(_04017_));
 sg13g2_a21o_1 _09667_ (.A2(_04008_),
    .A1(_04007_),
    .B1(_04017_),
    .X(_04018_));
 sg13g2_xnor2_1 _09668_ (.Y(_04019_),
    .A(_03989_),
    .B(_03990_));
 sg13g2_nand2b_1 _09669_ (.Y(_04020_),
    .B(_04018_),
    .A_N(_04019_));
 sg13g2_nor2_1 _09670_ (.A(_04012_),
    .B(_04015_),
    .Y(_04021_));
 sg13g2_xor2_1 _09671_ (.B(_04019_),
    .A(_04018_),
    .X(_04022_));
 sg13g2_o21ai_1 _09672_ (.B1(_04020_),
    .Y(_04023_),
    .A1(_04021_),
    .A2(_04022_));
 sg13g2_nand2_1 _09673_ (.Y(_04024_),
    .A(_04002_),
    .B(_04023_));
 sg13g2_nor2_1 _09674_ (.A(_04001_),
    .B(_04024_),
    .Y(_04025_));
 sg13g2_xor2_1 _09675_ (.B(_04023_),
    .A(_04002_),
    .X(_04026_));
 sg13g2_nor2_1 _09676_ (.A(_03876_),
    .B(_03900_),
    .Y(_04027_));
 sg13g2_and3_1 _09677_ (.X(_04028_),
    .A(net1590),
    .B(_03875_),
    .C(net1578));
 sg13g2_nand2_1 _09678_ (.Y(_04029_),
    .A(net1582),
    .B(_04028_));
 sg13g2_a22oi_1 _09679_ (.Y(_04030_),
    .B1(_04004_),
    .B2(_04005_),
    .A2(net1580),
    .A1(_03875_));
 sg13g2_or3_1 _09680_ (.A(_04006_),
    .B(_04029_),
    .C(_04030_),
    .X(_04031_));
 sg13g2_o21ai_1 _09681_ (.B1(_04029_),
    .Y(_04032_),
    .A1(_04006_),
    .A2(_04030_));
 sg13g2_nand2_1 _09682_ (.Y(_04033_),
    .A(_03870_),
    .B(net1576));
 sg13g2_nand2_1 _09683_ (.Y(_04034_),
    .A(net1588),
    .B(net1586));
 sg13g2_or2_1 _09684_ (.X(_04035_),
    .B(_04034_),
    .A(_04011_));
 sg13g2_xor2_1 _09685_ (.B(_04034_),
    .A(_04011_),
    .X(_04036_));
 sg13g2_nand2b_1 _09686_ (.Y(_04037_),
    .B(_04036_),
    .A_N(_04033_));
 sg13g2_xnor2_1 _09687_ (.Y(_04038_),
    .A(_04033_),
    .B(_04036_));
 sg13g2_nand3_1 _09688_ (.B(_04032_),
    .C(_04038_),
    .A(_04031_),
    .Y(_04039_));
 sg13g2_nand2_1 _09689_ (.Y(_04040_),
    .A(_04031_),
    .B(_04039_));
 sg13g2_xnor2_1 _09690_ (.Y(_04041_),
    .A(_04009_),
    .B(_04016_));
 sg13g2_nand2_1 _09691_ (.Y(_04042_),
    .A(_04040_),
    .B(_04041_));
 sg13g2_and2_1 _09692_ (.A(_04035_),
    .B(_04037_),
    .X(_04043_));
 sg13g2_nand2b_1 _09693_ (.Y(_04044_),
    .B(_03878_),
    .A_N(_04043_));
 sg13g2_xnor2_1 _09694_ (.Y(_04045_),
    .A(_03879_),
    .B(_04043_));
 sg13g2_xnor2_1 _09695_ (.Y(_04046_),
    .A(_04040_),
    .B(_04041_));
 sg13g2_o21ai_1 _09696_ (.B1(_04042_),
    .Y(_04047_),
    .A1(_04045_),
    .A2(_04046_));
 sg13g2_xor2_1 _09697_ (.B(_04022_),
    .A(_04021_),
    .X(_04048_));
 sg13g2_nand2_1 _09698_ (.Y(_04049_),
    .A(_04047_),
    .B(_04048_));
 sg13g2_xnor2_1 _09699_ (.Y(_04050_),
    .A(_04047_),
    .B(_04048_));
 sg13g2_o21ai_1 _09700_ (.B1(_04049_),
    .Y(_04051_),
    .A1(_04044_),
    .A2(_04050_));
 sg13g2_nand2_1 _09701_ (.Y(_04052_),
    .A(_04026_),
    .B(_04051_));
 sg13g2_nand2_1 _09702_ (.Y(_04053_),
    .A(_03870_),
    .B(net1575));
 sg13g2_and4_1 _09703_ (.A(net1593),
    .B(net1589),
    .C(net1585),
    .D(net1579),
    .X(_04054_));
 sg13g2_a22oi_1 _09704_ (.Y(_04055_),
    .B1(net1579),
    .B2(net1589),
    .A2(net1585),
    .A1(net1593));
 sg13g2_o21ai_1 _09705_ (.B1(_04053_),
    .Y(_04056_),
    .A1(_04054_),
    .A2(_04055_));
 sg13g2_or3_1 _09706_ (.A(_04053_),
    .B(_04054_),
    .C(_04055_),
    .X(_04057_));
 sg13g2_a22oi_1 _09707_ (.Y(_04058_),
    .B1(net1578),
    .B2(net1590),
    .A2(net1582),
    .A1(_03875_));
 sg13g2_a21oi_1 _09708_ (.A1(net1582),
    .A2(_04028_),
    .Y(_04059_),
    .B1(_04058_));
 sg13g2_and3_2 _09709_ (.X(_04060_),
    .A(_04056_),
    .B(_04057_),
    .C(_04059_));
 sg13g2_a21o_1 _09710_ (.A2(_04032_),
    .A1(_04031_),
    .B1(_04038_),
    .X(_04061_));
 sg13g2_and2_1 _09711_ (.A(_04039_),
    .B(_04061_),
    .X(_04062_));
 sg13g2_nand3_1 _09712_ (.B(_04060_),
    .C(_04061_),
    .A(_04039_),
    .Y(_04063_));
 sg13g2_a21o_1 _09713_ (.A2(_04061_),
    .A1(_04039_),
    .B1(_04060_),
    .X(_04064_));
 sg13g2_nor2b_1 _09714_ (.A(_04054_),
    .B_N(_04057_),
    .Y(_04065_));
 sg13g2_nor2b_1 _09715_ (.A(_03879_),
    .B_N(net1584),
    .Y(_04066_));
 sg13g2_nor2b_1 _09716_ (.A(_04065_),
    .B_N(_04066_),
    .Y(_04067_));
 sg13g2_xnor2_1 _09717_ (.Y(_04068_),
    .A(_04065_),
    .B(_04066_));
 sg13g2_xor2_1 _09718_ (.B(_04068_),
    .A(net1587),
    .X(_04069_));
 sg13g2_and3_1 _09719_ (.X(_04070_),
    .A(_04063_),
    .B(_04064_),
    .C(_04069_));
 sg13g2_a21oi_1 _09720_ (.A1(_04060_),
    .A2(_04062_),
    .Y(_04071_),
    .B1(_04070_));
 sg13g2_xnor2_1 _09721_ (.Y(_04072_),
    .A(_04045_),
    .B(_04046_));
 sg13g2_nor2_1 _09722_ (.A(_04071_),
    .B(_04072_),
    .Y(_04073_));
 sg13g2_a21o_1 _09723_ (.A2(_04068_),
    .A1(net1587),
    .B1(_04067_),
    .X(_04074_));
 sg13g2_xor2_1 _09724_ (.B(_04072_),
    .A(_04071_),
    .X(_04075_));
 sg13g2_a21oi_1 _09725_ (.A1(_04074_),
    .A2(_04075_),
    .Y(_04076_),
    .B1(_04073_));
 sg13g2_xor2_1 _09726_ (.B(_04050_),
    .A(_04044_),
    .X(_04077_));
 sg13g2_nor2b_1 _09727_ (.A(_04076_),
    .B_N(_04077_),
    .Y(_04078_));
 sg13g2_a21oi_1 _09728_ (.A1(_04056_),
    .A2(_04057_),
    .Y(_04079_),
    .B1(_04059_));
 sg13g2_nand2_1 _09729_ (.Y(_04080_),
    .A(_03870_),
    .B(net1585));
 sg13g2_nand2_1 _09730_ (.Y(_04081_),
    .A(net1592),
    .B(net1581));
 sg13g2_and4_1 _09731_ (.A(net1592),
    .B(net1588),
    .C(net1583),
    .D(net1579),
    .X(_04082_));
 sg13g2_nand4_1 _09732_ (.B(net1588),
    .C(net1581),
    .A(net1592),
    .Y(_04083_),
    .D(net1579));
 sg13g2_a22oi_1 _09733_ (.Y(_04084_),
    .B1(net1579),
    .B2(net1592),
    .A2(net1581),
    .A1(net1588));
 sg13g2_o21ai_1 _09734_ (.B1(_04080_),
    .Y(_04085_),
    .A1(_04082_),
    .A2(_04084_));
 sg13g2_or3_1 _09735_ (.A(_04080_),
    .B(_04082_),
    .C(_04084_),
    .X(_04086_));
 sg13g2_nand3_1 _09736_ (.B(_04085_),
    .C(_04086_),
    .A(_04027_),
    .Y(_04087_));
 sg13g2_nor3_1 _09737_ (.A(_04060_),
    .B(_04079_),
    .C(_04087_),
    .Y(_04088_));
 sg13g2_or3_1 _09738_ (.A(_04060_),
    .B(_04079_),
    .C(_04087_),
    .X(_04089_));
 sg13g2_o21ai_1 _09739_ (.B1(_04087_),
    .Y(_04090_),
    .A1(_04060_),
    .A2(_04079_));
 sg13g2_nand2_1 _09740_ (.Y(_04091_),
    .A(_03872_),
    .B(net1584));
 sg13g2_o21ai_1 _09741_ (.B1(_04083_),
    .Y(_04092_),
    .A1(_04080_),
    .A2(_04084_));
 sg13g2_nor2b_1 _09742_ (.A(_03879_),
    .B_N(net1576),
    .Y(_04093_));
 sg13g2_nand2_1 _09743_ (.Y(_04094_),
    .A(_04092_),
    .B(_04093_));
 sg13g2_xnor2_1 _09744_ (.Y(_04095_),
    .A(_04092_),
    .B(_04093_));
 sg13g2_xor2_1 _09745_ (.B(_04095_),
    .A(_04091_),
    .X(_04096_));
 sg13g2_and3_1 _09746_ (.X(_04097_),
    .A(_04089_),
    .B(_04090_),
    .C(_04096_));
 sg13g2_nor2_1 _09747_ (.A(_04088_),
    .B(_04097_),
    .Y(_04098_));
 sg13g2_a21oi_1 _09748_ (.A1(_04063_),
    .A2(_04064_),
    .Y(_04099_),
    .B1(_04069_));
 sg13g2_nor3_1 _09749_ (.A(_04070_),
    .B(_04098_),
    .C(_04099_),
    .Y(_04100_));
 sg13g2_or3_1 _09750_ (.A(_04070_),
    .B(_04098_),
    .C(_04099_),
    .X(_04101_));
 sg13g2_o21ai_1 _09751_ (.B1(_04094_),
    .Y(_04102_),
    .A1(_04091_),
    .A2(_04095_));
 sg13g2_o21ai_1 _09752_ (.B1(_04098_),
    .Y(_04103_),
    .A1(_04070_),
    .A2(_04099_));
 sg13g2_and3_1 _09753_ (.X(_04104_),
    .A(_04101_),
    .B(_04102_),
    .C(_04103_));
 sg13g2_nor2_1 _09754_ (.A(_04100_),
    .B(_04104_),
    .Y(_04105_));
 sg13g2_xnor2_1 _09755_ (.Y(_04106_),
    .A(_04074_),
    .B(_04075_));
 sg13g2_or2_1 _09756_ (.X(_04107_),
    .B(_04106_),
    .A(_04105_));
 sg13g2_nand2_1 _09757_ (.Y(_04108_),
    .A(net1587),
    .B(net1576));
 sg13g2_nand2_1 _09758_ (.Y(_04109_),
    .A(net1592),
    .B(net1577));
 sg13g2_nand2_1 _09759_ (.Y(_04110_),
    .A(net1588),
    .B(net1577));
 sg13g2_nand4_1 _09760_ (.B(net1588),
    .C(net1581),
    .A(net1592),
    .Y(_04111_),
    .D(net1577));
 sg13g2_nand2_1 _09761_ (.Y(_04112_),
    .A(_03870_),
    .B(net1579));
 sg13g2_a22oi_1 _09762_ (.Y(_04113_),
    .B1(net1577),
    .B2(net1588),
    .A2(net1581),
    .A1(net1592));
 sg13g2_xnor2_1 _09763_ (.Y(_04114_),
    .A(_04081_),
    .B(_04110_));
 sg13g2_o21ai_1 _09764_ (.B1(_04111_),
    .Y(_04115_),
    .A1(_04112_),
    .A2(_04113_));
 sg13g2_nor2b_1 _09765_ (.A(_03879_),
    .B_N(net1575),
    .Y(_04116_));
 sg13g2_nand2_1 _09766_ (.Y(_04117_),
    .A(_04115_),
    .B(_04116_));
 sg13g2_xnor2_1 _09767_ (.Y(_04118_),
    .A(_04115_),
    .B(_04116_));
 sg13g2_xor2_1 _09768_ (.B(_04118_),
    .A(_04108_),
    .X(_04119_));
 sg13g2_a21o_1 _09769_ (.A2(_04086_),
    .A1(_04085_),
    .B1(_04027_),
    .X(_04120_));
 sg13g2_and2_1 _09770_ (.A(_04087_),
    .B(_04120_),
    .X(_04121_));
 sg13g2_nand2_1 _09771_ (.Y(_04122_),
    .A(_04119_),
    .B(_04121_));
 sg13g2_a21oi_1 _09772_ (.A1(_04089_),
    .A2(_04090_),
    .Y(_04123_),
    .B1(_04096_));
 sg13g2_nor3_1 _09773_ (.A(_04097_),
    .B(_04122_),
    .C(_04123_),
    .Y(_04124_));
 sg13g2_or3_1 _09774_ (.A(_04097_),
    .B(_04122_),
    .C(_04123_),
    .X(_04125_));
 sg13g2_o21ai_1 _09775_ (.B1(_04117_),
    .Y(_04126_),
    .A1(_04108_),
    .A2(_04118_));
 sg13g2_inv_1 _09776_ (.Y(_04127_),
    .A(_04126_));
 sg13g2_o21ai_1 _09777_ (.B1(_04122_),
    .Y(_04128_),
    .A1(_04097_),
    .A2(_04123_));
 sg13g2_and2_1 _09778_ (.A(_04125_),
    .B(_04128_),
    .X(_04129_));
 sg13g2_a21oi_1 _09779_ (.A1(_04126_),
    .A2(_04128_),
    .Y(_04130_),
    .B1(_04124_));
 sg13g2_a21o_1 _09780_ (.A2(_04128_),
    .A1(_04126_),
    .B1(_04124_),
    .X(_04131_));
 sg13g2_a21oi_1 _09781_ (.A1(_04101_),
    .A2(_04103_),
    .Y(_04132_),
    .B1(_04102_));
 sg13g2_nor3_1 _09782_ (.A(_04104_),
    .B(_04130_),
    .C(_04132_),
    .Y(_04133_));
 sg13g2_o21ai_1 _09783_ (.B1(_04131_),
    .Y(_04134_),
    .A1(_04104_),
    .A2(_04132_));
 sg13g2_or3_1 _09784_ (.A(_04104_),
    .B(_04131_),
    .C(_04132_),
    .X(_04135_));
 sg13g2_nand2_1 _09785_ (.Y(_04136_),
    .A(net1587),
    .B(net1575));
 sg13g2_nand2_1 _09786_ (.Y(_04137_),
    .A(_03870_),
    .B(net1581));
 sg13g2_nor2_1 _09787_ (.A(_03871_),
    .B(_03900_),
    .Y(_04138_));
 sg13g2_nand2b_1 _09788_ (.Y(_04139_),
    .B(_04138_),
    .A_N(_04081_));
 sg13g2_nor2b_1 _09789_ (.A(_03879_),
    .B_N(net1585),
    .Y(_04140_));
 sg13g2_nand2b_1 _09790_ (.Y(_04141_),
    .B(_04140_),
    .A_N(_04139_));
 sg13g2_xnor2_1 _09791_ (.Y(_04142_),
    .A(_04139_),
    .B(_04140_));
 sg13g2_nand2b_1 _09792_ (.Y(_04143_),
    .B(_04142_),
    .A_N(_04136_));
 sg13g2_xnor2_1 _09793_ (.Y(_04144_),
    .A(_04136_),
    .B(_04142_));
 sg13g2_xnor2_1 _09794_ (.Y(_04145_),
    .A(_04112_),
    .B(_04114_));
 sg13g2_inv_1 _09795_ (.Y(_04146_),
    .A(_04145_));
 sg13g2_nand2_1 _09796_ (.Y(_04147_),
    .A(_04144_),
    .B(_04146_));
 sg13g2_xnor2_1 _09797_ (.Y(_04148_),
    .A(_04119_),
    .B(_04121_));
 sg13g2_nor2_1 _09798_ (.A(_04147_),
    .B(_04148_),
    .Y(_04149_));
 sg13g2_nand2_1 _09799_ (.Y(_04150_),
    .A(_04141_),
    .B(_04143_));
 sg13g2_xor2_1 _09800_ (.B(_04148_),
    .A(_04147_),
    .X(_04151_));
 sg13g2_a21oi_1 _09801_ (.A1(_04150_),
    .A2(_04151_),
    .Y(_04152_),
    .B1(_04149_));
 sg13g2_nand3_1 _09802_ (.B(_04127_),
    .C(_04128_),
    .A(_04125_),
    .Y(_04153_));
 sg13g2_a21oi_1 _09803_ (.A1(_04125_),
    .A2(_04128_),
    .Y(_04154_),
    .B1(_04127_));
 sg13g2_xnor2_1 _09804_ (.Y(_04155_),
    .A(_04127_),
    .B(_04129_));
 sg13g2_nand2b_1 _09805_ (.Y(_04156_),
    .B(_04155_),
    .A_N(_04152_));
 sg13g2_and2_1 _09806_ (.A(net1587),
    .B(net1579),
    .X(_04157_));
 sg13g2_nor2b_1 _09807_ (.A(_03879_),
    .B_N(net1579),
    .Y(_04158_));
 sg13g2_and2_1 _09808_ (.A(_04140_),
    .B(_04157_),
    .X(_04159_));
 sg13g2_xnor2_1 _09809_ (.Y(_04160_),
    .A(_04144_),
    .B(_04145_));
 sg13g2_nand2_1 _09810_ (.Y(_04161_),
    .A(_04159_),
    .B(_04160_));
 sg13g2_xnor2_1 _09811_ (.Y(_04162_),
    .A(_04150_),
    .B(_04151_));
 sg13g2_a21oi_1 _09812_ (.A1(net1587),
    .A2(net1585),
    .Y(_04163_),
    .B1(_04158_));
 sg13g2_or2_1 _09813_ (.X(_04164_),
    .B(_04163_),
    .A(_04159_));
 sg13g2_xnor2_1 _09814_ (.Y(_04165_),
    .A(_04109_),
    .B(_04137_));
 sg13g2_nor2_1 _09815_ (.A(_04164_),
    .B(_04165_),
    .Y(_04166_));
 sg13g2_a22oi_1 _09816_ (.Y(_04167_),
    .B1(_04138_),
    .B2(_04157_),
    .A2(net1581),
    .A1(_03878_));
 sg13g2_nor2_1 _09817_ (.A(net1577),
    .B(_04157_),
    .Y(_04168_));
 sg13g2_nor3_1 _09818_ (.A(_03873_),
    .B(_04167_),
    .C(_04168_),
    .Y(_04169_));
 sg13g2_nand4_1 _09819_ (.B(net1581),
    .C(net1577),
    .A(net1587),
    .Y(_04170_),
    .D(_04158_));
 sg13g2_a21oi_1 _09820_ (.A1(_03871_),
    .A2(_04157_),
    .Y(_04171_),
    .B1(_04170_));
 sg13g2_nand2_1 _09821_ (.Y(_04172_),
    .A(_04164_),
    .B(_04165_));
 sg13g2_o21ai_1 _09822_ (.B1(_04169_),
    .Y(_04173_),
    .A1(_04171_),
    .A2(_04172_));
 sg13g2_nor2b_1 _09823_ (.A(_04166_),
    .B_N(_04173_),
    .Y(_04174_));
 sg13g2_o21ai_1 _09824_ (.B1(_04161_),
    .Y(_04175_),
    .A1(_04162_),
    .A2(_04174_));
 sg13g2_nand2_1 _09825_ (.Y(_04176_),
    .A(_04166_),
    .B(_04171_));
 sg13g2_nor2_1 _09826_ (.A(_04159_),
    .B(_04160_),
    .Y(_04177_));
 sg13g2_o21ai_1 _09827_ (.B1(_04176_),
    .Y(_04178_),
    .A1(_04162_),
    .A2(_04177_));
 sg13g2_nand3b_1 _09828_ (.B(_04152_),
    .C(_04153_),
    .Y(_04179_),
    .A_N(_04154_));
 sg13g2_nand3_1 _09829_ (.B(_04178_),
    .C(_04179_),
    .A(_04175_),
    .Y(_04180_));
 sg13g2_a22oi_1 _09830_ (.Y(_04181_),
    .B1(_04156_),
    .B2(_04180_),
    .A2(_04135_),
    .A1(_04134_));
 sg13g2_nor2_1 _09831_ (.A(_04133_),
    .B(_04181_),
    .Y(_04182_));
 sg13g2_xor2_1 _09832_ (.B(_04106_),
    .A(_04105_),
    .X(_04183_));
 sg13g2_o21ai_1 _09833_ (.B1(_04183_),
    .Y(_04184_),
    .A1(_04133_),
    .A2(_04181_));
 sg13g2_xor2_1 _09834_ (.B(_04077_),
    .A(_04076_),
    .X(_04185_));
 sg13g2_a21oi_2 _09835_ (.B1(_04185_),
    .Y(_04186_),
    .A2(_04184_),
    .A1(_04107_));
 sg13g2_nor2_1 _09836_ (.A(_04078_),
    .B(_04186_),
    .Y(_04187_));
 sg13g2_xor2_1 _09837_ (.B(_04051_),
    .A(_04026_),
    .X(_04188_));
 sg13g2_o21ai_1 _09838_ (.B1(_04188_),
    .Y(_04189_),
    .A1(_04078_),
    .A2(_04186_));
 sg13g2_xnor2_1 _09839_ (.Y(_04190_),
    .A(_04001_),
    .B(_04024_));
 sg13g2_a21oi_1 _09840_ (.A1(_04052_),
    .A2(_04189_),
    .Y(_04191_),
    .B1(_04190_));
 sg13g2_xnor2_1 _09841_ (.Y(_04192_),
    .A(_03997_),
    .B(_03998_));
 sg13g2_o21ai_1 _09842_ (.B1(_04192_),
    .Y(_04193_),
    .A1(_04025_),
    .A2(_04191_));
 sg13g2_xor2_1 _09843_ (.B(_03974_),
    .A(_03967_),
    .X(_04194_));
 sg13g2_a21o_1 _09844_ (.A2(_04193_),
    .A1(_03999_),
    .B1(_04194_),
    .X(_04195_));
 sg13g2_nand2_1 _09845_ (.Y(_04196_),
    .A(_03975_),
    .B(_04195_));
 sg13g2_nand2_1 _09846_ (.Y(_04197_),
    .A(_03928_),
    .B(_03969_));
 sg13g2_and4_1 _09847_ (.A(_03928_),
    .B(_03936_),
    .C(_03969_),
    .D(_03973_),
    .X(_04198_));
 sg13g2_xnor2_1 _09848_ (.Y(_04199_),
    .A(_03936_),
    .B(_04197_));
 sg13g2_xnor2_1 _09849_ (.Y(_04200_),
    .A(_03973_),
    .B(_04199_));
 sg13g2_nand3_1 _09850_ (.B(_04195_),
    .C(_04198_),
    .A(_03975_),
    .Y(_04201_));
 sg13g2_and2_1 _09851_ (.A(_03858_),
    .B(_04201_),
    .X(_04202_));
 sg13g2_xor2_1 _09852_ (.B(net1464),
    .A(_03858_),
    .X(_04203_));
 sg13g2_a21oi_1 _09853_ (.A1(_03887_),
    .A2(_04203_),
    .Y(_04204_),
    .B1(_04202_));
 sg13g2_nor2_1 _09854_ (.A(_03855_),
    .B(_03883_),
    .Y(_04205_));
 sg13g2_xor2_1 _09855_ (.B(_03883_),
    .A(_03855_),
    .X(_04206_));
 sg13g2_o21ai_1 _09856_ (.B1(_03927_),
    .Y(_04207_),
    .A1(_04204_),
    .A2(_04205_));
 sg13g2_xor2_1 _09857_ (.B(_03888_),
    .A(_03862_),
    .X(_04208_));
 sg13g2_a21oi_1 _09858_ (.A1(_04207_),
    .A2(_04208_),
    .Y(_04209_),
    .B1(_03926_));
 sg13g2_a221oi_1 _09859_ (.B2(_04208_),
    .C1(_03926_),
    .B1(_04207_),
    .A1(_03856_),
    .Y(_04210_),
    .A2(_03890_));
 sg13g2_nor3_2 _09860_ (.A(_03924_),
    .B(_03925_),
    .C(_04210_),
    .Y(_04211_));
 sg13g2_nor2_1 _09861_ (.A(_03923_),
    .B(_04211_),
    .Y(_04212_));
 sg13g2_o21ai_1 _09862_ (.B1(_03921_),
    .Y(_04213_),
    .A1(_03923_),
    .A2(_04211_));
 sg13g2_a21oi_1 _09863_ (.A1(_03922_),
    .A2(_04213_),
    .Y(_04214_),
    .B1(_03920_));
 sg13g2_a21oi_2 _09864_ (.B1(_04214_),
    .Y(_04215_),
    .A2(_03889_),
    .A1(_03861_));
 sg13g2_o21ai_1 _09865_ (.B1(_03919_),
    .Y(_04216_),
    .A1(_03918_),
    .A2(_04215_));
 sg13g2_nand3_1 _09866_ (.B(_03922_),
    .C(_04213_),
    .A(_03920_),
    .Y(_04217_));
 sg13g2_nor2b_1 _09867_ (.A(_04214_),
    .B_N(_04217_),
    .Y(_04218_));
 sg13g2_o21ai_1 _09868_ (.B1(_03924_),
    .Y(_04219_),
    .A1(_03925_),
    .A2(_04210_));
 sg13g2_nor2b_1 _09869_ (.A(_04211_),
    .B_N(_04219_),
    .Y(_04220_));
 sg13g2_xnor2_1 _09870_ (.Y(_04221_),
    .A(_04204_),
    .B(_04206_));
 sg13g2_xor2_1 _09871_ (.B(_04203_),
    .A(_03887_),
    .X(_04222_));
 sg13g2_nand2_1 _09872_ (.Y(_04223_),
    .A(_04221_),
    .B(_04222_));
 sg13g2_xnor2_1 _09873_ (.Y(_04224_),
    .A(_04207_),
    .B(_04208_));
 sg13g2_nor2_1 _09874_ (.A(_04223_),
    .B(_04224_),
    .Y(_04225_));
 sg13g2_xor2_1 _09875_ (.B(_03890_),
    .A(_03856_),
    .X(_04226_));
 sg13g2_xnor2_1 _09876_ (.Y(_04227_),
    .A(_04209_),
    .B(_04226_));
 sg13g2_nand2_1 _09877_ (.Y(_04228_),
    .A(_04225_),
    .B(_04227_));
 sg13g2_and3_1 _09878_ (.X(_04229_),
    .A(_04220_),
    .B(_04225_),
    .C(_04227_));
 sg13g2_nand2_1 _09879_ (.Y(_04230_),
    .A(_03921_),
    .B(_03922_));
 sg13g2_xor2_1 _09880_ (.B(_04230_),
    .A(_04212_),
    .X(_04231_));
 sg13g2_and3_2 _09881_ (.X(_04232_),
    .A(_04218_),
    .B(_04229_),
    .C(_04231_));
 sg13g2_nor2b_1 _09882_ (.A(_03918_),
    .B_N(_03919_),
    .Y(_04233_));
 sg13g2_xnor2_1 _09883_ (.Y(_04234_),
    .A(_04215_),
    .B(_04233_));
 sg13g2_o21ai_1 _09884_ (.B1(_04216_),
    .Y(_04235_),
    .A1(_04232_),
    .A2(_04234_));
 sg13g2_nand2b_1 _09885_ (.Y(_04236_),
    .B(_03911_),
    .A_N(_03904_));
 sg13g2_o21ai_1 _09886_ (.B1(_04236_),
    .Y(_04237_),
    .A1(_03880_),
    .A2(_03915_));
 sg13g2_inv_1 _09887_ (.Y(_04238_),
    .A(_04237_));
 sg13g2_nand2b_1 _09888_ (.Y(_04239_),
    .B(_03882_),
    .A_N(_03865_));
 sg13g2_o21ai_1 _09889_ (.B1(_04239_),
    .Y(_04240_),
    .A1(_03893_),
    .A2(_03906_));
 sg13g2_a21oi_2 _09890_ (.B1(_04240_),
    .Y(_04241_),
    .A2(_04215_),
    .A1(_03918_));
 sg13g2_inv_1 _09891_ (.Y(_04242_),
    .A(_04241_));
 sg13g2_a21oi_1 _09892_ (.A1(_04229_),
    .A2(_04231_),
    .Y(_04243_),
    .B1(_04218_));
 sg13g2_nor2_1 _09893_ (.A(_04232_),
    .B(_04243_),
    .Y(_04244_));
 sg13g2_xnor2_1 _09894_ (.Y(_04245_),
    .A(_04220_),
    .B(_04228_));
 sg13g2_nand2b_1 _09895_ (.Y(_04246_),
    .B(_04221_),
    .A_N(_04222_));
 sg13g2_nor2_1 _09896_ (.A(_04224_),
    .B(_04246_),
    .Y(_04247_));
 sg13g2_nand4_1 _09897_ (.B(_04231_),
    .C(_04245_),
    .A(_04227_),
    .Y(_04248_),
    .D(_04247_));
 sg13g2_or4_1 _09898_ (.A(_04232_),
    .B(_04234_),
    .C(_04243_),
    .D(_04248_),
    .X(_04249_));
 sg13g2_xnor2_1 _09899_ (.Y(_04250_),
    .A(_04232_),
    .B(_04234_));
 sg13g2_and4_2 _09900_ (.A(_04235_),
    .B(_04238_),
    .C(_04241_),
    .D(_04249_),
    .X(_04251_));
 sg13g2_nand4_1 _09901_ (.B(_04135_),
    .C(_04156_),
    .A(_04134_),
    .Y(_04252_),
    .D(_04180_));
 sg13g2_nor2b_1 _09902_ (.A(_04181_),
    .B_N(_04252_),
    .Y(_04253_));
 sg13g2_xnor2_1 _09903_ (.Y(_04254_),
    .A(_04182_),
    .B(_04183_));
 sg13g2_mux2_1 _09904_ (.A0(_04253_),
    .A1(_04254_),
    .S(net1464),
    .X(_04255_));
 sg13g2_nand2_1 _09905_ (.Y(_04256_),
    .A(_04251_),
    .B(_04255_));
 sg13g2_a22oi_1 _09906_ (.Y(_00350_),
    .B1(net1484),
    .B2(_04256_),
    .A2(net1646),
    .A1(_00741_));
 sg13g2_nand3_1 _09907_ (.B(_04184_),
    .C(_04185_),
    .A(_04107_),
    .Y(_04257_));
 sg13g2_nor2b_1 _09908_ (.A(_04186_),
    .B_N(_04257_),
    .Y(_04258_));
 sg13g2_mux2_1 _09909_ (.A0(_04254_),
    .A1(_04258_),
    .S(net1464),
    .X(_04259_));
 sg13g2_nand2_1 _09910_ (.Y(_04260_),
    .A(_04251_),
    .B(_04259_));
 sg13g2_a22oi_1 _09911_ (.Y(_00351_),
    .B1(net1484),
    .B2(_04260_),
    .A2(net1646),
    .A1(_00740_));
 sg13g2_xnor2_1 _09912_ (.Y(_04261_),
    .A(_04187_),
    .B(_04188_));
 sg13g2_mux2_1 _09913_ (.A0(_04258_),
    .A1(_04261_),
    .S(net1464),
    .X(_04262_));
 sg13g2_nand2_1 _09914_ (.Y(_04263_),
    .A(_04251_),
    .B(_04262_));
 sg13g2_a22oi_1 _09915_ (.Y(_00352_),
    .B1(net1484),
    .B2(_04263_),
    .A2(net1646),
    .A1(_00743_));
 sg13g2_nand3_1 _09916_ (.B(_04189_),
    .C(_04190_),
    .A(_04052_),
    .Y(_04264_));
 sg13g2_nor2b_1 _09917_ (.A(_04191_),
    .B_N(_04264_),
    .Y(_04265_));
 sg13g2_mux2_1 _09918_ (.A0(_04261_),
    .A1(_04265_),
    .S(net1464),
    .X(_04266_));
 sg13g2_nand2_1 _09919_ (.Y(_04267_),
    .A(_04251_),
    .B(_04266_));
 sg13g2_a22oi_1 _09920_ (.Y(_00353_),
    .B1(net1484),
    .B2(_04267_),
    .A2(net1646),
    .A1(_00742_));
 sg13g2_or3_1 _09921_ (.A(_04025_),
    .B(_04191_),
    .C(_04192_),
    .X(_04268_));
 sg13g2_and2_1 _09922_ (.A(_04193_),
    .B(_04268_),
    .X(_04269_));
 sg13g2_mux2_1 _09923_ (.A0(_04265_),
    .A1(_04269_),
    .S(net1464),
    .X(_04270_));
 sg13g2_nand2_1 _09924_ (.Y(_04271_),
    .A(_04251_),
    .B(_04270_));
 sg13g2_a22oi_1 _09925_ (.Y(_00354_),
    .B1(net1484),
    .B2(_04271_),
    .A2(net1646),
    .A1(_00746_));
 sg13g2_nand3_1 _09926_ (.B(_04193_),
    .C(_04194_),
    .A(_03999_),
    .Y(_04272_));
 sg13g2_and2_1 _09927_ (.A(_04195_),
    .B(_04272_),
    .X(_04273_));
 sg13g2_mux2_1 _09928_ (.A0(_04269_),
    .A1(_04273_),
    .S(net1464),
    .X(_04274_));
 sg13g2_nand2_1 _09929_ (.Y(_04275_),
    .A(_04251_),
    .B(_04274_));
 sg13g2_a22oi_1 _09930_ (.Y(_00355_),
    .B1(net1484),
    .B2(_04275_),
    .A2(net1646),
    .A1(_00745_));
 sg13g2_xnor2_1 _09931_ (.Y(_04276_),
    .A(_04196_),
    .B(_04200_));
 sg13g2_o21ai_1 _09932_ (.B1(_04276_),
    .Y(_04277_),
    .A1(net1464),
    .A2(_04273_));
 sg13g2_nand2b_1 _09933_ (.Y(_04278_),
    .B(_04251_),
    .A_N(_04277_));
 sg13g2_a22oi_1 _09934_ (.Y(_00356_),
    .B1(net1484),
    .B2(_04278_),
    .A2(net1648),
    .A1(_00744_));
 sg13g2_nand3b_1 _09935_ (.B(_04215_),
    .C(_03918_),
    .Y(_04279_),
    .A_N(_04232_));
 sg13g2_nand3_1 _09936_ (.B(_04238_),
    .C(_04279_),
    .A(_04235_),
    .Y(_04280_));
 sg13g2_nor2b_1 _09937_ (.A(_04280_),
    .B_N(_04249_),
    .Y(_04281_));
 sg13g2_a21o_1 _09938_ (.A2(_04281_),
    .A1(_04222_),
    .B1(_04242_),
    .X(_04282_));
 sg13g2_a22oi_1 _09939_ (.Y(_00357_),
    .B1(net1485),
    .B2(_04282_),
    .A2(net1649),
    .A1(_00749_));
 sg13g2_xnor2_1 _09940_ (.Y(_04283_),
    .A(_04221_),
    .B(_04222_));
 sg13g2_a21o_1 _09941_ (.A2(_04283_),
    .A1(_04281_),
    .B1(_04242_),
    .X(_04284_));
 sg13g2_a22oi_1 _09942_ (.Y(_00358_),
    .B1(net1485),
    .B2(_04284_),
    .A2(net1649),
    .A1(_00748_));
 sg13g2_xnor2_1 _09943_ (.Y(_04285_),
    .A(_04223_),
    .B(_04224_));
 sg13g2_a21o_1 _09944_ (.A2(_04285_),
    .A1(_04281_),
    .B1(_04242_),
    .X(_04286_));
 sg13g2_a22oi_1 _09945_ (.Y(_00359_),
    .B1(net1485),
    .B2(_04286_),
    .A2(net1644),
    .A1(_00751_));
 sg13g2_xnor2_1 _09946_ (.Y(_04287_),
    .A(_04225_),
    .B(_04227_));
 sg13g2_a21o_1 _09947_ (.A2(_04287_),
    .A1(_04281_),
    .B1(_04242_),
    .X(_04288_));
 sg13g2_a22oi_1 _09948_ (.Y(_00360_),
    .B1(net1485),
    .B2(_04288_),
    .A2(net1644),
    .A1(_00750_));
 sg13g2_o21ai_1 _09949_ (.B1(_04241_),
    .Y(_04289_),
    .A1(_04245_),
    .A2(_04280_));
 sg13g2_a22oi_1 _09950_ (.Y(_00361_),
    .B1(net1485),
    .B2(_04289_),
    .A2(net1645),
    .A1(_00753_));
 sg13g2_xor2_1 _09951_ (.B(_04231_),
    .A(_04229_),
    .X(_04290_));
 sg13g2_o21ai_1 _09952_ (.B1(_04241_),
    .Y(_04291_),
    .A1(_04280_),
    .A2(_04290_));
 sg13g2_a22oi_1 _09953_ (.Y(_00362_),
    .B1(net1485),
    .B2(_04291_),
    .A2(net1649),
    .A1(_00752_));
 sg13g2_o21ai_1 _09954_ (.B1(_04241_),
    .Y(_04292_),
    .A1(_04244_),
    .A2(_04280_));
 sg13g2_a22oi_1 _09955_ (.Y(_00363_),
    .B1(net1485),
    .B2(_04292_),
    .A2(net1645),
    .A1(_00755_));
 sg13g2_o21ai_1 _09956_ (.B1(_04241_),
    .Y(_04293_),
    .A1(_04250_),
    .A2(_04280_));
 sg13g2_a22oi_1 _09957_ (.Y(_00364_),
    .B1(net1485),
    .B2(_04293_),
    .A2(net1645),
    .A1(_00754_));
 sg13g2_xor2_1 _09958_ (.B(_03905_),
    .A(_03881_),
    .X(_04294_));
 sg13g2_nand2_1 _09959_ (.Y(_04295_),
    .A(_04241_),
    .B(_04294_));
 sg13g2_a22oi_1 _09960_ (.Y(_00365_),
    .B1(net1484),
    .B2(_04295_),
    .A2(net1646),
    .A1(_00747_));
 sg13g2_mux2_2 _09961_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[0][8] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[1][8] ),
    .S(net1715),
    .X(_04296_));
 sg13g2_mux2_2 _09962_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[0][10] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[1][10] ),
    .S(net1710),
    .X(_04297_));
 sg13g2_mux2_2 _09963_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[0][14] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[1][14] ),
    .S(net1715),
    .X(_04298_));
 sg13g2_mux2_2 _09964_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[0][9] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[1][9] ),
    .S(net1710),
    .X(_04299_));
 sg13g2_mux2_2 _09965_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[0][11] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[1][11] ),
    .S(net1714),
    .X(_04300_));
 sg13g2_mux2_1 _09966_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[0][12] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[1][12] ),
    .S(net1714),
    .X(_04301_));
 sg13g2_mux2_2 _09967_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[0][13] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[1][13] ),
    .S(net1710),
    .X(_04302_));
 sg13g2_nand2b_1 _09968_ (.Y(_04303_),
    .B(net1713),
    .A_N(\u_tiny_nn_top.u_core.param_val_op_q[1][7] ));
 sg13g2_mux2_1 _09969_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[0][7] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[1][7] ),
    .S(net1713),
    .X(_04304_));
 sg13g2_o21ai_1 _09970_ (.B1(_04303_),
    .Y(_04305_),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[0][7] ),
    .A2(net1713));
 sg13g2_nor4_1 _09971_ (.A(_04297_),
    .B(_04299_),
    .C(_04301_),
    .D(_04304_),
    .Y(_04306_));
 sg13g2_nor4_1 _09972_ (.A(_04296_),
    .B(_04298_),
    .C(_04300_),
    .D(_04302_),
    .Y(_04307_));
 sg13g2_nand2_1 _09973_ (.Y(_04308_),
    .A(_04306_),
    .B(_04307_));
 sg13g2_mux2_2 _09974_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[0][5] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[1][5] ),
    .S(net1712),
    .X(_04309_));
 sg13g2_nand2_1 _09975_ (.Y(_04310_),
    .A(_00041_),
    .B(net1712));
 sg13g2_mux2_1 _09976_ (.A0(_00681_),
    .A1(_00682_),
    .S(net1712),
    .X(_04311_));
 sg13g2_o21ai_1 _09977_ (.B1(_04310_),
    .Y(_04312_),
    .A1(_00681_),
    .A2(net1712));
 sg13g2_mux2_2 _09978_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[0][0] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[1][0] ),
    .S(net1712),
    .X(_04313_));
 sg13g2_nor3_1 _09979_ (.A(net1574),
    .B(net1573),
    .C(net1571),
    .Y(_04314_));
 sg13g2_mux2_1 _09980_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[0][6] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[1][6] ),
    .S(net1713),
    .X(_04315_));
 sg13g2_mux2_2 _09981_ (.A0(_00040_),
    .A1(_00039_),
    .S(net1712),
    .X(_04316_));
 sg13g2_inv_2 _09982_ (.Y(_04317_),
    .A(_04316_));
 sg13g2_mux2_1 _09983_ (.A0(_00679_),
    .A1(_00680_),
    .S(net1712),
    .X(_04318_));
 sg13g2_mux2_1 _09984_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[0][3] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[1][3] ),
    .S(net1712),
    .X(_04319_));
 sg13g2_nor4_2 _09985_ (.A(net1570),
    .B(_04317_),
    .C(net1569),
    .Y(_04320_),
    .D(net1568));
 sg13g2_mux2_2 _09986_ (.A0(\u_tiny_nn_top.u_core.param_val_op_q[0][15] ),
    .A1(\u_tiny_nn_top.u_core.param_val_op_q[1][15] ),
    .S(net1716),
    .X(_04321_));
 sg13g2_nand3b_1 _09987_ (.B(_04320_),
    .C(_04314_),
    .Y(_04322_),
    .A_N(_04321_));
 sg13g2_or4_1 _09988_ (.A(net1573),
    .B(net1570),
    .C(_04317_),
    .D(net1569),
    .X(_04323_));
 sg13g2_nor4_2 _09989_ (.A(net1574),
    .B(net1571),
    .C(net1568),
    .Y(_04324_),
    .D(_04323_));
 sg13g2_nand2b_1 _09990_ (.Y(_04325_),
    .B(_04322_),
    .A_N(_04308_));
 sg13g2_mux2_2 _09991_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][8] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][8] ),
    .S(net1710),
    .X(_04326_));
 sg13g2_mux2_2 _09992_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][13] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][13] ),
    .S(net1711),
    .X(_04327_));
 sg13g2_mux2_2 _09993_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][10] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][10] ),
    .S(net1709),
    .X(_04328_));
 sg13g2_mux2_2 _09994_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][12] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][12] ),
    .S(net1697),
    .X(_04329_));
 sg13g2_mux2_2 _09995_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][7] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][7] ),
    .S(net1709),
    .X(_04330_));
 sg13g2_mux2_2 _09996_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][9] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][9] ),
    .S(net1697),
    .X(_04331_));
 sg13g2_mux2_2 _09997_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][14] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][14] ),
    .S(net1715),
    .X(_04332_));
 sg13g2_mux2_2 _09998_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][11] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][11] ),
    .S(net1709),
    .X(_04333_));
 sg13g2_nor4_1 _09999_ (.A(_04326_),
    .B(_04328_),
    .C(_04330_),
    .D(_04332_),
    .Y(_04334_));
 sg13g2_nor4_1 _10000_ (.A(_04327_),
    .B(_04329_),
    .C(_04331_),
    .D(_04333_),
    .Y(_04335_));
 sg13g2_and2_1 _10001_ (.A(_04334_),
    .B(_04335_),
    .X(_04336_));
 sg13g2_mux2_1 _10002_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][3] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][3] ),
    .S(net1695),
    .X(_04337_));
 sg13g2_mux2_1 _10003_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][2] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][2] ),
    .S(net1694),
    .X(_04338_));
 sg13g2_mux2_2 _10004_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][4] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][4] ),
    .S(net1706),
    .X(_04339_));
 sg13g2_nor3_1 _10005_ (.A(net1565),
    .B(net1563),
    .C(net1561),
    .Y(_04340_));
 sg13g2_mux2_1 _10006_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][1] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][1] ),
    .S(net1706),
    .X(_04341_));
 sg13g2_mux2_2 _10007_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][6] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][6] ),
    .S(net1706),
    .X(_04342_));
 sg13g2_mux2_2 _10008_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][0] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][0] ),
    .S(net1706),
    .X(_04343_));
 sg13g2_inv_1 _10009_ (.Y(_04344_),
    .A(_04343_));
 sg13g2_mux2_2 _10010_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][5] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][5] ),
    .S(net1694),
    .X(_04345_));
 sg13g2_inv_1 _10011_ (.Y(_04346_),
    .A(net1556));
 sg13g2_nor4_1 _10012_ (.A(net1560),
    .B(net1558),
    .C(net1557),
    .D(net1556),
    .Y(_04347_));
 sg13g2_nand2_2 _10013_ (.Y(_04348_),
    .A(_04340_),
    .B(_04347_));
 sg13g2_inv_1 _10014_ (.Y(_04349_),
    .A(_04348_));
 sg13g2_mux2_2 _10015_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[0][15] ),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][15] ),
    .S(net1711),
    .X(_04350_));
 sg13g2_o21ai_1 _10016_ (.B1(_04336_),
    .Y(_04351_),
    .A1(_04348_),
    .A2(_04350_));
 sg13g2_nand4_1 _10017_ (.B(_04297_),
    .C(_04300_),
    .A(_04296_),
    .Y(_04352_),
    .D(_04301_));
 sg13g2_nand4_1 _10018_ (.B(_04299_),
    .C(_04302_),
    .A(_04298_),
    .Y(_04353_),
    .D(_04304_));
 sg13g2_nor2_1 _10019_ (.A(_04352_),
    .B(_04353_),
    .Y(_04354_));
 sg13g2_nor2b_1 _10020_ (.A(_04324_),
    .B_N(_04354_),
    .Y(_04355_));
 sg13g2_nand4_1 _10021_ (.B(_04328_),
    .C(_04330_),
    .A(_04326_),
    .Y(_04356_),
    .D(_04332_));
 sg13g2_nand4_1 _10022_ (.B(_04329_),
    .C(_04331_),
    .A(_04327_),
    .Y(_04357_),
    .D(_04333_));
 sg13g2_nor2_1 _10023_ (.A(_04356_),
    .B(_04357_),
    .Y(_04358_));
 sg13g2_nand2_1 _10024_ (.Y(_04359_),
    .A(_04348_),
    .B(_04358_));
 sg13g2_nand3_1 _10025_ (.B(_04351_),
    .C(_04359_),
    .A(_04325_),
    .Y(_04360_));
 sg13g2_nor3_2 _10026_ (.A(net1650),
    .B(_04355_),
    .C(_04360_),
    .Y(_04361_));
 sg13g2_nor2_1 _10027_ (.A(_04298_),
    .B(_04332_),
    .Y(_04362_));
 sg13g2_nand2_1 _10028_ (.Y(_04363_),
    .A(_04298_),
    .B(_04332_));
 sg13g2_and2_1 _10029_ (.A(_04302_),
    .B(_04327_),
    .X(_04364_));
 sg13g2_or2_1 _10030_ (.X(_04365_),
    .B(_04327_),
    .A(_04302_));
 sg13g2_nand2b_1 _10031_ (.Y(_04366_),
    .B(_04365_),
    .A_N(_04364_));
 sg13g2_nor2_1 _10032_ (.A(_04301_),
    .B(_04329_),
    .Y(_04367_));
 sg13g2_nand2_1 _10033_ (.Y(_04368_),
    .A(_04301_),
    .B(_04329_));
 sg13g2_xnor2_1 _10034_ (.Y(_04369_),
    .A(_04300_),
    .B(_04333_));
 sg13g2_nor2_1 _10035_ (.A(_04297_),
    .B(_04328_),
    .Y(_04370_));
 sg13g2_and2_1 _10036_ (.A(_04299_),
    .B(_04331_),
    .X(_04371_));
 sg13g2_nand2_1 _10037_ (.Y(_04372_),
    .A(_04296_),
    .B(_04326_));
 sg13g2_and2_2 _10038_ (.A(net1570),
    .B(net1558),
    .X(_04373_));
 sg13g2_nand2_2 _10039_ (.Y(_04374_),
    .A(net1568),
    .B(net1558));
 sg13g2_nor2_1 _10040_ (.A(_04312_),
    .B(_04374_),
    .Y(_04375_));
 sg13g2_nand2_1 _10041_ (.Y(_04376_),
    .A(_04311_),
    .B(net1561));
 sg13g2_o21ai_1 _10042_ (.B1(_04376_),
    .Y(_04377_),
    .A1(_04312_),
    .A2(_04374_));
 sg13g2_nand2_1 _10043_ (.Y(_04378_),
    .A(net1574),
    .B(_04373_));
 sg13g2_xnor2_1 _10044_ (.Y(_04379_),
    .A(net1574),
    .B(_04373_));
 sg13g2_xnor2_1 _10045_ (.Y(_04380_),
    .A(_04346_),
    .B(_04377_));
 sg13g2_nor2b_1 _10046_ (.A(_04379_),
    .B_N(_04380_),
    .Y(_04381_));
 sg13g2_a21o_1 _10047_ (.A2(_04377_),
    .A1(net1556),
    .B1(_04381_),
    .X(_04382_));
 sg13g2_xnor2_1 _10048_ (.Y(_04383_),
    .A(net1570),
    .B(net1558));
 sg13g2_nor2b_1 _10049_ (.A(_04383_),
    .B_N(_04382_),
    .Y(_04384_));
 sg13g2_nor2_2 _10050_ (.A(_04373_),
    .B(_04384_),
    .Y(_04385_));
 sg13g2_inv_1 _10051_ (.Y(_04386_),
    .A(_04385_));
 sg13g2_a21oi_1 _10052_ (.A1(net1573),
    .A2(net1558),
    .Y(_04387_),
    .B1(net1568));
 sg13g2_a21oi_1 _10053_ (.A1(_04346_),
    .A2(_04375_),
    .Y(_04388_),
    .B1(_04387_));
 sg13g2_nand2_1 _10054_ (.Y(_04389_),
    .A(net1565),
    .B(_04388_));
 sg13g2_nand2_1 _10055_ (.Y(_04390_),
    .A(net1573),
    .B(_04374_));
 sg13g2_xor2_1 _10056_ (.B(_04390_),
    .A(net1561),
    .X(_04391_));
 sg13g2_nor2_1 _10057_ (.A(_04389_),
    .B(_04391_),
    .Y(_04392_));
 sg13g2_a22oi_1 _10058_ (.Y(_04393_),
    .B1(net1556),
    .B2(net1570),
    .A2(net1558),
    .A1(net1574));
 sg13g2_and2_2 _10059_ (.A(net1574),
    .B(net1556),
    .X(_04394_));
 sg13g2_nand2_1 _10060_ (.Y(_04395_),
    .A(_04373_),
    .B(_04394_));
 sg13g2_a21oi_1 _10061_ (.A1(_04373_),
    .A2(_04394_),
    .Y(_04396_),
    .B1(_04393_));
 sg13g2_xor2_1 _10062_ (.B(_04391_),
    .A(_04389_),
    .X(_04397_));
 sg13g2_a21oi_1 _10063_ (.A1(_04396_),
    .A2(_04397_),
    .Y(_04398_),
    .B1(_04392_));
 sg13g2_xnor2_1 _10064_ (.Y(_04399_),
    .A(_04379_),
    .B(_04380_));
 sg13g2_nand2b_1 _10065_ (.Y(_04400_),
    .B(_04399_),
    .A_N(_04398_));
 sg13g2_xnor2_1 _10066_ (.Y(_04401_),
    .A(_04398_),
    .B(_04399_));
 sg13g2_inv_1 _10067_ (.Y(_04402_),
    .A(_04401_));
 sg13g2_o21ai_1 _10068_ (.B1(_04400_),
    .Y(_04403_),
    .A1(_04395_),
    .A2(_04402_));
 sg13g2_nand2_1 _10069_ (.Y(_04404_),
    .A(_04378_),
    .B(_04383_));
 sg13g2_xor2_1 _10070_ (.B(_04404_),
    .A(_04382_),
    .X(_04405_));
 sg13g2_and2_1 _10071_ (.A(_04403_),
    .B(_04405_),
    .X(_04406_));
 sg13g2_xnor2_1 _10072_ (.Y(_04407_),
    .A(net1565),
    .B(_04388_));
 sg13g2_nand2_1 _10073_ (.Y(_04408_),
    .A(_04311_),
    .B(net1556));
 sg13g2_nand2_1 _10074_ (.Y(_04409_),
    .A(net1568),
    .B(net1556));
 sg13g2_nor2_1 _10075_ (.A(_04376_),
    .B(_04409_),
    .Y(_04410_));
 sg13g2_xor2_1 _10076_ (.B(_04409_),
    .A(_04376_),
    .X(_04411_));
 sg13g2_a21oi_1 _10077_ (.A1(net1569),
    .A2(_04411_),
    .Y(_04412_),
    .B1(_04410_));
 sg13g2_xor2_1 _10078_ (.B(_04408_),
    .A(_04374_),
    .X(_04413_));
 sg13g2_nand2b_1 _10079_ (.Y(_04414_),
    .B(_04413_),
    .A_N(_04412_));
 sg13g2_nor2b_2 _10080_ (.A(_04316_),
    .B_N(net1562),
    .Y(_04415_));
 sg13g2_nand2_1 _10081_ (.Y(_04416_),
    .A(_04317_),
    .B(net1563));
 sg13g2_xor2_1 _10082_ (.B(net1563),
    .A(_04316_),
    .X(_04417_));
 sg13g2_xor2_1 _10083_ (.B(_04413_),
    .A(_04412_),
    .X(_04418_));
 sg13g2_o21ai_1 _10084_ (.B1(_04414_),
    .Y(_04419_),
    .A1(_04417_),
    .A2(_04418_));
 sg13g2_nor2b_1 _10085_ (.A(_04407_),
    .B_N(_04419_),
    .Y(_04420_));
 sg13g2_nand2_1 _10086_ (.Y(_04421_),
    .A(_04315_),
    .B(net1563));
 sg13g2_nand2_2 _10087_ (.Y(_04422_),
    .A(_04317_),
    .B(_04339_));
 sg13g2_nand2_1 _10088_ (.Y(_04423_),
    .A(_04315_),
    .B(net1561));
 sg13g2_nor2_1 _10089_ (.A(_04421_),
    .B(_04422_),
    .Y(_04424_));
 sg13g2_xnor2_1 _10090_ (.Y(_04425_),
    .A(_04415_),
    .B(_04423_));
 sg13g2_xor2_1 _10091_ (.B(_04425_),
    .A(_04394_),
    .X(_04426_));
 sg13g2_xor2_1 _10092_ (.B(_04419_),
    .A(_04407_),
    .X(_04427_));
 sg13g2_inv_1 _10093_ (.Y(_04428_),
    .A(_04427_));
 sg13g2_a21oi_1 _10094_ (.A1(_04426_),
    .A2(_04428_),
    .Y(_04429_),
    .B1(_04420_));
 sg13g2_xnor2_1 _10095_ (.Y(_04430_),
    .A(_04396_),
    .B(_04397_));
 sg13g2_a21oi_1 _10096_ (.A1(_04394_),
    .A2(_04425_),
    .Y(_04431_),
    .B1(_04424_));
 sg13g2_xor2_1 _10097_ (.B(_04430_),
    .A(_04429_),
    .X(_04432_));
 sg13g2_nand2b_1 _10098_ (.Y(_04433_),
    .B(_04432_),
    .A_N(_04431_));
 sg13g2_o21ai_1 _10099_ (.B1(_04433_),
    .Y(_04434_),
    .A1(_04429_),
    .A2(_04430_));
 sg13g2_xnor2_1 _10100_ (.Y(_04435_),
    .A(_04395_),
    .B(_04401_));
 sg13g2_nand2_1 _10101_ (.Y(_04436_),
    .A(_04434_),
    .B(_04435_));
 sg13g2_and4_1 _10102_ (.A(net1573),
    .B(net1568),
    .C(net1565),
    .D(_04339_),
    .X(_04437_));
 sg13g2_nand2_1 _10103_ (.Y(_04438_),
    .A(net1569),
    .B(_04342_));
 sg13g2_a22oi_1 _10104_ (.Y(_04439_),
    .B1(net1561),
    .B2(net1568),
    .A2(net1565),
    .A1(net1573));
 sg13g2_or3_1 _10105_ (.A(_04437_),
    .B(_04438_),
    .C(_04439_),
    .X(_04440_));
 sg13g2_nand2b_1 _10106_ (.Y(_04441_),
    .B(_04440_),
    .A_N(_04437_));
 sg13g2_xor2_1 _10107_ (.B(_04411_),
    .A(net1569),
    .X(_04442_));
 sg13g2_nand2_1 _10108_ (.Y(_04443_),
    .A(_04317_),
    .B(net1559));
 sg13g2_nor2b_1 _10109_ (.A(_04316_),
    .B_N(net1558),
    .Y(_04444_));
 sg13g2_nand2_1 _10110_ (.Y(_04445_),
    .A(net1560),
    .B(_04444_));
 sg13g2_xnor2_1 _10111_ (.Y(_04446_),
    .A(net1560),
    .B(_04444_));
 sg13g2_xor2_1 _10112_ (.B(_04442_),
    .A(_04441_),
    .X(_04447_));
 sg13g2_nor2b_1 _10113_ (.A(_04446_),
    .B_N(_04447_),
    .Y(_04448_));
 sg13g2_a21o_1 _10114_ (.A2(_04442_),
    .A1(_04441_),
    .B1(_04448_),
    .X(_04449_));
 sg13g2_xnor2_1 _10115_ (.Y(_04450_),
    .A(_04417_),
    .B(_04418_));
 sg13g2_nand2b_1 _10116_ (.Y(_04451_),
    .B(_04449_),
    .A_N(_04450_));
 sg13g2_nand2_1 _10117_ (.Y(_04452_),
    .A(_04309_),
    .B(net1561));
 sg13g2_nand2_1 _10118_ (.Y(_04453_),
    .A(net1570),
    .B(net1564));
 sg13g2_xor2_1 _10119_ (.B(_04453_),
    .A(_04445_),
    .X(_04454_));
 sg13g2_nand2b_1 _10120_ (.Y(_04455_),
    .B(_04454_),
    .A_N(_04452_));
 sg13g2_xnor2_1 _10121_ (.Y(_04456_),
    .A(_04452_),
    .B(_04454_));
 sg13g2_inv_1 _10122_ (.Y(_04457_),
    .A(_04456_));
 sg13g2_xor2_1 _10123_ (.B(_04450_),
    .A(_04449_),
    .X(_04458_));
 sg13g2_o21ai_1 _10124_ (.B1(_04451_),
    .Y(_04459_),
    .A1(_04457_),
    .A2(_04458_));
 sg13g2_xor2_1 _10125_ (.B(_04427_),
    .A(_04426_),
    .X(_04460_));
 sg13g2_nand2b_1 _10126_ (.Y(_04461_),
    .B(_04459_),
    .A_N(_04460_));
 sg13g2_o21ai_1 _10127_ (.B1(_04455_),
    .Y(_04462_),
    .A1(_04445_),
    .A2(_04453_));
 sg13g2_inv_1 _10128_ (.Y(_04463_),
    .A(_04462_));
 sg13g2_xor2_1 _10129_ (.B(_04460_),
    .A(_04459_),
    .X(_04464_));
 sg13g2_o21ai_1 _10130_ (.B1(_04461_),
    .Y(_04465_),
    .A1(_04463_),
    .A2(_04464_));
 sg13g2_xnor2_1 _10131_ (.Y(_04466_),
    .A(_04431_),
    .B(_04432_));
 sg13g2_and2_1 _10132_ (.A(_04465_),
    .B(_04466_),
    .X(_04467_));
 sg13g2_and4_1 _10133_ (.A(net1573),
    .B(net1567),
    .C(net1564),
    .D(net1562),
    .X(_04468_));
 sg13g2_nand4_1 _10134_ (.B(net1567),
    .C(net1564),
    .A(net1572),
    .Y(_04469_),
    .D(net1562));
 sg13g2_nand2_1 _10135_ (.Y(_04470_),
    .A(_04318_),
    .B(_04345_));
 sg13g2_a22oi_1 _10136_ (.Y(_04471_),
    .B1(net1562),
    .B2(net1572),
    .A2(net1564),
    .A1(net1567));
 sg13g2_or3_1 _10137_ (.A(_04468_),
    .B(_04470_),
    .C(_04471_),
    .X(_04472_));
 sg13g2_o21ai_1 _10138_ (.B1(_04469_),
    .Y(_04473_),
    .A1(_04470_),
    .A2(_04471_));
 sg13g2_o21ai_1 _10139_ (.B1(_04438_),
    .Y(_04474_),
    .A1(_04437_),
    .A2(_04439_));
 sg13g2_and3_1 _10140_ (.X(_04475_),
    .A(_04440_),
    .B(_04473_),
    .C(_04474_));
 sg13g2_a21oi_1 _10141_ (.A1(_04440_),
    .A2(_04474_),
    .Y(_04476_),
    .B1(_04473_));
 sg13g2_nor2b_1 _10142_ (.A(_04316_),
    .B_N(net1556),
    .Y(_04477_));
 sg13g2_nand2_1 _10143_ (.Y(_04478_),
    .A(_04313_),
    .B(_04477_));
 sg13g2_xnor2_1 _10144_ (.Y(_04479_),
    .A(_04313_),
    .B(_04477_));
 sg13g2_xnor2_1 _10145_ (.Y(_04480_),
    .A(_04344_),
    .B(_04479_));
 sg13g2_or3_1 _10146_ (.A(_04475_),
    .B(_04476_),
    .C(_04480_),
    .X(_04481_));
 sg13g2_nand2b_1 _10147_ (.Y(_04482_),
    .B(_04481_),
    .A_N(_04475_));
 sg13g2_xnor2_1 _10148_ (.Y(_04483_),
    .A(_04446_),
    .B(_04447_));
 sg13g2_xnor2_1 _10149_ (.Y(_04484_),
    .A(_04482_),
    .B(_04483_));
 sg13g2_nand2_1 _10150_ (.Y(_04485_),
    .A(_04309_),
    .B(net1565));
 sg13g2_o21ai_1 _10151_ (.B1(_04478_),
    .Y(_04486_),
    .A1(_04344_),
    .A2(_04479_));
 sg13g2_nand2b_1 _10152_ (.Y(_04487_),
    .B(_04486_),
    .A_N(_04421_));
 sg13g2_xor2_1 _10153_ (.B(_04486_),
    .A(_04421_),
    .X(_04488_));
 sg13g2_xor2_1 _10154_ (.B(_04488_),
    .A(_04485_),
    .X(_04489_));
 sg13g2_nor2b_1 _10155_ (.A(_04484_),
    .B_N(_04489_),
    .Y(_04490_));
 sg13g2_a21o_1 _10156_ (.A2(_04483_),
    .A1(_04482_),
    .B1(_04490_),
    .X(_04491_));
 sg13g2_xnor2_1 _10157_ (.Y(_04492_),
    .A(_04457_),
    .B(_04458_));
 sg13g2_nand2b_1 _10158_ (.Y(_04493_),
    .B(_04491_),
    .A_N(_04492_));
 sg13g2_o21ai_1 _10159_ (.B1(_04487_),
    .Y(_04494_),
    .A1(_04485_),
    .A2(_04488_));
 sg13g2_inv_1 _10160_ (.Y(_04495_),
    .A(_04494_));
 sg13g2_xor2_1 _10161_ (.B(_04492_),
    .A(_04491_),
    .X(_04496_));
 sg13g2_o21ai_1 _10162_ (.B1(_04493_),
    .Y(_04497_),
    .A1(_04495_),
    .A2(_04496_));
 sg13g2_xnor2_1 _10163_ (.Y(_04498_),
    .A(_04463_),
    .B(_04464_));
 sg13g2_nor2b_1 _10164_ (.A(_04498_),
    .B_N(_04497_),
    .Y(_04499_));
 sg13g2_and4_1 _10165_ (.A(net1572),
    .B(net1566),
    .C(net1562),
    .D(net1559),
    .X(_04500_));
 sg13g2_nand4_1 _10166_ (.B(net1566),
    .C(net1562),
    .A(net1572),
    .Y(_04501_),
    .D(net1559));
 sg13g2_nand2_1 _10167_ (.Y(_04502_),
    .A(_04318_),
    .B(net1561));
 sg13g2_a22oi_1 _10168_ (.Y(_04503_),
    .B1(net1559),
    .B2(net1572),
    .A2(net1562),
    .A1(net1566));
 sg13g2_or3_1 _10169_ (.A(_04500_),
    .B(_04502_),
    .C(_04503_),
    .X(_04504_));
 sg13g2_o21ai_1 _10170_ (.B1(_04501_),
    .Y(_04505_),
    .A1(_04502_),
    .A2(_04503_));
 sg13g2_o21ai_1 _10171_ (.B1(_04470_),
    .Y(_04506_),
    .A1(_04468_),
    .A2(_04471_));
 sg13g2_and3_1 _10172_ (.X(_04507_),
    .A(_04472_),
    .B(_04505_),
    .C(_04506_));
 sg13g2_nand3_1 _10173_ (.B(_04505_),
    .C(_04506_),
    .A(_04472_),
    .Y(_04508_));
 sg13g2_nand2_1 _10174_ (.Y(_04509_),
    .A(net1571),
    .B(net1558));
 sg13g2_nand2_1 _10175_ (.Y(_04510_),
    .A(_04313_),
    .B(net1561));
 sg13g2_or2_1 _10176_ (.X(_04511_),
    .B(_04509_),
    .A(_04422_));
 sg13g2_xnor2_1 _10177_ (.Y(_04512_),
    .A(_04422_),
    .B(_04509_));
 sg13g2_a21oi_1 _10178_ (.A1(_04472_),
    .A2(_04506_),
    .Y(_04513_),
    .B1(_04505_));
 sg13g2_or3_1 _10179_ (.A(_04507_),
    .B(_04512_),
    .C(_04513_),
    .X(_04514_));
 sg13g2_o21ai_1 _10180_ (.B1(_04508_),
    .Y(_04515_),
    .A1(_04512_),
    .A2(_04513_));
 sg13g2_o21ai_1 _10181_ (.B1(_04480_),
    .Y(_04516_),
    .A1(_04475_),
    .A2(_04476_));
 sg13g2_nand3_1 _10182_ (.B(_04515_),
    .C(_04516_),
    .A(_04481_),
    .Y(_04517_));
 sg13g2_a21o_1 _10183_ (.A2(_04516_),
    .A1(_04481_),
    .B1(_04515_),
    .X(_04518_));
 sg13g2_nand2_1 _10184_ (.Y(_04519_),
    .A(_04309_),
    .B(net1563));
 sg13g2_inv_1 _10185_ (.Y(_04520_),
    .A(_04519_));
 sg13g2_nand2_1 _10186_ (.Y(_04521_),
    .A(net1570),
    .B(net1560));
 sg13g2_nor2_1 _10187_ (.A(_04511_),
    .B(_04521_),
    .Y(_04522_));
 sg13g2_xor2_1 _10188_ (.B(_04521_),
    .A(_04511_),
    .X(_04523_));
 sg13g2_xnor2_1 _10189_ (.Y(_04524_),
    .A(_04519_),
    .B(_04523_));
 sg13g2_nand3_1 _10190_ (.B(_04518_),
    .C(_04524_),
    .A(_04517_),
    .Y(_04525_));
 sg13g2_nand2_1 _10191_ (.Y(_04526_),
    .A(_04517_),
    .B(_04525_));
 sg13g2_xnor2_1 _10192_ (.Y(_04527_),
    .A(_04484_),
    .B(_04489_));
 sg13g2_nand2_1 _10193_ (.Y(_04528_),
    .A(_04526_),
    .B(_04527_));
 sg13g2_a21oi_2 _10194_ (.B1(_04522_),
    .Y(_04529_),
    .A2(_04523_),
    .A1(_04520_));
 sg13g2_xnor2_1 _10195_ (.Y(_04530_),
    .A(_04526_),
    .B(_04527_));
 sg13g2_o21ai_1 _10196_ (.B1(_04528_),
    .Y(_04531_),
    .A1(_04529_),
    .A2(_04530_));
 sg13g2_xnor2_1 _10197_ (.Y(_04532_),
    .A(_04495_),
    .B(_04496_));
 sg13g2_nand2b_1 _10198_ (.Y(_04533_),
    .B(_04531_),
    .A_N(_04532_));
 sg13g2_and4_1 _10199_ (.A(net1572),
    .B(net1566),
    .C(net1559),
    .D(net1557),
    .X(_04534_));
 sg13g2_nand4_1 _10200_ (.B(net1566),
    .C(net1559),
    .A(net1572),
    .Y(_04535_),
    .D(net1557));
 sg13g2_nand2_1 _10201_ (.Y(_04536_),
    .A(_04318_),
    .B(net1564));
 sg13g2_a22oi_1 _10202_ (.Y(_04537_),
    .B1(net1557),
    .B2(net1572),
    .A2(net1559),
    .A1(net1566));
 sg13g2_or3_1 _10203_ (.A(_04534_),
    .B(_04536_),
    .C(_04537_),
    .X(_04538_));
 sg13g2_o21ai_1 _10204_ (.B1(_04535_),
    .Y(_04539_),
    .A1(_04536_),
    .A2(_04537_));
 sg13g2_o21ai_1 _10205_ (.B1(_04502_),
    .Y(_04540_),
    .A1(_04500_),
    .A2(_04503_));
 sg13g2_and3_1 _10206_ (.X(_04541_),
    .A(_04504_),
    .B(_04539_),
    .C(_04540_));
 sg13g2_nand3_1 _10207_ (.B(_04539_),
    .C(_04540_),
    .A(_04504_),
    .Y(_04542_));
 sg13g2_a22oi_1 _10208_ (.Y(_04543_),
    .B1(_04345_),
    .B2(net1571),
    .A2(net1564),
    .A1(_04317_));
 sg13g2_nand2_1 _10209_ (.Y(_04544_),
    .A(net1571),
    .B(net1564));
 sg13g2_nand3_1 _10210_ (.B(net1564),
    .C(_04477_),
    .A(net1571),
    .Y(_04545_));
 sg13g2_nor2b_1 _10211_ (.A(_04543_),
    .B_N(_04545_),
    .Y(_04546_));
 sg13g2_nand2b_1 _10212_ (.Y(_04547_),
    .B(_04545_),
    .A_N(_04543_));
 sg13g2_a21oi_1 _10213_ (.A1(_04504_),
    .A2(_04540_),
    .Y(_04548_),
    .B1(_04539_));
 sg13g2_a21o_1 _10214_ (.A2(_04540_),
    .A1(_04504_),
    .B1(_04539_),
    .X(_04549_));
 sg13g2_nand3_1 _10215_ (.B(_04546_),
    .C(_04549_),
    .A(_04542_),
    .Y(_04550_));
 sg13g2_a21oi_1 _10216_ (.A1(_04546_),
    .A2(_04549_),
    .Y(_04551_),
    .B1(_04541_));
 sg13g2_o21ai_1 _10217_ (.B1(_04542_),
    .Y(_04552_),
    .A1(_04547_),
    .A2(_04548_));
 sg13g2_o21ai_1 _10218_ (.B1(_04512_),
    .Y(_04553_),
    .A1(_04507_),
    .A2(_04513_));
 sg13g2_nand3_1 _10219_ (.B(_04552_),
    .C(_04553_),
    .A(_04514_),
    .Y(_04554_));
 sg13g2_nand2_1 _10220_ (.Y(_04555_),
    .A(net1574),
    .B(net1559));
 sg13g2_inv_1 _10221_ (.Y(_04556_),
    .A(_04555_));
 sg13g2_nand2_1 _10222_ (.Y(_04557_),
    .A(net1570),
    .B(net1557));
 sg13g2_nor2_1 _10223_ (.A(_04545_),
    .B(_04557_),
    .Y(_04558_));
 sg13g2_xor2_1 _10224_ (.B(_04557_),
    .A(_04545_),
    .X(_04559_));
 sg13g2_xnor2_1 _10225_ (.Y(_04560_),
    .A(_04556_),
    .B(_04559_));
 sg13g2_a21oi_1 _10226_ (.A1(_04514_),
    .A2(_04553_),
    .Y(_04561_),
    .B1(_04552_));
 sg13g2_a21o_1 _10227_ (.A2(_04553_),
    .A1(_04514_),
    .B1(_04551_),
    .X(_04562_));
 sg13g2_nand4_1 _10228_ (.B(_04542_),
    .C(_04550_),
    .A(_04514_),
    .Y(_04563_),
    .D(_04553_));
 sg13g2_a21oi_1 _10229_ (.A1(_04562_),
    .A2(_04563_),
    .Y(_04564_),
    .B1(_04560_));
 sg13g2_o21ai_1 _10230_ (.B1(_04554_),
    .Y(_04565_),
    .A1(_04560_),
    .A2(_04561_));
 sg13g2_a21o_1 _10231_ (.A2(_04518_),
    .A1(_04517_),
    .B1(_04524_),
    .X(_04566_));
 sg13g2_and3_1 _10232_ (.X(_04567_),
    .A(_04525_),
    .B(_04565_),
    .C(_04566_));
 sg13g2_a21oi_1 _10233_ (.A1(_04556_),
    .A2(_04559_),
    .Y(_04568_),
    .B1(_04558_));
 sg13g2_a21oi_1 _10234_ (.A1(_04525_),
    .A2(_04566_),
    .Y(_04569_),
    .B1(_04565_));
 sg13g2_or3_1 _10235_ (.A(_04567_),
    .B(_04568_),
    .C(_04569_),
    .X(_04570_));
 sg13g2_nand2b_1 _10236_ (.Y(_04571_),
    .B(_04570_),
    .A_N(_04567_));
 sg13g2_xor2_1 _10237_ (.B(_04530_),
    .A(_04529_),
    .X(_04572_));
 sg13g2_and2_1 _10238_ (.A(_04571_),
    .B(_04572_),
    .X(_04573_));
 sg13g2_and3_1 _10239_ (.X(_04574_),
    .A(_04560_),
    .B(_04562_),
    .C(_04563_));
 sg13g2_nand4_1 _10240_ (.B(net1566),
    .C(net1563),
    .A(net1569),
    .Y(_04575_),
    .D(net1557));
 sg13g2_inv_1 _10241_ (.Y(_04576_),
    .A(_04575_));
 sg13g2_o21ai_1 _10242_ (.B1(_04536_),
    .Y(_04577_),
    .A1(_04534_),
    .A2(_04537_));
 sg13g2_and3_1 _10243_ (.X(_04578_),
    .A(_04538_),
    .B(_04576_),
    .C(_04577_));
 sg13g2_nand3_1 _10244_ (.B(_04576_),
    .C(_04577_),
    .A(_04538_),
    .Y(_04579_));
 sg13g2_a21oi_1 _10245_ (.A1(_04538_),
    .A2(_04577_),
    .Y(_04580_),
    .B1(_04576_));
 sg13g2_nor2_1 _10246_ (.A(_04578_),
    .B(_04580_),
    .Y(_04581_));
 sg13g2_nand2_1 _10247_ (.Y(_04582_),
    .A(net1571),
    .B(net1563));
 sg13g2_or2_2 _10248_ (.X(_04583_),
    .B(_04582_),
    .A(_04422_));
 sg13g2_xnor2_1 _10249_ (.Y(_04584_),
    .A(_04415_),
    .B(_04510_));
 sg13g2_inv_1 _10250_ (.Y(_04585_),
    .A(_04584_));
 sg13g2_o21ai_1 _10251_ (.B1(_04579_),
    .Y(_04586_),
    .A1(_04580_),
    .A2(_04585_));
 sg13g2_o21ai_1 _10252_ (.B1(_04547_),
    .Y(_04587_),
    .A1(_04541_),
    .A2(_04548_));
 sg13g2_and3_1 _10253_ (.X(_04588_),
    .A(_04550_),
    .B(_04586_),
    .C(_04587_));
 sg13g2_nand2_2 _10254_ (.Y(_04589_),
    .A(net1574),
    .B(net1557));
 sg13g2_nor2_1 _10255_ (.A(_04583_),
    .B(_04589_),
    .Y(_04590_));
 sg13g2_xor2_1 _10256_ (.B(_04589_),
    .A(_04583_),
    .X(_04591_));
 sg13g2_xnor2_1 _10257_ (.Y(_04592_),
    .A(_04583_),
    .B(_04589_));
 sg13g2_a21oi_1 _10258_ (.A1(_04550_),
    .A2(_04587_),
    .Y(_04593_),
    .B1(_04586_));
 sg13g2_a21o_1 _10259_ (.A2(_04587_),
    .A1(_04550_),
    .B1(_04586_),
    .X(_04594_));
 sg13g2_nor3_1 _10260_ (.A(_04588_),
    .B(_04592_),
    .C(_04593_),
    .Y(_04595_));
 sg13g2_a21oi_1 _10261_ (.A1(_04591_),
    .A2(_04594_),
    .Y(_04596_),
    .B1(_04588_));
 sg13g2_nor3_1 _10262_ (.A(_04564_),
    .B(_04574_),
    .C(_04596_),
    .Y(_04597_));
 sg13g2_or3_1 _10263_ (.A(_04564_),
    .B(_04574_),
    .C(_04596_),
    .X(_04598_));
 sg13g2_o21ai_1 _10264_ (.B1(_04596_),
    .Y(_04599_),
    .A1(_04564_),
    .A2(_04574_));
 sg13g2_nand3_1 _10265_ (.B(_04598_),
    .C(_04599_),
    .A(_04590_),
    .Y(_04600_));
 sg13g2_a21o_1 _10266_ (.A2(_04599_),
    .A1(_04590_),
    .B1(_04597_),
    .X(_04601_));
 sg13g2_o21ai_1 _10267_ (.B1(_04568_),
    .Y(_04602_),
    .A1(_04567_),
    .A2(_04569_));
 sg13g2_and3_1 _10268_ (.X(_04603_),
    .A(_04570_),
    .B(_04601_),
    .C(_04602_));
 sg13g2_nand3_1 _10269_ (.B(_04601_),
    .C(_04602_),
    .A(_04570_),
    .Y(_04604_));
 sg13g2_a21o_1 _10270_ (.A2(_04599_),
    .A1(_04598_),
    .B1(_04590_),
    .X(_04605_));
 sg13g2_o21ai_1 _10271_ (.B1(_04592_),
    .Y(_04606_),
    .A1(_04588_),
    .A2(_04593_));
 sg13g2_nand2_1 _10272_ (.Y(_04607_),
    .A(net1569),
    .B(net1560));
 sg13g2_nand2_1 _10273_ (.Y(_04608_),
    .A(net1571),
    .B(net1557));
 sg13g2_nor2_1 _10274_ (.A(_04607_),
    .B(_04608_),
    .Y(_04609_));
 sg13g2_nand2_1 _10275_ (.Y(_04610_),
    .A(_04415_),
    .B(_04609_));
 sg13g2_o21ai_1 _10276_ (.B1(_04582_),
    .Y(_04611_),
    .A1(_04316_),
    .A2(_04344_));
 sg13g2_o21ai_1 _10277_ (.B1(_04607_),
    .Y(_04612_),
    .A1(_04416_),
    .A2(_04608_));
 sg13g2_a22oi_1 _10278_ (.Y(_04613_),
    .B1(_04611_),
    .B2(_04612_),
    .A2(_04609_),
    .A1(_04417_));
 sg13g2_nor2_1 _10279_ (.A(_04443_),
    .B(_04544_),
    .Y(_04614_));
 sg13g2_xor2_1 _10280_ (.B(_04544_),
    .A(_04443_),
    .X(_04615_));
 sg13g2_a22oi_1 _10281_ (.Y(_04616_),
    .B1(_04343_),
    .B2(net1566),
    .A2(net1562),
    .A1(net1569));
 sg13g2_nor2_1 _10282_ (.A(_04576_),
    .B(_04616_),
    .Y(_04617_));
 sg13g2_nand2_1 _10283_ (.Y(_04618_),
    .A(_04615_),
    .B(_04617_));
 sg13g2_xnor2_1 _10284_ (.Y(_04619_),
    .A(_04615_),
    .B(_04617_));
 sg13g2_o21ai_1 _10285_ (.B1(_04610_),
    .Y(_04620_),
    .A1(_04613_),
    .A2(_04619_));
 sg13g2_xnor2_1 _10286_ (.Y(_04621_),
    .A(_04581_),
    .B(_04584_));
 sg13g2_or2_1 _10287_ (.X(_04622_),
    .B(_04621_),
    .A(_04618_));
 sg13g2_nor2_1 _10288_ (.A(_04614_),
    .B(_04620_),
    .Y(_04623_));
 sg13g2_a22oi_1 _10289_ (.Y(_04624_),
    .B1(_04620_),
    .B2(_04614_),
    .A2(_04617_),
    .A1(_04615_));
 sg13g2_a221oi_1 _10290_ (.B2(_04621_),
    .C1(_04595_),
    .B1(_04624_),
    .A1(_04622_),
    .Y(_04625_),
    .A2(_04623_));
 sg13g2_nand4_1 _10291_ (.B(_04605_),
    .C(_04606_),
    .A(_04600_),
    .Y(_04626_),
    .D(_04625_));
 sg13g2_a21oi_1 _10292_ (.A1(_04570_),
    .A2(_04602_),
    .Y(_04627_),
    .B1(_04601_));
 sg13g2_nor2_1 _10293_ (.A(_04603_),
    .B(_04627_),
    .Y(_04628_));
 sg13g2_o21ai_1 _10294_ (.B1(_04604_),
    .Y(_04629_),
    .A1(_04626_),
    .A2(_04627_));
 sg13g2_or2_1 _10295_ (.X(_04630_),
    .B(_04572_),
    .A(_04571_));
 sg13g2_nand2b_1 _10296_ (.Y(_04631_),
    .B(_04630_),
    .A_N(_04573_));
 sg13g2_a21oi_1 _10297_ (.A1(_04629_),
    .A2(_04630_),
    .Y(_04632_),
    .B1(_04573_));
 sg13g2_xor2_1 _10298_ (.B(_04532_),
    .A(_04531_),
    .X(_04633_));
 sg13g2_o21ai_1 _10299_ (.B1(_04533_),
    .Y(_04634_),
    .A1(_04632_),
    .A2(_04633_));
 sg13g2_nand2b_1 _10300_ (.Y(_04635_),
    .B(_04498_),
    .A_N(_04497_));
 sg13g2_nand2b_1 _10301_ (.Y(_04636_),
    .B(_04635_),
    .A_N(_04499_));
 sg13g2_a21o_1 _10302_ (.A2(_04635_),
    .A1(_04634_),
    .B1(_04499_),
    .X(_04637_));
 sg13g2_xor2_1 _10303_ (.B(_04466_),
    .A(_04465_),
    .X(_04638_));
 sg13g2_a21oi_1 _10304_ (.A1(_04637_),
    .A2(_04638_),
    .Y(_04639_),
    .B1(_04467_));
 sg13g2_xnor2_1 _10305_ (.Y(_04640_),
    .A(_04434_),
    .B(_04435_));
 sg13g2_o21ai_1 _10306_ (.B1(_04436_),
    .Y(_04641_),
    .A1(_04639_),
    .A2(_04640_));
 sg13g2_xnor2_1 _10307_ (.Y(_04642_),
    .A(_04403_),
    .B(_04405_));
 sg13g2_inv_1 _10308_ (.Y(_04643_),
    .A(_04642_));
 sg13g2_a21oi_2 _10309_ (.B1(_04406_),
    .Y(_04644_),
    .A2(_04643_),
    .A1(_04641_));
 sg13g2_and2_2 _10310_ (.A(_04385_),
    .B(_04644_),
    .X(_04645_));
 sg13g2_a21oi_1 _10311_ (.A1(_04385_),
    .A2(_04644_),
    .Y(_04646_),
    .B1(_04305_));
 sg13g2_nand3_1 _10312_ (.B(_04385_),
    .C(_04644_),
    .A(_04305_),
    .Y(_04647_));
 sg13g2_nor2b_1 _10313_ (.A(_04646_),
    .B_N(_04647_),
    .Y(_04648_));
 sg13g2_a21oi_1 _10314_ (.A1(_04330_),
    .A2(_04647_),
    .Y(_04649_),
    .B1(_04646_));
 sg13g2_nor2_1 _10315_ (.A(_04296_),
    .B(_04326_),
    .Y(_04650_));
 sg13g2_xor2_1 _10316_ (.B(_04326_),
    .A(_04296_),
    .X(_04651_));
 sg13g2_o21ai_1 _10317_ (.B1(_04372_),
    .Y(_04652_),
    .A1(_04649_),
    .A2(_04650_));
 sg13g2_xnor2_1 _10318_ (.Y(_04653_),
    .A(_04299_),
    .B(_04331_));
 sg13g2_inv_1 _10319_ (.Y(_04654_),
    .A(_04653_));
 sg13g2_a21oi_1 _10320_ (.A1(_04652_),
    .A2(_04654_),
    .Y(_04655_),
    .B1(_04371_));
 sg13g2_a221oi_1 _10321_ (.B2(_04654_),
    .C1(_04371_),
    .B1(_04652_),
    .A1(_04297_),
    .Y(_04656_),
    .A2(_04328_));
 sg13g2_nor3_1 _10322_ (.A(_04369_),
    .B(_04370_),
    .C(_04656_),
    .Y(_04657_));
 sg13g2_a21oi_1 _10323_ (.A1(_04300_),
    .A2(_04333_),
    .Y(_04658_),
    .B1(_04657_));
 sg13g2_o21ai_1 _10324_ (.B1(_04368_),
    .Y(_04659_),
    .A1(_04367_),
    .A2(_04658_));
 sg13g2_a21oi_1 _10325_ (.A1(_04365_),
    .A2(_04659_),
    .Y(_04660_),
    .B1(_04364_));
 sg13g2_o21ai_1 _10326_ (.B1(_04363_),
    .Y(_04661_),
    .A1(_04362_),
    .A2(_04660_));
 sg13g2_and2_1 _10327_ (.A(_04362_),
    .B(_04660_),
    .X(_04662_));
 sg13g2_or2_1 _10328_ (.X(_04663_),
    .B(_04660_),
    .A(_04363_));
 sg13g2_a21oi_2 _10329_ (.B1(_04662_),
    .Y(_04664_),
    .A2(_04663_),
    .A1(_04661_));
 sg13g2_xnor2_1 _10330_ (.Y(_04665_),
    .A(_04366_),
    .B(_04659_));
 sg13g2_o21ai_1 _10331_ (.B1(_04369_),
    .Y(_04666_),
    .A1(_04370_),
    .A2(_04656_));
 sg13g2_nor2b_1 _10332_ (.A(_04657_),
    .B_N(_04666_),
    .Y(_04667_));
 sg13g2_xor2_1 _10333_ (.B(_04651_),
    .A(_04649_),
    .X(_04668_));
 sg13g2_xnor2_1 _10334_ (.Y(_04669_),
    .A(_04330_),
    .B(_04648_));
 sg13g2_nor2_1 _10335_ (.A(_04668_),
    .B(_04669_),
    .Y(_04670_));
 sg13g2_xnor2_1 _10336_ (.Y(_04671_),
    .A(_04652_),
    .B(_04653_));
 sg13g2_nand2_1 _10337_ (.Y(_04672_),
    .A(_04670_),
    .B(_04671_));
 sg13g2_xor2_1 _10338_ (.B(_04328_),
    .A(_04297_),
    .X(_04673_));
 sg13g2_xor2_1 _10339_ (.B(_04673_),
    .A(_04655_),
    .X(_04674_));
 sg13g2_inv_1 _10340_ (.Y(_04675_),
    .A(_04674_));
 sg13g2_nor2_1 _10341_ (.A(_04672_),
    .B(_04674_),
    .Y(_04676_));
 sg13g2_and2_1 _10342_ (.A(_04667_),
    .B(_04676_),
    .X(_04677_));
 sg13g2_nand2b_1 _10343_ (.Y(_04678_),
    .B(_04368_),
    .A_N(_04367_));
 sg13g2_xor2_1 _10344_ (.B(_04678_),
    .A(_04658_),
    .X(_04679_));
 sg13g2_and3_1 _10345_ (.X(_04680_),
    .A(_04665_),
    .B(_04677_),
    .C(_04679_));
 sg13g2_o21ai_1 _10346_ (.B1(_04661_),
    .Y(_04681_),
    .A1(_04664_),
    .A2(_04680_));
 sg13g2_nand2b_1 _10347_ (.Y(_04682_),
    .B(_04662_),
    .A_N(_04680_));
 sg13g2_a22oi_1 _10348_ (.Y(_04683_),
    .B1(_04358_),
    .B2(_04349_),
    .A2(_04354_),
    .A1(_04324_));
 sg13g2_and3_1 _10349_ (.X(_04684_),
    .A(_04681_),
    .B(_04682_),
    .C(_04683_));
 sg13g2_nand3b_1 _10350_ (.B(_04349_),
    .C(_04336_),
    .Y(_04685_),
    .A_N(_04350_));
 sg13g2_o21ai_1 _10351_ (.B1(_04685_),
    .Y(_04686_),
    .A1(_04308_),
    .A2(_04322_));
 sg13g2_or2_2 _10352_ (.X(_04687_),
    .B(_04686_),
    .A(_04662_));
 sg13g2_inv_1 _10353_ (.Y(_04688_),
    .A(_04687_));
 sg13g2_xnor2_1 _10354_ (.Y(_04689_),
    .A(_04667_),
    .B(_04676_));
 sg13g2_nor2b_1 _10355_ (.A(_04668_),
    .B_N(_04669_),
    .Y(_04690_));
 sg13g2_nand4_1 _10356_ (.B(_04675_),
    .C(_04679_),
    .A(_04671_),
    .Y(_04691_),
    .D(_04690_));
 sg13g2_a21oi_1 _10357_ (.A1(_04677_),
    .A2(_04679_),
    .Y(_04692_),
    .B1(_04665_));
 sg13g2_or2_1 _10358_ (.X(_04693_),
    .B(_04692_),
    .A(_04680_));
 sg13g2_or4_1 _10359_ (.A(_04664_),
    .B(_04689_),
    .C(_04691_),
    .D(_04693_),
    .X(_04694_));
 sg13g2_and3_2 _10360_ (.X(_04695_),
    .A(net1417),
    .B(_04688_),
    .C(_04694_));
 sg13g2_xnor2_1 _10361_ (.Y(_04696_),
    .A(_04626_),
    .B(_04628_));
 sg13g2_xnor2_1 _10362_ (.Y(_04697_),
    .A(_04629_),
    .B(_04631_));
 sg13g2_mux2_1 _10363_ (.A0(_04697_),
    .A1(_04696_),
    .S(_04645_),
    .X(_04698_));
 sg13g2_nand2_1 _10364_ (.Y(_04699_),
    .A(_04695_),
    .B(_04698_));
 sg13g2_a22oi_1 _10365_ (.Y(_00366_),
    .B1(net1482),
    .B2(_04699_),
    .A2(net1647),
    .A1(_00725_));
 sg13g2_xor2_1 _10366_ (.B(_04633_),
    .A(_04632_),
    .X(_04700_));
 sg13g2_mux2_1 _10367_ (.A0(_04700_),
    .A1(_04697_),
    .S(_04645_),
    .X(_04701_));
 sg13g2_nand2_1 _10368_ (.Y(_04702_),
    .A(_04695_),
    .B(_04701_));
 sg13g2_a22oi_1 _10369_ (.Y(_00367_),
    .B1(net1482),
    .B2(_04702_),
    .A2(net1647),
    .A1(_00724_));
 sg13g2_xnor2_1 _10370_ (.Y(_04703_),
    .A(_04634_),
    .B(_04636_));
 sg13g2_mux2_1 _10371_ (.A0(_04703_),
    .A1(_04700_),
    .S(_04645_),
    .X(_04704_));
 sg13g2_nand2_1 _10372_ (.Y(_04705_),
    .A(_04695_),
    .B(_04704_));
 sg13g2_a22oi_1 _10373_ (.Y(_00368_),
    .B1(net1482),
    .B2(_04705_),
    .A2(net1647),
    .A1(_00727_));
 sg13g2_xor2_1 _10374_ (.B(_04638_),
    .A(_04637_),
    .X(_04706_));
 sg13g2_mux2_1 _10375_ (.A0(_04706_),
    .A1(_04703_),
    .S(_04645_),
    .X(_04707_));
 sg13g2_nand2_1 _10376_ (.Y(_04708_),
    .A(_04695_),
    .B(_04707_));
 sg13g2_a22oi_1 _10377_ (.Y(_00369_),
    .B1(net1482),
    .B2(_04708_),
    .A2(net1647),
    .A1(_00726_));
 sg13g2_xor2_1 _10378_ (.B(_04640_),
    .A(_04639_),
    .X(_04709_));
 sg13g2_mux2_1 _10379_ (.A0(_04709_),
    .A1(_04706_),
    .S(_04645_),
    .X(_04710_));
 sg13g2_nand2_1 _10380_ (.Y(_04711_),
    .A(_04695_),
    .B(_04710_));
 sg13g2_a22oi_1 _10381_ (.Y(_00370_),
    .B1(net1482),
    .B2(_04711_),
    .A2(net1647),
    .A1(_00730_));
 sg13g2_xnor2_1 _10382_ (.Y(_04712_),
    .A(_04641_),
    .B(_04642_));
 sg13g2_mux2_1 _10383_ (.A0(_04712_),
    .A1(_04709_),
    .S(_04645_),
    .X(_04713_));
 sg13g2_nand2_1 _10384_ (.Y(_04714_),
    .A(_04695_),
    .B(_04713_));
 sg13g2_a22oi_1 _10385_ (.Y(_00371_),
    .B1(net1482),
    .B2(_04714_),
    .A2(net1647),
    .A1(_00729_));
 sg13g2_nor2_1 _10386_ (.A(_04386_),
    .B(_04712_),
    .Y(_04715_));
 sg13g2_nand2_1 _10387_ (.Y(_04716_),
    .A(_04377_),
    .B(_04394_));
 sg13g2_a21oi_1 _10388_ (.A1(_04373_),
    .A2(_04716_),
    .Y(_04717_),
    .B1(_04384_));
 sg13g2_xnor2_1 _10389_ (.Y(_04718_),
    .A(_04644_),
    .B(_04717_));
 sg13g2_nand3b_1 _10390_ (.B(_04718_),
    .C(_04695_),
    .Y(_04719_),
    .A_N(_04715_));
 sg13g2_a22oi_1 _10391_ (.Y(_00372_),
    .B1(net1482),
    .B2(_04719_),
    .A2(net1647),
    .A1(_00728_));
 sg13g2_nand2b_1 _10392_ (.Y(_04720_),
    .B(net1417),
    .A_N(_04669_));
 sg13g2_nand2_1 _10393_ (.Y(_04721_),
    .A(_04688_),
    .B(_04720_));
 sg13g2_a22oi_1 _10394_ (.Y(_00373_),
    .B1(_04361_),
    .B2(_04721_),
    .A2(net1648),
    .A1(_00732_));
 sg13g2_xnor2_1 _10395_ (.Y(_04722_),
    .A(_04668_),
    .B(_04669_));
 sg13g2_a21o_1 _10396_ (.A2(_04722_),
    .A1(_04684_),
    .B1(_04687_),
    .X(_04723_));
 sg13g2_a22oi_1 _10397_ (.Y(_00374_),
    .B1(net1483),
    .B2(_04723_),
    .A2(net1646),
    .A1(_00733_));
 sg13g2_xnor2_1 _10398_ (.Y(_04724_),
    .A(_04670_),
    .B(_04671_));
 sg13g2_a21o_1 _10399_ (.A2(_04724_),
    .A1(net1417),
    .B1(_04687_),
    .X(_04725_));
 sg13g2_a22oi_1 _10400_ (.Y(_00375_),
    .B1(net1483),
    .B2(_04725_),
    .A2(net1644),
    .A1(_00734_));
 sg13g2_xnor2_1 _10401_ (.Y(_04726_),
    .A(_04672_),
    .B(_04674_));
 sg13g2_a21o_1 _10402_ (.A2(_04726_),
    .A1(net1417),
    .B1(_04687_),
    .X(_04727_));
 sg13g2_a22oi_1 _10403_ (.Y(_00376_),
    .B1(net1483),
    .B2(_04727_),
    .A2(net1644),
    .A1(_00735_));
 sg13g2_a21o_1 _10404_ (.A2(_04689_),
    .A1(net1417),
    .B1(_04687_),
    .X(_04728_));
 sg13g2_a22oi_1 _10405_ (.Y(_00377_),
    .B1(net1483),
    .B2(_04728_),
    .A2(net1644),
    .A1(_00736_));
 sg13g2_xnor2_1 _10406_ (.Y(_04729_),
    .A(_04677_),
    .B(_04679_));
 sg13g2_a21o_1 _10407_ (.A2(_04729_),
    .A1(net1417),
    .B1(_04687_),
    .X(_04730_));
 sg13g2_a22oi_1 _10408_ (.Y(_00378_),
    .B1(net1483),
    .B2(_04730_),
    .A2(net1644),
    .A1(_00737_));
 sg13g2_a21o_1 _10409_ (.A2(_04693_),
    .A1(net1417),
    .B1(_04687_),
    .X(_04731_));
 sg13g2_a22oi_1 _10410_ (.Y(_00379_),
    .B1(net1483),
    .B2(_04731_),
    .A2(net1644),
    .A1(_00738_));
 sg13g2_xor2_1 _10411_ (.B(_04680_),
    .A(_04664_),
    .X(_04732_));
 sg13g2_a21o_1 _10412_ (.A2(_04732_),
    .A1(net1417),
    .B1(_04687_),
    .X(_04733_));
 sg13g2_a22oi_1 _10413_ (.Y(_00380_),
    .B1(net1483),
    .B2(_04733_),
    .A2(net1644),
    .A1(_00739_));
 sg13g2_xor2_1 _10414_ (.B(_04350_),
    .A(_04321_),
    .X(_04734_));
 sg13g2_nand2_1 _10415_ (.Y(_04735_),
    .A(_04688_),
    .B(_04734_));
 sg13g2_a22oi_1 _10416_ (.Y(_00381_),
    .B1(net1482),
    .B2(_04735_),
    .A2(net1647),
    .A1(_00731_));
 sg13g2_nor2_2 _10417_ (.A(\u_tiny_nn_top.state_q[16] ),
    .B(\u_tiny_nn_top.state_q[2] ),
    .Y(_04736_));
 sg13g2_and2_1 _10418_ (.A(net1766),
    .B(net1745),
    .X(_04737_));
 sg13g2_nand2_1 _10419_ (.Y(_04738_),
    .A(net1766),
    .B(net1745));
 sg13g2_nor4_1 _10420_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[12] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[11] ),
    .C(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[14] ),
    .D(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[13] ),
    .Y(_04739_));
 sg13g2_nor4_1 _10421_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[8] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[7] ),
    .C(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[10] ),
    .D(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[9] ),
    .Y(_04740_));
 sg13g2_and2_1 _10422_ (.A(_04739_),
    .B(_04740_),
    .X(_04741_));
 sg13g2_nor4_1 _10423_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[11] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[12] ),
    .C(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[13] ),
    .D(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[14] ),
    .Y(_04742_));
 sg13g2_nor4_1 _10424_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[7] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[8] ),
    .C(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[9] ),
    .D(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[10] ),
    .Y(_04743_));
 sg13g2_and2_1 _10425_ (.A(_04742_),
    .B(_04743_),
    .X(_04744_));
 sg13g2_a22oi_1 _10426_ (.Y(_04745_),
    .B1(_04744_),
    .B2(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[15] ),
    .A2(_04741_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[15] ));
 sg13g2_nand4_1 _10427_ (.B(_00743_),
    .C(_00745_),
    .A(_00742_),
    .Y(_04746_),
    .D(_00746_));
 sg13g2_nor3_1 _10428_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[1] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[0] ),
    .C(_04746_),
    .Y(_04747_));
 sg13g2_nand2_1 _10429_ (.Y(_04748_),
    .A(_00116_),
    .B(_04747_));
 sg13g2_nand4_1 _10430_ (.B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[11] ),
    .C(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[14] ),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[12] ),
    .Y(_04749_),
    .D(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[13] ));
 sg13g2_nand3_1 _10431_ (.B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[7] ),
    .C(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[10] ),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[8] ),
    .Y(_04750_));
 sg13g2_nor3_1 _10432_ (.A(_00751_),
    .B(_04749_),
    .C(_04750_),
    .Y(_04751_));
 sg13g2_o21ai_1 _10433_ (.B1(_04748_),
    .Y(_04752_),
    .A1(_04741_),
    .A2(_04751_));
 sg13g2_nand4_1 _10434_ (.B(_00727_),
    .C(_00729_),
    .A(_00726_),
    .Y(_04753_),
    .D(_00730_));
 sg13g2_nor3_1 _10435_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[1] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[0] ),
    .C(_04753_),
    .Y(_04754_));
 sg13g2_nand2_1 _10436_ (.Y(_04755_),
    .A(_00115_),
    .B(_04754_));
 sg13g2_nand4_1 _10437_ (.B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[12] ),
    .C(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[13] ),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[11] ),
    .Y(_04756_),
    .D(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[14] ));
 sg13g2_nand3_1 _10438_ (.B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[8] ),
    .C(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[9] ),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[7] ),
    .Y(_04757_));
 sg13g2_nor3_1 _10439_ (.A(_00735_),
    .B(_04756_),
    .C(_04757_),
    .Y(_04758_));
 sg13g2_o21ai_1 _10440_ (.B1(_04755_),
    .Y(_04759_),
    .A1(_04744_),
    .A2(_04758_));
 sg13g2_nand4_1 _10441_ (.B(_04745_),
    .C(_04752_),
    .A(net1743),
    .Y(_04760_),
    .D(_04759_));
 sg13g2_and2_1 _10442_ (.A(_00728_),
    .B(_04754_),
    .X(_04761_));
 sg13g2_nand2_1 _10443_ (.Y(_04762_),
    .A(_04758_),
    .B(_04761_));
 sg13g2_and2_1 _10444_ (.A(_00744_),
    .B(_04747_),
    .X(_04763_));
 sg13g2_and2_1 _10445_ (.A(_04751_),
    .B(_04763_),
    .X(_04764_));
 sg13g2_a21oi_1 _10446_ (.A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[15] ),
    .A2(_04764_),
    .Y(_04765_),
    .B1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[15] ));
 sg13g2_nor2_1 _10447_ (.A(_04762_),
    .B(_04765_),
    .Y(_04766_));
 sg13g2_a21o_1 _10448_ (.A2(_04764_),
    .A1(_00747_),
    .B1(_00731_),
    .X(_04767_));
 sg13g2_a21oi_2 _10449_ (.B1(_04760_),
    .Y(_04768_),
    .A2(_04767_),
    .A1(_04766_));
 sg13g2_and2_1 _10450_ (.A(net1732),
    .B(_04768_),
    .X(_04769_));
 sg13g2_and3_2 _10451_ (.X(_04770_),
    .A(_00747_),
    .B(_04741_),
    .C(_04763_));
 sg13g2_nor2_2 _10452_ (.A(_00739_),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[14] ),
    .Y(_04771_));
 sg13g2_nand2_2 _10453_ (.Y(_04772_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[14] ),
    .B(_00754_));
 sg13g2_nor2_1 _10454_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[12] ),
    .B(_00752_),
    .Y(_04773_));
 sg13g2_nand2_1 _10455_ (.Y(_04774_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[11] ),
    .B(_00753_));
 sg13g2_nand2b_1 _10456_ (.Y(_04775_),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[8] ),
    .A_N(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[8] ));
 sg13g2_nor2b_1 _10457_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[7] ),
    .B_N(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[7] ),
    .Y(_04776_));
 sg13g2_nor2b_1 _10458_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[8] ),
    .B_N(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[8] ),
    .Y(_04777_));
 sg13g2_a221oi_1 _10459_ (.B2(_04776_),
    .C1(_04777_),
    .B1(_04775_),
    .A1(_00734_),
    .Y(_04778_),
    .A2(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[9] ));
 sg13g2_nand2b_1 _10460_ (.Y(_04779_),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[10] ),
    .A_N(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[10] ));
 sg13g2_o21ai_1 _10461_ (.B1(_04779_),
    .Y(_04780_),
    .A1(_00734_),
    .A2(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[9] ));
 sg13g2_a22oi_1 _10462_ (.Y(_04781_),
    .B1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[11] ),
    .B2(_00736_),
    .A2(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[10] ),
    .A1(_00735_));
 sg13g2_o21ai_1 _10463_ (.B1(_04781_),
    .Y(_04782_),
    .A1(_04778_),
    .A2(_04780_));
 sg13g2_a21o_1 _10464_ (.A2(_04782_),
    .A1(_04774_),
    .B1(_04773_),
    .X(_04783_));
 sg13g2_nand2_1 _10465_ (.Y(_04784_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[13] ),
    .B(_00755_));
 sg13g2_a22oi_1 _10466_ (.Y(_04785_),
    .B1(_00755_),
    .B2(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[13] ),
    .A2(_00752_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[12] ));
 sg13g2_nand2_2 _10467_ (.Y(_04786_),
    .A(_00739_),
    .B(_00754_));
 sg13g2_xnor2_1 _10468_ (.Y(_04787_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[14] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[14] ));
 sg13g2_nand2_1 _10469_ (.Y(_04788_),
    .A(_00738_),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[13] ));
 sg13g2_nand2_1 _10470_ (.Y(_04789_),
    .A(_04787_),
    .B(_04788_));
 sg13g2_a21oi_2 _10471_ (.B1(_04789_),
    .Y(_04790_),
    .A2(_04785_),
    .A1(_04783_));
 sg13g2_a21o_1 _10472_ (.A2(_04785_),
    .A1(_04783_),
    .B1(_04789_),
    .X(_04791_));
 sg13g2_nand2_1 _10473_ (.Y(_04792_),
    .A(net1731),
    .B(net1532));
 sg13g2_nand2b_1 _10474_ (.Y(_04793_),
    .B(net1520),
    .A_N(_00124_));
 sg13g2_mux2_2 _10475_ (.A0(_00123_),
    .A1(_00124_),
    .S(net1520),
    .X(_04794_));
 sg13g2_o21ai_1 _10476_ (.B1(_04793_),
    .Y(_04795_),
    .A1(_00123_),
    .A2(net1520));
 sg13g2_nand2b_1 _10477_ (.Y(_04796_),
    .B(net1520),
    .A_N(_00123_));
 sg13g2_mux2_2 _10478_ (.A0(_00124_),
    .A1(_00123_),
    .S(net1520),
    .X(_04797_));
 sg13g2_o21ai_1 _10479_ (.B1(_04796_),
    .Y(_04798_),
    .A1(_00124_),
    .A2(net1518));
 sg13g2_xnor2_1 _10480_ (.Y(_04799_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[10] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[10] ));
 sg13g2_xor2_1 _10481_ (.B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[10] ),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[10] ),
    .X(_04800_));
 sg13g2_xor2_1 _10482_ (.B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[11] ),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[11] ),
    .X(_04801_));
 sg13g2_xor2_1 _10483_ (.B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[9] ),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[9] ),
    .X(_04802_));
 sg13g2_inv_1 _10484_ (.Y(_04803_),
    .A(_04802_));
 sg13g2_xnor2_1 _10485_ (.Y(_04804_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[8] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[8] ));
 sg13g2_and3_1 _10486_ (.X(_04805_),
    .A(_00120_),
    .B(_04772_),
    .C(_04791_));
 sg13g2_a21oi_2 _10487_ (.B1(_00756_),
    .Y(_04806_),
    .A2(_04791_),
    .A1(_04772_));
 sg13g2_or2_1 _10488_ (.X(_04807_),
    .B(_04806_),
    .A(_04805_));
 sg13g2_nor2_2 _10489_ (.A(_04805_),
    .B(_04806_),
    .Y(_04808_));
 sg13g2_nand2_1 _10490_ (.Y(_04809_),
    .A(_00119_),
    .B(_00120_));
 sg13g2_o21ai_1 _10491_ (.B1(_04809_),
    .Y(_04810_),
    .A1(_04805_),
    .A2(_04806_));
 sg13g2_a21o_1 _10492_ (.A2(net1532),
    .A1(net1731),
    .B1(_00127_),
    .X(_04811_));
 sg13g2_nand3b_1 _10493_ (.B(_04772_),
    .C(_04791_),
    .Y(_04812_),
    .A_N(_00128_));
 sg13g2_nand2_1 _10494_ (.Y(_04813_),
    .A(_04811_),
    .B(_04812_));
 sg13g2_a22oi_1 _10495_ (.Y(_04814_),
    .B1(_04812_),
    .B2(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[8] ),
    .A2(_04811_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[8] ));
 sg13g2_a22oi_1 _10496_ (.Y(_04815_),
    .B1(net1505),
    .B2(_04814_),
    .A2(_04810_),
    .A1(_04804_));
 sg13g2_a221oi_1 _10497_ (.B2(_04814_),
    .C1(_04802_),
    .B1(net1505),
    .A1(_04804_),
    .Y(_04816_),
    .A2(_04810_));
 sg13g2_o21ai_1 _10498_ (.B1(_04799_),
    .Y(_04817_),
    .A1(_04801_),
    .A2(_04816_));
 sg13g2_nand3_1 _10499_ (.B(net1731),
    .C(net1532),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[10] ),
    .Y(_04818_));
 sg13g2_o21ai_1 _10500_ (.B1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[10] ),
    .Y(_04819_),
    .A1(_04771_),
    .A2(_04790_));
 sg13g2_nand2_1 _10501_ (.Y(_04820_),
    .A(_04818_),
    .B(_04819_));
 sg13g2_and2_2 _10502_ (.A(_04818_),
    .B(_04819_),
    .X(_04821_));
 sg13g2_nand3_1 _10503_ (.B(net1731),
    .C(net1532),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[12] ),
    .Y(_04822_));
 sg13g2_o21ai_1 _10504_ (.B1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[12] ),
    .Y(_04823_),
    .A1(_04771_),
    .A2(_04790_));
 sg13g2_nand2_1 _10505_ (.Y(_04824_),
    .A(_04822_),
    .B(_04823_));
 sg13g2_and2_1 _10506_ (.A(_04822_),
    .B(_04823_),
    .X(_04825_));
 sg13g2_o21ai_1 _10507_ (.B1(_00736_),
    .Y(_04826_),
    .A1(_04771_),
    .A2(_04790_));
 sg13g2_nand3_1 _10508_ (.B(net1731),
    .C(net1532),
    .A(_00753_),
    .Y(_04827_));
 sg13g2_and2_1 _10509_ (.A(_04826_),
    .B(_04827_),
    .X(_04828_));
 sg13g2_nand2_1 _10510_ (.Y(_04829_),
    .A(_04826_),
    .B(_04827_));
 sg13g2_xnor2_1 _10511_ (.Y(_04830_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[12] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[12] ));
 sg13g2_a21oi_1 _10512_ (.A1(_04826_),
    .A2(_04827_),
    .Y(_04831_),
    .B1(_04830_));
 sg13g2_a221oi_1 _10513_ (.B2(_04827_),
    .C1(_04830_),
    .B1(_04826_),
    .A1(_04822_),
    .Y(_04832_),
    .A2(_04823_));
 sg13g2_nand2_1 _10514_ (.Y(_04833_),
    .A(_04784_),
    .B(_04788_));
 sg13g2_and3_1 _10515_ (.X(_04834_),
    .A(_04826_),
    .B(_04827_),
    .C(_04830_));
 sg13g2_nor3_1 _10516_ (.A(_04832_),
    .B(_04833_),
    .C(_04834_),
    .Y(_04835_));
 sg13g2_o21ai_1 _10517_ (.B1(_04801_),
    .Y(_04836_),
    .A1(_04820_),
    .A2(_04835_));
 sg13g2_nor2_1 _10518_ (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[13] ),
    .B(net1521),
    .Y(_04837_));
 sg13g2_a21oi_1 _10519_ (.A1(_00738_),
    .A2(net1521),
    .Y(_04838_),
    .B1(_04837_));
 sg13g2_mux2_1 _10520_ (.A0(_00755_),
    .A1(_00738_),
    .S(net1521),
    .X(_04839_));
 sg13g2_a21oi_1 _10521_ (.A1(_04833_),
    .A2(_04839_),
    .Y(_04840_),
    .B1(_04787_));
 sg13g2_a22oi_1 _10522_ (.Y(_04841_),
    .B1(_04825_),
    .B2(_04831_),
    .A2(_04788_),
    .A1(_04784_));
 sg13g2_nand3_1 _10523_ (.B(net1731),
    .C(net1532),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[9] ),
    .Y(_04842_));
 sg13g2_o21ai_1 _10524_ (.B1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[9] ),
    .Y(_04843_),
    .A1(_04771_),
    .A2(_04790_));
 sg13g2_nand2_2 _10525_ (.Y(_04844_),
    .A(_04842_),
    .B(_04843_));
 sg13g2_and2_1 _10526_ (.A(_04842_),
    .B(_04843_),
    .X(_04845_));
 sg13g2_and3_1 _10527_ (.X(_04846_),
    .A(_04800_),
    .B(_04842_),
    .C(_04843_));
 sg13g2_a21oi_1 _10528_ (.A1(_04842_),
    .A2(_04843_),
    .Y(_04847_),
    .B1(_04800_));
 sg13g2_nor3_1 _10529_ (.A(_04803_),
    .B(_04846_),
    .C(_04847_),
    .Y(_04848_));
 sg13g2_nand3_1 _10530_ (.B(_04818_),
    .C(_04819_),
    .A(_04800_),
    .Y(_04849_));
 sg13g2_a21oi_1 _10531_ (.A1(_04830_),
    .A2(_04849_),
    .Y(_04850_),
    .B1(_04801_));
 sg13g2_nor4_1 _10532_ (.A(_04840_),
    .B(_04841_),
    .C(_04848_),
    .D(_04850_),
    .Y(_04851_));
 sg13g2_or3_1 _10533_ (.A(_04799_),
    .B(_04802_),
    .C(_04815_),
    .X(_04852_));
 sg13g2_nand4_1 _10534_ (.B(_04836_),
    .C(_04851_),
    .A(_04817_),
    .Y(_04853_),
    .D(_04852_));
 sg13g2_nor2_1 _10535_ (.A(_04797_),
    .B(_04853_),
    .Y(_04854_));
 sg13g2_nor2_2 _10536_ (.A(_04795_),
    .B(_04854_),
    .Y(_04855_));
 sg13g2_xnor2_1 _10537_ (.Y(_04856_),
    .A(_04794_),
    .B(_04854_));
 sg13g2_xnor2_1 _10538_ (.Y(_04857_),
    .A(_04802_),
    .B(_04815_));
 sg13g2_xnor2_1 _10539_ (.Y(_04858_),
    .A(_04803_),
    .B(_04815_));
 sg13g2_nor2_2 _10540_ (.A(_04853_),
    .B(_04858_),
    .Y(_04859_));
 sg13g2_a21oi_2 _10541_ (.B1(_04853_),
    .Y(_04860_),
    .A2(_04858_),
    .A1(_04797_));
 sg13g2_inv_1 _10542_ (.Y(_04861_),
    .A(_04860_));
 sg13g2_xor2_1 _10543_ (.B(_04810_),
    .A(_04804_),
    .X(_04862_));
 sg13g2_xnor2_1 _10544_ (.Y(_04863_),
    .A(_04804_),
    .B(_04810_));
 sg13g2_xnor2_1 _10545_ (.Y(_04864_),
    .A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[7] ),
    .B(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[7] ));
 sg13g2_nand3_1 _10546_ (.B(net1731),
    .C(net1532),
    .A(_00118_),
    .Y(_04865_));
 sg13g2_o21ai_1 _10547_ (.B1(_00117_),
    .Y(_04866_),
    .A1(_04771_),
    .A2(_04790_));
 sg13g2_nand2_2 _10548_ (.Y(_04867_),
    .A(_04865_),
    .B(_04866_));
 sg13g2_inv_1 _10549_ (.Y(_04868_),
    .A(_04867_));
 sg13g2_nand3_1 _10550_ (.B(net1731),
    .C(net1532),
    .A(_00126_),
    .Y(_04869_));
 sg13g2_o21ai_1 _10551_ (.B1(_00125_),
    .Y(_04870_),
    .A1(_04771_),
    .A2(_04790_));
 sg13g2_nand2_2 _10552_ (.Y(_04871_),
    .A(_04869_),
    .B(_04870_));
 sg13g2_a22oi_1 _10553_ (.Y(_04872_),
    .B1(_04869_),
    .B2(_04870_),
    .A2(_04866_),
    .A1(_04865_));
 sg13g2_mux2_2 _10554_ (.A0(_00122_),
    .A1(_00121_),
    .S(net1518),
    .X(_04873_));
 sg13g2_nor2_1 _10555_ (.A(_04797_),
    .B(_04872_),
    .Y(_04874_));
 sg13g2_xnor2_1 _10556_ (.Y(_04875_),
    .A(_04873_),
    .B(_04874_));
 sg13g2_nand2_1 _10557_ (.Y(_04876_),
    .A(_04872_),
    .B(_04873_));
 sg13g2_mux2_1 _10558_ (.A0(_00132_),
    .A1(_00131_),
    .S(net1518),
    .X(_04877_));
 sg13g2_inv_1 _10559_ (.Y(_04878_),
    .A(_04877_));
 sg13g2_mux2_1 _10560_ (.A0(_00130_),
    .A1(_00129_),
    .S(net1518),
    .X(_04879_));
 sg13g2_nand4_1 _10561_ (.B(_04873_),
    .C(_04877_),
    .A(_04872_),
    .Y(_04880_),
    .D(_04879_));
 sg13g2_mux2_1 _10562_ (.A0(_00134_),
    .A1(_00133_),
    .S(net1519),
    .X(_04881_));
 sg13g2_inv_1 _10563_ (.Y(_04882_),
    .A(_04881_));
 sg13g2_a21oi_1 _10564_ (.A1(_04872_),
    .A2(_04873_),
    .Y(_04883_),
    .B1(_04797_));
 sg13g2_a21oi_1 _10565_ (.A1(_04798_),
    .A2(_04878_),
    .Y(_04884_),
    .B1(_04883_));
 sg13g2_nand2_1 _10566_ (.Y(_04885_),
    .A(_04798_),
    .B(_04880_));
 sg13g2_o21ai_1 _10567_ (.B1(_04798_),
    .Y(_04886_),
    .A1(_04880_),
    .A2(_04882_));
 sg13g2_mux2_1 _10568_ (.A0(_00115_),
    .A1(_00116_),
    .S(net1519),
    .X(_04887_));
 sg13g2_a21o_1 _10569_ (.A2(_04887_),
    .A1(_04886_),
    .B1(_04797_),
    .X(_04888_));
 sg13g2_nor2_1 _10570_ (.A(_04797_),
    .B(net1742),
    .Y(_04889_));
 sg13g2_a21oi_1 _10571_ (.A1(net1742),
    .A2(_04888_),
    .Y(_04890_),
    .B1(_04889_));
 sg13g2_mux2_1 _10572_ (.A0(_04797_),
    .A1(_04890_),
    .S(_04863_),
    .X(_04891_));
 sg13g2_a21oi_1 _10573_ (.A1(_04857_),
    .A2(_04891_),
    .Y(_04892_),
    .B1(_04861_));
 sg13g2_mux2_2 _10574_ (.A0(_00117_),
    .A1(_00118_),
    .S(net1520),
    .X(_04893_));
 sg13g2_mux2_1 _10575_ (.A0(_00125_),
    .A1(_00126_),
    .S(net1520),
    .X(_04894_));
 sg13g2_nor2_1 _10576_ (.A(_04794_),
    .B(_04893_),
    .Y(_04895_));
 sg13g2_a21oi_1 _10577_ (.A1(_04893_),
    .A2(_04894_),
    .Y(_04896_),
    .B1(_04794_));
 sg13g2_mux2_1 _10578_ (.A0(_00121_),
    .A1(_00122_),
    .S(net1518),
    .X(_04897_));
 sg13g2_nand2b_1 _10579_ (.Y(_04898_),
    .B(_04897_),
    .A_N(_04896_));
 sg13g2_nand2_1 _10580_ (.Y(_04899_),
    .A(_04795_),
    .B(_04898_));
 sg13g2_nand2b_1 _10581_ (.Y(_04900_),
    .B(net1518),
    .A_N(_00132_));
 sg13g2_o21ai_1 _10582_ (.B1(_04900_),
    .Y(_04901_),
    .A1(_00131_),
    .A2(net1518));
 sg13g2_o21ai_1 _10583_ (.B1(_04795_),
    .Y(_04902_),
    .A1(_04898_),
    .A2(_04901_));
 sg13g2_mux2_1 _10584_ (.A0(_00129_),
    .A1(_00130_),
    .S(net1518),
    .X(_04903_));
 sg13g2_mux2_1 _10585_ (.A0(_00133_),
    .A1(_00134_),
    .S(net1519),
    .X(_04904_));
 sg13g2_a21o_1 _10586_ (.A2(_04903_),
    .A1(_04902_),
    .B1(_04794_),
    .X(_04905_));
 sg13g2_o21ai_1 _10587_ (.B1(_04905_),
    .Y(_04906_),
    .A1(_04794_),
    .A2(_04904_));
 sg13g2_nand2b_1 _10588_ (.Y(_04907_),
    .B(net1520),
    .A_N(_00115_));
 sg13g2_o21ai_1 _10589_ (.B1(_04907_),
    .Y(_04908_),
    .A1(_00116_),
    .A2(net1521));
 sg13g2_a21oi_1 _10590_ (.A1(_04795_),
    .A2(_04908_),
    .Y(_04909_),
    .B1(_04906_));
 sg13g2_and2_1 _10591_ (.A(_04892_),
    .B(_04909_),
    .X(_04910_));
 sg13g2_xor2_1 _10592_ (.B(_04887_),
    .A(_04886_),
    .X(_04911_));
 sg13g2_mux2_1 _10593_ (.A0(_04888_),
    .A1(_04911_),
    .S(net1742),
    .X(_04912_));
 sg13g2_mux2_1 _10594_ (.A0(_04798_),
    .A1(_04912_),
    .S(_04863_),
    .X(_04913_));
 sg13g2_o21ai_1 _10595_ (.B1(_04860_),
    .Y(_04914_),
    .A1(_04858_),
    .A2(_04913_));
 sg13g2_xor2_1 _10596_ (.B(_04908_),
    .A(_04906_),
    .X(_04915_));
 sg13g2_nor2b_1 _10597_ (.A(_04914_),
    .B_N(_04915_),
    .Y(_04916_));
 sg13g2_xor2_1 _10598_ (.B(_04915_),
    .A(_04914_),
    .X(_04917_));
 sg13g2_inv_1 _10599_ (.Y(_04918_),
    .A(_04917_));
 sg13g2_xnor2_1 _10600_ (.Y(_04919_),
    .A(_04882_),
    .B(_04885_));
 sg13g2_mux4_1 _10601_ (.S0(net1742),
    .A0(_04798_),
    .A1(_04888_),
    .A2(_04911_),
    .A3(_04919_),
    .S1(_04863_),
    .X(_04920_));
 sg13g2_o21ai_1 _10602_ (.B1(_04860_),
    .Y(_04921_),
    .A1(_04858_),
    .A2(_04920_));
 sg13g2_xor2_1 _10603_ (.B(_04905_),
    .A(_04904_),
    .X(_04922_));
 sg13g2_nor2b_1 _10604_ (.A(_04921_),
    .B_N(_04922_),
    .Y(_04923_));
 sg13g2_nand2b_1 _10605_ (.Y(_04924_),
    .B(_04919_),
    .A_N(net1741));
 sg13g2_xor2_1 _10606_ (.B(_04884_),
    .A(_04879_),
    .X(_04925_));
 sg13g2_nand2_1 _10607_ (.Y(_04926_),
    .A(net1742),
    .B(_04925_));
 sg13g2_mux4_1 _10608_ (.S0(net1742),
    .A0(_04888_),
    .A1(_04911_),
    .A2(_04919_),
    .A3(_04925_),
    .S1(_04863_),
    .X(_04927_));
 sg13g2_o21ai_1 _10609_ (.B1(_04860_),
    .Y(_04928_),
    .A1(_04858_),
    .A2(_04927_));
 sg13g2_xnor2_1 _10610_ (.Y(_04929_),
    .A(_04902_),
    .B(_04903_));
 sg13g2_nor2_1 _10611_ (.A(_04928_),
    .B(_04929_),
    .Y(_04930_));
 sg13g2_xor2_1 _10612_ (.B(_04929_),
    .A(_04928_),
    .X(_04931_));
 sg13g2_nor2_2 _10613_ (.A(_04853_),
    .B(_04857_),
    .Y(_04932_));
 sg13g2_nor2b_1 _10614_ (.A(_04891_),
    .B_N(_04932_),
    .Y(_04933_));
 sg13g2_xnor2_1 _10615_ (.Y(_04934_),
    .A(_04877_),
    .B(_04883_));
 sg13g2_mux4_1 _10616_ (.S0(net1741),
    .A0(_04911_),
    .A1(_04919_),
    .A2(_04925_),
    .A3(_04934_),
    .S1(_04863_),
    .X(_04935_));
 sg13g2_a21o_1 _10617_ (.A2(_04935_),
    .A1(_04859_),
    .B1(_04933_),
    .X(_04936_));
 sg13g2_xnor2_1 _10618_ (.Y(_04937_),
    .A(_04899_),
    .B(_04901_));
 sg13g2_and2_1 _10619_ (.A(_04936_),
    .B(_04937_),
    .X(_04938_));
 sg13g2_nand3_1 _10620_ (.B(_04924_),
    .C(_04926_),
    .A(_04862_),
    .Y(_04939_));
 sg13g2_and2_1 _10621_ (.A(net1741),
    .B(_04875_),
    .X(_04940_));
 sg13g2_nor2b_1 _10622_ (.A(net1741),
    .B_N(_04934_),
    .Y(_04941_));
 sg13g2_nor3_1 _10623_ (.A(_04862_),
    .B(_04940_),
    .C(_04941_),
    .Y(_04942_));
 sg13g2_nor2b_1 _10624_ (.A(_04942_),
    .B_N(_04859_),
    .Y(_04943_));
 sg13g2_a22oi_1 _10625_ (.Y(_04944_),
    .B1(_04939_),
    .B2(_04943_),
    .A2(_04932_),
    .A1(_04913_));
 sg13g2_xor2_1 _10626_ (.B(_04897_),
    .A(_04896_),
    .X(_04945_));
 sg13g2_nor2_1 _10627_ (.A(_04944_),
    .B(_04945_),
    .Y(_04946_));
 sg13g2_nor2_1 _10628_ (.A(_04797_),
    .B(_04867_),
    .Y(_04947_));
 sg13g2_xnor2_1 _10629_ (.Y(_04948_),
    .A(_04871_),
    .B(_04947_));
 sg13g2_mux2_1 _10630_ (.A0(_04875_),
    .A1(_04948_),
    .S(net1741),
    .X(_04949_));
 sg13g2_mux4_1 _10631_ (.S0(_04862_),
    .A0(_04875_),
    .A1(_04925_),
    .A2(_04948_),
    .A3(_04934_),
    .S1(net1741),
    .X(_04950_));
 sg13g2_a22oi_1 _10632_ (.Y(_04951_),
    .B1(_04950_),
    .B2(_04859_),
    .A2(_04932_),
    .A1(_04920_));
 sg13g2_xnor2_1 _10633_ (.Y(_04952_),
    .A(_04894_),
    .B(_04895_));
 sg13g2_nor2b_1 _10634_ (.A(_04951_),
    .B_N(_04952_),
    .Y(_04953_));
 sg13g2_mux4_1 _10635_ (.S0(_04862_),
    .A0(_04948_),
    .A1(_04934_),
    .A2(_04868_),
    .A3(_04875_),
    .S1(net1741),
    .X(_04954_));
 sg13g2_a22oi_1 _10636_ (.Y(_04955_),
    .B1(_04954_),
    .B2(_04859_),
    .A2(_04932_),
    .A1(_04927_));
 sg13g2_nor2_1 _10637_ (.A(_04893_),
    .B(_04955_),
    .Y(_04956_));
 sg13g2_xnor2_1 _10638_ (.Y(_04957_),
    .A(_04951_),
    .B(_04952_));
 sg13g2_a21o_1 _10639_ (.A2(_04957_),
    .A1(_04956_),
    .B1(_04953_),
    .X(_04958_));
 sg13g2_xor2_1 _10640_ (.B(_04945_),
    .A(_04944_),
    .X(_04959_));
 sg13g2_a21o_1 _10641_ (.A2(_04959_),
    .A1(_04958_),
    .B1(_04946_),
    .X(_04960_));
 sg13g2_xor2_1 _10642_ (.B(_04937_),
    .A(_04936_),
    .X(_04961_));
 sg13g2_a21o_1 _10643_ (.A2(_04961_),
    .A1(_04960_),
    .B1(_04938_),
    .X(_04962_));
 sg13g2_a21o_1 _10644_ (.A2(_04962_),
    .A1(_04931_),
    .B1(_04930_),
    .X(_04963_));
 sg13g2_xnor2_1 _10645_ (.Y(_04964_),
    .A(_04921_),
    .B(_04922_));
 sg13g2_a21o_1 _10646_ (.A2(_04964_),
    .A1(_04963_),
    .B1(_04923_),
    .X(_04965_));
 sg13g2_a21o_1 _10647_ (.A2(_04965_),
    .A1(_04918_),
    .B1(_04916_),
    .X(_04966_));
 sg13g2_xnor2_1 _10648_ (.Y(_04967_),
    .A(_04892_),
    .B(_04909_));
 sg13g2_inv_1 _10649_ (.Y(_04968_),
    .A(_04967_));
 sg13g2_a21o_2 _10650_ (.A2(_04968_),
    .A1(_04966_),
    .B1(_04910_),
    .X(_04969_));
 sg13g2_xor2_1 _10651_ (.B(_04969_),
    .A(_04856_),
    .X(_04970_));
 sg13g2_xnor2_1 _10652_ (.Y(_04971_),
    .A(_04918_),
    .B(_04965_));
 sg13g2_xor2_1 _10653_ (.B(_04962_),
    .A(_04931_),
    .X(_04972_));
 sg13g2_xnor2_1 _10654_ (.Y(_04973_),
    .A(_04960_),
    .B(_04961_));
 sg13g2_xor2_1 _10655_ (.B(_04959_),
    .A(_04958_),
    .X(_04974_));
 sg13g2_xnor2_1 _10656_ (.Y(_04975_),
    .A(_04956_),
    .B(_04957_));
 sg13g2_nand2_1 _10657_ (.Y(_04976_),
    .A(_04932_),
    .B(_04935_));
 sg13g2_nor2_1 _10658_ (.A(_04863_),
    .B(_04949_),
    .Y(_04977_));
 sg13g2_o21ai_1 _10659_ (.B1(_04863_),
    .Y(_04978_),
    .A1(net1741),
    .A2(_04867_));
 sg13g2_nand2_1 _10660_ (.Y(_04979_),
    .A(_04859_),
    .B(_04978_));
 sg13g2_o21ai_1 _10661_ (.B1(_04976_),
    .Y(_04980_),
    .A1(_04977_),
    .A2(_04979_));
 sg13g2_inv_1 _10662_ (.Y(_04981_),
    .A(_04980_));
 sg13g2_xor2_1 _10663_ (.B(_04955_),
    .A(_04893_),
    .X(_04982_));
 sg13g2_nor2_1 _10664_ (.A(_04980_),
    .B(_04982_),
    .Y(_04983_));
 sg13g2_nand2_1 _10665_ (.Y(_04984_),
    .A(_04975_),
    .B(_04983_));
 sg13g2_nor2_1 _10666_ (.A(_04974_),
    .B(_04984_),
    .Y(_04985_));
 sg13g2_nand2_1 _10667_ (.Y(_04986_),
    .A(_04973_),
    .B(_04985_));
 sg13g2_nor2_1 _10668_ (.A(_04972_),
    .B(_04986_),
    .Y(_04987_));
 sg13g2_xnor2_1 _10669_ (.Y(_04988_),
    .A(_04963_),
    .B(_04964_));
 sg13g2_nand2_1 _10670_ (.Y(_04989_),
    .A(_04987_),
    .B(_04988_));
 sg13g2_nand2b_1 _10671_ (.Y(_04990_),
    .B(_04971_),
    .A_N(_04989_));
 sg13g2_xnor2_1 _10672_ (.Y(_04991_),
    .A(_04966_),
    .B(_04968_));
 sg13g2_nand2b_1 _10673_ (.Y(_04992_),
    .B(_04991_),
    .A_N(_04990_));
 sg13g2_nor2_1 _10674_ (.A(_04970_),
    .B(_04992_),
    .Y(_04993_));
 sg13g2_nor2_1 _10675_ (.A(net1533),
    .B(_04993_),
    .Y(_04994_));
 sg13g2_nand2_1 _10676_ (.Y(_04995_),
    .A(_04808_),
    .B(net1505));
 sg13g2_a21oi_2 _10677_ (.B1(_04855_),
    .Y(_04996_),
    .A2(_04969_),
    .A1(_04856_));
 sg13g2_nor2_1 _10678_ (.A(_04862_),
    .B(_04941_),
    .Y(_04997_));
 sg13g2_nor2_1 _10679_ (.A(_04925_),
    .B(_04934_),
    .Y(_04998_));
 sg13g2_a21oi_1 _10680_ (.A1(_04924_),
    .A2(_04998_),
    .Y(_04999_),
    .B1(_04997_));
 sg13g2_o21ai_1 _10681_ (.B1(_04867_),
    .Y(_05000_),
    .A1(net1742),
    .A2(_04871_));
 sg13g2_nand2_1 _10682_ (.Y(_05001_),
    .A(_04862_),
    .B(_05000_));
 sg13g2_a21oi_1 _10683_ (.A1(_04857_),
    .A2(_05001_),
    .Y(_05002_),
    .B1(_04853_));
 sg13g2_o21ai_1 _10684_ (.B1(_05002_),
    .Y(_05003_),
    .A1(_04876_),
    .A2(_04999_));
 sg13g2_inv_2 _10685_ (.Y(_05004_),
    .A(_05003_));
 sg13g2_o21ai_1 _10686_ (.B1(_04996_),
    .Y(_05005_),
    .A1(_04989_),
    .A2(_05004_));
 sg13g2_xor2_1 _10687_ (.B(_05005_),
    .A(_04971_),
    .X(_05006_));
 sg13g2_inv_2 _10688_ (.Y(_05007_),
    .A(_05006_));
 sg13g2_a221oi_1 _10689_ (.B2(_05003_),
    .C1(_04855_),
    .B1(_04987_),
    .A1(_04856_),
    .Y(_05008_),
    .A2(_04969_));
 sg13g2_xnor2_1 _10690_ (.Y(_05009_),
    .A(_04988_),
    .B(_05008_));
 sg13g2_nand2_1 _10691_ (.Y(_05010_),
    .A(_05007_),
    .B(net1453));
 sg13g2_a221oi_1 _10692_ (.B2(_05003_),
    .C1(_04855_),
    .B1(_04985_),
    .A1(_04856_),
    .Y(_05011_),
    .A2(_04969_));
 sg13g2_xor2_1 _10693_ (.B(_05011_),
    .A(_04973_),
    .X(_05012_));
 sg13g2_xnor2_1 _10694_ (.Y(_05013_),
    .A(_04973_),
    .B(_05011_));
 sg13g2_nand2_1 _10695_ (.Y(_05014_),
    .A(_04996_),
    .B(_05004_));
 sg13g2_xnor2_1 _10696_ (.Y(_05015_),
    .A(_04981_),
    .B(_05014_));
 sg13g2_nand3_1 _10697_ (.B(_04983_),
    .C(_05003_),
    .A(_04975_),
    .Y(_05016_));
 sg13g2_and2_1 _10698_ (.A(_04996_),
    .B(_05016_),
    .X(_05017_));
 sg13g2_xnor2_1 _10699_ (.Y(_05018_),
    .A(_04974_),
    .B(_05017_));
 sg13g2_xor2_1 _10700_ (.B(_05017_),
    .A(_04974_),
    .X(_05019_));
 sg13g2_o21ai_1 _10701_ (.B1(_05012_),
    .Y(_05020_),
    .A1(_05015_),
    .A2(_05019_));
 sg13g2_o21ai_1 _10702_ (.B1(_04996_),
    .Y(_05021_),
    .A1(_04986_),
    .A2(_05004_));
 sg13g2_xor2_1 _10703_ (.B(_05021_),
    .A(_04972_),
    .X(_05022_));
 sg13g2_a221oi_1 _10704_ (.B2(_05003_),
    .C1(_04855_),
    .B1(_04981_),
    .A1(_04856_),
    .Y(_05023_),
    .A2(_04969_));
 sg13g2_xnor2_1 _10705_ (.Y(_05024_),
    .A(_04982_),
    .B(_05023_));
 sg13g2_nor2_1 _10706_ (.A(_05013_),
    .B(_05024_),
    .Y(_05025_));
 sg13g2_nor2b_1 _10707_ (.A(_05025_),
    .B_N(net1440),
    .Y(_05026_));
 sg13g2_nand2b_1 _10708_ (.Y(_05027_),
    .B(net1441),
    .A_N(_05025_));
 sg13g2_a221oi_1 _10709_ (.B2(_05003_),
    .C1(_04855_),
    .B1(_04983_),
    .A1(_04856_),
    .Y(_05028_),
    .A2(_04969_));
 sg13g2_xnor2_1 _10710_ (.Y(_05029_),
    .A(_04975_),
    .B(_05028_));
 sg13g2_and2_1 _10711_ (.A(net1441),
    .B(_05029_),
    .X(_05030_));
 sg13g2_a22oi_1 _10712_ (.Y(_05031_),
    .B1(_05030_),
    .B2(_05018_),
    .A2(_05026_),
    .A1(_05020_));
 sg13g2_a221oi_1 _10713_ (.B2(_05018_),
    .C1(net1454),
    .B1(_05030_),
    .A1(_05020_),
    .Y(_05032_),
    .A2(_05026_));
 sg13g2_nor2_2 _10714_ (.A(net1442),
    .B(_05032_),
    .Y(_05033_));
 sg13g2_nand2_1 _10715_ (.Y(_05034_),
    .A(_04995_),
    .B(_05033_));
 sg13g2_or2_2 _10716_ (.X(_05035_),
    .B(net1454),
    .A(_05006_));
 sg13g2_inv_1 _10717_ (.Y(_05036_),
    .A(_05035_));
 sg13g2_nand2_1 _10718_ (.Y(_05037_),
    .A(_05012_),
    .B(net1441));
 sg13g2_nand2_1 _10719_ (.Y(_05038_),
    .A(_05015_),
    .B(_05024_));
 sg13g2_nor2_1 _10720_ (.A(_05019_),
    .B(_05029_),
    .Y(_05039_));
 sg13g2_a21oi_1 _10721_ (.A1(_05038_),
    .A2(_05039_),
    .Y(_05040_),
    .B1(_05037_));
 sg13g2_o21ai_1 _10722_ (.B1(_04813_),
    .Y(_05041_),
    .A1(_05035_),
    .A2(_05040_));
 sg13g2_inv_1 _10723_ (.Y(_05042_),
    .A(_05041_));
 sg13g2_nand2b_1 _10724_ (.Y(_05043_),
    .B(_05039_),
    .A_N(_05038_));
 sg13g2_nor2_1 _10725_ (.A(_05035_),
    .B(_05037_),
    .Y(_05044_));
 sg13g2_nand3_1 _10726_ (.B(_05043_),
    .C(_05044_),
    .A(_04845_),
    .Y(_05045_));
 sg13g2_nor2b_1 _10727_ (.A(_05041_),
    .B_N(_05045_),
    .Y(_05046_));
 sg13g2_a21o_1 _10728_ (.A2(_05044_),
    .A1(_05043_),
    .B1(_04845_),
    .X(_05047_));
 sg13g2_nand2_1 _10729_ (.Y(_05048_),
    .A(_04821_),
    .B(_05047_));
 sg13g2_a21oi_1 _10730_ (.A1(_05034_),
    .A2(_05046_),
    .Y(_05049_),
    .B1(_05048_));
 sg13g2_nor3_1 _10731_ (.A(net1505),
    .B(_05035_),
    .C(_05040_),
    .Y(_05050_));
 sg13g2_nand2b_1 _10732_ (.Y(_05051_),
    .B(_05050_),
    .A_N(_05031_));
 sg13g2_a221oi_1 _10733_ (.B2(_04820_),
    .C1(_05051_),
    .B1(_05045_),
    .A1(_04808_),
    .Y(_05052_),
    .A2(_05033_));
 sg13g2_o21ai_1 _10734_ (.B1(_04996_),
    .Y(_05053_),
    .A1(_04990_),
    .A2(_05004_));
 sg13g2_xor2_1 _10735_ (.B(_05053_),
    .A(_04991_),
    .X(_05054_));
 sg13g2_xnor2_1 _10736_ (.Y(_05055_),
    .A(_04991_),
    .B(_05053_));
 sg13g2_o21ai_1 _10737_ (.B1(_04996_),
    .Y(_05056_),
    .A1(_04992_),
    .A2(_05004_));
 sg13g2_xnor2_1 _10738_ (.Y(_05057_),
    .A(_04970_),
    .B(_05056_));
 sg13g2_xor2_1 _10739_ (.B(_05056_),
    .A(_04970_),
    .X(_05058_));
 sg13g2_nor2_1 _10740_ (.A(_04824_),
    .B(_04828_),
    .Y(_05059_));
 sg13g2_nand2_1 _10741_ (.Y(_05060_),
    .A(_04839_),
    .B(_05059_));
 sg13g2_inv_1 _10742_ (.Y(_05061_),
    .A(_05060_));
 sg13g2_nor4_1 _10743_ (.A(_04786_),
    .B(net1438),
    .C(net1437),
    .D(_05060_),
    .Y(_05062_));
 sg13g2_o21ai_1 _10744_ (.B1(_05062_),
    .Y(_05063_),
    .A1(_05049_),
    .A2(_05052_));
 sg13g2_and2_1 _10745_ (.A(_04994_),
    .B(_05063_),
    .X(_05064_));
 sg13g2_nor2_1 _10746_ (.A(_04825_),
    .B(_04839_),
    .Y(_05065_));
 sg13g2_nand4_1 _10747_ (.B(net1505),
    .C(_04828_),
    .A(_04807_),
    .Y(_05066_),
    .D(_04844_));
 sg13g2_nand3_1 _10748_ (.B(_04820_),
    .C(_05065_),
    .A(_04786_),
    .Y(_05067_));
 sg13g2_nor3_1 _10749_ (.A(net1435),
    .B(_05066_),
    .C(_05067_),
    .Y(_05068_));
 sg13g2_nor2b_2 _10750_ (.A(_05068_),
    .B_N(net1419),
    .Y(_05069_));
 sg13g2_nor2_1 _10751_ (.A(_05029_),
    .B(net1436),
    .Y(_05070_));
 sg13g2_nor2_1 _10752_ (.A(_05015_),
    .B(net1439),
    .Y(_05071_));
 sg13g2_o21ai_1 _10753_ (.B1(net1436),
    .Y(_05072_),
    .A1(_05024_),
    .A2(_05055_));
 sg13g2_a21oi_1 _10754_ (.A1(net1442),
    .A2(_05071_),
    .Y(_05073_),
    .B1(_05072_));
 sg13g2_nor2_1 _10755_ (.A(_05070_),
    .B(_05073_),
    .Y(_05074_));
 sg13g2_and3_1 _10756_ (.X(_05075_),
    .A(_00731_),
    .B(_04744_),
    .C(_04761_));
 sg13g2_nor2_1 _10757_ (.A(_04764_),
    .B(_05075_),
    .Y(_05076_));
 sg13g2_or2_1 _10758_ (.X(_05077_),
    .B(_05075_),
    .A(_04764_));
 sg13g2_a221oi_1 _10759_ (.B2(_05074_),
    .C1(net1516),
    .B1(_05069_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[0] ),
    .Y(_05078_),
    .A2(net1533));
 sg13g2_o21ai_1 _10760_ (.B1(net1535),
    .Y(_05079_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[0] ),
    .A2(_05076_));
 sg13g2_o21ai_1 _10761_ (.B1(_04769_),
    .Y(_05080_),
    .A1(_05078_),
    .A2(_05079_));
 sg13g2_nor2_2 _10762_ (.A(\u_tiny_nn_top.data_i_q[0] ),
    .B(net1744),
    .Y(_05081_));
 sg13g2_o21ai_1 _10763_ (.B1(_05080_),
    .Y(_05082_),
    .A1(net982),
    .A2(net1733));
 sg13g2_nor2_1 _10764_ (.A(_05081_),
    .B(_05082_),
    .Y(_00382_));
 sg13g2_nor2_1 _10765_ (.A(_05010_),
    .B(_05015_),
    .Y(_05083_));
 sg13g2_nor2_1 _10766_ (.A(_05007_),
    .B(_05024_),
    .Y(_05084_));
 sg13g2_o21ai_1 _10767_ (.B1(_05055_),
    .Y(_05085_),
    .A1(_05083_),
    .A2(_05084_));
 sg13g2_a21oi_1 _10768_ (.A1(_05029_),
    .A2(net1439),
    .Y(_05086_),
    .B1(_05057_));
 sg13g2_a22oi_1 _10769_ (.Y(_05087_),
    .B1(_05085_),
    .B2(_05086_),
    .A2(_05057_),
    .A1(_05018_));
 sg13g2_a221oi_1 _10770_ (.B2(_05087_),
    .C1(net1516),
    .B1(_05069_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[1] ),
    .Y(_05088_),
    .A2(net1533));
 sg13g2_o21ai_1 _10771_ (.B1(net1535),
    .Y(_05089_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[1] ),
    .A2(net1517));
 sg13g2_o21ai_1 _10772_ (.B1(_04769_),
    .Y(_05090_),
    .A1(_05088_),
    .A2(_05089_));
 sg13g2_nor2_1 _10773_ (.A(net1851),
    .B(net1743),
    .Y(_05091_));
 sg13g2_o21ai_1 _10774_ (.B1(_05090_),
    .Y(_05092_),
    .A1(net975),
    .A2(net1733));
 sg13g2_nor2_1 _10775_ (.A(_05091_),
    .B(_05092_),
    .Y(_00383_));
 sg13g2_nand2_1 _10776_ (.Y(_05093_),
    .A(_05018_),
    .B(net1439));
 sg13g2_nor2_1 _10777_ (.A(_05015_),
    .B(_05035_),
    .Y(_05094_));
 sg13g2_nor3_1 _10778_ (.A(_05015_),
    .B(net1440),
    .C(_05035_),
    .Y(_05095_));
 sg13g2_a21oi_1 _10779_ (.A1(net1442),
    .A2(_05029_),
    .Y(_05096_),
    .B1(net1439));
 sg13g2_o21ai_1 _10780_ (.B1(_05096_),
    .Y(_05097_),
    .A1(_05010_),
    .A2(_05024_));
 sg13g2_o21ai_1 _10781_ (.B1(_05093_),
    .Y(_05098_),
    .A1(_05095_),
    .A2(_05097_));
 sg13g2_nand2_1 _10782_ (.Y(_05099_),
    .A(net1436),
    .B(_05098_));
 sg13g2_o21ai_1 _10783_ (.B1(_05099_),
    .Y(_05100_),
    .A1(_05013_),
    .A2(net1436));
 sg13g2_inv_1 _10784_ (.Y(_05101_),
    .A(_05100_));
 sg13g2_a221oi_1 _10785_ (.B2(_05101_),
    .C1(net1516),
    .B1(_05069_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[2] ),
    .Y(_05102_),
    .A2(net1533));
 sg13g2_o21ai_1 _10786_ (.B1(net1535),
    .Y(_05103_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[2] ),
    .A2(net1517));
 sg13g2_o21ai_1 _10787_ (.B1(_04769_),
    .Y(_05104_),
    .A1(_05102_),
    .A2(_05103_));
 sg13g2_nor2_2 _10788_ (.A(\u_tiny_nn_top.data_i_q[2] ),
    .B(net1744),
    .Y(_05105_));
 sg13g2_o21ai_1 _10789_ (.B1(_05104_),
    .Y(_05106_),
    .A1(net985),
    .A2(net1733));
 sg13g2_nor2_1 _10790_ (.A(_05105_),
    .B(_05106_),
    .Y(_00384_));
 sg13g2_a21o_1 _10791_ (.A2(_05094_),
    .A1(net1440),
    .B1(net1439),
    .X(_05107_));
 sg13g2_nor2_1 _10792_ (.A(net1454),
    .B(_05024_),
    .Y(_05108_));
 sg13g2_nor3_1 _10793_ (.A(net1440),
    .B(_05024_),
    .C(_05035_),
    .Y(_05109_));
 sg13g2_nand3_1 _10794_ (.B(net1453),
    .C(_05029_),
    .A(_05007_),
    .Y(_05110_));
 sg13g2_o21ai_1 _10795_ (.B1(_05110_),
    .Y(_05111_),
    .A1(_05007_),
    .A2(_05018_));
 sg13g2_o21ai_1 _10796_ (.B1(_05055_),
    .Y(_05112_),
    .A1(_05109_),
    .A2(_05111_));
 sg13g2_a21oi_1 _10797_ (.A1(_05013_),
    .A2(_05107_),
    .Y(_05113_),
    .B1(_05057_));
 sg13g2_a22oi_1 _10798_ (.Y(_05114_),
    .B1(_05112_),
    .B2(_05113_),
    .A2(net1437),
    .A1(net1440));
 sg13g2_a221oi_1 _10799_ (.B2(_05114_),
    .C1(net1516),
    .B1(_05069_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[3] ),
    .Y(_05115_),
    .A2(net1533));
 sg13g2_o21ai_1 _10800_ (.B1(net1535),
    .Y(_05116_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[3] ),
    .A2(net1517));
 sg13g2_o21ai_1 _10801_ (.B1(_04768_),
    .Y(_05117_),
    .A1(_05115_),
    .A2(_05116_));
 sg13g2_o21ai_1 _10802_ (.B1(net1733),
    .Y(_05118_),
    .A1(net1848),
    .A2(net1743));
 sg13g2_nor2b_1 _10803_ (.A(_05118_),
    .B_N(_05117_),
    .Y(_05119_));
 sg13g2_a21o_1 _10804_ (.A2(net1734),
    .A1(net941),
    .B1(_05119_),
    .X(_00385_));
 sg13g2_nor2_1 _10805_ (.A(net1454),
    .B(net1436),
    .Y(_05120_));
 sg13g2_nor2_1 _10806_ (.A(_05015_),
    .B(_05037_),
    .Y(_05121_));
 sg13g2_nor2_1 _10807_ (.A(net1442),
    .B(_05018_),
    .Y(_05122_));
 sg13g2_o21ai_1 _10808_ (.B1(_05122_),
    .Y(_05123_),
    .A1(net1453),
    .A2(_05121_));
 sg13g2_a21oi_1 _10809_ (.A1(net1441),
    .A2(_05108_),
    .Y(_05124_),
    .B1(net1442));
 sg13g2_o21ai_1 _10810_ (.B1(_05123_),
    .Y(_05125_),
    .A1(_05012_),
    .A2(_05124_));
 sg13g2_a21oi_1 _10811_ (.A1(_05029_),
    .A2(_05036_),
    .Y(_05126_),
    .B1(net1438));
 sg13g2_o21ai_1 _10812_ (.B1(net1436),
    .Y(_05127_),
    .A1(net1440),
    .A2(_05126_));
 sg13g2_a21oi_1 _10813_ (.A1(_05055_),
    .A2(_05125_),
    .Y(_05128_),
    .B1(_05127_));
 sg13g2_nor2_1 _10814_ (.A(_05120_),
    .B(_05128_),
    .Y(_05129_));
 sg13g2_a221oi_1 _10815_ (.B2(_05129_),
    .C1(net1516),
    .B1(_05069_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[4] ),
    .Y(_05130_),
    .A2(net1533));
 sg13g2_o21ai_1 _10816_ (.B1(net1535),
    .Y(_05131_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[4] ),
    .A2(net1517));
 sg13g2_o21ai_1 _10817_ (.B1(_04768_),
    .Y(_05132_),
    .A1(_05130_),
    .A2(_05131_));
 sg13g2_o21ai_1 _10818_ (.B1(net1732),
    .Y(_05133_),
    .A1(net1845),
    .A2(net1743));
 sg13g2_nor2b_1 _10819_ (.A(_05133_),
    .B_N(_05132_),
    .Y(_05134_));
 sg13g2_a21o_1 _10820_ (.A2(net1734),
    .A1(net953),
    .B1(_05134_),
    .X(_00386_));
 sg13g2_nand3_1 _10821_ (.B(net1453),
    .C(_05012_),
    .A(_05007_),
    .Y(_05135_));
 sg13g2_a21oi_1 _10822_ (.A1(net1442),
    .A2(net1440),
    .Y(_05136_),
    .B1(net1438));
 sg13g2_a221oi_1 _10823_ (.B2(_05136_),
    .C1(net1437),
    .B1(_05135_),
    .A1(net1453),
    .Y(_05137_),
    .A2(net1438));
 sg13g2_a221oi_1 _10824_ (.B2(_05020_),
    .C1(net1453),
    .B1(_05030_),
    .A1(_05019_),
    .Y(_05138_),
    .A2(_05027_));
 sg13g2_o21ai_1 _10825_ (.B1(_05007_),
    .Y(_05139_),
    .A1(net1437),
    .A2(_05138_));
 sg13g2_nor2b_1 _10826_ (.A(_05137_),
    .B_N(_05139_),
    .Y(_05140_));
 sg13g2_a221oi_1 _10827_ (.B2(_05140_),
    .C1(net1516),
    .B1(_05069_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[5] ),
    .Y(_05141_),
    .A2(net1533));
 sg13g2_o21ai_1 _10828_ (.B1(net1535),
    .Y(_05142_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[5] ),
    .A2(net1517));
 sg13g2_o21ai_1 _10829_ (.B1(_04768_),
    .Y(_05143_),
    .A1(_05141_),
    .A2(_05142_));
 sg13g2_o21ai_1 _10830_ (.B1(net1733),
    .Y(_05144_),
    .A1(net1842),
    .A2(net1743));
 sg13g2_nor2b_1 _10831_ (.A(_05144_),
    .B_N(_05143_),
    .Y(_05145_));
 sg13g2_a21o_1 _10832_ (.A2(net1734),
    .A1(net958),
    .B1(_05145_),
    .X(_00387_));
 sg13g2_o21ai_1 _10833_ (.B1(net1436),
    .Y(_05146_),
    .A1(_05007_),
    .A2(net1454));
 sg13g2_nand3b_1 _10834_ (.B(_05018_),
    .C(net1441),
    .Y(_05147_),
    .A_N(_05015_));
 sg13g2_nor3_1 _10835_ (.A(net1453),
    .B(_05013_),
    .C(_05030_),
    .Y(_05148_));
 sg13g2_a22oi_1 _10836_ (.Y(_05149_),
    .B1(_05147_),
    .B2(_05148_),
    .A2(net1440),
    .A1(net1453));
 sg13g2_nand2_1 _10837_ (.Y(_05150_),
    .A(_05018_),
    .B(_05026_));
 sg13g2_nand3_1 _10838_ (.B(_05149_),
    .C(_05150_),
    .A(_05055_),
    .Y(_05151_));
 sg13g2_nor2_1 _10839_ (.A(net1442),
    .B(net1437),
    .Y(_05152_));
 sg13g2_a22oi_1 _10840_ (.Y(_05153_),
    .B1(_05151_),
    .B2(_05152_),
    .A2(_05146_),
    .A1(_05055_));
 sg13g2_a221oi_1 _10841_ (.B2(_05153_),
    .C1(net1516),
    .B1(_05069_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[6] ),
    .Y(_05154_),
    .A2(net1534));
 sg13g2_o21ai_1 _10842_ (.B1(net1535),
    .Y(_05155_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[6] ),
    .A2(net1517));
 sg13g2_o21ai_1 _10843_ (.B1(_04768_),
    .Y(_05156_),
    .A1(_05154_),
    .A2(_05155_));
 sg13g2_o21ai_1 _10844_ (.B1(_04738_),
    .Y(_05157_),
    .A1(net1839),
    .A2(net1743));
 sg13g2_nor2b_1 _10845_ (.A(_05157_),
    .B_N(_05156_),
    .Y(_05158_));
 sg13g2_a21o_1 _10846_ (.A2(net1734),
    .A1(net1006),
    .B1(_05158_),
    .X(_00388_));
 sg13g2_nand2_1 _10847_ (.Y(_05159_),
    .A(net1062),
    .B(net1734));
 sg13g2_o21ai_1 _10848_ (.B1(net1435),
    .Y(_05160_),
    .A1(_05033_),
    .A2(net1438));
 sg13g2_xnor2_1 _10849_ (.Y(_05161_),
    .A(_04807_),
    .B(_05160_));
 sg13g2_a221oi_1 _10850_ (.B2(_05161_),
    .C1(net1516),
    .B1(net1419),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[7] ),
    .Y(_05162_),
    .A2(net1534));
 sg13g2_a21oi_1 _10851_ (.A1(_00749_),
    .A2(net1515),
    .Y(_05163_),
    .B1(_05162_));
 sg13g2_nand2_2 _10852_ (.Y(_05164_),
    .A(_04762_),
    .B(_04768_));
 sg13g2_nor2_1 _10853_ (.A(net1836),
    .B(net1745),
    .Y(_05165_));
 sg13g2_o21ai_1 _10854_ (.B1(net1732),
    .Y(_05166_),
    .A1(_05163_),
    .A2(_05164_));
 sg13g2_o21ai_1 _10855_ (.B1(_05159_),
    .Y(_00389_),
    .A1(_05165_),
    .A2(_05166_));
 sg13g2_nor2_1 _10856_ (.A(_04807_),
    .B(_05033_),
    .Y(_05167_));
 sg13g2_o21ai_1 _10857_ (.B1(_04808_),
    .Y(_05168_),
    .A1(net1442),
    .A2(_05032_));
 sg13g2_nor2_1 _10858_ (.A(_05042_),
    .B(_05050_),
    .Y(_05169_));
 sg13g2_xnor2_1 _10859_ (.Y(_05170_),
    .A(_04808_),
    .B(net1505));
 sg13g2_o21ai_1 _10860_ (.B1(_05055_),
    .Y(_05171_),
    .A1(_05167_),
    .A2(_05169_));
 sg13g2_a21o_1 _10861_ (.A2(_05169_),
    .A1(_05167_),
    .B1(_05171_),
    .X(_05172_));
 sg13g2_a21oi_1 _10862_ (.A1(net1505),
    .A2(net1438),
    .Y(_05173_),
    .B1(net1437));
 sg13g2_a22oi_1 _10863_ (.Y(_05174_),
    .B1(_05172_),
    .B2(_05173_),
    .A2(_05170_),
    .A1(net1437));
 sg13g2_a221oi_1 _10864_ (.B2(_05174_),
    .C1(net1513),
    .B1(net1419),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[8] ),
    .Y(_05175_),
    .A2(net1534));
 sg13g2_a21oi_1 _10865_ (.A1(_00748_),
    .A2(net1513),
    .Y(_05176_),
    .B1(_05175_));
 sg13g2_nor2_1 _10866_ (.A(net1832),
    .B(net1743),
    .Y(_05177_));
 sg13g2_o21ai_1 _10867_ (.B1(net1732),
    .Y(_05178_),
    .A1(_05164_),
    .A2(_05176_));
 sg13g2_nand2_1 _10868_ (.Y(_05179_),
    .A(net1066),
    .B(net1734));
 sg13g2_o21ai_1 _10869_ (.B1(_05179_),
    .Y(_00390_),
    .A1(_05177_),
    .A2(_05178_));
 sg13g2_nand2_1 _10870_ (.Y(_05180_),
    .A(net1045),
    .B(net1735));
 sg13g2_and2_1 _10871_ (.A(_05045_),
    .B(_05047_),
    .X(_05181_));
 sg13g2_o21ai_1 _10872_ (.B1(_05041_),
    .Y(_05182_),
    .A1(_05050_),
    .A2(_05168_));
 sg13g2_a21oi_1 _10873_ (.A1(_05181_),
    .A2(_05182_),
    .Y(_05183_),
    .B1(net1438));
 sg13g2_o21ai_1 _10874_ (.B1(_05183_),
    .Y(_05184_),
    .A1(_05181_),
    .A2(_05182_));
 sg13g2_a21oi_1 _10875_ (.A1(_04844_),
    .A2(net1438),
    .Y(_05185_),
    .B1(net1437));
 sg13g2_nand3_1 _10876_ (.B(net1505),
    .C(_04844_),
    .A(_04808_),
    .Y(_05186_));
 sg13g2_xnor2_1 _10877_ (.Y(_05187_),
    .A(_04844_),
    .B(_04995_));
 sg13g2_o21ai_1 _10878_ (.B1(net1419),
    .Y(_05188_),
    .A1(net1435),
    .A2(_05187_));
 sg13g2_a21o_1 _10879_ (.A2(_05185_),
    .A1(_05184_),
    .B1(_05188_),
    .X(_05189_));
 sg13g2_a21oi_1 _10880_ (.A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[9] ),
    .A2(net1534),
    .Y(_05190_),
    .B1(net1515));
 sg13g2_a22oi_1 _10881_ (.Y(_05191_),
    .B1(_05189_),
    .B2(_05190_),
    .A2(net1513),
    .A1(_00751_));
 sg13g2_nor2_2 _10882_ (.A(\u_tiny_nn_top.data_i_q[9] ),
    .B(net1744),
    .Y(_05192_));
 sg13g2_o21ai_1 _10883_ (.B1(net1732),
    .Y(_05193_),
    .A1(_05164_),
    .A2(_05191_));
 sg13g2_o21ai_1 _10884_ (.B1(_05180_),
    .Y(_00391_),
    .A1(_05192_),
    .A2(_05193_));
 sg13g2_nand2_1 _10885_ (.Y(_05194_),
    .A(net1785),
    .B(net1735));
 sg13g2_nand3_1 _10886_ (.B(net1435),
    .C(_05183_),
    .A(_05047_),
    .Y(_05195_));
 sg13g2_o21ai_1 _10887_ (.B1(_05195_),
    .Y(_05196_),
    .A1(net1435),
    .A2(_05186_));
 sg13g2_xnor2_1 _10888_ (.Y(_05197_),
    .A(_04821_),
    .B(_05196_));
 sg13g2_a221oi_1 _10889_ (.B2(_05197_),
    .C1(_05077_),
    .B1(_05064_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[10] ),
    .Y(_05198_),
    .A2(_04770_));
 sg13g2_a21oi_1 _10890_ (.A1(_00750_),
    .A2(net1513),
    .Y(_05199_),
    .B1(_05198_));
 sg13g2_nor2_2 _10891_ (.A(\u_tiny_nn_top.data_i_q[10] ),
    .B(net1744),
    .Y(_05200_));
 sg13g2_o21ai_1 _10892_ (.B1(net1733),
    .Y(_05201_),
    .A1(_05164_),
    .A2(_05199_));
 sg13g2_o21ai_1 _10893_ (.B1(_05194_),
    .Y(_00392_),
    .A1(_05200_),
    .A2(_05201_));
 sg13g2_nand2_1 _10894_ (.Y(_05202_),
    .A(net1028),
    .B(net1735));
 sg13g2_nor3_1 _10895_ (.A(_04821_),
    .B(net1435),
    .C(_05186_),
    .Y(_05203_));
 sg13g2_and4_1 _10896_ (.A(_04821_),
    .B(_05047_),
    .C(net1435),
    .D(_05183_),
    .X(_05204_));
 sg13g2_nor2_1 _10897_ (.A(_05203_),
    .B(_05204_),
    .Y(_05205_));
 sg13g2_xnor2_1 _10898_ (.Y(_05206_),
    .A(_04828_),
    .B(_05205_));
 sg13g2_a221oi_1 _10899_ (.B2(_05206_),
    .C1(net1514),
    .B1(net1419),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[11] ),
    .Y(_05207_),
    .A2(net1534));
 sg13g2_a21oi_1 _10900_ (.A1(_00753_),
    .A2(net1514),
    .Y(_05208_),
    .B1(_05207_));
 sg13g2_nor2_2 _10901_ (.A(\u_tiny_nn_top.data_i_q[11] ),
    .B(net1744),
    .Y(_05209_));
 sg13g2_o21ai_1 _10902_ (.B1(net1732),
    .Y(_05210_),
    .A1(_05164_),
    .A2(_05208_));
 sg13g2_o21ai_1 _10903_ (.B1(_05202_),
    .Y(_00393_),
    .A1(_05209_),
    .A2(_05210_));
 sg13g2_nand2_1 _10904_ (.Y(_05211_),
    .A(net1035),
    .B(net1735));
 sg13g2_nor4_2 _10905_ (.A(_04821_),
    .B(_04829_),
    .C(net1435),
    .Y(_05212_),
    .D(_05186_));
 sg13g2_a21oi_1 _10906_ (.A1(_04829_),
    .A2(_05204_),
    .Y(_05213_),
    .B1(_05212_));
 sg13g2_xnor2_1 _10907_ (.Y(_05214_),
    .A(_04824_),
    .B(_05213_));
 sg13g2_a221oi_1 _10908_ (.B2(_05214_),
    .C1(net1514),
    .B1(net1419),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[12] ),
    .Y(_05215_),
    .A2(net1534));
 sg13g2_a21oi_1 _10909_ (.A1(_00752_),
    .A2(net1513),
    .Y(_05216_),
    .B1(_05215_));
 sg13g2_nor2_2 _10910_ (.A(net1828),
    .B(net1744),
    .Y(_05217_));
 sg13g2_o21ai_1 _10911_ (.B1(net1732),
    .Y(_05218_),
    .A1(_05164_),
    .A2(_05216_));
 sg13g2_o21ai_1 _10912_ (.B1(_05211_),
    .Y(_00394_),
    .A1(_05217_),
    .A2(_05218_));
 sg13g2_a22oi_1 _10913_ (.Y(_05219_),
    .B1(_05212_),
    .B2(_04824_),
    .A2(_05204_),
    .A1(_05059_));
 sg13g2_xnor2_1 _10914_ (.Y(_05220_),
    .A(_04838_),
    .B(_05219_));
 sg13g2_a22oi_1 _10915_ (.Y(_05221_),
    .B1(net1419),
    .B2(_05220_),
    .A2(net1534),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[13] ));
 sg13g2_a21oi_1 _10916_ (.A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[13] ),
    .A2(net1513),
    .Y(_05222_),
    .B1(_05164_));
 sg13g2_o21ai_1 _10917_ (.B1(_05222_),
    .Y(_05223_),
    .A1(net1513),
    .A2(_05221_));
 sg13g2_nor2_2 _10918_ (.A(\u_tiny_nn_top.data_i_q[13] ),
    .B(net1744),
    .Y(_05224_));
 sg13g2_nor2_1 _10919_ (.A(net1735),
    .B(_05224_),
    .Y(_05225_));
 sg13g2_a22oi_1 _10920_ (.Y(_05226_),
    .B1(_05223_),
    .B2(_05225_),
    .A2(net1734),
    .A1(net1023));
 sg13g2_inv_1 _10921_ (.Y(_00395_),
    .A(_05226_));
 sg13g2_nand2_1 _10922_ (.Y(_05227_),
    .A(net1058),
    .B(net1735));
 sg13g2_a22oi_1 _10923_ (.Y(_05228_),
    .B1(_05212_),
    .B2(_05065_),
    .A2(_05204_),
    .A1(_05061_));
 sg13g2_xnor2_1 _10924_ (.Y(_05229_),
    .A(_04786_),
    .B(_05228_));
 sg13g2_a221oi_1 _10925_ (.B2(_05229_),
    .C1(net1514),
    .B1(net1419),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[14] ),
    .Y(_05230_),
    .A2(net1534));
 sg13g2_a21oi_1 _10926_ (.A1(_00754_),
    .A2(net1513),
    .Y(_05231_),
    .B1(_05230_));
 sg13g2_nor2_2 _10927_ (.A(net1827),
    .B(net1744),
    .Y(_05232_));
 sg13g2_o21ai_1 _10928_ (.B1(net1732),
    .Y(_05233_),
    .A1(_05164_),
    .A2(_05231_));
 sg13g2_o21ai_1 _10929_ (.B1(_05227_),
    .Y(_00396_),
    .A1(_05232_),
    .A2(_05233_));
 sg13g2_nand2_1 _10930_ (.Y(_05234_),
    .A(net1010),
    .B(net1734));
 sg13g2_nor2b_1 _10931_ (.A(net1533),
    .B_N(_04996_),
    .Y(_05235_));
 sg13g2_a22oi_1 _10932_ (.Y(_05236_),
    .B1(_05063_),
    .B2(_05235_),
    .A2(_04770_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[15] ));
 sg13g2_o21ai_1 _10933_ (.B1(net1535),
    .Y(_05237_),
    .A1(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[15] ),
    .A2(net1517));
 sg13g2_a21oi_1 _10934_ (.A1(net1517),
    .A2(_05236_),
    .Y(_05238_),
    .B1(_05237_));
 sg13g2_nor3_2 _10935_ (.A(_04760_),
    .B(_04766_),
    .C(_05238_),
    .Y(_05239_));
 sg13g2_o21ai_1 _10936_ (.B1(net1733),
    .Y(_05240_),
    .A1(net1826),
    .A2(net1743));
 sg13g2_o21ai_1 _10937_ (.B1(_05234_),
    .Y(_00397_),
    .A1(_05239_),
    .A2(_05240_));
 sg13g2_nand2_1 _10938_ (.Y(_05241_),
    .A(net670),
    .B(net1750));
 sg13g2_o21ai_1 _10939_ (.B1(_05241_),
    .Y(_00398_),
    .A1(net1769),
    .A2(net1750));
 sg13g2_mux2_1 _10940_ (.A0(net1850),
    .A1(net872),
    .S(net1750),
    .X(_00399_));
 sg13g2_nand2_1 _10941_ (.Y(_05242_),
    .A(net562),
    .B(net1751));
 sg13g2_o21ai_1 _10942_ (.B1(_05242_),
    .Y(_00400_),
    .A1(net1771),
    .A2(net1751));
 sg13g2_mux2_1 _10943_ (.A0(net1846),
    .A1(net899),
    .S(net1751),
    .X(_00401_));
 sg13g2_mux2_1 _10944_ (.A0(net1843),
    .A1(net900),
    .S(net1751),
    .X(_00402_));
 sg13g2_mux2_1 _10945_ (.A0(net1840),
    .A1(net944),
    .S(net1750),
    .X(_00403_));
 sg13g2_mux2_1 _10946_ (.A0(net1838),
    .A1(net845),
    .S(net1752),
    .X(_00404_));
 sg13g2_mux2_1 _10947_ (.A0(net1835),
    .A1(net914),
    .S(net1753),
    .X(_00405_));
 sg13g2_mux2_1 _10948_ (.A0(net1831),
    .A1(net950),
    .S(net1761),
    .X(_00406_));
 sg13g2_nand2_1 _10949_ (.Y(_05243_),
    .A(net747),
    .B(net1755));
 sg13g2_o21ai_1 _10950_ (.B1(_05243_),
    .Y(_00407_),
    .A1(net1773),
    .A2(net1755));
 sg13g2_nand2_1 _10951_ (.Y(_05244_),
    .A(net649),
    .B(net1753));
 sg13g2_o21ai_1 _10952_ (.B1(_05244_),
    .Y(_00408_),
    .A1(net1775),
    .A2(net1753));
 sg13g2_nand2_1 _10953_ (.Y(_05245_),
    .A(net483),
    .B(net1753));
 sg13g2_o21ai_1 _10954_ (.B1(_05245_),
    .Y(_00409_),
    .A1(net1777),
    .A2(net1753));
 sg13g2_nand2_1 _10955_ (.Y(_05246_),
    .A(net606),
    .B(net1753));
 sg13g2_o21ai_1 _10956_ (.B1(_05246_),
    .Y(_00410_),
    .A1(net1779),
    .A2(net1755));
 sg13g2_nand2_1 _10957_ (.Y(_05247_),
    .A(net777),
    .B(net1761));
 sg13g2_o21ai_1 _10958_ (.B1(_05247_),
    .Y(_00411_),
    .A1(net1782),
    .A2(net1761));
 sg13g2_nand2_1 _10959_ (.Y(_05248_),
    .A(net589),
    .B(net1761));
 sg13g2_o21ai_1 _10960_ (.B1(_05248_),
    .Y(_00412_),
    .A1(net1783),
    .A2(net1761));
 sg13g2_mux2_1 _10961_ (.A0(net1825),
    .A1(net938),
    .S(net1762),
    .X(_00413_));
 sg13g2_nor2_1 _10962_ (.A(net1794),
    .B(net695),
    .Y(_05249_));
 sg13g2_a21oi_1 _10963_ (.A1(net1769),
    .A2(net1794),
    .Y(_00414_),
    .B1(_05249_));
 sg13g2_mux2_1 _10964_ (.A0(net733),
    .A1(net1849),
    .S(net1794),
    .X(_00415_));
 sg13g2_nor2_1 _10965_ (.A(net1794),
    .B(net609),
    .Y(_05250_));
 sg13g2_a21oi_1 _10966_ (.A1(net1771),
    .A2(net1794),
    .Y(_00416_),
    .B1(_05250_));
 sg13g2_mux2_1 _10967_ (.A0(net535),
    .A1(net1847),
    .S(net1796),
    .X(_00417_));
 sg13g2_mux2_1 _10968_ (.A0(net536),
    .A1(net1844),
    .S(net1796),
    .X(_00418_));
 sg13g2_mux2_1 _10969_ (.A0(net537),
    .A1(net1841),
    .S(net1796),
    .X(_00419_));
 sg13g2_mux2_1 _10970_ (.A0(net735),
    .A1(net1837),
    .S(net1794),
    .X(_00420_));
 sg13g2_mux2_1 _10971_ (.A0(net708),
    .A1(net1833),
    .S(net1797),
    .X(_00421_));
 sg13g2_mux2_1 _10972_ (.A0(net699),
    .A1(net1830),
    .S(net1795),
    .X(_00422_));
 sg13g2_nor2_1 _10973_ (.A(net1795),
    .B(net616),
    .Y(_05251_));
 sg13g2_a21oi_1 _10974_ (.A1(net1774),
    .A2(net1795),
    .Y(_00423_),
    .B1(_05251_));
 sg13g2_nor2_1 _10975_ (.A(net1796),
    .B(net628),
    .Y(_05252_));
 sg13g2_a21oi_1 _10976_ (.A1(net1776),
    .A2(net1795),
    .Y(_00424_),
    .B1(_05252_));
 sg13g2_nor2_1 _10977_ (.A(net1795),
    .B(net683),
    .Y(_05253_));
 sg13g2_a21oi_1 _10978_ (.A1(net1777),
    .A2(net1795),
    .Y(_00425_),
    .B1(_05253_));
 sg13g2_nor2_1 _10979_ (.A(net1794),
    .B(net577),
    .Y(_05254_));
 sg13g2_a21oi_1 _10980_ (.A1(net1779),
    .A2(net1794),
    .Y(_00426_),
    .B1(_05254_));
 sg13g2_nor2_1 _10981_ (.A(net1795),
    .B(net605),
    .Y(_05255_));
 sg13g2_a21oi_1 _10982_ (.A1(net1782),
    .A2(net1795),
    .Y(_00427_),
    .B1(_05255_));
 sg13g2_nor2_1 _10983_ (.A(net1797),
    .B(net671),
    .Y(_05256_));
 sg13g2_a21oi_1 _10984_ (.A1(net1783),
    .A2(net1797),
    .Y(_00428_),
    .B1(net672));
 sg13g2_mux2_1 _10985_ (.A0(net764),
    .A1(net1823),
    .S(net1797),
    .X(_00429_));
 sg13g2_mux2_1 _10986_ (.A0(net670),
    .A1(net854),
    .S(net1750),
    .X(_00430_));
 sg13g2_mux2_1 _10987_ (.A0(net872),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][1] ),
    .S(net1751),
    .X(_00431_));
 sg13g2_mux2_1 _10988_ (.A0(net562),
    .A1(net824),
    .S(net1751),
    .X(_00432_));
 sg13g2_mux2_1 _10989_ (.A0(net899),
    .A1(net861),
    .S(net1751),
    .X(_00433_));
 sg13g2_mux2_1 _10990_ (.A0(net900),
    .A1(net866),
    .S(net1756),
    .X(_00434_));
 sg13g2_mux2_1 _10991_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[7][5] ),
    .A1(net925),
    .S(net1750),
    .X(_00435_));
 sg13g2_mux2_1 _10992_ (.A0(net845),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][6] ),
    .S(net1752),
    .X(_00436_));
 sg13g2_mux2_1 _10993_ (.A0(net914),
    .A1(net948),
    .S(net1754),
    .X(_00437_));
 sg13g2_mux2_1 _10994_ (.A0(net950),
    .A1(net951),
    .S(net1761),
    .X(_00438_));
 sg13g2_mux2_1 _10995_ (.A0(net747),
    .A1(net911),
    .S(net1754),
    .X(_00439_));
 sg13g2_mux2_1 _10996_ (.A0(net649),
    .A1(net881),
    .S(net1754),
    .X(_00440_));
 sg13g2_mux2_1 _10997_ (.A0(net483),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[5][11] ),
    .S(net1753),
    .X(_00441_));
 sg13g2_mux2_1 _10998_ (.A0(net606),
    .A1(net879),
    .S(net1753),
    .X(_00442_));
 sg13g2_mux2_1 _10999_ (.A0(net777),
    .A1(net920),
    .S(net1754),
    .X(_00443_));
 sg13g2_mux2_1 _11000_ (.A0(net589),
    .A1(net842),
    .S(net1762),
    .X(_00444_));
 sg13g2_mux2_1 _11001_ (.A0(net938),
    .A1(net896),
    .S(net1759),
    .X(_00445_));
 sg13g2_nor2_1 _11002_ (.A(net684),
    .B(net1800),
    .Y(_05257_));
 sg13g2_a21oi_1 _11003_ (.A1(net1769),
    .A2(net1800),
    .Y(_00446_),
    .B1(_05257_));
 sg13g2_mux2_1 _11004_ (.A0(net712),
    .A1(net1850),
    .S(net1800),
    .X(_00447_));
 sg13g2_nor2_1 _11005_ (.A(net819),
    .B(net1800),
    .Y(_05258_));
 sg13g2_a21oi_1 _11006_ (.A1(net1771),
    .A2(net1800),
    .Y(_00448_),
    .B1(_05258_));
 sg13g2_mux2_1 _11007_ (.A0(net540),
    .A1(net1846),
    .S(net1799),
    .X(_00449_));
 sg13g2_mux2_1 _11008_ (.A0(net529),
    .A1(net1843),
    .S(net1800),
    .X(_00450_));
 sg13g2_mux2_1 _11009_ (.A0(net550),
    .A1(net1840),
    .S(net1799),
    .X(_00451_));
 sg13g2_mux2_1 _11010_ (.A0(net720),
    .A1(net1838),
    .S(net1800),
    .X(_00452_));
 sg13g2_mux2_1 _11011_ (.A0(net821),
    .A1(net1835),
    .S(net1801),
    .X(_00453_));
 sg13g2_mux2_1 _11012_ (.A0(net723),
    .A1(net1831),
    .S(net1801),
    .X(_00454_));
 sg13g2_nor2_1 _11013_ (.A(net679),
    .B(net1798),
    .Y(_05259_));
 sg13g2_a21oi_1 _11014_ (.A1(net1773),
    .A2(net1798),
    .Y(_00455_),
    .B1(_05259_));
 sg13g2_nor2_1 _11015_ (.A(net680),
    .B(net1798),
    .Y(_05260_));
 sg13g2_a21oi_1 _11016_ (.A1(net1775),
    .A2(net1799),
    .Y(_00456_),
    .B1(_05260_));
 sg13g2_nor2_1 _11017_ (.A(net790),
    .B(net1798),
    .Y(_05261_));
 sg13g2_a21oi_1 _11018_ (.A1(net1777),
    .A2(net1798),
    .Y(_00457_),
    .B1(_05261_));
 sg13g2_nor2_1 _11019_ (.A(net772),
    .B(net1799),
    .Y(_05262_));
 sg13g2_a21oi_1 _11020_ (.A1(net1779),
    .A2(net1799),
    .Y(_00458_),
    .B1(_05262_));
 sg13g2_nor2_1 _11021_ (.A(net714),
    .B(net1799),
    .Y(_05263_));
 sg13g2_a21oi_1 _11022_ (.A1(net1782),
    .A2(net1799),
    .Y(_00459_),
    .B1(_05263_));
 sg13g2_nor2_1 _11023_ (.A(net713),
    .B(net1798),
    .Y(_05264_));
 sg13g2_a21oi_1 _11024_ (.A1(net1783),
    .A2(net1798),
    .Y(_00460_),
    .B1(_05264_));
 sg13g2_mux2_1 _11025_ (.A0(net685),
    .A1(net1825),
    .S(net1798),
    .X(_00461_));
 sg13g2_nor2_2 _11026_ (.A(net854),
    .B(net1750),
    .Y(_05265_));
 sg13g2_a21oi_1 _11027_ (.A1(_00684_),
    .A2(net1757),
    .Y(_00462_),
    .B1(_05265_));
 sg13g2_mux2_1 _11028_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[5][1] ),
    .A1(net933),
    .S(net1752),
    .X(_00463_));
 sg13g2_mux2_1 _11029_ (.A0(net824),
    .A1(net940),
    .S(net1752),
    .X(_00464_));
 sg13g2_mux2_1 _11030_ (.A0(net861),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][3] ),
    .S(net1752),
    .X(_00465_));
 sg13g2_mux2_1 _11031_ (.A0(net866),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][4] ),
    .S(net1752),
    .X(_00466_));
 sg13g2_mux2_1 _11032_ (.A0(net925),
    .A1(net931),
    .S(net1750),
    .X(_00467_));
 sg13g2_mux2_1 _11033_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[5][6] ),
    .A1(net923),
    .S(net1757),
    .X(_00468_));
 sg13g2_mux2_1 _11034_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[5][7] ),
    .A1(net907),
    .S(net1758),
    .X(_00469_));
 sg13g2_mux2_1 _11035_ (.A0(net951),
    .A1(net967),
    .S(net1761),
    .X(_00470_));
 sg13g2_mux2_1 _11036_ (.A0(net911),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][9] ),
    .S(net1754),
    .X(_00471_));
 sg13g2_mux2_1 _11037_ (.A0(net881),
    .A1(net859),
    .S(net1758),
    .X(_00472_));
 sg13g2_mux2_1 _11038_ (.A0(net921),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][11] ),
    .S(net1754),
    .X(_00473_));
 sg13g2_mux2_1 _11039_ (.A0(net879),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[3][12] ),
    .S(net1754),
    .X(_00474_));
 sg13g2_mux2_1 _11040_ (.A0(net920),
    .A1(net677),
    .S(net1758),
    .X(_00475_));
 sg13g2_mux2_1 _11041_ (.A0(net842),
    .A1(net917),
    .S(net1762),
    .X(_00476_));
 sg13g2_mux2_1 _11042_ (.A0(net896),
    .A1(net847),
    .S(net1758),
    .X(_00477_));
 sg13g2_nor2_1 _11043_ (.A(net1806),
    .B(net659),
    .Y(_05266_));
 sg13g2_a21oi_1 _11044_ (.A1(net1770),
    .A2(net1806),
    .Y(_00478_),
    .B1(net660));
 sg13g2_mux2_1 _11045_ (.A0(net548),
    .A1(net1851),
    .S(net1806),
    .X(_00479_));
 sg13g2_nor2_1 _11046_ (.A(net1806),
    .B(net507),
    .Y(_05267_));
 sg13g2_a21oi_1 _11047_ (.A1(net1772),
    .A2(net1806),
    .Y(_00480_),
    .B1(net508));
 sg13g2_mux2_1 _11048_ (.A0(net731),
    .A1(net1848),
    .S(net1806),
    .X(_00481_));
 sg13g2_mux2_1 _11049_ (.A0(net541),
    .A1(\u_tiny_nn_top.data_i_q[4] ),
    .S(\u_tiny_nn_top.param_write_q[3] ),
    .X(_00482_));
 sg13g2_mux2_1 _11050_ (.A0(net527),
    .A1(net1842),
    .S(net1806),
    .X(_00483_));
 sg13g2_mux2_1 _11051_ (.A0(net689),
    .A1(net1839),
    .S(net1806),
    .X(_00484_));
 sg13g2_mux2_1 _11052_ (.A0(net697),
    .A1(net1836),
    .S(net1807),
    .X(_00485_));
 sg13g2_mux2_1 _11053_ (.A0(net702),
    .A1(net1832),
    .S(net1808),
    .X(_00486_));
 sg13g2_nor2_1 _11054_ (.A(net1809),
    .B(net629),
    .Y(_05268_));
 sg13g2_a21oi_1 _11055_ (.A1(net1773),
    .A2(net1809),
    .Y(_00487_),
    .B1(net630));
 sg13g2_nor2_1 _11056_ (.A(net1807),
    .B(net722),
    .Y(_05269_));
 sg13g2_a21oi_1 _11057_ (.A1(net1775),
    .A2(net1807),
    .Y(_00488_),
    .B1(_05269_));
 sg13g2_nor2_1 _11058_ (.A(net1807),
    .B(net663),
    .Y(_05270_));
 sg13g2_a21oi_1 _11059_ (.A1(net1778),
    .A2(net1807),
    .Y(_00489_),
    .B1(_05270_));
 sg13g2_nor2_1 _11060_ (.A(net1807),
    .B(net667),
    .Y(_05271_));
 sg13g2_a21oi_1 _11061_ (.A1(net1780),
    .A2(net1807),
    .Y(_00490_),
    .B1(_05271_));
 sg13g2_nor2_1 _11062_ (.A(net1808),
    .B(net627),
    .Y(_05272_));
 sg13g2_a21oi_1 _11063_ (.A1(net1781),
    .A2(net1807),
    .Y(_00491_),
    .B1(_05272_));
 sg13g2_nor2_1 _11064_ (.A(net1808),
    .B(net700),
    .Y(_05273_));
 sg13g2_a21oi_1 _11065_ (.A1(net1784),
    .A2(net1808),
    .Y(_00492_),
    .B1(_05273_));
 sg13g2_mux2_1 _11066_ (.A0(net715),
    .A1(net1826),
    .S(net1808),
    .X(_00493_));
 sg13g2_nand2_1 _11067_ (.Y(_05274_),
    .A(net560),
    .B(net1757));
 sg13g2_o21ai_1 _11068_ (.B1(_05274_),
    .Y(_00494_),
    .A1(_00684_),
    .A2(net1757));
 sg13g2_mux2_1 _11069_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[3][1] ),
    .A1(net870),
    .S(net1760),
    .X(_00495_));
 sg13g2_mux2_1 _11070_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[3][2] ),
    .A1(net833),
    .S(net1757),
    .X(_00496_));
 sg13g2_mux2_1 _11071_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[3][3] ),
    .A1(net915),
    .S(net1752),
    .X(_00497_));
 sg13g2_mux2_1 _11072_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[3][4] ),
    .A1(net882),
    .S(net1757),
    .X(_00498_));
 sg13g2_mux2_1 _11073_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[3][5] ),
    .A1(net888),
    .S(net1752),
    .X(_00499_));
 sg13g2_mux2_1 _11074_ (.A0(net923),
    .A1(net927),
    .S(net1757),
    .X(_00500_));
 sg13g2_mux2_1 _11075_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[3][7] ),
    .A1(net837),
    .S(net1758),
    .X(_00501_));
 sg13g2_mux2_1 _11076_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[3][8] ),
    .A1(net817),
    .S(net1759),
    .X(_00502_));
 sg13g2_mux2_1 _11077_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[3][9] ),
    .A1(net897),
    .S(net1758),
    .X(_00503_));
 sg13g2_mux2_1 _11078_ (.A0(net859),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][10] ),
    .S(net1758),
    .X(_00504_));
 sg13g2_mux2_1 _11079_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[3][11] ),
    .A1(net825),
    .S(net1757),
    .X(_00505_));
 sg13g2_mux2_1 _11080_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[3][12] ),
    .A1(net850),
    .S(net1758),
    .X(_00506_));
 sg13g2_mux2_1 _11081_ (.A0(net677),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][13] ),
    .S(net1759),
    .X(_00507_));
 sg13g2_mux2_1 _11082_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[3][14] ),
    .A1(net894),
    .S(net1762),
    .X(_00508_));
 sg13g2_mux2_1 _11083_ (.A0(net847),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[1][15] ),
    .S(net1759),
    .X(_00509_));
 sg13g2_nor2_1 _11084_ (.A(net1814),
    .B(net658),
    .Y(_05275_));
 sg13g2_a21oi_1 _11085_ (.A1(net1769),
    .A2(net1814),
    .Y(_00510_),
    .B1(_05275_));
 sg13g2_mux2_1 _11086_ (.A0(net555),
    .A1(net1851),
    .S(net1814),
    .X(_00511_));
 sg13g2_nor2_1 _11087_ (.A(net1814),
    .B(net501),
    .Y(_05276_));
 sg13g2_a21oi_1 _11088_ (.A1(net1771),
    .A2(net1814),
    .Y(_00512_),
    .B1(_05276_));
 sg13g2_mux2_1 _11089_ (.A0(net692),
    .A1(net1848),
    .S(net1814),
    .X(_00513_));
 sg13g2_mux2_1 _11090_ (.A0(net539),
    .A1(net1845),
    .S(net1815),
    .X(_00514_));
 sg13g2_mux2_1 _11091_ (.A0(net814),
    .A1(net1842),
    .S(net1814),
    .X(_00515_));
 sg13g2_mux2_1 _11092_ (.A0(net681),
    .A1(net1839),
    .S(net1814),
    .X(_00516_));
 sg13g2_mux2_1 _11093_ (.A0(net856),
    .A1(net1836),
    .S(net1815),
    .X(_00517_));
 sg13g2_mux2_1 _11094_ (.A0(net710),
    .A1(net1832),
    .S(net1817),
    .X(_00518_));
 sg13g2_nor2_1 _11095_ (.A(net1817),
    .B(net634),
    .Y(_05277_));
 sg13g2_a21oi_1 _11096_ (.A1(net1773),
    .A2(net1817),
    .Y(_00519_),
    .B1(_05277_));
 sg13g2_nor2_1 _11097_ (.A(net1816),
    .B(net725),
    .Y(_05278_));
 sg13g2_a21oi_1 _11098_ (.A1(net1775),
    .A2(net1816),
    .Y(_00520_),
    .B1(net726));
 sg13g2_nor2_1 _11099_ (.A(net1815),
    .B(net612),
    .Y(_05279_));
 sg13g2_a21oi_1 _11100_ (.A1(net1778),
    .A2(net1815),
    .Y(_00521_),
    .B1(_05279_));
 sg13g2_nor2_1 _11101_ (.A(net1817),
    .B(net651),
    .Y(_05280_));
 sg13g2_a21oi_1 _11102_ (.A1(net1780),
    .A2(net1817),
    .Y(_00522_),
    .B1(_05280_));
 sg13g2_nor2_1 _11103_ (.A(net1817),
    .B(net666),
    .Y(_05281_));
 sg13g2_a21oi_1 _11104_ (.A1(net1781),
    .A2(net1817),
    .Y(_00523_),
    .B1(_05281_));
 sg13g2_nor2_1 _11105_ (.A(net1818),
    .B(net736),
    .Y(_05282_));
 sg13g2_a21oi_1 _11106_ (.A1(net1784),
    .A2(net1818),
    .Y(_00524_),
    .B1(net737));
 sg13g2_mux2_1 _11107_ (.A0(net755),
    .A1(net1826),
    .S(net1818),
    .X(_00525_));
 sg13g2_nor2b_1 _11108_ (.A(\u_tiny_nn_top.state_q[15] ),
    .B_N(net1854),
    .Y(_05283_));
 sg13g2_a221oi_1 _11109_ (.B2(net1765),
    .C1(_05283_),
    .B1(_02867_),
    .A1(_00163_),
    .Y(_05284_),
    .A2(_01063_));
 sg13g2_nor2_1 _11110_ (.A(net778),
    .B(net1676),
    .Y(_05285_));
 sg13g2_a21oi_1 _11111_ (.A1(net1769),
    .A2(net1676),
    .Y(_00526_),
    .B1(_05285_));
 sg13g2_mux2_1 _11112_ (.A0(net840),
    .A1(net1850),
    .S(net1676),
    .X(_00527_));
 sg13g2_nor2_1 _11113_ (.A(net858),
    .B(net1677),
    .Y(_05286_));
 sg13g2_a21oi_1 _11114_ (.A1(net1771),
    .A2(net1677),
    .Y(_00528_),
    .B1(_05286_));
 sg13g2_mux2_1 _11115_ (.A0(net803),
    .A1(net1846),
    .S(net1679),
    .X(_00529_));
 sg13g2_mux2_1 _11116_ (.A0(net780),
    .A1(net1843),
    .S(net1678),
    .X(_00530_));
 sg13g2_mux2_1 _11117_ (.A0(net810),
    .A1(net1840),
    .S(net1676),
    .X(_00531_));
 sg13g2_mux2_1 _11118_ (.A0(net797),
    .A1(net1838),
    .S(net1678),
    .X(_00532_));
 sg13g2_mux2_1 _11119_ (.A0(net781),
    .A1(net1835),
    .S(net1680),
    .X(_00533_));
 sg13g2_mux2_1 _11120_ (.A0(net693),
    .A1(net1831),
    .S(net1680),
    .X(_00534_));
 sg13g2_nor2_1 _11121_ (.A(net792),
    .B(net1680),
    .Y(_05287_));
 sg13g2_a21oi_1 _11122_ (.A1(net1773),
    .A2(net1680),
    .Y(_00535_),
    .B1(_05287_));
 sg13g2_nor2_1 _11123_ (.A(net804),
    .B(net1677),
    .Y(_05288_));
 sg13g2_a21oi_1 _11124_ (.A1(net1775),
    .A2(net1677),
    .Y(_00536_),
    .B1(_05288_));
 sg13g2_nor2_1 _11125_ (.A(net886),
    .B(net1677),
    .Y(_05289_));
 sg13g2_a21oi_1 _11126_ (.A1(net1777),
    .A2(net1679),
    .Y(_00537_),
    .B1(_05289_));
 sg13g2_nor2_1 _11127_ (.A(net762),
    .B(net1680),
    .Y(_05290_));
 sg13g2_a21oi_1 _11128_ (.A1(net1779),
    .A2(net1680),
    .Y(_00538_),
    .B1(_05290_));
 sg13g2_nor2_1 _11129_ (.A(net701),
    .B(net1686),
    .Y(_05291_));
 sg13g2_a21oi_1 _11130_ (.A1(net1781),
    .A2(net1686),
    .Y(_00539_),
    .B1(_05291_));
 sg13g2_nor2_1 _11131_ (.A(net495),
    .B(net1686),
    .Y(_05292_));
 sg13g2_a21oi_1 _11132_ (.A1(net1783),
    .A2(net1686),
    .Y(_00540_),
    .B1(_05292_));
 sg13g2_mux2_1 _11133_ (.A0(net816),
    .A1(net1825),
    .S(net1685),
    .X(_00541_));
 sg13g2_nor2_1 _11134_ (.A(net1862),
    .B(net504),
    .Y(_05293_));
 sg13g2_a21oi_1 _11135_ (.A1(net1769),
    .A2(net1862),
    .Y(_00542_),
    .B1(_05293_));
 sg13g2_mux2_1 _11136_ (.A0(net591),
    .A1(net1849),
    .S(net1862),
    .X(_00543_));
 sg13g2_nor2_1 _11137_ (.A(net1862),
    .B(net497),
    .Y(_05294_));
 sg13g2_a21oi_1 _11138_ (.A1(net1771),
    .A2(net1862),
    .Y(_00544_),
    .B1(_05294_));
 sg13g2_mux2_1 _11139_ (.A0(net565),
    .A1(net1847),
    .S(net1862),
    .X(_00545_));
 sg13g2_mux2_1 _11140_ (.A0(net519),
    .A1(net1843),
    .S(net1863),
    .X(_00546_));
 sg13g2_mux2_1 _11141_ (.A0(net563),
    .A1(net1840),
    .S(net1865),
    .X(_00547_));
 sg13g2_mux2_1 _11142_ (.A0(net574),
    .A1(net1837),
    .S(net1862),
    .X(_00548_));
 sg13g2_mux2_1 _11143_ (.A0(net662),
    .A1(net1833),
    .S(net1864),
    .X(_00549_));
 sg13g2_mux2_1 _11144_ (.A0(net583),
    .A1(net1830),
    .S(net1864),
    .X(_00550_));
 sg13g2_nor2_1 _11145_ (.A(net1863),
    .B(net498),
    .Y(_05295_));
 sg13g2_a21oi_1 _11146_ (.A1(net1774),
    .A2(net1865),
    .Y(_00551_),
    .B1(_05295_));
 sg13g2_nor2_1 _11147_ (.A(net1864),
    .B(net493),
    .Y(_05296_));
 sg13g2_a21oi_1 _11148_ (.A1(net1776),
    .A2(net1864),
    .Y(_00552_),
    .B1(_05296_));
 sg13g2_nor2_1 _11149_ (.A(net1863),
    .B(net520),
    .Y(_05297_));
 sg13g2_a21oi_1 _11150_ (.A1(net1777),
    .A2(net1863),
    .Y(_00553_),
    .B1(_05297_));
 sg13g2_nor2_1 _11151_ (.A(net1863),
    .B(net513),
    .Y(_05298_));
 sg13g2_a21oi_1 _11152_ (.A1(net1779),
    .A2(net1862),
    .Y(_00554_),
    .B1(_05298_));
 sg13g2_nor2_1 _11153_ (.A(net1863),
    .B(net646),
    .Y(_05299_));
 sg13g2_a21oi_1 _11154_ (.A1(net1782),
    .A2(net1863),
    .Y(_00555_),
    .B1(_05299_));
 sg13g2_nor2_1 _11155_ (.A(net1864),
    .B(net503),
    .Y(_05300_));
 sg13g2_a21oi_1 _11156_ (.A1(net1783),
    .A2(net1864),
    .Y(_00556_),
    .B1(_05300_));
 sg13g2_mux2_1 _11157_ (.A0(net635),
    .A1(net1823),
    .S(net1864),
    .X(_00557_));
 sg13g2_mux2_1 _11158_ (.A0(net909),
    .A1(net778),
    .S(net1676),
    .X(_00558_));
 sg13g2_mux2_1 _11159_ (.A0(net893),
    .A1(net840),
    .S(net1679),
    .X(_00559_));
 sg13g2_mux2_1 _11160_ (.A0(net929),
    .A1(net858),
    .S(net1677),
    .X(_00560_));
 sg13g2_mux2_1 _11161_ (.A0(net775),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[6][3] ),
    .S(net1678),
    .X(_00561_));
 sg13g2_mux2_1 _11162_ (.A0(net796),
    .A1(net780),
    .S(net1678),
    .X(_00562_));
 sg13g2_mux2_1 _11163_ (.A0(net782),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[6][5] ),
    .S(net1676),
    .X(_00563_));
 sg13g2_mux2_1 _11164_ (.A0(net801),
    .A1(net797),
    .S(net1683),
    .X(_00564_));
 sg13g2_mux2_1 _11165_ (.A0(net831),
    .A1(net781),
    .S(net1680),
    .X(_00565_));
 sg13g2_mux2_1 _11166_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][8] ),
    .A1(net693),
    .S(net1680),
    .X(_00566_));
 sg13g2_mux2_1 _11167_ (.A0(net753),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[6][9] ),
    .S(net1681),
    .X(_00567_));
 sg13g2_mux2_1 _11168_ (.A0(net757),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[6][10] ),
    .S(net1677),
    .X(_00568_));
 sg13g2_mux2_1 _11169_ (.A0(net843),
    .A1(net886),
    .S(net1677),
    .X(_00569_));
 sg13g2_mux2_1 _11170_ (.A0(net791),
    .A1(net762),
    .S(net1681),
    .X(_00570_));
 sg13g2_mux2_1 _11171_ (.A0(net789),
    .A1(net701),
    .S(net1685),
    .X(_00571_));
 sg13g2_mux2_1 _11172_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[4][14] ),
    .A1(net495),
    .S(net1685),
    .X(_00572_));
 sg13g2_mux2_1 _11173_ (.A0(net739),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[6][15] ),
    .S(net1687),
    .X(_00573_));
 sg13g2_nor2_1 _11174_ (.A(net1804),
    .B(net524),
    .Y(_05301_));
 sg13g2_a21oi_1 _11175_ (.A1(net1769),
    .A2(net1804),
    .Y(_00574_),
    .B1(net525));
 sg13g2_mux2_1 _11176_ (.A0(net717),
    .A1(net1850),
    .S(net1804),
    .X(_00575_));
 sg13g2_nor2_1 _11177_ (.A(net1804),
    .B(net728),
    .Y(_05302_));
 sg13g2_a21oi_1 _11178_ (.A1(net1771),
    .A2(net1804),
    .Y(_00576_),
    .B1(net729));
 sg13g2_mux2_1 _11179_ (.A0(net559),
    .A1(net1846),
    .S(net1803),
    .X(_00577_));
 sg13g2_mux2_1 _11180_ (.A0(net553),
    .A1(net1843),
    .S(net1804),
    .X(_00578_));
 sg13g2_mux2_1 _11181_ (.A0(net551),
    .A1(net1840),
    .S(net1804),
    .X(_00579_));
 sg13g2_mux2_1 _11182_ (.A0(net581),
    .A1(net1838),
    .S(net1804),
    .X(_00580_));
 sg13g2_mux2_1 _11183_ (.A0(net721),
    .A1(net1835),
    .S(net1802),
    .X(_00581_));
 sg13g2_mux2_1 _11184_ (.A0(net648),
    .A1(net1831),
    .S(net1802),
    .X(_00582_));
 sg13g2_nor2_1 _11185_ (.A(net1803),
    .B(net534),
    .Y(_05303_));
 sg13g2_a21oi_1 _11186_ (.A1(net1773),
    .A2(net1803),
    .Y(_00583_),
    .B1(_05303_));
 sg13g2_nor2_1 _11187_ (.A(net1802),
    .B(net568),
    .Y(_05304_));
 sg13g2_a21oi_1 _11188_ (.A1(net1775),
    .A2(net1805),
    .Y(_00584_),
    .B1(_05304_));
 sg13g2_nor2_1 _11189_ (.A(net1802),
    .B(net590),
    .Y(_05305_));
 sg13g2_a21oi_1 _11190_ (.A1(net1777),
    .A2(net1802),
    .Y(_00585_),
    .B1(_05305_));
 sg13g2_nor2_1 _11191_ (.A(net1803),
    .B(net502),
    .Y(_05306_));
 sg13g2_a21oi_1 _11192_ (.A1(net1779),
    .A2(net1803),
    .Y(_00586_),
    .B1(_05306_));
 sg13g2_nor2_1 _11193_ (.A(net1803),
    .B(net494),
    .Y(_05307_));
 sg13g2_a21oi_1 _11194_ (.A1(net1782),
    .A2(net1803),
    .Y(_00587_),
    .B1(_05307_));
 sg13g2_nor2_1 _11195_ (.A(net1805),
    .B(net586),
    .Y(_05308_));
 sg13g2_a21oi_1 _11196_ (.A1(net1783),
    .A2(net1805),
    .Y(_00588_),
    .B1(net587));
 sg13g2_mux2_1 _11197_ (.A0(net636),
    .A1(net1825),
    .S(net1802),
    .X(_00589_));
 sg13g2_nand2_2 _11198_ (.Y(_05309_),
    .A(net909),
    .B(net1676));
 sg13g2_o21ai_1 _11199_ (.B1(_05309_),
    .Y(_00590_),
    .A1(_00683_),
    .A2(net1682));
 sg13g2_mux2_1 _11200_ (.A0(net913),
    .A1(net893),
    .S(net1678),
    .X(_00591_));
 sg13g2_mux2_1 _11201_ (.A0(net748),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[4][2] ),
    .S(net1683),
    .X(_00592_));
 sg13g2_mux2_1 _11202_ (.A0(net793),
    .A1(net775),
    .S(net1678),
    .X(_00593_));
 sg13g2_mux2_1 _11203_ (.A0(net769),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[4][4] ),
    .S(net1682),
    .X(_00594_));
 sg13g2_mux2_1 _11204_ (.A0(net741),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[4][5] ),
    .S(net1676),
    .X(_00595_));
 sg13g2_mux2_1 _11205_ (.A0(net813),
    .A1(net801),
    .S(net1682),
    .X(_00596_));
 sg13g2_mux2_1 _11206_ (.A0(net751),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[4][7] ),
    .S(net1685),
    .X(_00597_));
 sg13g2_mux2_1 _11207_ (.A0(net863),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[4][8] ),
    .S(net1687),
    .X(_00598_));
 sg13g2_mux2_1 _11208_ (.A0(net743),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[4][9] ),
    .S(net1685),
    .X(_00599_));
 sg13g2_mux2_1 _11209_ (.A0(net812),
    .A1(net757),
    .S(net1683),
    .X(_00600_));
 sg13g2_mux2_1 _11210_ (.A0(\u_tiny_nn_top.u_core.mul_val_op_q[2][11] ),
    .A1(net843),
    .S(net1683),
    .X(_00601_));
 sg13g2_mux2_1 _11211_ (.A0(net745),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[4][12] ),
    .S(net1685),
    .X(_00602_));
 sg13g2_mux2_1 _11212_ (.A0(net849),
    .A1(net789),
    .S(net1687),
    .X(_00603_));
 sg13g2_mux2_1 _11213_ (.A0(net787),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[4][14] ),
    .S(net1688),
    .X(_00604_));
 sg13g2_mux2_1 _11214_ (.A0(net865),
    .A1(net739),
    .S(net1687),
    .X(_00605_));
 sg13g2_nor2_1 _11215_ (.A(net1810),
    .B(net545),
    .Y(_05310_));
 sg13g2_a21oi_1 _11216_ (.A1(net1770),
    .A2(net1810),
    .Y(_00606_),
    .B1(_05310_));
 sg13g2_mux2_1 _11217_ (.A0(net543),
    .A1(net1851),
    .S(net1810),
    .X(_00607_));
 sg13g2_nor2_1 _11218_ (.A(net1810),
    .B(net516),
    .Y(_05311_));
 sg13g2_a21oi_1 _11219_ (.A1(net1772),
    .A2(net1810),
    .Y(_00608_),
    .B1(_05311_));
 sg13g2_mux2_1 _11220_ (.A0(net584),
    .A1(net1848),
    .S(net1810),
    .X(_00609_));
 sg13g2_mux2_1 _11221_ (.A0(net523),
    .A1(net1845),
    .S(net1810),
    .X(_00610_));
 sg13g2_mux2_1 _11222_ (.A0(net546),
    .A1(\u_tiny_nn_top.data_i_q[5] ),
    .S(net1810),
    .X(_00611_));
 sg13g2_mux2_1 _11223_ (.A0(net621),
    .A1(net1839),
    .S(net1811),
    .X(_00612_));
 sg13g2_mux2_1 _11224_ (.A0(net637),
    .A1(net1836),
    .S(net1812),
    .X(_00613_));
 sg13g2_mux2_1 _11225_ (.A0(net623),
    .A1(net1832),
    .S(net1812),
    .X(_00614_));
 sg13g2_nor2_1 _11226_ (.A(net1813),
    .B(net596),
    .Y(_05312_));
 sg13g2_a21oi_1 _11227_ (.A1(net1773),
    .A2(net1813),
    .Y(_00615_),
    .B1(net597));
 sg13g2_nor2_1 _11228_ (.A(net1811),
    .B(net652),
    .Y(_05313_));
 sg13g2_a21oi_1 _11229_ (.A1(net1775),
    .A2(net1811),
    .Y(_00616_),
    .B1(net653));
 sg13g2_nor2_1 _11230_ (.A(net1812),
    .B(net522),
    .Y(_05314_));
 sg13g2_a21oi_1 _11231_ (.A1(net1778),
    .A2(net1812),
    .Y(_00617_),
    .B1(_05314_));
 sg13g2_nor2_1 _11232_ (.A(net1812),
    .B(net538),
    .Y(_05315_));
 sg13g2_a21oi_1 _11233_ (.A1(net1780),
    .A2(net1812),
    .Y(_00618_),
    .B1(_05315_));
 sg13g2_nor2_1 _11234_ (.A(net1813),
    .B(net505),
    .Y(_05316_));
 sg13g2_a21oi_1 _11235_ (.A1(net1781),
    .A2(net1812),
    .Y(_00619_),
    .B1(net506));
 sg13g2_nor2_1 _11236_ (.A(net1813),
    .B(net510),
    .Y(_05317_));
 sg13g2_a21oi_1 _11237_ (.A1(net1784),
    .A2(net1813),
    .Y(_00620_),
    .B1(net511));
 sg13g2_mux2_1 _11238_ (.A0(net575),
    .A1(net1826),
    .S(net1812),
    .X(_00621_));
 sg13g2_nor2_1 _11239_ (.A(net668),
    .B(net1684),
    .Y(_05318_));
 sg13g2_a21oi_1 _11240_ (.A1(_00683_),
    .A2(net1682),
    .Y(_00622_),
    .B1(_05318_));
 sg13g2_mux2_1 _11241_ (.A0(net642),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][1] ),
    .S(net1684),
    .X(_00623_));
 sg13g2_mux2_1 _11242_ (.A0(net625),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][2] ),
    .S(net1682),
    .X(_00624_));
 sg13g2_mux2_1 _11243_ (.A0(net592),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][3] ),
    .S(net1682),
    .X(_00625_));
 sg13g2_mux2_1 _11244_ (.A0(net706),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][4] ),
    .S(net1682),
    .X(_00626_));
 sg13g2_mux2_1 _11245_ (.A0(net557),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][5] ),
    .S(net1678),
    .X(_00627_));
 sg13g2_mux2_1 _11246_ (.A0(net572),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][6] ),
    .S(net1684),
    .X(_00628_));
 sg13g2_mux2_1 _11247_ (.A0(net570),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][7] ),
    .S(net1687),
    .X(_00629_));
 sg13g2_mux2_1 _11248_ (.A0(net632),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][8] ),
    .S(net1687),
    .X(_00630_));
 sg13g2_mux2_1 _11249_ (.A0(net618),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][9] ),
    .S(net1685),
    .X(_00631_));
 sg13g2_mux2_1 _11250_ (.A0(net607),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][10] ),
    .S(net1684),
    .X(_00632_));
 sg13g2_mux2_1 _11251_ (.A0(net686),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][11] ),
    .S(net1682),
    .X(_00633_));
 sg13g2_mux2_1 _11252_ (.A0(net566),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][12] ),
    .S(net1685),
    .X(_00634_));
 sg13g2_mux2_1 _11253_ (.A0(net579),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][13] ),
    .S(net1687),
    .X(_00635_));
 sg13g2_mux2_1 _11254_ (.A0(net644),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][14] ),
    .S(net1688),
    .X(_00636_));
 sg13g2_mux2_1 _11255_ (.A0(net614),
    .A1(\u_tiny_nn_top.u_core.mul_val_op_q[2][15] ),
    .S(net1687),
    .X(_00637_));
 sg13g2_dfrbp_1 _11256_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net68),
    .D(net904),
    .Q_N(_05626_),
    .Q(\u_tiny_nn_top.relu_q ));
 sg13g2_dfrbp_1 _11257_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net414),
    .D(_00189_),
    .Q_N(_05625_),
    .Q(\u_tiny_nn_top.param_write_q[6] ));
 sg13g2_dfrbp_1 _11258_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net413),
    .D(_00190_),
    .Q_N(_00100_),
    .Q(\u_tiny_nn_top.start_count_q[0] ));
 sg13g2_dfrbp_1 _11259_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net412),
    .D(net785),
    .Q_N(_00102_),
    .Q(\u_tiny_nn_top.start_count_q[1] ));
 sg13g2_dfrbp_1 _11260_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net411),
    .D(_00192_),
    .Q_N(_00104_),
    .Q(\u_tiny_nn_top.start_count_q[2] ));
 sg13g2_dfrbp_1 _11261_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net410),
    .D(net828),
    .Q_N(_00106_),
    .Q(\u_tiny_nn_top.start_count_q[3] ));
 sg13g2_dfrbp_1 _11262_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net409),
    .D(_00194_),
    .Q_N(_00108_),
    .Q(\u_tiny_nn_top.start_count_q[4] ));
 sg13g2_dfrbp_1 _11263_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net408),
    .D(_00195_),
    .Q_N(_00110_),
    .Q(\u_tiny_nn_top.start_count_q[5] ));
 sg13g2_dfrbp_1 _11264_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net407),
    .D(net800),
    .Q_N(_00112_),
    .Q(\u_tiny_nn_top.start_count_q[6] ));
 sg13g2_dfrbp_1 _11265_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net406),
    .D(net809),
    .Q_N(_00114_),
    .Q(\u_tiny_nn_top.start_count_q[7] ));
 sg13g2_dfrbp_1 _11266_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net405),
    .D(_00198_),
    .Q_N(_00099_),
    .Q(\u_tiny_nn_top.counter_q[0] ));
 sg13g2_dfrbp_1 _11267_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net404),
    .D(net1081),
    .Q_N(_05624_),
    .Q(\u_tiny_nn_top.counter_q[1] ));
 sg13g2_dfrbp_1 _11268_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net403),
    .D(_00200_),
    .Q_N(_00103_),
    .Q(\u_tiny_nn_top.counter_q[2] ));
 sg13g2_dfrbp_1 _11269_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net402),
    .D(net1032),
    .Q_N(_00105_),
    .Q(\u_tiny_nn_top.counter_q[3] ));
 sg13g2_dfrbp_1 _11270_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net401),
    .D(net1054),
    .Q_N(_00107_),
    .Q(\u_tiny_nn_top.counter_q[4] ));
 sg13g2_dfrbp_1 _11271_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net400),
    .D(net1025),
    .Q_N(_00109_),
    .Q(\u_tiny_nn_top.counter_q[5] ));
 sg13g2_dfrbp_1 _11272_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net399),
    .D(net1040),
    .Q_N(_00111_),
    .Q(\u_tiny_nn_top.counter_q[6] ));
 sg13g2_dfrbp_1 _11273_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net398),
    .D(net1009),
    .Q_N(_00113_),
    .Q(\u_tiny_nn_top.counter_q[7] ));
 sg13g2_dfrbp_1 _11274_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net397),
    .D(net492),
    .Q_N(_00169_),
    .Q(\u_tiny_nn_top.phase_q ));
 sg13g2_dfrbp_1 _11275_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net396),
    .D(net705),
    .Q_N(_05623_),
    .Q(\u_tiny_nn_top.max_val_skid_q[0] ));
 sg13g2_dfrbp_1 _11276_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net395),
    .D(net878),
    .Q_N(_05622_),
    .Q(\u_tiny_nn_top.max_val_skid_q[1] ));
 sg13g2_dfrbp_1 _11277_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net394),
    .D(net902),
    .Q_N(_05621_),
    .Q(\u_tiny_nn_top.max_val_skid_q[2] ));
 sg13g2_dfrbp_1 _11278_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net393),
    .D(net836),
    .Q_N(_05620_),
    .Q(\u_tiny_nn_top.max_val_skid_q[3] ));
 sg13g2_dfrbp_1 _11279_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net392),
    .D(net830),
    .Q_N(_05619_),
    .Q(\u_tiny_nn_top.max_val_skid_q[4] ));
 sg13g2_dfrbp_1 _11280_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net391),
    .D(net774),
    .Q_N(_05618_),
    .Q(\u_tiny_nn_top.max_val_skid_q[5] ));
 sg13g2_dfrbp_1 _11281_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net390),
    .D(net853),
    .Q_N(_05617_),
    .Q(\u_tiny_nn_top.max_val_skid_q[6] ));
 sg13g2_dfrbp_1 _11282_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net389),
    .D(net937),
    .Q_N(_05616_),
    .Q(\u_tiny_nn_top.max_val_skid_q[7] ));
 sg13g2_dfrbp_1 _11283_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1868),
    .D(_00179_),
    .Q_N(uo_out[0]),
    .Q(_00170_));
 sg13g2_dfrbp_1 _11284_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1866),
    .D(_00180_),
    .Q_N(uo_out[1]),
    .Q(_00171_));
 sg13g2_dfrbp_1 _11285_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1866),
    .D(_00181_),
    .Q_N(uo_out[2]),
    .Q(_00172_));
 sg13g2_dfrbp_1 _11286_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1866),
    .D(_00182_),
    .Q_N(uo_out[3]),
    .Q(_00173_));
 sg13g2_dfrbp_1 _11287_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1866),
    .D(_00183_),
    .Q_N(uo_out[4]),
    .Q(_00174_));
 sg13g2_dfrbp_1 _11288_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1866),
    .D(_00184_),
    .Q_N(uo_out[5]),
    .Q(_00175_));
 sg13g2_dfrbp_1 _11289_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1866),
    .D(_00185_),
    .Q_N(uo_out[6]),
    .Q(_00176_));
 sg13g2_dfrbp_1 _11290_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1866),
    .D(net919),
    .Q_N(uo_out[7]),
    .Q(_00177_));
 sg13g2_dfrbp_1 _11291_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1867),
    .D(net9),
    .Q_N(_05627_),
    .Q(\u_tiny_nn_top.data_i_q[0] ));
 sg13g2_dfrbp_1 _11292_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1867),
    .D(net10),
    .Q_N(_00101_),
    .Q(\u_tiny_nn_top.data_i_q[1] ));
 sg13g2_dfrbp_1 _11293_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1867),
    .D(net11),
    .Q_N(_05628_),
    .Q(\u_tiny_nn_top.data_i_q[2] ));
 sg13g2_dfrbp_1 _11294_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1867),
    .D(net12),
    .Q_N(_05629_),
    .Q(\u_tiny_nn_top.data_i_q[3] ));
 sg13g2_dfrbp_1 _11295_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1867),
    .D(net13),
    .Q_N(_05630_),
    .Q(\u_tiny_nn_top.data_i_q[4] ));
 sg13g2_dfrbp_1 _11296_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1867),
    .D(net14),
    .Q_N(_05631_),
    .Q(\u_tiny_nn_top.data_i_q[5] ));
 sg13g2_dfrbp_1 _11297_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1867),
    .D(net15),
    .Q_N(_00017_),
    .Q(\u_tiny_nn_top.data_i_q[6] ));
 sg13g2_dfrbp_1 _11298_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1866),
    .D(net16),
    .Q_N(_05632_),
    .Q(\u_tiny_nn_top.data_i_q[7] ));
 sg13g2_dfrbp_1 _11299_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1871),
    .D(net1),
    .Q_N(_05633_),
    .Q(\u_tiny_nn_top.data_i_q[8] ));
 sg13g2_dfrbp_1 _11300_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1871),
    .D(net2),
    .Q_N(_05634_),
    .Q(\u_tiny_nn_top.data_i_q[9] ));
 sg13g2_dfrbp_1 _11301_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1871),
    .D(net3),
    .Q_N(_05635_),
    .Q(\u_tiny_nn_top.data_i_q[10] ));
 sg13g2_dfrbp_1 _11302_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1871),
    .D(net4),
    .Q_N(_05636_),
    .Q(\u_tiny_nn_top.data_i_q[11] ));
 sg13g2_dfrbp_1 _11303_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1872),
    .D(net5),
    .Q_N(_05637_),
    .Q(\u_tiny_nn_top.data_i_q[12] ));
 sg13g2_dfrbp_1 _11304_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1872),
    .D(net6),
    .Q_N(_05638_),
    .Q(\u_tiny_nn_top.data_i_q[13] ));
 sg13g2_dfrbp_1 _11305_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1868),
    .D(net7),
    .Q_N(_05639_),
    .Q(\u_tiny_nn_top.data_i_q[14] ));
 sg13g2_dfrbp_1 _11306_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1867),
    .D(net8),
    .Q_N(_00168_),
    .Q(\u_tiny_nn_top.data_i_q[15] ));
 sg13g2_dfrbp_1 _11307_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net380),
    .D(_00215_),
    .Q_N(_00083_),
    .Q(\u_tiny_nn_top.core_accumulate_result[0] ));
 sg13g2_dfrbp_1 _11308_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net379),
    .D(_00216_),
    .Q_N(_00085_),
    .Q(\u_tiny_nn_top.core_accumulate_result[1] ));
 sg13g2_dfrbp_1 _11309_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net378),
    .D(_00217_),
    .Q_N(_00087_),
    .Q(\u_tiny_nn_top.core_accumulate_result[2] ));
 sg13g2_dfrbp_1 _11310_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net377),
    .D(_00218_),
    .Q_N(_00089_),
    .Q(\u_tiny_nn_top.core_accumulate_result[3] ));
 sg13g2_dfrbp_1 _11311_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net376),
    .D(_00219_),
    .Q_N(_00091_),
    .Q(\u_tiny_nn_top.core_accumulate_result[4] ));
 sg13g2_dfrbp_1 _11312_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net375),
    .D(_00220_),
    .Q_N(_00093_),
    .Q(\u_tiny_nn_top.core_accumulate_result[5] ));
 sg13g2_dfrbp_1 _11313_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net374),
    .D(_00221_),
    .Q_N(_00095_),
    .Q(\u_tiny_nn_top.core_accumulate_result[6] ));
 sg13g2_dfrbp_1 _11314_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net373),
    .D(_00222_),
    .Q_N(_00097_),
    .Q(\u_tiny_nn_top.core_accumulate_result[7] ));
 sg13g2_dfrbp_1 _11315_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net372),
    .D(_00223_),
    .Q_N(_00084_),
    .Q(\u_tiny_nn_top.core_accumulate_result[8] ));
 sg13g2_dfrbp_1 _11316_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net371),
    .D(_00224_),
    .Q_N(_00086_),
    .Q(\u_tiny_nn_top.core_accumulate_result[9] ));
 sg13g2_dfrbp_1 _11317_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net370),
    .D(_00225_),
    .Q_N(_00088_),
    .Q(\u_tiny_nn_top.core_accumulate_result[10] ));
 sg13g2_dfrbp_1 _11318_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net369),
    .D(_00226_),
    .Q_N(_00090_),
    .Q(\u_tiny_nn_top.core_accumulate_result[11] ));
 sg13g2_dfrbp_1 _11319_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net368),
    .D(_00227_),
    .Q_N(_00092_),
    .Q(\u_tiny_nn_top.core_accumulate_result[12] ));
 sg13g2_dfrbp_1 _11320_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net367),
    .D(_00228_),
    .Q_N(_00094_),
    .Q(\u_tiny_nn_top.core_accumulate_result[13] ));
 sg13g2_dfrbp_1 _11321_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net366),
    .D(_00229_),
    .Q_N(_00096_),
    .Q(\u_tiny_nn_top.core_accumulate_result[14] ));
 sg13g2_dfrbp_1 _11322_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net365),
    .D(_00230_),
    .Q_N(_00098_),
    .Q(\u_tiny_nn_top.core_accumulate_result[15] ));
 sg13g2_dfrbp_1 _11323_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net364),
    .D(net675),
    .Q_N(_05615_),
    .Q(\u_tiny_nn_top.param_write_q[0] ));
 sg13g2_dfrbp_1 _11324_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net362),
    .D(net1027),
    .Q_N(_05614_),
    .Q(\u_tiny_nn_top.param_write_q[1] ));
 sg13g2_dfrbp_1 _11325_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net360),
    .D(_00233_),
    .Q_N(_05613_),
    .Q(\u_tiny_nn_top.param_write_q[2] ));
 sg13g2_dfrbp_1 _11326_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net358),
    .D(net1092),
    .Q_N(_05612_),
    .Q(\u_tiny_nn_top.param_write_q[3] ));
 sg13g2_dfrbp_1 _11327_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net356),
    .D(_00235_),
    .Q_N(_05611_),
    .Q(\u_tiny_nn_top.param_write_q[4] ));
 sg13g2_dfrbp_1 _11328_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net354),
    .D(_00236_),
    .Q_N(_05610_),
    .Q(\u_tiny_nn_top.param_write_q[5] ));
 sg13g2_dfrbp_1 _11329_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net352),
    .D(net1060),
    .Q_N(_05609_),
    .Q(\u_tiny_nn_top.param_write_q[7] ));
 sg13g2_dfrbp_1 _11330_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net350),
    .D(_00238_),
    .Q_N(_05608_),
    .Q(\u_tiny_nn_top.max_val_q[0] ));
 sg13g2_dfrbp_1 _11331_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net348),
    .D(_00239_),
    .Q_N(_05607_),
    .Q(\u_tiny_nn_top.max_val_q[1] ));
 sg13g2_dfrbp_1 _11332_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net346),
    .D(_00240_),
    .Q_N(_05606_),
    .Q(\u_tiny_nn_top.max_val_q[2] ));
 sg13g2_dfrbp_1 _11333_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net344),
    .D(_00241_),
    .Q_N(_05605_),
    .Q(\u_tiny_nn_top.max_val_q[3] ));
 sg13g2_dfrbp_1 _11334_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net342),
    .D(_00242_),
    .Q_N(_05604_),
    .Q(\u_tiny_nn_top.max_val_q[4] ));
 sg13g2_dfrbp_1 _11335_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net340),
    .D(_00243_),
    .Q_N(_05603_),
    .Q(\u_tiny_nn_top.max_val_q[5] ));
 sg13g2_dfrbp_1 _11336_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net338),
    .D(_00244_),
    .Q_N(_05602_),
    .Q(\u_tiny_nn_top.max_val_q[6] ));
 sg13g2_dfrbp_1 _11337_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net336),
    .D(_00245_),
    .Q_N(_05601_),
    .Q(\u_tiny_nn_top.max_val_q[7] ));
 sg13g2_dfrbp_1 _11338_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net334),
    .D(_00246_),
    .Q_N(_05600_),
    .Q(\u_tiny_nn_top.max_val_q[8] ));
 sg13g2_dfrbp_1 _11339_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net332),
    .D(net955),
    .Q_N(_05599_),
    .Q(\u_tiny_nn_top.max_val_q[9] ));
 sg13g2_dfrbp_1 _11340_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net330),
    .D(_00248_),
    .Q_N(_05598_),
    .Q(\u_tiny_nn_top.max_val_q[10] ));
 sg13g2_dfrbp_1 _11341_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net328),
    .D(net996),
    .Q_N(_05597_),
    .Q(\u_tiny_nn_top.max_val_q[11] ));
 sg13g2_dfrbp_1 _11342_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net326),
    .D(net961),
    .Q_N(_05596_),
    .Q(\u_tiny_nn_top.max_val_q[12] ));
 sg13g2_dfrbp_1 _11343_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net324),
    .D(net974),
    .Q_N(_05595_),
    .Q(\u_tiny_nn_top.max_val_q[13] ));
 sg13g2_dfrbp_1 _11344_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net322),
    .D(_00252_),
    .Q_N(_05594_),
    .Q(\u_tiny_nn_top.max_val_q[14] ));
 sg13g2_dfrbp_1 _11345_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net320),
    .D(_00253_),
    .Q_N(_05593_),
    .Q(\u_tiny_nn_top.max_val_q[15] ));
 sg13g2_dfrbp_1 _11346_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1870),
    .D(net1004),
    .Q_N(\u_tiny_nn_top.state_q[0] ),
    .Q(_00178_));
 sg13g2_dfrbp_1 _11347_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1869),
    .D(net977),
    .Q_N(_05640_),
    .Q(\u_tiny_nn_top.state_q[1] ));
 sg13g2_dfrbp_1 _11348_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1869),
    .D(net1089),
    .Q_N(_05641_),
    .Q(\u_tiny_nn_top.state_q[2] ));
 sg13g2_dfrbp_1 _11349_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1869),
    .D(net990),
    .Q_N(_00036_),
    .Q(\u_tiny_nn_top.state_q[3] ));
 sg13g2_dfrbp_1 _11350_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1870),
    .D(net994),
    .Q_N(_00164_),
    .Q(\u_tiny_nn_top.state_q[4] ));
 sg13g2_dfrbp_1 _11351_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1870),
    .D(_00001_),
    .Q_N(_05642_),
    .Q(\u_tiny_nn_top.state_q[5] ));
 sg13g2_dfrbp_1 _11352_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1869),
    .D(_00014_),
    .Q_N(_05643_),
    .Q(\u_tiny_nn_top.state_q[6] ));
 sg13g2_dfrbp_1 _11353_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1870),
    .D(_00002_),
    .Q_N(_05644_),
    .Q(\u_tiny_nn_top.state_q[7] ));
 sg13g2_dfrbp_1 _11354_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1871),
    .D(net488),
    .Q_N(_00167_),
    .Q(\u_tiny_nn_top.state_q[8] ));
 sg13g2_dfrbp_1 _11355_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1870),
    .D(_00016_),
    .Q_N(_05645_),
    .Q(\u_tiny_nn_top.state_q[9] ));
 sg13g2_dfrbp_1 _11356_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1869),
    .D(net807),
    .Q_N(_00166_),
    .Q(\u_tiny_nn_top.state_q[10] ));
 sg13g2_dfrbp_1 _11357_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1869),
    .D(_00005_),
    .Q_N(_00161_),
    .Q(\u_tiny_nn_top.core_mul_add_op_b_en ));
 sg13g2_dfrbp_1 _11358_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1871),
    .D(_00006_),
    .Q_N(_05646_),
    .Q(\u_tiny_nn_top.state_q[12] ));
 sg13g2_dfrbp_1 _11359_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1871),
    .D(net486),
    .Q_N(_00165_),
    .Q(\u_tiny_nn_top.state_q[13] ));
 sg13g2_dfrbp_1 _11360_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1870),
    .D(net490),
    .Q_N(_05647_),
    .Q(\u_tiny_nn_top.state_q[14] ));
 sg13g2_dfrbp_1 _11361_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1869),
    .D(net885),
    .Q_N(_00163_),
    .Q(\u_tiny_nn_top.state_q[15] ));
 sg13g2_dfrbp_1 _11362_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1869),
    .D(_00003_),
    .Q_N(_05648_),
    .Q(\u_tiny_nn_top.state_q[16] ));
 sg13g2_dfrbp_1 _11363_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1871),
    .D(_00010_),
    .Q_N(_00162_),
    .Q(\u_tiny_nn_top.state_q[17] ));
 sg13g2_dfrbp_1 _11364_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net317),
    .D(_00254_),
    .Q_N(_05592_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][0] ));
 sg13g2_dfrbp_1 _11365_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net316),
    .D(net533),
    .Q_N(_00038_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][1] ));
 sg13g2_dfrbp_1 _11366_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net315),
    .D(_00256_),
    .Q_N(_00040_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][2] ));
 sg13g2_dfrbp_1 _11367_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net314),
    .D(net665),
    .Q_N(_05591_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][3] ));
 sg13g2_dfrbp_1 _11368_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net313),
    .D(_00258_),
    .Q_N(_00042_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][4] ));
 sg13g2_dfrbp_1 _11369_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net312),
    .D(_00259_),
    .Q_N(_05590_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][5] ));
 sg13g2_dfrbp_1 _11370_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net311),
    .D(net595),
    .Q_N(_05589_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][6] ));
 sg13g2_dfrbp_1 _11371_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net310),
    .D(net767),
    .Q_N(_05588_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][7] ));
 sg13g2_dfrbp_1 _11372_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net309),
    .D(net657),
    .Q_N(_05587_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][8] ));
 sg13g2_dfrbp_1 _11373_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net308),
    .D(_00263_),
    .Q_N(_05586_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][9] ));
 sg13g2_dfrbp_1 _11374_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net307),
    .D(_00264_),
    .Q_N(_05585_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][10] ));
 sg13g2_dfrbp_1 _11375_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net306),
    .D(_00265_),
    .Q_N(_05584_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][11] ));
 sg13g2_dfrbp_1 _11376_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net305),
    .D(_00266_),
    .Q_N(_05583_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][12] ));
 sg13g2_dfrbp_1 _11377_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net304),
    .D(_00267_),
    .Q_N(_05582_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][13] ));
 sg13g2_dfrbp_1 _11378_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net303),
    .D(net601),
    .Q_N(_05581_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][14] ));
 sg13g2_dfrbp_1 _11379_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net302),
    .D(net640),
    .Q_N(_05580_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[0][15] ));
 sg13g2_dfrbp_1 _11380_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net301),
    .D(_00270_),
    .Q_N(_00143_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][0] ));
 sg13g2_dfrbp_1 _11381_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net300),
    .D(_00271_),
    .Q_N(_00151_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][1] ));
 sg13g2_dfrbp_1 _11382_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net299),
    .D(_00272_),
    .Q_N(_00147_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][2] ));
 sg13g2_dfrbp_1 _11383_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net298),
    .D(_00273_),
    .Q_N(_00157_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][3] ));
 sg13g2_dfrbp_1 _11384_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net297),
    .D(_00274_),
    .Q_N(_00155_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][4] ));
 sg13g2_dfrbp_1 _11385_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net296),
    .D(_00275_),
    .Q_N(_00159_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][5] ));
 sg13g2_dfrbp_1 _11386_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net295),
    .D(_00276_),
    .Q_N(_00142_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][6] ));
 sg13g2_dfrbp_1 _11387_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net294),
    .D(_00277_),
    .Q_N(_00145_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][7] ));
 sg13g2_dfrbp_1 _11388_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net293),
    .D(_00278_),
    .Q_N(_00153_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][8] ));
 sg13g2_dfrbp_1 _11389_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net292),
    .D(_00279_),
    .Q_N(_05579_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][9] ));
 sg13g2_dfrbp_1 _11390_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net291),
    .D(_00280_),
    .Q_N(_05578_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][10] ));
 sg13g2_dfrbp_1 _11391_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net290),
    .D(_00281_),
    .Q_N(_05577_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][11] ));
 sg13g2_dfrbp_1 _11392_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net289),
    .D(_00282_),
    .Q_N(_05576_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][12] ));
 sg13g2_dfrbp_1 _11393_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net288),
    .D(_00283_),
    .Q_N(_05575_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][13] ));
 sg13g2_dfrbp_1 _11394_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net287),
    .D(_00284_),
    .Q_N(_05574_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][14] ));
 sg13g2_dfrbp_1 _11395_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net286),
    .D(_00285_),
    .Q_N(_00150_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][15] ));
 sg13g2_dfrbp_1 _11396_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net285),
    .D(_00286_),
    .Q_N(_00144_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][0] ));
 sg13g2_dfrbp_1 _11397_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net284),
    .D(_00287_),
    .Q_N(_00152_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][1] ));
 sg13g2_dfrbp_1 _11398_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net283),
    .D(_00288_),
    .Q_N(_00148_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][2] ));
 sg13g2_dfrbp_1 _11399_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net282),
    .D(_00289_),
    .Q_N(_00158_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][3] ));
 sg13g2_dfrbp_1 _11400_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net281),
    .D(_00290_),
    .Q_N(_00156_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][4] ));
 sg13g2_dfrbp_1 _11401_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net280),
    .D(_00291_),
    .Q_N(_00160_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][5] ));
 sg13g2_dfrbp_1 _11402_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net279),
    .D(_00292_),
    .Q_N(_00141_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][6] ));
 sg13g2_dfrbp_1 _11403_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net278),
    .D(_00293_),
    .Q_N(_00146_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][7] ));
 sg13g2_dfrbp_1 _11404_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net277),
    .D(_00294_),
    .Q_N(_00154_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][8] ));
 sg13g2_dfrbp_1 _11405_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net276),
    .D(_00295_),
    .Q_N(_05573_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][9] ));
 sg13g2_dfrbp_1 _11406_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net275),
    .D(_00296_),
    .Q_N(_05572_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][10] ));
 sg13g2_dfrbp_1 _11407_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net274),
    .D(_00297_),
    .Q_N(_05571_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][11] ));
 sg13g2_dfrbp_1 _11408_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net273),
    .D(_00298_),
    .Q_N(_05570_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][12] ));
 sg13g2_dfrbp_1 _11409_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net272),
    .D(_00299_),
    .Q_N(_05569_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][13] ));
 sg13g2_dfrbp_1 _11410_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net271),
    .D(_00300_),
    .Q_N(_05568_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][14] ));
 sg13g2_dfrbp_1 _11411_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net270),
    .D(_00301_),
    .Q_N(_00149_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][15] ));
 sg13g2_dfrbp_1 _11412_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net269),
    .D(_00302_),
    .Q_N(_00034_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][0] ));
 sg13g2_dfrbp_1 _11413_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net268),
    .D(_00303_),
    .Q_N(_00032_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][1] ));
 sg13g2_dfrbp_1 _11414_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net267),
    .D(_00304_),
    .Q_N(_00030_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][2] ));
 sg13g2_dfrbp_1 _11415_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net266),
    .D(_00305_),
    .Q_N(_00028_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][3] ));
 sg13g2_dfrbp_1 _11416_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net265),
    .D(_00306_),
    .Q_N(_00026_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][4] ));
 sg13g2_dfrbp_1 _11417_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net264),
    .D(_00307_),
    .Q_N(_00024_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][5] ));
 sg13g2_dfrbp_1 _11418_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net263),
    .D(_00308_),
    .Q_N(_00019_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][6] ));
 sg13g2_dfrbp_1 _11419_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net262),
    .D(_00309_),
    .Q_N(_00022_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][7] ));
 sg13g2_dfrbp_1 _11420_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net261),
    .D(_00310_),
    .Q_N(_00057_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][8] ));
 sg13g2_dfrbp_1 _11421_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net260),
    .D(_00311_),
    .Q_N(_00061_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][9] ));
 sg13g2_dfrbp_1 _11422_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net259),
    .D(_00312_),
    .Q_N(_00059_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][10] ));
 sg13g2_dfrbp_1 _11423_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net258),
    .D(_00313_),
    .Q_N(_00065_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][11] ));
 sg13g2_dfrbp_1 _11424_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net257),
    .D(_00314_),
    .Q_N(_00063_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][12] ));
 sg13g2_dfrbp_1 _11425_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net256),
    .D(_00315_),
    .Q_N(_00069_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][13] ));
 sg13g2_dfrbp_1 _11426_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net255),
    .D(_00316_),
    .Q_N(_00067_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][14] ));
 sg13g2_dfrbp_1 _11427_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net254),
    .D(_00317_),
    .Q_N(_00021_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][15] ));
 sg13g2_dfrbp_1 _11428_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net253),
    .D(_00318_),
    .Q_N(_05567_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][0] ));
 sg13g2_dfrbp_1 _11429_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net251),
    .D(_00319_),
    .Q_N(_05566_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][1] ));
 sg13g2_dfrbp_1 _11430_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net249),
    .D(_00320_),
    .Q_N(_05565_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][2] ));
 sg13g2_dfrbp_1 _11431_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net247),
    .D(_00321_),
    .Q_N(_05564_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][3] ));
 sg13g2_dfrbp_1 _11432_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net245),
    .D(_00322_),
    .Q_N(_05563_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][4] ));
 sg13g2_dfrbp_1 _11433_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net243),
    .D(_00323_),
    .Q_N(_05562_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][5] ));
 sg13g2_dfrbp_1 _11434_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net241),
    .D(_00324_),
    .Q_N(_05561_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][6] ));
 sg13g2_dfrbp_1 _11435_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net239),
    .D(_00325_),
    .Q_N(_05560_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][7] ));
 sg13g2_dfrbp_1 _11436_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net237),
    .D(_00326_),
    .Q_N(_00058_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][8] ));
 sg13g2_dfrbp_1 _11437_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net235),
    .D(_00327_),
    .Q_N(_00062_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][9] ));
 sg13g2_dfrbp_1 _11438_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net233),
    .D(_00328_),
    .Q_N(_00060_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][10] ));
 sg13g2_dfrbp_1 _11439_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net231),
    .D(_00329_),
    .Q_N(_00066_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][11] ));
 sg13g2_dfrbp_1 _11440_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net229),
    .D(_00330_),
    .Q_N(_00064_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][12] ));
 sg13g2_dfrbp_1 _11441_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net227),
    .D(_00331_),
    .Q_N(_00070_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][13] ));
 sg13g2_dfrbp_1 _11442_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net225),
    .D(_00332_),
    .Q_N(_00068_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][14] ));
 sg13g2_dfrbp_1 _11443_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net223),
    .D(_00333_),
    .Q_N(_05559_),
    .Q(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][15] ));
 sg13g2_dfrbp_1 _11444_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net221),
    .D(_00334_),
    .Q_N(_05558_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[0] ));
 sg13g2_dfrbp_1 _11445_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net220),
    .D(_00335_),
    .Q_N(_05557_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[1] ));
 sg13g2_dfrbp_1 _11446_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net219),
    .D(_00336_),
    .Q_N(_05556_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[2] ));
 sg13g2_dfrbp_1 _11447_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net218),
    .D(_00337_),
    .Q_N(_05555_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[3] ));
 sg13g2_dfrbp_1 _11448_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net217),
    .D(_00338_),
    .Q_N(_00078_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[4] ));
 sg13g2_dfrbp_1 _11449_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net216),
    .D(_00339_),
    .Q_N(_00079_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[5] ));
 sg13g2_dfrbp_1 _11450_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net215),
    .D(_00340_),
    .Q_N(_00071_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[6] ));
 sg13g2_dfrbp_1 _11451_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net214),
    .D(_00341_),
    .Q_N(_00074_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[7] ));
 sg13g2_dfrbp_1 _11452_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net213),
    .D(_00342_),
    .Q_N(_00077_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[8] ));
 sg13g2_dfrbp_1 _11453_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net212),
    .D(_00343_),
    .Q_N(_00073_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[9] ));
 sg13g2_dfrbp_1 _11454_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net211),
    .D(_00344_),
    .Q_N(_00080_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[10] ));
 sg13g2_dfrbp_1 _11455_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net210),
    .D(_00345_),
    .Q_N(_00082_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[11] ));
 sg13g2_dfrbp_1 _11456_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net209),
    .D(_00346_),
    .Q_N(_00081_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[12] ));
 sg13g2_dfrbp_1 _11457_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net208),
    .D(_00347_),
    .Q_N(_00072_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[13] ));
 sg13g2_dfrbp_1 _11458_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net207),
    .D(_00348_),
    .Q_N(_00075_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[14] ));
 sg13g2_dfrbp_1 _11459_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net206),
    .D(_00349_),
    .Q_N(_00076_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[15] ));
 sg13g2_dfrbp_1 _11460_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net205),
    .D(_00350_),
    .Q_N(_00117_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[0] ));
 sg13g2_dfrbp_1 _11461_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net203),
    .D(_00351_),
    .Q_N(_00125_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[1] ));
 sg13g2_dfrbp_1 _11462_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net201),
    .D(_00352_),
    .Q_N(_00121_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[2] ));
 sg13g2_dfrbp_1 _11463_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net199),
    .D(_00353_),
    .Q_N(_00131_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[3] ));
 sg13g2_dfrbp_1 _11464_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net197),
    .D(_00354_),
    .Q_N(_00129_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[4] ));
 sg13g2_dfrbp_1 _11465_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net195),
    .D(_00355_),
    .Q_N(_00133_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[5] ));
 sg13g2_dfrbp_1 _11466_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net193),
    .D(_00356_),
    .Q_N(_00116_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[6] ));
 sg13g2_dfrbp_1 _11467_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net191),
    .D(_00357_),
    .Q_N(_00120_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[7] ));
 sg13g2_dfrbp_1 _11468_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net189),
    .D(_00358_),
    .Q_N(_00128_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[8] ));
 sg13g2_dfrbp_1 _11469_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net187),
    .D(_00359_),
    .Q_N(_05554_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[9] ));
 sg13g2_dfrbp_1 _11470_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net185),
    .D(_00360_),
    .Q_N(_05553_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[10] ));
 sg13g2_dfrbp_1 _11471_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net183),
    .D(_00361_),
    .Q_N(_05552_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[11] ));
 sg13g2_dfrbp_1 _11472_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net181),
    .D(_00362_),
    .Q_N(_05551_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[12] ));
 sg13g2_dfrbp_1 _11473_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net179),
    .D(_00363_),
    .Q_N(_05550_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[13] ));
 sg13g2_dfrbp_1 _11474_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net177),
    .D(_00364_),
    .Q_N(_05549_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[14] ));
 sg13g2_dfrbp_1 _11475_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net175),
    .D(_00365_),
    .Q_N(_00123_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[15] ));
 sg13g2_dfrbp_1 _11476_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net173),
    .D(_00366_),
    .Q_N(_00118_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[0] ));
 sg13g2_dfrbp_1 _11477_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net171),
    .D(_00367_),
    .Q_N(_00126_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[1] ));
 sg13g2_dfrbp_1 _11478_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net169),
    .D(_00368_),
    .Q_N(_00122_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[2] ));
 sg13g2_dfrbp_1 _11479_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net167),
    .D(_00369_),
    .Q_N(_00132_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[3] ));
 sg13g2_dfrbp_1 _11480_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net165),
    .D(_00370_),
    .Q_N(_00130_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[4] ));
 sg13g2_dfrbp_1 _11481_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net163),
    .D(_00371_),
    .Q_N(_00134_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[5] ));
 sg13g2_dfrbp_1 _11482_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net161),
    .D(_00372_),
    .Q_N(_00115_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[6] ));
 sg13g2_dfrbp_1 _11483_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net159),
    .D(_00373_),
    .Q_N(_00119_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[7] ));
 sg13g2_dfrbp_1 _11484_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net157),
    .D(_00374_),
    .Q_N(_00127_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[8] ));
 sg13g2_dfrbp_1 _11485_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net155),
    .D(_00375_),
    .Q_N(_05548_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[9] ));
 sg13g2_dfrbp_1 _11486_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net153),
    .D(_00376_),
    .Q_N(_05547_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[10] ));
 sg13g2_dfrbp_1 _11487_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net151),
    .D(_00377_),
    .Q_N(_05546_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[11] ));
 sg13g2_dfrbp_1 _11488_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net149),
    .D(_00378_),
    .Q_N(_05545_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[12] ));
 sg13g2_dfrbp_1 _11489_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net147),
    .D(_00379_),
    .Q_N(_05544_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[13] ));
 sg13g2_dfrbp_1 _11490_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net145),
    .D(_00380_),
    .Q_N(_05543_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[14] ));
 sg13g2_dfrbp_1 _11491_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net143),
    .D(_00381_),
    .Q_N(_00124_),
    .Q(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[15] ));
 sg13g2_dfrbp_1 _11492_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net142),
    .D(_00382_),
    .Q_N(_00035_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][0] ));
 sg13g2_dfrbp_1 _11493_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net141),
    .D(_00383_),
    .Q_N(_00033_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][1] ));
 sg13g2_dfrbp_1 _11494_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net140),
    .D(_00384_),
    .Q_N(_00031_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][2] ));
 sg13g2_dfrbp_1 _11495_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net139),
    .D(_00385_),
    .Q_N(_00029_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][3] ));
 sg13g2_dfrbp_1 _11496_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net138),
    .D(_00386_),
    .Q_N(_00027_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][4] ));
 sg13g2_dfrbp_1 _11497_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net137),
    .D(_00387_),
    .Q_N(_00025_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][5] ));
 sg13g2_dfrbp_1 _11498_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net136),
    .D(_00388_),
    .Q_N(_00018_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][6] ));
 sg13g2_dfrbp_1 _11499_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net135),
    .D(_00389_),
    .Q_N(_00023_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][7] ));
 sg13g2_dfrbp_1 _11500_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net134),
    .D(_00390_),
    .Q_N(_05542_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][8] ));
 sg13g2_dfrbp_1 _11501_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net133),
    .D(_00391_),
    .Q_N(_05541_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][9] ));
 sg13g2_dfrbp_1 _11502_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net132),
    .D(_00392_),
    .Q_N(_05540_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][10] ));
 sg13g2_dfrbp_1 _11503_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net131),
    .D(_00393_),
    .Q_N(_05539_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][11] ));
 sg13g2_dfrbp_1 _11504_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net130),
    .D(_00394_),
    .Q_N(_05538_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][12] ));
 sg13g2_dfrbp_1 _11505_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net129),
    .D(_00395_),
    .Q_N(_05537_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][13] ));
 sg13g2_dfrbp_1 _11506_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net128),
    .D(_00396_),
    .Q_N(_05536_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][14] ));
 sg13g2_dfrbp_1 _11507_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net127),
    .D(_00397_),
    .Q_N(_00020_),
    .Q(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][15] ));
 sg13g2_dfrbp_1 _11508_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net126),
    .D(_00398_),
    .Q_N(_05535_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][0] ));
 sg13g2_dfrbp_1 _11509_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net125),
    .D(_00399_),
    .Q_N(_05534_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][1] ));
 sg13g2_dfrbp_1 _11510_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net124),
    .D(_00400_),
    .Q_N(_05533_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][2] ));
 sg13g2_dfrbp_1 _11511_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net123),
    .D(_00401_),
    .Q_N(_05532_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][3] ));
 sg13g2_dfrbp_1 _11512_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net122),
    .D(_00402_),
    .Q_N(_05531_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][4] ));
 sg13g2_dfrbp_1 _11513_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net121),
    .D(_00403_),
    .Q_N(_05530_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][5] ));
 sg13g2_dfrbp_1 _11514_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net120),
    .D(_00404_),
    .Q_N(_05529_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][6] ));
 sg13g2_dfrbp_1 _11515_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net119),
    .D(_00405_),
    .Q_N(_05528_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][7] ));
 sg13g2_dfrbp_1 _11516_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net118),
    .D(_00406_),
    .Q_N(_05527_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][8] ));
 sg13g2_dfrbp_1 _11517_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net117),
    .D(_00407_),
    .Q_N(_05526_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][9] ));
 sg13g2_dfrbp_1 _11518_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net116),
    .D(_00408_),
    .Q_N(_05525_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][10] ));
 sg13g2_dfrbp_1 _11519_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net115),
    .D(_00409_),
    .Q_N(_05524_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][11] ));
 sg13g2_dfrbp_1 _11520_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net114),
    .D(_00410_),
    .Q_N(_05523_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][12] ));
 sg13g2_dfrbp_1 _11521_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net113),
    .D(_00411_),
    .Q_N(_05522_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][13] ));
 sg13g2_dfrbp_1 _11522_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net112),
    .D(_00412_),
    .Q_N(_05521_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][14] ));
 sg13g2_dfrbp_1 _11523_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net111),
    .D(_00413_),
    .Q_N(_05520_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[7][15] ));
 sg13g2_dfrbp_1 _11524_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net110),
    .D(_00414_),
    .Q_N(_05519_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][0] ));
 sg13g2_dfrbp_1 _11525_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net109),
    .D(_00415_),
    .Q_N(_05518_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][1] ));
 sg13g2_dfrbp_1 _11526_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net108),
    .D(_00416_),
    .Q_N(_05517_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][2] ));
 sg13g2_dfrbp_1 _11527_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net107),
    .D(_00417_),
    .Q_N(_00135_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][3] ));
 sg13g2_dfrbp_1 _11528_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net106),
    .D(_00418_),
    .Q_N(_00139_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][4] ));
 sg13g2_dfrbp_1 _11529_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net105),
    .D(_00419_),
    .Q_N(_00137_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][5] ));
 sg13g2_dfrbp_1 _11530_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net104),
    .D(_00420_),
    .Q_N(_05516_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][6] ));
 sg13g2_dfrbp_1 _11531_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net103),
    .D(net709),
    .Q_N(_05515_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][7] ));
 sg13g2_dfrbp_1 _11532_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net102),
    .D(_00422_),
    .Q_N(_05514_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][8] ));
 sg13g2_dfrbp_1 _11533_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net101),
    .D(_00423_),
    .Q_N(_05513_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][9] ));
 sg13g2_dfrbp_1 _11534_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net100),
    .D(_00424_),
    .Q_N(_05512_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][10] ));
 sg13g2_dfrbp_1 _11535_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net99),
    .D(_00425_),
    .Q_N(_05511_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][11] ));
 sg13g2_dfrbp_1 _11536_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net98),
    .D(_00426_),
    .Q_N(_05510_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][12] ));
 sg13g2_dfrbp_1 _11537_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net97),
    .D(_00427_),
    .Q_N(_05509_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][13] ));
 sg13g2_dfrbp_1 _11538_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net96),
    .D(net673),
    .Q_N(_05508_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][14] ));
 sg13g2_dfrbp_1 _11539_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net95),
    .D(net765),
    .Q_N(_05507_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[7][15] ));
 sg13g2_dfrbp_1 _11540_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net94),
    .D(_00430_),
    .Q_N(_05506_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][0] ));
 sg13g2_dfrbp_1 _11541_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net93),
    .D(net873),
    .Q_N(_05505_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][1] ));
 sg13g2_dfrbp_1 _11542_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net92),
    .D(_00432_),
    .Q_N(_05504_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][2] ));
 sg13g2_dfrbp_1 _11543_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net91),
    .D(_00433_),
    .Q_N(_05503_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][3] ));
 sg13g2_dfrbp_1 _11544_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net90),
    .D(_00434_),
    .Q_N(_05502_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][4] ));
 sg13g2_dfrbp_1 _11545_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net89),
    .D(net926),
    .Q_N(_05501_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][5] ));
 sg13g2_dfrbp_1 _11546_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net88),
    .D(net846),
    .Q_N(_05500_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][6] ));
 sg13g2_dfrbp_1 _11547_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net87),
    .D(_00437_),
    .Q_N(_05499_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][7] ));
 sg13g2_dfrbp_1 _11548_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net86),
    .D(_00438_),
    .Q_N(_05498_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][8] ));
 sg13g2_dfrbp_1 _11549_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net85),
    .D(_00439_),
    .Q_N(_05497_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][9] ));
 sg13g2_dfrbp_1 _11550_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net84),
    .D(_00440_),
    .Q_N(_05496_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][10] ));
 sg13g2_dfrbp_1 _11551_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net83),
    .D(net484),
    .Q_N(_05495_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][11] ));
 sg13g2_dfrbp_1 _11552_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net82),
    .D(_00442_),
    .Q_N(_05494_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][12] ));
 sg13g2_dfrbp_1 _11553_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net81),
    .D(_00443_),
    .Q_N(_05493_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][13] ));
 sg13g2_dfrbp_1 _11554_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net80),
    .D(_00444_),
    .Q_N(_05492_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][14] ));
 sg13g2_dfrbp_1 _11555_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net79),
    .D(_00445_),
    .Q_N(_05491_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[5][15] ));
 sg13g2_dfrbp_1 _11556_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net78),
    .D(_00446_),
    .Q_N(_05490_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][0] ));
 sg13g2_dfrbp_1 _11557_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net77),
    .D(_00447_),
    .Q_N(_05489_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][1] ));
 sg13g2_dfrbp_1 _11558_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net76),
    .D(_00448_),
    .Q_N(_05488_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][2] ));
 sg13g2_dfrbp_1 _11559_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net75),
    .D(_00449_),
    .Q_N(_00051_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][3] ));
 sg13g2_dfrbp_1 _11560_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net74),
    .D(_00450_),
    .Q_N(_00055_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][4] ));
 sg13g2_dfrbp_1 _11561_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net73),
    .D(_00451_),
    .Q_N(_00053_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][5] ));
 sg13g2_dfrbp_1 _11562_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net72),
    .D(_00452_),
    .Q_N(_05487_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][6] ));
 sg13g2_dfrbp_1 _11563_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net71),
    .D(net822),
    .Q_N(_05486_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][7] ));
 sg13g2_dfrbp_1 _11564_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net70),
    .D(net724),
    .Q_N(_05485_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][8] ));
 sg13g2_dfrbp_1 _11565_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net69),
    .D(_00455_),
    .Q_N(_05484_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][9] ));
 sg13g2_dfrbp_1 _11566_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net67),
    .D(_00456_),
    .Q_N(_05483_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][10] ));
 sg13g2_dfrbp_1 _11567_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net66),
    .D(_00457_),
    .Q_N(_05482_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][11] ));
 sg13g2_dfrbp_1 _11568_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net65),
    .D(_00458_),
    .Q_N(_05481_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][12] ));
 sg13g2_dfrbp_1 _11569_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net64),
    .D(_00459_),
    .Q_N(_05480_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][13] ));
 sg13g2_dfrbp_1 _11570_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net63),
    .D(_00460_),
    .Q_N(_05479_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][14] ));
 sg13g2_dfrbp_1 _11571_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net62),
    .D(_00461_),
    .Q_N(_05478_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[5][15] ));
 sg13g2_dfrbp_1 _11572_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net61),
    .D(_00462_),
    .Q_N(_05477_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][0] ));
 sg13g2_dfrbp_1 _11573_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net60),
    .D(net934),
    .Q_N(_05476_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][1] ));
 sg13g2_dfrbp_1 _11574_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net59),
    .D(_00464_),
    .Q_N(_05475_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][2] ));
 sg13g2_dfrbp_1 _11575_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net58),
    .D(net862),
    .Q_N(_05474_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][3] ));
 sg13g2_dfrbp_1 _11576_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net57),
    .D(net867),
    .Q_N(_05473_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][4] ));
 sg13g2_dfrbp_1 _11577_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net56),
    .D(_00467_),
    .Q_N(_05472_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][5] ));
 sg13g2_dfrbp_1 _11578_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net55),
    .D(net924),
    .Q_N(_05471_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][6] ));
 sg13g2_dfrbp_1 _11579_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net54),
    .D(net908),
    .Q_N(_05470_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][7] ));
 sg13g2_dfrbp_1 _11580_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net53),
    .D(_00470_),
    .Q_N(_05469_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][8] ));
 sg13g2_dfrbp_1 _11581_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net52),
    .D(net912),
    .Q_N(_05468_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][9] ));
 sg13g2_dfrbp_1 _11582_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net51),
    .D(_00472_),
    .Q_N(_05467_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][10] ));
 sg13g2_dfrbp_1 _11583_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net50),
    .D(net922),
    .Q_N(_05466_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][11] ));
 sg13g2_dfrbp_1 _11584_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net49),
    .D(net880),
    .Q_N(_05465_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][12] ));
 sg13g2_dfrbp_1 _11585_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net48),
    .D(_00475_),
    .Q_N(_05464_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][13] ));
 sg13g2_dfrbp_1 _11586_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net47),
    .D(_00476_),
    .Q_N(_05463_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][14] ));
 sg13g2_dfrbp_1 _11587_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net46),
    .D(_00477_),
    .Q_N(_05462_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[3][15] ));
 sg13g2_dfrbp_1 _11588_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net45),
    .D(net661),
    .Q_N(_05461_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][0] ));
 sg13g2_dfrbp_1 _11589_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net44),
    .D(net549),
    .Q_N(_00043_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][1] ));
 sg13g2_dfrbp_1 _11590_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net43),
    .D(net509),
    .Q_N(_00045_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][2] ));
 sg13g2_dfrbp_1 _11591_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net42),
    .D(net732),
    .Q_N(_05460_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][3] ));
 sg13g2_dfrbp_1 _11592_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net41),
    .D(net542),
    .Q_N(_00047_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][4] ));
 sg13g2_dfrbp_1 _11593_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net40),
    .D(net528),
    .Q_N(_00049_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][5] ));
 sg13g2_dfrbp_1 _11594_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net39),
    .D(net690),
    .Q_N(_05459_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][6] ));
 sg13g2_dfrbp_1 _11595_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net38),
    .D(net698),
    .Q_N(_05458_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][7] ));
 sg13g2_dfrbp_1 _11596_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net37),
    .D(net703),
    .Q_N(_05457_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][8] ));
 sg13g2_dfrbp_1 _11597_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net36),
    .D(net631),
    .Q_N(_05456_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][9] ));
 sg13g2_dfrbp_1 _11598_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net35),
    .D(_00488_),
    .Q_N(_05455_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][10] ));
 sg13g2_dfrbp_1 _11599_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net34),
    .D(_00489_),
    .Q_N(_05454_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][11] ));
 sg13g2_dfrbp_1 _11600_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net33),
    .D(_00490_),
    .Q_N(_05453_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][12] ));
 sg13g2_dfrbp_1 _11601_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net482),
    .D(_00491_),
    .Q_N(_05452_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][13] ));
 sg13g2_dfrbp_1 _11602_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net481),
    .D(_00492_),
    .Q_N(_05451_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][14] ));
 sg13g2_dfrbp_1 _11603_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net480),
    .D(net716),
    .Q_N(_05450_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[3][15] ));
 sg13g2_dfrbp_1 _11604_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net479),
    .D(net561),
    .Q_N(_05449_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][0] ));
 sg13g2_dfrbp_1 _11605_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net478),
    .D(net871),
    .Q_N(_05448_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][1] ));
 sg13g2_dfrbp_1 _11606_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net477),
    .D(net834),
    .Q_N(_05447_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][2] ));
 sg13g2_dfrbp_1 _11607_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net476),
    .D(net916),
    .Q_N(_05446_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][3] ));
 sg13g2_dfrbp_1 _11608_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net475),
    .D(net883),
    .Q_N(_05445_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][4] ));
 sg13g2_dfrbp_1 _11609_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net474),
    .D(net889),
    .Q_N(_05444_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][5] ));
 sg13g2_dfrbp_1 _11610_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net473),
    .D(_00500_),
    .Q_N(_05443_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][6] ));
 sg13g2_dfrbp_1 _11611_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net472),
    .D(net838),
    .Q_N(_05442_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][7] ));
 sg13g2_dfrbp_1 _11612_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net471),
    .D(net818),
    .Q_N(_05441_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][8] ));
 sg13g2_dfrbp_1 _11613_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net470),
    .D(net898),
    .Q_N(_05440_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][9] ));
 sg13g2_dfrbp_1 _11614_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net469),
    .D(net860),
    .Q_N(_05439_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][10] ));
 sg13g2_dfrbp_1 _11615_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net468),
    .D(net826),
    .Q_N(_05438_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][11] ));
 sg13g2_dfrbp_1 _11616_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net467),
    .D(net851),
    .Q_N(_05437_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][12] ));
 sg13g2_dfrbp_1 _11617_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net466),
    .D(net678),
    .Q_N(_05436_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][13] ));
 sg13g2_dfrbp_1 _11618_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net465),
    .D(net895),
    .Q_N(_05435_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][14] ));
 sg13g2_dfrbp_1 _11619_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net464),
    .D(net848),
    .Q_N(_05434_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[1][15] ));
 sg13g2_dfrbp_1 _11620_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net463),
    .D(_00510_),
    .Q_N(_05433_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][0] ));
 sg13g2_dfrbp_1 _11621_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net462),
    .D(net556),
    .Q_N(_00037_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][1] ));
 sg13g2_dfrbp_1 _11622_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net461),
    .D(_00512_),
    .Q_N(_00039_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][2] ));
 sg13g2_dfrbp_1 _11623_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net460),
    .D(_00513_),
    .Q_N(_05432_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][3] ));
 sg13g2_dfrbp_1 _11624_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net459),
    .D(_00514_),
    .Q_N(_00041_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][4] ));
 sg13g2_dfrbp_1 _11625_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net458),
    .D(_00515_),
    .Q_N(_05431_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][5] ));
 sg13g2_dfrbp_1 _11626_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net457),
    .D(net682),
    .Q_N(_05430_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][6] ));
 sg13g2_dfrbp_1 _11627_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net456),
    .D(net857),
    .Q_N(_05429_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][7] ));
 sg13g2_dfrbp_1 _11628_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net455),
    .D(net711),
    .Q_N(_05428_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][8] ));
 sg13g2_dfrbp_1 _11629_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net454),
    .D(_00519_),
    .Q_N(_05427_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][9] ));
 sg13g2_dfrbp_1 _11630_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net453),
    .D(net727),
    .Q_N(_05426_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][10] ));
 sg13g2_dfrbp_1 _11631_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net452),
    .D(_00521_),
    .Q_N(_05425_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][11] ));
 sg13g2_dfrbp_1 _11632_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net451),
    .D(_00522_),
    .Q_N(_05424_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][12] ));
 sg13g2_dfrbp_1 _11633_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net450),
    .D(_00523_),
    .Q_N(_05423_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][13] ));
 sg13g2_dfrbp_1 _11634_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net449),
    .D(net738),
    .Q_N(_05422_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][14] ));
 sg13g2_dfrbp_1 _11635_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net448),
    .D(net756),
    .Q_N(_05421_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[1][15] ));
 sg13g2_dfrbp_1 _11636_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net447),
    .D(_00526_),
    .Q_N(_05420_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][0] ));
 sg13g2_dfrbp_1 _11637_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net446),
    .D(_00527_),
    .Q_N(_05419_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][1] ));
 sg13g2_dfrbp_1 _11638_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net445),
    .D(_00528_),
    .Q_N(_05418_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][2] ));
 sg13g2_dfrbp_1 _11639_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net444),
    .D(_00529_),
    .Q_N(_05417_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][3] ));
 sg13g2_dfrbp_1 _11640_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net443),
    .D(_00530_),
    .Q_N(_05416_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][4] ));
 sg13g2_dfrbp_1 _11641_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net442),
    .D(_00531_),
    .Q_N(_05415_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][5] ));
 sg13g2_dfrbp_1 _11642_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net441),
    .D(_00532_),
    .Q_N(_05414_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][6] ));
 sg13g2_dfrbp_1 _11643_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net440),
    .D(_00533_),
    .Q_N(_05413_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][7] ));
 sg13g2_dfrbp_1 _11644_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net439),
    .D(_00534_),
    .Q_N(_05412_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][8] ));
 sg13g2_dfrbp_1 _11645_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net438),
    .D(_00535_),
    .Q_N(_05411_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][9] ));
 sg13g2_dfrbp_1 _11646_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net437),
    .D(_00536_),
    .Q_N(_05410_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][10] ));
 sg13g2_dfrbp_1 _11647_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net436),
    .D(_00537_),
    .Q_N(_05409_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][11] ));
 sg13g2_dfrbp_1 _11648_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net435),
    .D(_00538_),
    .Q_N(_05408_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][12] ));
 sg13g2_dfrbp_1 _11649_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net434),
    .D(_00539_),
    .Q_N(_05407_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][13] ));
 sg13g2_dfrbp_1 _11650_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net433),
    .D(_00540_),
    .Q_N(_05406_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][14] ));
 sg13g2_dfrbp_1 _11651_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net432),
    .D(_00541_),
    .Q_N(_05405_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[6][15] ));
 sg13g2_dfrbp_1 _11652_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net431),
    .D(_00542_),
    .Q_N(_05404_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][0] ));
 sg13g2_dfrbp_1 _11653_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net430),
    .D(_00543_),
    .Q_N(_05403_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][1] ));
 sg13g2_dfrbp_1 _11654_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net429),
    .D(_00544_),
    .Q_N(_05402_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][2] ));
 sg13g2_dfrbp_1 _11655_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net428),
    .D(_00545_),
    .Q_N(_00136_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][3] ));
 sg13g2_dfrbp_1 _11656_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net427),
    .D(_00546_),
    .Q_N(_00140_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][4] ));
 sg13g2_dfrbp_1 _11657_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net426),
    .D(net564),
    .Q_N(_00138_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][5] ));
 sg13g2_dfrbp_1 _11658_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net425),
    .D(_00548_),
    .Q_N(_05401_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][6] ));
 sg13g2_dfrbp_1 _11659_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net424),
    .D(_00549_),
    .Q_N(_05400_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][7] ));
 sg13g2_dfrbp_1 _11660_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net423),
    .D(_00550_),
    .Q_N(_05399_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][8] ));
 sg13g2_dfrbp_1 _11661_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net422),
    .D(net499),
    .Q_N(_05398_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][9] ));
 sg13g2_dfrbp_1 _11662_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net421),
    .D(_00552_),
    .Q_N(_05397_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][10] ));
 sg13g2_dfrbp_1 _11663_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net420),
    .D(_00553_),
    .Q_N(_05396_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][11] ));
 sg13g2_dfrbp_1 _11664_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net419),
    .D(_00554_),
    .Q_N(_05395_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][12] ));
 sg13g2_dfrbp_1 _11665_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net418),
    .D(_00555_),
    .Q_N(_05394_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][13] ));
 sg13g2_dfrbp_1 _11666_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net417),
    .D(_00556_),
    .Q_N(_05393_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][14] ));
 sg13g2_dfrbp_1 _11667_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net416),
    .D(_00557_),
    .Q_N(_05392_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[6][15] ));
 sg13g2_dfrbp_1 _11668_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net415),
    .D(_00558_),
    .Q_N(_05391_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][0] ));
 sg13g2_dfrbp_1 _11669_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net388),
    .D(_00559_),
    .Q_N(_05390_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][1] ));
 sg13g2_dfrbp_1 _11670_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net387),
    .D(_00560_),
    .Q_N(_05389_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][2] ));
 sg13g2_dfrbp_1 _11671_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net386),
    .D(net776),
    .Q_N(_05388_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][3] ));
 sg13g2_dfrbp_1 _11672_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net385),
    .D(_00562_),
    .Q_N(_05387_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][4] ));
 sg13g2_dfrbp_1 _11673_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net384),
    .D(net783),
    .Q_N(_05386_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][5] ));
 sg13g2_dfrbp_1 _11674_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net383),
    .D(_00564_),
    .Q_N(_05385_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][6] ));
 sg13g2_dfrbp_1 _11675_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net382),
    .D(_00565_),
    .Q_N(_05384_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][7] ));
 sg13g2_dfrbp_1 _11676_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net381),
    .D(net694),
    .Q_N(_05383_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][8] ));
 sg13g2_dfrbp_1 _11677_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net363),
    .D(net754),
    .Q_N(_05382_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][9] ));
 sg13g2_dfrbp_1 _11678_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net361),
    .D(net758),
    .Q_N(_05381_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][10] ));
 sg13g2_dfrbp_1 _11679_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net359),
    .D(_00569_),
    .Q_N(_05380_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][11] ));
 sg13g2_dfrbp_1 _11680_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net357),
    .D(_00570_),
    .Q_N(_05379_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][12] ));
 sg13g2_dfrbp_1 _11681_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net355),
    .D(_00571_),
    .Q_N(_05378_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][13] ));
 sg13g2_dfrbp_1 _11682_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net353),
    .D(net496),
    .Q_N(_05377_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][14] ));
 sg13g2_dfrbp_1 _11683_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net351),
    .D(net740),
    .Q_N(_05376_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[4][15] ));
 sg13g2_dfrbp_1 _11684_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net349),
    .D(net526),
    .Q_N(_05375_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][0] ));
 sg13g2_dfrbp_1 _11685_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net347),
    .D(net718),
    .Q_N(_05374_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][1] ));
 sg13g2_dfrbp_1 _11686_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net345),
    .D(net730),
    .Q_N(_05373_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][2] ));
 sg13g2_dfrbp_1 _11687_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net343),
    .D(_00577_),
    .Q_N(_00052_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][3] ));
 sg13g2_dfrbp_1 _11688_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net341),
    .D(net554),
    .Q_N(_00056_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][4] ));
 sg13g2_dfrbp_1 _11689_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net339),
    .D(net552),
    .Q_N(_00054_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][5] ));
 sg13g2_dfrbp_1 _11690_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net337),
    .D(net582),
    .Q_N(_05372_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][6] ));
 sg13g2_dfrbp_1 _11691_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net335),
    .D(_00581_),
    .Q_N(_05371_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][7] ));
 sg13g2_dfrbp_1 _11692_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net333),
    .D(_00582_),
    .Q_N(_05370_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][8] ));
 sg13g2_dfrbp_1 _11693_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net331),
    .D(_00583_),
    .Q_N(_05369_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][9] ));
 sg13g2_dfrbp_1 _11694_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net329),
    .D(net569),
    .Q_N(_05368_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][10] ));
 sg13g2_dfrbp_1 _11695_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net327),
    .D(_00585_),
    .Q_N(_05367_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][11] ));
 sg13g2_dfrbp_1 _11696_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net325),
    .D(_00586_),
    .Q_N(_05366_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][12] ));
 sg13g2_dfrbp_1 _11697_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net323),
    .D(_00587_),
    .Q_N(_05365_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][13] ));
 sg13g2_dfrbp_1 _11698_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net321),
    .D(net588),
    .Q_N(_05364_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][14] ));
 sg13g2_dfrbp_1 _11699_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net319),
    .D(_00589_),
    .Q_N(_05363_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[4][15] ));
 sg13g2_dfrbp_1 _11700_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net318),
    .D(net910),
    .Q_N(_05362_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][0] ));
 sg13g2_dfrbp_1 _11701_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net252),
    .D(_00591_),
    .Q_N(_05361_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][1] ));
 sg13g2_dfrbp_1 _11702_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net250),
    .D(net749),
    .Q_N(_05360_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][2] ));
 sg13g2_dfrbp_1 _11703_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net248),
    .D(_00593_),
    .Q_N(_05359_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][3] ));
 sg13g2_dfrbp_1 _11704_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net246),
    .D(net770),
    .Q_N(_05358_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][4] ));
 sg13g2_dfrbp_1 _11705_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net244),
    .D(net742),
    .Q_N(_05357_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][5] ));
 sg13g2_dfrbp_1 _11706_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net242),
    .D(_00596_),
    .Q_N(_05356_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][6] ));
 sg13g2_dfrbp_1 _11707_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net240),
    .D(net752),
    .Q_N(_05355_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][7] ));
 sg13g2_dfrbp_1 _11708_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net238),
    .D(net864),
    .Q_N(_05354_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][8] ));
 sg13g2_dfrbp_1 _11709_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net236),
    .D(net744),
    .Q_N(_05353_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][9] ));
 sg13g2_dfrbp_1 _11710_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net234),
    .D(_00600_),
    .Q_N(_05352_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][10] ));
 sg13g2_dfrbp_1 _11711_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net232),
    .D(net844),
    .Q_N(_05351_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][11] ));
 sg13g2_dfrbp_1 _11712_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net230),
    .D(net746),
    .Q_N(_05350_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][12] ));
 sg13g2_dfrbp_1 _11713_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net228),
    .D(_00603_),
    .Q_N(_05349_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][13] ));
 sg13g2_dfrbp_1 _11714_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net226),
    .D(net788),
    .Q_N(_05348_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][14] ));
 sg13g2_dfrbp_1 _11715_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net224),
    .D(_00605_),
    .Q_N(_05347_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[2][15] ));
 sg13g2_dfrbp_1 _11716_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net222),
    .D(_00606_),
    .Q_N(_05346_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][0] ));
 sg13g2_dfrbp_1 _11717_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net204),
    .D(net544),
    .Q_N(_00044_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][1] ));
 sg13g2_dfrbp_1 _11718_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net202),
    .D(_00608_),
    .Q_N(_00046_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][2] ));
 sg13g2_dfrbp_1 _11719_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net200),
    .D(net585),
    .Q_N(_05345_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][3] ));
 sg13g2_dfrbp_1 _11720_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net198),
    .D(_00610_),
    .Q_N(_00048_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][4] ));
 sg13g2_dfrbp_1 _11721_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net196),
    .D(net547),
    .Q_N(_00050_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][5] ));
 sg13g2_dfrbp_1 _11722_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net194),
    .D(net622),
    .Q_N(_05344_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][6] ));
 sg13g2_dfrbp_1 _11723_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net192),
    .D(net638),
    .Q_N(_05343_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][7] ));
 sg13g2_dfrbp_1 _11724_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net190),
    .D(net624),
    .Q_N(_05342_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][8] ));
 sg13g2_dfrbp_1 _11725_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net188),
    .D(net598),
    .Q_N(_05341_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][9] ));
 sg13g2_dfrbp_1 _11726_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net186),
    .D(net654),
    .Q_N(_05340_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][10] ));
 sg13g2_dfrbp_1 _11727_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net184),
    .D(_00617_),
    .Q_N(_05339_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][11] ));
 sg13g2_dfrbp_1 _11728_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net182),
    .D(_00618_),
    .Q_N(_05338_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][12] ));
 sg13g2_dfrbp_1 _11729_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net180),
    .D(_00619_),
    .Q_N(_05337_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][13] ));
 sg13g2_dfrbp_1 _11730_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net178),
    .D(net512),
    .Q_N(_05336_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][14] ));
 sg13g2_dfrbp_1 _11731_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net176),
    .D(net576),
    .Q_N(_05335_),
    .Q(\u_tiny_nn_top.u_core.param_val_op_q[2][15] ));
 sg13g2_dfrbp_1 _11732_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net174),
    .D(net669),
    .Q_N(_05334_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][0] ));
 sg13g2_dfrbp_1 _11733_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net172),
    .D(net643),
    .Q_N(_05333_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][1] ));
 sg13g2_dfrbp_1 _11734_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net170),
    .D(net626),
    .Q_N(_05332_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][2] ));
 sg13g2_dfrbp_1 _11735_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net168),
    .D(net593),
    .Q_N(_05331_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][3] ));
 sg13g2_dfrbp_1 _11736_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net166),
    .D(net707),
    .Q_N(_05330_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][4] ));
 sg13g2_dfrbp_1 _11737_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net164),
    .D(net558),
    .Q_N(_05329_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][5] ));
 sg13g2_dfrbp_1 _11738_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net162),
    .D(net573),
    .Q_N(_05328_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][6] ));
 sg13g2_dfrbp_1 _11739_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net160),
    .D(net571),
    .Q_N(_05327_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][7] ));
 sg13g2_dfrbp_1 _11740_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net158),
    .D(net633),
    .Q_N(_05326_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][8] ));
 sg13g2_dfrbp_1 _11741_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net156),
    .D(net619),
    .Q_N(_05325_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][9] ));
 sg13g2_dfrbp_1 _11742_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net154),
    .D(net608),
    .Q_N(_05324_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][10] ));
 sg13g2_dfrbp_1 _11743_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net152),
    .D(net687),
    .Q_N(_05323_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][11] ));
 sg13g2_dfrbp_1 _11744_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net150),
    .D(net567),
    .Q_N(_05322_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][12] ));
 sg13g2_dfrbp_1 _11745_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net148),
    .D(net580),
    .Q_N(_05321_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][13] ));
 sg13g2_dfrbp_1 _11746_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net146),
    .D(net645),
    .Q_N(_05320_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][14] ));
 sg13g2_dfrbp_1 _11747_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net144),
    .D(net615),
    .Q_N(_05319_),
    .Q(\u_tiny_nn_top.u_core.mul_val_op_q[0][15] ));
 sg13g2_tiehi _11599__34 (.L_HI(net34));
 sg13g2_tiehi _11598__35 (.L_HI(net35));
 sg13g2_tiehi _11597__36 (.L_HI(net36));
 sg13g2_tiehi _11596__37 (.L_HI(net37));
 sg13g2_tiehi _11595__38 (.L_HI(net38));
 sg13g2_tiehi _11594__39 (.L_HI(net39));
 sg13g2_tiehi _11593__40 (.L_HI(net40));
 sg13g2_tiehi _11592__41 (.L_HI(net41));
 sg13g2_tiehi _11591__42 (.L_HI(net42));
 sg13g2_tiehi _11590__43 (.L_HI(net43));
 sg13g2_tiehi _11589__44 (.L_HI(net44));
 sg13g2_tiehi _11588__45 (.L_HI(net45));
 sg13g2_tiehi _11587__46 (.L_HI(net46));
 sg13g2_tiehi _11586__47 (.L_HI(net47));
 sg13g2_tiehi _11585__48 (.L_HI(net48));
 sg13g2_tiehi _11584__49 (.L_HI(net49));
 sg13g2_tiehi _11583__50 (.L_HI(net50));
 sg13g2_tiehi _11582__51 (.L_HI(net51));
 sg13g2_tiehi _11581__52 (.L_HI(net52));
 sg13g2_tiehi _11580__53 (.L_HI(net53));
 sg13g2_tiehi _11579__54 (.L_HI(net54));
 sg13g2_tiehi _11578__55 (.L_HI(net55));
 sg13g2_tiehi _11577__56 (.L_HI(net56));
 sg13g2_tiehi _11576__57 (.L_HI(net57));
 sg13g2_tiehi _11575__58 (.L_HI(net58));
 sg13g2_tiehi _11574__59 (.L_HI(net59));
 sg13g2_tiehi _11573__60 (.L_HI(net60));
 sg13g2_tiehi _11572__61 (.L_HI(net61));
 sg13g2_tiehi _11571__62 (.L_HI(net62));
 sg13g2_tiehi _11570__63 (.L_HI(net63));
 sg13g2_tiehi _11569__64 (.L_HI(net64));
 sg13g2_tiehi _11568__65 (.L_HI(net65));
 sg13g2_tiehi _11567__66 (.L_HI(net66));
 sg13g2_tiehi _11566__67 (.L_HI(net67));
 sg13g2_tiehi _11256__68 (.L_HI(net68));
 sg13g2_tiehi _11565__69 (.L_HI(net69));
 sg13g2_tiehi _11564__70 (.L_HI(net70));
 sg13g2_tiehi _11563__71 (.L_HI(net71));
 sg13g2_tiehi _11562__72 (.L_HI(net72));
 sg13g2_tiehi _11561__73 (.L_HI(net73));
 sg13g2_tiehi _11560__74 (.L_HI(net74));
 sg13g2_tiehi _11559__75 (.L_HI(net75));
 sg13g2_tiehi _11558__76 (.L_HI(net76));
 sg13g2_tiehi _11557__77 (.L_HI(net77));
 sg13g2_tiehi _11556__78 (.L_HI(net78));
 sg13g2_tiehi _11555__79 (.L_HI(net79));
 sg13g2_tiehi _11554__80 (.L_HI(net80));
 sg13g2_tiehi _11553__81 (.L_HI(net81));
 sg13g2_tiehi _11552__82 (.L_HI(net82));
 sg13g2_tiehi _11551__83 (.L_HI(net83));
 sg13g2_tiehi _11550__84 (.L_HI(net84));
 sg13g2_tiehi _11549__85 (.L_HI(net85));
 sg13g2_tiehi _11548__86 (.L_HI(net86));
 sg13g2_tiehi _11547__87 (.L_HI(net87));
 sg13g2_tiehi _11546__88 (.L_HI(net88));
 sg13g2_tiehi _11545__89 (.L_HI(net89));
 sg13g2_tiehi _11544__90 (.L_HI(net90));
 sg13g2_tiehi _11543__91 (.L_HI(net91));
 sg13g2_tiehi _11542__92 (.L_HI(net92));
 sg13g2_tiehi _11541__93 (.L_HI(net93));
 sg13g2_tiehi _11540__94 (.L_HI(net94));
 sg13g2_tiehi _11539__95 (.L_HI(net95));
 sg13g2_tiehi _11538__96 (.L_HI(net96));
 sg13g2_tiehi _11537__97 (.L_HI(net97));
 sg13g2_tiehi _11536__98 (.L_HI(net98));
 sg13g2_tiehi _11535__99 (.L_HI(net99));
 sg13g2_tiehi _11534__100 (.L_HI(net100));
 sg13g2_tiehi _11533__101 (.L_HI(net101));
 sg13g2_tiehi _11532__102 (.L_HI(net102));
 sg13g2_tiehi _11531__103 (.L_HI(net103));
 sg13g2_tiehi _11530__104 (.L_HI(net104));
 sg13g2_tiehi _11529__105 (.L_HI(net105));
 sg13g2_tiehi _11528__106 (.L_HI(net106));
 sg13g2_tiehi _11527__107 (.L_HI(net107));
 sg13g2_tiehi _11526__108 (.L_HI(net108));
 sg13g2_tiehi _11525__109 (.L_HI(net109));
 sg13g2_tiehi _11524__110 (.L_HI(net110));
 sg13g2_tiehi _11523__111 (.L_HI(net111));
 sg13g2_tiehi _11522__112 (.L_HI(net112));
 sg13g2_tiehi _11521__113 (.L_HI(net113));
 sg13g2_tiehi _11520__114 (.L_HI(net114));
 sg13g2_tiehi _11519__115 (.L_HI(net115));
 sg13g2_tiehi _11518__116 (.L_HI(net116));
 sg13g2_tiehi _11517__117 (.L_HI(net117));
 sg13g2_tiehi _11516__118 (.L_HI(net118));
 sg13g2_tiehi _11515__119 (.L_HI(net119));
 sg13g2_tiehi _11514__120 (.L_HI(net120));
 sg13g2_tiehi _11513__121 (.L_HI(net121));
 sg13g2_tiehi _11512__122 (.L_HI(net122));
 sg13g2_tiehi _11511__123 (.L_HI(net123));
 sg13g2_tiehi _11510__124 (.L_HI(net124));
 sg13g2_tiehi _11509__125 (.L_HI(net125));
 sg13g2_tiehi _11508__126 (.L_HI(net126));
 sg13g2_tiehi _11507__127 (.L_HI(net127));
 sg13g2_tiehi _11506__128 (.L_HI(net128));
 sg13g2_tiehi _11505__129 (.L_HI(net129));
 sg13g2_tiehi _11504__130 (.L_HI(net130));
 sg13g2_tiehi _11503__131 (.L_HI(net131));
 sg13g2_tiehi _11502__132 (.L_HI(net132));
 sg13g2_tiehi _11501__133 (.L_HI(net133));
 sg13g2_tiehi _11500__134 (.L_HI(net134));
 sg13g2_tiehi _11499__135 (.L_HI(net135));
 sg13g2_tiehi _11498__136 (.L_HI(net136));
 sg13g2_tiehi _11497__137 (.L_HI(net137));
 sg13g2_tiehi _11496__138 (.L_HI(net138));
 sg13g2_tiehi _11495__139 (.L_HI(net139));
 sg13g2_tiehi _11494__140 (.L_HI(net140));
 sg13g2_tiehi _11493__141 (.L_HI(net141));
 sg13g2_tiehi _11492__142 (.L_HI(net142));
 sg13g2_tiehi _11491__143 (.L_HI(net143));
 sg13g2_tiehi _11747__144 (.L_HI(net144));
 sg13g2_tiehi _11490__145 (.L_HI(net145));
 sg13g2_tiehi _11746__146 (.L_HI(net146));
 sg13g2_tiehi _11489__147 (.L_HI(net147));
 sg13g2_tiehi _11745__148 (.L_HI(net148));
 sg13g2_tiehi _11488__149 (.L_HI(net149));
 sg13g2_tiehi _11744__150 (.L_HI(net150));
 sg13g2_tiehi _11487__151 (.L_HI(net151));
 sg13g2_tiehi _11743__152 (.L_HI(net152));
 sg13g2_tiehi _11486__153 (.L_HI(net153));
 sg13g2_tiehi _11742__154 (.L_HI(net154));
 sg13g2_tiehi _11485__155 (.L_HI(net155));
 sg13g2_tiehi _11741__156 (.L_HI(net156));
 sg13g2_tiehi _11484__157 (.L_HI(net157));
 sg13g2_tiehi _11740__158 (.L_HI(net158));
 sg13g2_tiehi _11483__159 (.L_HI(net159));
 sg13g2_tiehi _11739__160 (.L_HI(net160));
 sg13g2_tiehi _11482__161 (.L_HI(net161));
 sg13g2_tiehi _11738__162 (.L_HI(net162));
 sg13g2_tiehi _11481__163 (.L_HI(net163));
 sg13g2_tiehi _11737__164 (.L_HI(net164));
 sg13g2_tiehi _11480__165 (.L_HI(net165));
 sg13g2_tiehi _11736__166 (.L_HI(net166));
 sg13g2_tiehi _11479__167 (.L_HI(net167));
 sg13g2_tiehi _11735__168 (.L_HI(net168));
 sg13g2_tiehi _11478__169 (.L_HI(net169));
 sg13g2_tiehi _11734__170 (.L_HI(net170));
 sg13g2_tiehi _11477__171 (.L_HI(net171));
 sg13g2_tiehi _11733__172 (.L_HI(net172));
 sg13g2_tiehi _11476__173 (.L_HI(net173));
 sg13g2_tiehi _11732__174 (.L_HI(net174));
 sg13g2_tiehi _11475__175 (.L_HI(net175));
 sg13g2_tiehi _11731__176 (.L_HI(net176));
 sg13g2_tiehi _11474__177 (.L_HI(net177));
 sg13g2_tiehi _11730__178 (.L_HI(net178));
 sg13g2_tiehi _11473__179 (.L_HI(net179));
 sg13g2_tiehi _11729__180 (.L_HI(net180));
 sg13g2_tiehi _11472__181 (.L_HI(net181));
 sg13g2_tiehi _11728__182 (.L_HI(net182));
 sg13g2_tiehi _11471__183 (.L_HI(net183));
 sg13g2_tiehi _11727__184 (.L_HI(net184));
 sg13g2_tiehi _11470__185 (.L_HI(net185));
 sg13g2_tiehi _11726__186 (.L_HI(net186));
 sg13g2_tiehi _11469__187 (.L_HI(net187));
 sg13g2_tiehi _11725__188 (.L_HI(net188));
 sg13g2_tiehi _11468__189 (.L_HI(net189));
 sg13g2_tiehi _11724__190 (.L_HI(net190));
 sg13g2_tiehi _11467__191 (.L_HI(net191));
 sg13g2_tiehi _11723__192 (.L_HI(net192));
 sg13g2_tiehi _11466__193 (.L_HI(net193));
 sg13g2_tiehi _11722__194 (.L_HI(net194));
 sg13g2_tiehi _11465__195 (.L_HI(net195));
 sg13g2_tiehi _11721__196 (.L_HI(net196));
 sg13g2_tiehi _11464__197 (.L_HI(net197));
 sg13g2_tiehi _11720__198 (.L_HI(net198));
 sg13g2_tiehi _11463__199 (.L_HI(net199));
 sg13g2_tiehi _11719__200 (.L_HI(net200));
 sg13g2_tiehi _11462__201 (.L_HI(net201));
 sg13g2_tiehi _11718__202 (.L_HI(net202));
 sg13g2_tiehi _11461__203 (.L_HI(net203));
 sg13g2_tiehi _11717__204 (.L_HI(net204));
 sg13g2_tiehi _11460__205 (.L_HI(net205));
 sg13g2_tiehi _11459__206 (.L_HI(net206));
 sg13g2_tiehi _11458__207 (.L_HI(net207));
 sg13g2_tiehi _11457__208 (.L_HI(net208));
 sg13g2_tiehi _11456__209 (.L_HI(net209));
 sg13g2_tiehi _11455__210 (.L_HI(net210));
 sg13g2_tiehi _11454__211 (.L_HI(net211));
 sg13g2_tiehi _11453__212 (.L_HI(net212));
 sg13g2_tiehi _11452__213 (.L_HI(net213));
 sg13g2_tiehi _11451__214 (.L_HI(net214));
 sg13g2_tiehi _11450__215 (.L_HI(net215));
 sg13g2_tiehi _11449__216 (.L_HI(net216));
 sg13g2_tiehi _11448__217 (.L_HI(net217));
 sg13g2_tiehi _11447__218 (.L_HI(net218));
 sg13g2_tiehi _11446__219 (.L_HI(net219));
 sg13g2_tiehi _11445__220 (.L_HI(net220));
 sg13g2_tiehi _11444__221 (.L_HI(net221));
 sg13g2_tiehi _11716__222 (.L_HI(net222));
 sg13g2_tiehi _11443__223 (.L_HI(net223));
 sg13g2_tiehi _11715__224 (.L_HI(net224));
 sg13g2_tiehi _11442__225 (.L_HI(net225));
 sg13g2_tiehi _11714__226 (.L_HI(net226));
 sg13g2_tiehi _11441__227 (.L_HI(net227));
 sg13g2_tiehi _11713__228 (.L_HI(net228));
 sg13g2_tiehi _11440__229 (.L_HI(net229));
 sg13g2_tiehi _11712__230 (.L_HI(net230));
 sg13g2_tiehi _11439__231 (.L_HI(net231));
 sg13g2_tiehi _11711__232 (.L_HI(net232));
 sg13g2_tiehi _11438__233 (.L_HI(net233));
 sg13g2_tiehi _11710__234 (.L_HI(net234));
 sg13g2_tiehi _11437__235 (.L_HI(net235));
 sg13g2_tiehi _11709__236 (.L_HI(net236));
 sg13g2_tiehi _11436__237 (.L_HI(net237));
 sg13g2_tiehi _11708__238 (.L_HI(net238));
 sg13g2_tiehi _11435__239 (.L_HI(net239));
 sg13g2_tiehi _11707__240 (.L_HI(net240));
 sg13g2_tiehi _11434__241 (.L_HI(net241));
 sg13g2_tiehi _11706__242 (.L_HI(net242));
 sg13g2_tiehi _11433__243 (.L_HI(net243));
 sg13g2_tiehi _11705__244 (.L_HI(net244));
 sg13g2_tiehi _11432__245 (.L_HI(net245));
 sg13g2_tiehi _11704__246 (.L_HI(net246));
 sg13g2_tiehi _11431__247 (.L_HI(net247));
 sg13g2_tiehi _11703__248 (.L_HI(net248));
 sg13g2_tiehi _11430__249 (.L_HI(net249));
 sg13g2_tiehi _11702__250 (.L_HI(net250));
 sg13g2_tiehi _11429__251 (.L_HI(net251));
 sg13g2_tiehi _11701__252 (.L_HI(net252));
 sg13g2_tiehi _11428__253 (.L_HI(net253));
 sg13g2_tiehi _11427__254 (.L_HI(net254));
 sg13g2_tiehi _11426__255 (.L_HI(net255));
 sg13g2_tiehi _11425__256 (.L_HI(net256));
 sg13g2_tiehi _11424__257 (.L_HI(net257));
 sg13g2_tiehi _11423__258 (.L_HI(net258));
 sg13g2_tiehi _11422__259 (.L_HI(net259));
 sg13g2_tiehi _11421__260 (.L_HI(net260));
 sg13g2_tiehi _11420__261 (.L_HI(net261));
 sg13g2_tiehi _11419__262 (.L_HI(net262));
 sg13g2_tiehi _11418__263 (.L_HI(net263));
 sg13g2_tiehi _11417__264 (.L_HI(net264));
 sg13g2_tiehi _11416__265 (.L_HI(net265));
 sg13g2_tiehi _11415__266 (.L_HI(net266));
 sg13g2_tiehi _11414__267 (.L_HI(net267));
 sg13g2_tiehi _11413__268 (.L_HI(net268));
 sg13g2_tiehi _11412__269 (.L_HI(net269));
 sg13g2_tiehi _11411__270 (.L_HI(net270));
 sg13g2_tiehi _11410__271 (.L_HI(net271));
 sg13g2_tiehi _11409__272 (.L_HI(net272));
 sg13g2_tiehi _11408__273 (.L_HI(net273));
 sg13g2_tiehi _11407__274 (.L_HI(net274));
 sg13g2_tiehi _11406__275 (.L_HI(net275));
 sg13g2_tiehi _11405__276 (.L_HI(net276));
 sg13g2_tiehi _11404__277 (.L_HI(net277));
 sg13g2_tiehi _11403__278 (.L_HI(net278));
 sg13g2_tiehi _11402__279 (.L_HI(net279));
 sg13g2_tiehi _11401__280 (.L_HI(net280));
 sg13g2_tiehi _11400__281 (.L_HI(net281));
 sg13g2_tiehi _11399__282 (.L_HI(net282));
 sg13g2_tiehi _11398__283 (.L_HI(net283));
 sg13g2_tiehi _11397__284 (.L_HI(net284));
 sg13g2_tiehi _11396__285 (.L_HI(net285));
 sg13g2_tiehi _11395__286 (.L_HI(net286));
 sg13g2_tiehi _11394__287 (.L_HI(net287));
 sg13g2_tiehi _11393__288 (.L_HI(net288));
 sg13g2_tiehi _11392__289 (.L_HI(net289));
 sg13g2_tiehi _11391__290 (.L_HI(net290));
 sg13g2_tiehi _11390__291 (.L_HI(net291));
 sg13g2_tiehi _11389__292 (.L_HI(net292));
 sg13g2_tiehi _11388__293 (.L_HI(net293));
 sg13g2_tiehi _11387__294 (.L_HI(net294));
 sg13g2_tiehi _11386__295 (.L_HI(net295));
 sg13g2_tiehi _11385__296 (.L_HI(net296));
 sg13g2_tiehi _11384__297 (.L_HI(net297));
 sg13g2_tiehi _11383__298 (.L_HI(net298));
 sg13g2_tiehi _11382__299 (.L_HI(net299));
 sg13g2_tiehi _11381__300 (.L_HI(net300));
 sg13g2_tiehi _11380__301 (.L_HI(net301));
 sg13g2_tiehi _11379__302 (.L_HI(net302));
 sg13g2_tiehi _11378__303 (.L_HI(net303));
 sg13g2_tiehi _11377__304 (.L_HI(net304));
 sg13g2_tiehi _11376__305 (.L_HI(net305));
 sg13g2_tiehi _11375__306 (.L_HI(net306));
 sg13g2_tiehi _11374__307 (.L_HI(net307));
 sg13g2_tiehi _11373__308 (.L_HI(net308));
 sg13g2_tiehi _11372__309 (.L_HI(net309));
 sg13g2_tiehi _11371__310 (.L_HI(net310));
 sg13g2_tiehi _11370__311 (.L_HI(net311));
 sg13g2_tiehi _11369__312 (.L_HI(net312));
 sg13g2_tiehi _11368__313 (.L_HI(net313));
 sg13g2_tiehi _11367__314 (.L_HI(net314));
 sg13g2_tiehi _11366__315 (.L_HI(net315));
 sg13g2_tiehi _11365__316 (.L_HI(net316));
 sg13g2_tiehi _11364__317 (.L_HI(net317));
 sg13g2_tiehi _11700__318 (.L_HI(net318));
 sg13g2_tiehi _11699__319 (.L_HI(net319));
 sg13g2_tiehi _11345__320 (.L_HI(net320));
 sg13g2_tiehi _11698__321 (.L_HI(net321));
 sg13g2_tiehi _11344__322 (.L_HI(net322));
 sg13g2_tiehi _11697__323 (.L_HI(net323));
 sg13g2_tiehi _11343__324 (.L_HI(net324));
 sg13g2_tiehi _11696__325 (.L_HI(net325));
 sg13g2_tiehi _11342__326 (.L_HI(net326));
 sg13g2_tiehi _11695__327 (.L_HI(net327));
 sg13g2_tiehi _11341__328 (.L_HI(net328));
 sg13g2_tiehi _11694__329 (.L_HI(net329));
 sg13g2_tiehi _11340__330 (.L_HI(net330));
 sg13g2_tiehi _11693__331 (.L_HI(net331));
 sg13g2_tiehi _11339__332 (.L_HI(net332));
 sg13g2_tiehi _11692__333 (.L_HI(net333));
 sg13g2_tiehi _11338__334 (.L_HI(net334));
 sg13g2_tiehi _11691__335 (.L_HI(net335));
 sg13g2_tiehi _11337__336 (.L_HI(net336));
 sg13g2_tiehi _11690__337 (.L_HI(net337));
 sg13g2_tiehi _11336__338 (.L_HI(net338));
 sg13g2_tiehi _11689__339 (.L_HI(net339));
 sg13g2_tiehi _11335__340 (.L_HI(net340));
 sg13g2_tiehi _11688__341 (.L_HI(net341));
 sg13g2_tiehi _11334__342 (.L_HI(net342));
 sg13g2_tiehi _11687__343 (.L_HI(net343));
 sg13g2_tiehi _11333__344 (.L_HI(net344));
 sg13g2_tiehi _11686__345 (.L_HI(net345));
 sg13g2_tiehi _11332__346 (.L_HI(net346));
 sg13g2_tiehi _11685__347 (.L_HI(net347));
 sg13g2_tiehi _11331__348 (.L_HI(net348));
 sg13g2_tiehi _11684__349 (.L_HI(net349));
 sg13g2_tiehi _11330__350 (.L_HI(net350));
 sg13g2_tiehi _11683__351 (.L_HI(net351));
 sg13g2_tiehi _11329__352 (.L_HI(net352));
 sg13g2_tiehi _11682__353 (.L_HI(net353));
 sg13g2_tiehi _11328__354 (.L_HI(net354));
 sg13g2_tiehi _11681__355 (.L_HI(net355));
 sg13g2_tiehi _11327__356 (.L_HI(net356));
 sg13g2_tiehi _11680__357 (.L_HI(net357));
 sg13g2_tiehi _11326__358 (.L_HI(net358));
 sg13g2_tiehi _11679__359 (.L_HI(net359));
 sg13g2_tiehi _11325__360 (.L_HI(net360));
 sg13g2_tiehi _11678__361 (.L_HI(net361));
 sg13g2_tiehi _11324__362 (.L_HI(net362));
 sg13g2_tiehi _11677__363 (.L_HI(net363));
 sg13g2_tiehi _11323__364 (.L_HI(net364));
 sg13g2_tiehi _11322__365 (.L_HI(net365));
 sg13g2_tiehi _11321__366 (.L_HI(net366));
 sg13g2_tiehi _11320__367 (.L_HI(net367));
 sg13g2_tiehi _11319__368 (.L_HI(net368));
 sg13g2_tiehi _11318__369 (.L_HI(net369));
 sg13g2_tiehi _11317__370 (.L_HI(net370));
 sg13g2_tiehi _11316__371 (.L_HI(net371));
 sg13g2_tiehi _11315__372 (.L_HI(net372));
 sg13g2_tiehi _11314__373 (.L_HI(net373));
 sg13g2_tiehi _11313__374 (.L_HI(net374));
 sg13g2_tiehi _11312__375 (.L_HI(net375));
 sg13g2_tiehi _11311__376 (.L_HI(net376));
 sg13g2_tiehi _11310__377 (.L_HI(net377));
 sg13g2_tiehi _11309__378 (.L_HI(net378));
 sg13g2_tiehi _11308__379 (.L_HI(net379));
 sg13g2_tiehi _11307__380 (.L_HI(net380));
 sg13g2_tiehi _11676__381 (.L_HI(net381));
 sg13g2_tiehi _11675__382 (.L_HI(net382));
 sg13g2_tiehi _11674__383 (.L_HI(net383));
 sg13g2_tiehi _11673__384 (.L_HI(net384));
 sg13g2_tiehi _11672__385 (.L_HI(net385));
 sg13g2_tiehi _11671__386 (.L_HI(net386));
 sg13g2_tiehi _11670__387 (.L_HI(net387));
 sg13g2_tiehi _11669__388 (.L_HI(net388));
 sg13g2_tiehi _11282__389 (.L_HI(net389));
 sg13g2_tiehi _11281__390 (.L_HI(net390));
 sg13g2_tiehi _11280__391 (.L_HI(net391));
 sg13g2_tiehi _11279__392 (.L_HI(net392));
 sg13g2_tiehi _11278__393 (.L_HI(net393));
 sg13g2_tiehi _11277__394 (.L_HI(net394));
 sg13g2_tiehi _11276__395 (.L_HI(net395));
 sg13g2_tiehi _11275__396 (.L_HI(net396));
 sg13g2_tiehi _11274__397 (.L_HI(net397));
 sg13g2_tiehi _11273__398 (.L_HI(net398));
 sg13g2_tiehi _11272__399 (.L_HI(net399));
 sg13g2_tiehi _11271__400 (.L_HI(net400));
 sg13g2_tiehi _11270__401 (.L_HI(net401));
 sg13g2_tiehi _11269__402 (.L_HI(net402));
 sg13g2_tiehi _11268__403 (.L_HI(net403));
 sg13g2_tiehi _11267__404 (.L_HI(net404));
 sg13g2_tiehi _11266__405 (.L_HI(net405));
 sg13g2_tiehi _11265__406 (.L_HI(net406));
 sg13g2_tiehi _11264__407 (.L_HI(net407));
 sg13g2_tiehi _11263__408 (.L_HI(net408));
 sg13g2_tiehi _11262__409 (.L_HI(net409));
 sg13g2_tiehi _11261__410 (.L_HI(net410));
 sg13g2_tiehi _11260__411 (.L_HI(net411));
 sg13g2_tiehi _11259__412 (.L_HI(net412));
 sg13g2_tiehi _11258__413 (.L_HI(net413));
 sg13g2_tiehi _11257__414 (.L_HI(net414));
 sg13g2_tiehi _11668__415 (.L_HI(net415));
 sg13g2_tiehi _11667__416 (.L_HI(net416));
 sg13g2_tiehi _11666__417 (.L_HI(net417));
 sg13g2_tiehi _11665__418 (.L_HI(net418));
 sg13g2_tiehi _11664__419 (.L_HI(net419));
 sg13g2_tiehi _11663__420 (.L_HI(net420));
 sg13g2_tiehi _11662__421 (.L_HI(net421));
 sg13g2_tiehi _11661__422 (.L_HI(net422));
 sg13g2_tiehi _11660__423 (.L_HI(net423));
 sg13g2_tiehi _11659__424 (.L_HI(net424));
 sg13g2_tiehi _11658__425 (.L_HI(net425));
 sg13g2_tiehi _11657__426 (.L_HI(net426));
 sg13g2_tiehi _11656__427 (.L_HI(net427));
 sg13g2_tiehi _11655__428 (.L_HI(net428));
 sg13g2_tiehi _11654__429 (.L_HI(net429));
 sg13g2_tiehi _11653__430 (.L_HI(net430));
 sg13g2_tiehi _11652__431 (.L_HI(net431));
 sg13g2_tiehi _11651__432 (.L_HI(net432));
 sg13g2_tiehi _11650__433 (.L_HI(net433));
 sg13g2_tiehi _11649__434 (.L_HI(net434));
 sg13g2_tiehi _11648__435 (.L_HI(net435));
 sg13g2_tiehi _11647__436 (.L_HI(net436));
 sg13g2_tiehi _11646__437 (.L_HI(net437));
 sg13g2_tiehi _11645__438 (.L_HI(net438));
 sg13g2_tiehi _11644__439 (.L_HI(net439));
 sg13g2_tiehi _11643__440 (.L_HI(net440));
 sg13g2_tiehi _11642__441 (.L_HI(net441));
 sg13g2_tiehi _11641__442 (.L_HI(net442));
 sg13g2_tiehi _11640__443 (.L_HI(net443));
 sg13g2_tiehi _11639__444 (.L_HI(net444));
 sg13g2_tiehi _11638__445 (.L_HI(net445));
 sg13g2_tiehi _11637__446 (.L_HI(net446));
 sg13g2_tiehi _11636__447 (.L_HI(net447));
 sg13g2_tiehi _11635__448 (.L_HI(net448));
 sg13g2_tiehi _11634__449 (.L_HI(net449));
 sg13g2_tiehi _11633__450 (.L_HI(net450));
 sg13g2_tiehi _11632__451 (.L_HI(net451));
 sg13g2_tiehi _11631__452 (.L_HI(net452));
 sg13g2_tiehi _11630__453 (.L_HI(net453));
 sg13g2_tiehi _11629__454 (.L_HI(net454));
 sg13g2_tiehi _11628__455 (.L_HI(net455));
 sg13g2_tiehi _11627__456 (.L_HI(net456));
 sg13g2_tiehi _11626__457 (.L_HI(net457));
 sg13g2_tiehi _11625__458 (.L_HI(net458));
 sg13g2_tiehi _11624__459 (.L_HI(net459));
 sg13g2_tiehi _11623__460 (.L_HI(net460));
 sg13g2_tiehi _11622__461 (.L_HI(net461));
 sg13g2_tiehi _11621__462 (.L_HI(net462));
 sg13g2_tiehi _11620__463 (.L_HI(net463));
 sg13g2_tiehi _11619__464 (.L_HI(net464));
 sg13g2_tiehi _11618__465 (.L_HI(net465));
 sg13g2_tiehi _11617__466 (.L_HI(net466));
 sg13g2_tiehi _11616__467 (.L_HI(net467));
 sg13g2_tiehi _11615__468 (.L_HI(net468));
 sg13g2_tiehi _11614__469 (.L_HI(net469));
 sg13g2_tiehi _11613__470 (.L_HI(net470));
 sg13g2_tiehi _11612__471 (.L_HI(net471));
 sg13g2_tiehi _11611__472 (.L_HI(net472));
 sg13g2_tiehi _11610__473 (.L_HI(net473));
 sg13g2_tiehi _11609__474 (.L_HI(net474));
 sg13g2_tiehi _11608__475 (.L_HI(net475));
 sg13g2_tiehi _11607__476 (.L_HI(net476));
 sg13g2_tiehi _11606__477 (.L_HI(net477));
 sg13g2_tiehi _11605__478 (.L_HI(net478));
 sg13g2_tiehi _11604__479 (.L_HI(net479));
 sg13g2_tiehi _11603__480 (.L_HI(net480));
 sg13g2_tiehi _11602__481 (.L_HI(net481));
 sg13g2_tiehi _11601__482 (.L_HI(net482));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_gregac_tiny_nn_18 (.L_LO(net18));
 sg13g2_tielo tt_um_gregac_tiny_nn_19 (.L_LO(net19));
 sg13g2_tielo tt_um_gregac_tiny_nn_20 (.L_LO(net20));
 sg13g2_tielo tt_um_gregac_tiny_nn_21 (.L_LO(net21));
 sg13g2_tielo tt_um_gregac_tiny_nn_22 (.L_LO(net22));
 sg13g2_tielo tt_um_gregac_tiny_nn_23 (.L_LO(net23));
 sg13g2_tielo tt_um_gregac_tiny_nn_24 (.L_LO(net24));
 sg13g2_tielo tt_um_gregac_tiny_nn_25 (.L_LO(net25));
 sg13g2_tielo tt_um_gregac_tiny_nn_26 (.L_LO(net26));
 sg13g2_tielo tt_um_gregac_tiny_nn_27 (.L_LO(net27));
 sg13g2_tielo tt_um_gregac_tiny_nn_28 (.L_LO(net28));
 sg13g2_tielo tt_um_gregac_tiny_nn_29 (.L_LO(net29));
 sg13g2_tielo tt_um_gregac_tiny_nn_30 (.L_LO(net30));
 sg13g2_tielo tt_um_gregac_tiny_nn_31 (.L_LO(net31));
 sg13g2_tielo tt_um_gregac_tiny_nn_32 (.L_LO(net32));
 sg13g2_tiehi _11600__33 (.L_HI(net33));
 sg13g2_buf_2 fanout1417 (.A(_04684_),
    .X(net1417));
 sg13g2_buf_2 fanout1418 (.A(_02320_),
    .X(net1418));
 sg13g2_buf_2 fanout1419 (.A(_05064_),
    .X(net1419));
 sg13g2_buf_2 fanout1420 (.A(_03750_),
    .X(net1420));
 sg13g2_buf_2 fanout1421 (.A(_03270_),
    .X(net1421));
 sg13g2_buf_2 fanout1422 (.A(_02298_),
    .X(net1422));
 sg13g2_buf_2 fanout1423 (.A(net1424),
    .X(net1423));
 sg13g2_buf_1 fanout1424 (.A(_01596_),
    .X(net1424));
 sg13g2_buf_2 fanout1425 (.A(net1426),
    .X(net1425));
 sg13g2_buf_2 fanout1426 (.A(_01596_),
    .X(net1426));
 sg13g2_buf_2 fanout1427 (.A(net1428),
    .X(net1427));
 sg13g2_buf_2 fanout1428 (.A(_01593_),
    .X(net1428));
 sg13g2_buf_2 fanout1429 (.A(_01561_),
    .X(net1429));
 sg13g2_buf_2 fanout1430 (.A(_01563_),
    .X(net1430));
 sg13g2_buf_2 fanout1431 (.A(_01560_),
    .X(net1431));
 sg13g2_buf_2 fanout1432 (.A(_01558_),
    .X(net1432));
 sg13g2_buf_1 fanout1433 (.A(_01558_),
    .X(net1433));
 sg13g2_buf_2 fanout1434 (.A(_01549_),
    .X(net1434));
 sg13g2_buf_2 fanout1435 (.A(_05058_),
    .X(net1435));
 sg13g2_buf_2 fanout1436 (.A(_05058_),
    .X(net1436));
 sg13g2_buf_2 fanout1437 (.A(_05057_),
    .X(net1437));
 sg13g2_buf_2 fanout1438 (.A(_05054_),
    .X(net1438));
 sg13g2_buf_1 fanout1439 (.A(_05054_),
    .X(net1439));
 sg13g2_buf_2 fanout1440 (.A(_05022_),
    .X(net1440));
 sg13g2_buf_1 fanout1441 (.A(_05022_),
    .X(net1441));
 sg13g2_buf_2 fanout1442 (.A(_05006_),
    .X(net1442));
 sg13g2_buf_2 fanout1443 (.A(net1444),
    .X(net1443));
 sg13g2_buf_2 fanout1444 (.A(_02293_),
    .X(net1444));
 sg13g2_buf_2 fanout1445 (.A(net1446),
    .X(net1445));
 sg13g2_buf_2 fanout1446 (.A(_02233_),
    .X(net1446));
 sg13g2_buf_2 fanout1447 (.A(net1448),
    .X(net1447));
 sg13g2_buf_2 fanout1448 (.A(_02233_),
    .X(net1448));
 sg13g2_buf_2 fanout1449 (.A(net1450),
    .X(net1449));
 sg13g2_buf_2 fanout1450 (.A(_01898_),
    .X(net1450));
 sg13g2_buf_2 fanout1451 (.A(net1452),
    .X(net1451));
 sg13g2_buf_2 fanout1452 (.A(_01897_),
    .X(net1452));
 sg13g2_buf_2 fanout1453 (.A(net1454),
    .X(net1453));
 sg13g2_buf_2 fanout1454 (.A(_05009_),
    .X(net1454));
 sg13g2_buf_2 fanout1455 (.A(_02248_),
    .X(net1455));
 sg13g2_buf_1 fanout1456 (.A(_02248_),
    .X(net1456));
 sg13g2_buf_2 fanout1457 (.A(_02245_),
    .X(net1457));
 sg13g2_buf_2 fanout1458 (.A(net1459),
    .X(net1458));
 sg13g2_buf_2 fanout1459 (.A(_02243_),
    .X(net1459));
 sg13g2_buf_2 fanout1460 (.A(net1461),
    .X(net1460));
 sg13g2_buf_2 fanout1461 (.A(_01945_),
    .X(net1461));
 sg13g2_buf_2 fanout1462 (.A(_01918_),
    .X(net1462));
 sg13g2_buf_2 fanout1463 (.A(_01498_),
    .X(net1463));
 sg13g2_buf_4 fanout1464 (.X(net1464),
    .A(_04201_));
 sg13g2_buf_2 fanout1465 (.A(net1466),
    .X(net1465));
 sg13g2_buf_1 fanout1466 (.A(_03715_),
    .X(net1466));
 sg13g2_buf_2 fanout1467 (.A(net1468),
    .X(net1467));
 sg13g2_buf_1 fanout1468 (.A(_03253_),
    .X(net1468));
 sg13g2_buf_2 fanout1469 (.A(_01922_),
    .X(net1469));
 sg13g2_buf_2 fanout1470 (.A(_02200_),
    .X(net1470));
 sg13g2_buf_2 fanout1471 (.A(_02826_),
    .X(net1471));
 sg13g2_buf_1 fanout1472 (.A(_02826_),
    .X(net1472));
 sg13g2_buf_2 fanout1473 (.A(net1474),
    .X(net1473));
 sg13g2_buf_2 fanout1474 (.A(_02826_),
    .X(net1474));
 sg13g2_buf_2 fanout1475 (.A(_02083_),
    .X(net1475));
 sg13g2_buf_2 fanout1476 (.A(_01359_),
    .X(net1476));
 sg13g2_buf_2 fanout1477 (.A(net1478),
    .X(net1477));
 sg13g2_buf_1 fanout1478 (.A(net1481),
    .X(net1478));
 sg13g2_buf_2 fanout1479 (.A(net1481),
    .X(net1479));
 sg13g2_buf_2 fanout1480 (.A(net1481),
    .X(net1480));
 sg13g2_buf_1 fanout1481 (.A(_00926_),
    .X(net1481));
 sg13g2_buf_4 fanout1482 (.X(net1482),
    .A(net1483));
 sg13g2_buf_4 fanout1483 (.X(net1483),
    .A(_04361_));
 sg13g2_buf_4 fanout1484 (.X(net1484),
    .A(_03917_));
 sg13g2_buf_4 fanout1485 (.X(net1485),
    .A(_03917_));
 sg13g2_buf_2 fanout1486 (.A(_01620_),
    .X(net1486));
 sg13g2_buf_2 fanout1487 (.A(net1489),
    .X(net1487));
 sg13g2_buf_2 fanout1488 (.A(net1489),
    .X(net1488));
 sg13g2_buf_2 fanout1489 (.A(_01619_),
    .X(net1489));
 sg13g2_buf_2 fanout1490 (.A(_01318_),
    .X(net1490));
 sg13g2_buf_2 fanout1491 (.A(net1492),
    .X(net1491));
 sg13g2_buf_2 fanout1492 (.A(_03440_),
    .X(net1492));
 sg13g2_buf_2 fanout1493 (.A(_02983_),
    .X(net1493));
 sg13g2_buf_2 fanout1494 (.A(_02983_),
    .X(net1494));
 sg13g2_buf_4 fanout1495 (.X(net1495),
    .A(_01315_));
 sg13g2_buf_2 fanout1496 (.A(_01315_),
    .X(net1496));
 sg13g2_buf_2 fanout1497 (.A(net1499),
    .X(net1497));
 sg13g2_buf_4 fanout1498 (.X(net1498),
    .A(net1499));
 sg13g2_buf_4 fanout1499 (.X(net1499),
    .A(_01314_));
 sg13g2_buf_2 fanout1500 (.A(net1501),
    .X(net1500));
 sg13g2_buf_1 fanout1501 (.A(_01264_),
    .X(net1501));
 sg13g2_buf_2 fanout1502 (.A(_02090_),
    .X(net1502));
 sg13g2_buf_2 fanout1503 (.A(_01067_),
    .X(net1503));
 sg13g2_buf_2 fanout1504 (.A(_01067_),
    .X(net1504));
 sg13g2_buf_2 fanout1505 (.A(_04813_),
    .X(net1505));
 sg13g2_buf_4 fanout1506 (.X(net1506),
    .A(_01736_));
 sg13g2_buf_2 fanout1507 (.A(net1508),
    .X(net1507));
 sg13g2_buf_2 fanout1508 (.A(net1509),
    .X(net1508));
 sg13g2_buf_1 fanout1509 (.A(net1511),
    .X(net1509));
 sg13g2_buf_2 fanout1510 (.A(net1511),
    .X(net1510));
 sg13g2_buf_1 fanout1511 (.A(net1512),
    .X(net1511));
 sg13g2_buf_2 fanout1512 (.A(_01189_),
    .X(net1512));
 sg13g2_buf_2 fanout1513 (.A(net1515),
    .X(net1513));
 sg13g2_buf_1 fanout1514 (.A(net1515),
    .X(net1514));
 sg13g2_buf_1 fanout1515 (.A(_05077_),
    .X(net1515));
 sg13g2_buf_2 fanout1516 (.A(_05077_),
    .X(net1516));
 sg13g2_buf_2 fanout1517 (.A(_05076_),
    .X(net1517));
 sg13g2_buf_4 fanout1518 (.X(net1518),
    .A(net1519));
 sg13g2_buf_2 fanout1519 (.A(net1521),
    .X(net1519));
 sg13g2_buf_2 fanout1520 (.A(net1521),
    .X(net1520));
 sg13g2_buf_2 fanout1521 (.A(_04792_),
    .X(net1521));
 sg13g2_buf_2 fanout1522 (.A(_02912_),
    .X(net1522));
 sg13g2_buf_1 fanout1523 (.A(_02912_),
    .X(net1523));
 sg13g2_buf_2 fanout1524 (.A(net1525),
    .X(net1524));
 sg13g2_buf_2 fanout1525 (.A(_02910_),
    .X(net1525));
 sg13g2_buf_2 fanout1526 (.A(_02081_),
    .X(net1526));
 sg13g2_buf_2 fanout1527 (.A(_02047_),
    .X(net1527));
 sg13g2_buf_4 fanout1528 (.X(net1528),
    .A(_02007_));
 sg13g2_buf_4 fanout1529 (.X(net1529),
    .A(_01366_));
 sg13g2_buf_2 fanout1530 (.A(net1531),
    .X(net1530));
 sg13g2_buf_2 fanout1531 (.A(_01182_),
    .X(net1531));
 sg13g2_buf_2 fanout1532 (.A(_04791_),
    .X(net1532));
 sg13g2_buf_2 fanout1533 (.A(_04770_),
    .X(net1533));
 sg13g2_buf_2 fanout1534 (.A(_04770_),
    .X(net1534));
 sg13g2_buf_2 fanout1535 (.A(_04762_),
    .X(net1535));
 sg13g2_buf_2 fanout1536 (.A(net1537),
    .X(net1536));
 sg13g2_buf_2 fanout1537 (.A(_03376_),
    .X(net1537));
 sg13g2_buf_2 fanout1538 (.A(net1539),
    .X(net1538));
 sg13g2_buf_2 fanout1539 (.A(_03375_),
    .X(net1539));
 sg13g2_buf_4 fanout1540 (.X(net1540),
    .A(net1542));
 sg13g2_buf_2 fanout1541 (.A(net1542),
    .X(net1541));
 sg13g2_buf_2 fanout1542 (.A(net1544),
    .X(net1542));
 sg13g2_buf_2 fanout1543 (.A(net1544),
    .X(net1543));
 sg13g2_buf_1 fanout1544 (.A(_02040_),
    .X(net1544));
 sg13g2_buf_2 fanout1545 (.A(_01968_),
    .X(net1545));
 sg13g2_buf_2 fanout1546 (.A(net1547),
    .X(net1546));
 sg13g2_buf_2 fanout1547 (.A(_01968_),
    .X(net1547));
 sg13g2_buf_2 fanout1548 (.A(_01967_),
    .X(net1548));
 sg13g2_buf_4 fanout1549 (.X(net1549),
    .A(_01689_));
 sg13g2_buf_2 fanout1550 (.A(_01689_),
    .X(net1550));
 sg13g2_buf_2 fanout1551 (.A(net1553),
    .X(net1551));
 sg13g2_buf_2 fanout1552 (.A(net1553),
    .X(net1552));
 sg13g2_buf_2 fanout1553 (.A(_01689_),
    .X(net1553));
 sg13g2_buf_4 fanout1554 (.X(net1554),
    .A(_01060_));
 sg13g2_buf_4 fanout1555 (.X(net1555),
    .A(_01022_));
 sg13g2_buf_2 fanout1556 (.A(_04345_),
    .X(net1556));
 sg13g2_buf_2 fanout1557 (.A(_04343_),
    .X(net1557));
 sg13g2_buf_2 fanout1558 (.A(_04342_),
    .X(net1558));
 sg13g2_buf_2 fanout1559 (.A(net1560),
    .X(net1559));
 sg13g2_buf_4 fanout1560 (.X(net1560),
    .A(_04341_));
 sg13g2_buf_4 fanout1561 (.X(net1561),
    .A(_04339_));
 sg13g2_buf_2 fanout1562 (.A(net1563),
    .X(net1562));
 sg13g2_buf_4 fanout1563 (.X(net1563),
    .A(_04338_));
 sg13g2_buf_2 fanout1564 (.A(net1565),
    .X(net1564));
 sg13g2_buf_4 fanout1565 (.X(net1565),
    .A(_04337_));
 sg13g2_buf_2 fanout1566 (.A(net1567),
    .X(net1566));
 sg13g2_buf_1 fanout1567 (.A(net1568),
    .X(net1567));
 sg13g2_buf_2 fanout1568 (.A(_04319_),
    .X(net1568));
 sg13g2_buf_2 fanout1569 (.A(_04318_),
    .X(net1569));
 sg13g2_buf_4 fanout1570 (.X(net1570),
    .A(_04315_));
 sg13g2_buf_2 fanout1571 (.A(_04313_),
    .X(net1571));
 sg13g2_buf_2 fanout1572 (.A(net1573),
    .X(net1572));
 sg13g2_buf_2 fanout1573 (.A(_04311_),
    .X(net1573));
 sg13g2_buf_4 fanout1574 (.X(net1574),
    .A(_04309_));
 sg13g2_buf_2 fanout1575 (.A(_03902_),
    .X(net1575));
 sg13g2_buf_2 fanout1576 (.A(_03901_),
    .X(net1576));
 sg13g2_buf_2 fanout1577 (.A(_03899_),
    .X(net1577));
 sg13g2_buf_1 fanout1578 (.A(_03899_),
    .X(net1578));
 sg13g2_buf_2 fanout1579 (.A(_03898_),
    .X(net1579));
 sg13g2_buf_2 fanout1580 (.A(_03898_),
    .X(net1580));
 sg13g2_buf_2 fanout1581 (.A(net1583),
    .X(net1581));
 sg13g2_buf_2 fanout1582 (.A(net1583),
    .X(net1582));
 sg13g2_buf_1 fanout1583 (.A(_03896_),
    .X(net1583));
 sg13g2_buf_2 fanout1584 (.A(_03895_),
    .X(net1584));
 sg13g2_buf_2 fanout1585 (.A(_03894_),
    .X(net1585));
 sg13g2_buf_1 fanout1586 (.A(_03894_),
    .X(net1586));
 sg13g2_buf_2 fanout1587 (.A(_03872_),
    .X(net1587));
 sg13g2_buf_2 fanout1588 (.A(net1589),
    .X(net1588));
 sg13g2_buf_2 fanout1589 (.A(_03868_),
    .X(net1589));
 sg13g2_buf_2 fanout1590 (.A(net1591),
    .X(net1590));
 sg13g2_buf_2 fanout1591 (.A(_03867_),
    .X(net1591));
 sg13g2_buf_2 fanout1592 (.A(net1593),
    .X(net1592));
 sg13g2_buf_2 fanout1593 (.A(_03866_),
    .X(net1593));
 sg13g2_buf_2 fanout1594 (.A(_03426_),
    .X(net1594));
 sg13g2_buf_2 fanout1595 (.A(_03426_),
    .X(net1595));
 sg13g2_buf_2 fanout1596 (.A(_03424_),
    .X(net1596));
 sg13g2_buf_2 fanout1597 (.A(_03423_),
    .X(net1597));
 sg13g2_buf_1 fanout1598 (.A(_03423_),
    .X(net1598));
 sg13g2_buf_2 fanout1599 (.A(_03422_),
    .X(net1599));
 sg13g2_buf_2 fanout1600 (.A(_03422_),
    .X(net1600));
 sg13g2_buf_2 fanout1601 (.A(_03421_),
    .X(net1601));
 sg13g2_buf_1 fanout1602 (.A(_03421_),
    .X(net1602));
 sg13g2_buf_2 fanout1603 (.A(_03420_),
    .X(net1603));
 sg13g2_buf_2 fanout1604 (.A(_03419_),
    .X(net1604));
 sg13g2_buf_1 fanout1605 (.A(_03419_),
    .X(net1605));
 sg13g2_buf_2 fanout1606 (.A(net1607),
    .X(net1606));
 sg13g2_buf_2 fanout1607 (.A(net1608),
    .X(net1607));
 sg13g2_buf_2 fanout1608 (.A(_03400_),
    .X(net1608));
 sg13g2_buf_2 fanout1609 (.A(_03399_),
    .X(net1609));
 sg13g2_buf_4 fanout1610 (.X(net1610),
    .A(_03398_));
 sg13g2_buf_1 fanout1611 (.A(_03398_),
    .X(net1611));
 sg13g2_buf_2 fanout1612 (.A(_03396_),
    .X(net1612));
 sg13g2_buf_2 fanout1613 (.A(_03393_),
    .X(net1613));
 sg13g2_buf_2 fanout1614 (.A(_03391_),
    .X(net1614));
 sg13g2_buf_2 fanout1615 (.A(_03391_),
    .X(net1615));
 sg13g2_buf_2 fanout1616 (.A(net1617),
    .X(net1616));
 sg13g2_buf_2 fanout1617 (.A(_03390_),
    .X(net1617));
 sg13g2_buf_2 fanout1618 (.A(net1619),
    .X(net1618));
 sg13g2_buf_2 fanout1619 (.A(net1620),
    .X(net1619));
 sg13g2_buf_2 fanout1620 (.A(_02955_),
    .X(net1620));
 sg13g2_buf_2 fanout1621 (.A(_02954_),
    .X(net1621));
 sg13g2_buf_2 fanout1622 (.A(_02952_),
    .X(net1622));
 sg13g2_buf_1 fanout1623 (.A(_02952_),
    .X(net1623));
 sg13g2_buf_2 fanout1624 (.A(_02950_),
    .X(net1624));
 sg13g2_buf_2 fanout1625 (.A(net1626),
    .X(net1625));
 sg13g2_buf_2 fanout1626 (.A(_02948_),
    .X(net1626));
 sg13g2_buf_2 fanout1627 (.A(_02943_),
    .X(net1627));
 sg13g2_buf_1 fanout1628 (.A(_02943_),
    .X(net1628));
 sg13g2_buf_2 fanout1629 (.A(_02925_),
    .X(net1629));
 sg13g2_buf_2 fanout1630 (.A(_02925_),
    .X(net1630));
 sg13g2_buf_2 fanout1631 (.A(_02923_),
    .X(net1631));
 sg13g2_buf_2 fanout1632 (.A(_02923_),
    .X(net1632));
 sg13g2_buf_2 fanout1633 (.A(_02922_),
    .X(net1633));
 sg13g2_buf_2 fanout1634 (.A(_02922_),
    .X(net1634));
 sg13g2_buf_2 fanout1635 (.A(net1636),
    .X(net1635));
 sg13g2_buf_2 fanout1636 (.A(_02921_),
    .X(net1636));
 sg13g2_buf_2 fanout1637 (.A(net1639),
    .X(net1637));
 sg13g2_buf_1 fanout1638 (.A(net1639),
    .X(net1638));
 sg13g2_buf_2 fanout1639 (.A(_02919_),
    .X(net1639));
 sg13g2_buf_2 fanout1640 (.A(net1641),
    .X(net1640));
 sg13g2_buf_2 fanout1641 (.A(_02918_),
    .X(net1641));
 sg13g2_buf_2 fanout1642 (.A(net1643),
    .X(net1642));
 sg13g2_buf_2 fanout1643 (.A(_02916_),
    .X(net1643));
 sg13g2_buf_2 fanout1644 (.A(net1645),
    .X(net1644));
 sg13g2_buf_1 fanout1645 (.A(net1650),
    .X(net1645));
 sg13g2_buf_2 fanout1646 (.A(net1648),
    .X(net1646));
 sg13g2_buf_2 fanout1647 (.A(net1648),
    .X(net1647));
 sg13g2_buf_1 fanout1648 (.A(net1649),
    .X(net1648));
 sg13g2_buf_1 fanout1649 (.A(_02909_),
    .X(net1649));
 sg13g2_buf_4 fanout1650 (.X(net1650),
    .A(_02909_));
 sg13g2_buf_2 fanout1651 (.A(net1652),
    .X(net1651));
 sg13g2_buf_2 fanout1652 (.A(net1653),
    .X(net1652));
 sg13g2_buf_2 fanout1653 (.A(_02900_),
    .X(net1653));
 sg13g2_buf_2 fanout1654 (.A(net1657),
    .X(net1654));
 sg13g2_buf_2 fanout1655 (.A(net1657),
    .X(net1655));
 sg13g2_buf_1 fanout1656 (.A(net1657),
    .X(net1656));
 sg13g2_buf_2 fanout1657 (.A(net1658),
    .X(net1657));
 sg13g2_buf_2 fanout1658 (.A(_02884_),
    .X(net1658));
 sg13g2_buf_2 fanout1659 (.A(net1660),
    .X(net1659));
 sg13g2_buf_2 fanout1660 (.A(net1663),
    .X(net1660));
 sg13g2_buf_2 fanout1661 (.A(net1663),
    .X(net1661));
 sg13g2_buf_2 fanout1662 (.A(net1663),
    .X(net1662));
 sg13g2_buf_2 fanout1663 (.A(_02870_),
    .X(net1663));
 sg13g2_buf_2 fanout1664 (.A(net1665),
    .X(net1664));
 sg13g2_buf_1 fanout1665 (.A(net1666),
    .X(net1665));
 sg13g2_buf_2 fanout1666 (.A(_02305_),
    .X(net1666));
 sg13g2_buf_2 fanout1667 (.A(_01688_),
    .X(net1667));
 sg13g2_buf_2 fanout1668 (.A(_01648_),
    .X(net1668));
 sg13g2_buf_2 fanout1669 (.A(net1670),
    .X(net1669));
 sg13g2_buf_2 fanout1670 (.A(_01270_),
    .X(net1670));
 sg13g2_buf_2 fanout1671 (.A(net1673),
    .X(net1671));
 sg13g2_buf_2 fanout1672 (.A(net1673),
    .X(net1672));
 sg13g2_buf_2 fanout1673 (.A(_01208_),
    .X(net1673));
 sg13g2_buf_2 fanout1674 (.A(_01188_),
    .X(net1674));
 sg13g2_buf_1 fanout1675 (.A(_01188_),
    .X(net1675));
 sg13g2_buf_4 fanout1676 (.X(net1676),
    .A(net1679));
 sg13g2_buf_2 fanout1677 (.A(net1678),
    .X(net1677));
 sg13g2_buf_4 fanout1678 (.X(net1678),
    .A(net1679));
 sg13g2_buf_2 fanout1679 (.A(net1681),
    .X(net1679));
 sg13g2_buf_4 fanout1680 (.X(net1680),
    .A(net1681));
 sg13g2_buf_2 fanout1681 (.A(_05284_),
    .X(net1681));
 sg13g2_buf_4 fanout1682 (.X(net1682),
    .A(net1684));
 sg13g2_buf_2 fanout1683 (.A(net1684),
    .X(net1683));
 sg13g2_buf_4 fanout1684 (.X(net1684),
    .A(_05284_));
 sg13g2_buf_4 fanout1685 (.X(net1685),
    .A(net1688));
 sg13g2_buf_1 fanout1686 (.A(net1688),
    .X(net1686));
 sg13g2_buf_4 fanout1687 (.X(net1687),
    .A(net1688));
 sg13g2_buf_2 fanout1688 (.A(_05284_),
    .X(net1688));
 sg13g2_buf_4 fanout1689 (.X(net1689),
    .A(net1691));
 sg13g2_buf_2 fanout1690 (.A(net1691),
    .X(net1690));
 sg13g2_buf_2 fanout1691 (.A(net1699),
    .X(net1691));
 sg13g2_buf_4 fanout1692 (.X(net1692),
    .A(net1699));
 sg13g2_buf_1 fanout1693 (.A(net1699),
    .X(net1693));
 sg13g2_buf_4 fanout1694 (.X(net1694),
    .A(net1698));
 sg13g2_buf_2 fanout1695 (.A(net1698),
    .X(net1695));
 sg13g2_buf_4 fanout1696 (.X(net1696),
    .A(net1697));
 sg13g2_buf_4 fanout1697 (.X(net1697),
    .A(net1698));
 sg13g2_buf_2 fanout1698 (.A(net1699),
    .X(net1698));
 sg13g2_buf_2 fanout1699 (.A(net1716),
    .X(net1699));
 sg13g2_buf_4 fanout1700 (.X(net1700),
    .A(net1705));
 sg13g2_buf_2 fanout1701 (.A(net1705),
    .X(net1701));
 sg13g2_buf_4 fanout1702 (.X(net1702),
    .A(net1705));
 sg13g2_buf_4 fanout1703 (.X(net1703),
    .A(net1705));
 sg13g2_buf_2 fanout1704 (.A(net1705),
    .X(net1704));
 sg13g2_buf_2 fanout1705 (.A(net1716),
    .X(net1705));
 sg13g2_buf_4 fanout1706 (.X(net1706),
    .A(net1708));
 sg13g2_buf_2 fanout1707 (.A(net1708),
    .X(net1707));
 sg13g2_buf_2 fanout1708 (.A(net1714),
    .X(net1708));
 sg13g2_buf_4 fanout1709 (.X(net1709),
    .A(net1711));
 sg13g2_buf_4 fanout1710 (.X(net1710),
    .A(net1711));
 sg13g2_buf_2 fanout1711 (.A(net1714),
    .X(net1711));
 sg13g2_buf_4 fanout1712 (.X(net1712),
    .A(net1713));
 sg13g2_buf_4 fanout1713 (.X(net1713),
    .A(net1714));
 sg13g2_buf_2 fanout1714 (.A(net1716),
    .X(net1714));
 sg13g2_buf_4 fanout1715 (.X(net1715),
    .A(net1716));
 sg13g2_buf_4 fanout1716 (.X(net1716),
    .A(_02914_));
 sg13g2_buf_4 fanout1717 (.X(net1717),
    .A(net1718));
 sg13g2_buf_4 fanout1718 (.X(net1718),
    .A(_02816_));
 sg13g2_buf_2 fanout1719 (.A(net1721),
    .X(net1719));
 sg13g2_buf_1 fanout1720 (.A(net1721),
    .X(net1720));
 sg13g2_buf_2 fanout1721 (.A(_02239_),
    .X(net1721));
 sg13g2_buf_2 fanout1722 (.A(net1723),
    .X(net1722));
 sg13g2_buf_2 fanout1723 (.A(_01955_),
    .X(net1723));
 sg13g2_buf_2 fanout1724 (.A(net1725),
    .X(net1724));
 sg13g2_buf_2 fanout1725 (.A(net1726),
    .X(net1725));
 sg13g2_buf_2 fanout1726 (.A(_00928_),
    .X(net1726));
 sg13g2_buf_2 fanout1727 (.A(net1728),
    .X(net1727));
 sg13g2_buf_2 fanout1728 (.A(net1729),
    .X(net1728));
 sg13g2_buf_2 fanout1729 (.A(_00828_),
    .X(net1729));
 sg13g2_buf_2 fanout1730 (.A(_00823_),
    .X(net1730));
 sg13g2_buf_2 fanout1731 (.A(_04772_),
    .X(net1731));
 sg13g2_buf_2 fanout1732 (.A(net1733),
    .X(net1732));
 sg13g2_buf_2 fanout1733 (.A(_04738_),
    .X(net1733));
 sg13g2_buf_2 fanout1734 (.A(_04737_),
    .X(net1734));
 sg13g2_buf_2 fanout1735 (.A(_04737_),
    .X(net1735));
 sg13g2_buf_4 fanout1736 (.X(net1736),
    .A(_00783_));
 sg13g2_buf_1 fanout1737 (.A(_00783_),
    .X(net1737));
 sg13g2_buf_2 fanout1738 (.A(net1739),
    .X(net1738));
 sg13g2_buf_2 fanout1739 (.A(net1740),
    .X(net1739));
 sg13g2_buf_2 fanout1740 (.A(_00782_),
    .X(net1740));
 sg13g2_buf_2 fanout1741 (.A(net1742),
    .X(net1741));
 sg13g2_buf_4 fanout1742 (.X(net1742),
    .A(_04864_));
 sg13g2_buf_2 fanout1743 (.A(net1745),
    .X(net1743));
 sg13g2_buf_4 fanout1744 (.X(net1744),
    .A(_04736_));
 sg13g2_buf_1 fanout1745 (.A(_04736_),
    .X(net1745));
 sg13g2_buf_4 fanout1746 (.X(net1746),
    .A(_02036_));
 sg13g2_buf_1 fanout1747 (.A(_02036_),
    .X(net1747));
 sg13g2_buf_4 fanout1748 (.X(net1748),
    .A(net1749));
 sg13g2_buf_1 fanout1749 (.A(_01676_),
    .X(net1749));
 sg13g2_buf_4 fanout1750 (.X(net1750),
    .A(net1751));
 sg13g2_buf_4 fanout1751 (.X(net1751),
    .A(net1756));
 sg13g2_buf_4 fanout1752 (.X(net1752),
    .A(net1756));
 sg13g2_buf_2 fanout1753 (.A(net1754),
    .X(net1753));
 sg13g2_buf_4 fanout1754 (.X(net1754),
    .A(net1755));
 sg13g2_buf_2 fanout1755 (.A(net1756),
    .X(net1755));
 sg13g2_buf_2 fanout1756 (.A(net1760),
    .X(net1756));
 sg13g2_buf_4 fanout1757 (.X(net1757),
    .A(net1760));
 sg13g2_buf_4 fanout1758 (.X(net1758),
    .A(net1759));
 sg13g2_buf_2 fanout1759 (.A(net1760),
    .X(net1759));
 sg13g2_buf_4 fanout1760 (.X(net1760),
    .A(_01184_));
 sg13g2_buf_4 fanout1761 (.X(net1761),
    .A(_01184_));
 sg13g2_buf_4 fanout1762 (.X(net1762),
    .A(_01184_));
 sg13g2_buf_4 fanout1763 (.X(net1763),
    .A(_00825_));
 sg13g2_buf_4 fanout1764 (.X(net1764),
    .A(_00788_));
 sg13g2_buf_4 fanout1765 (.X(net1765),
    .A(net1766));
 sg13g2_buf_4 fanout1766 (.X(net1766),
    .A(_00787_));
 sg13g2_buf_2 fanout1767 (.A(net1768),
    .X(net1767));
 sg13g2_buf_4 fanout1768 (.X(net1768),
    .A(_00661_));
 sg13g2_buf_8 fanout1769 (.A(_00646_),
    .X(net1769));
 sg13g2_buf_4 fanout1770 (.X(net1770),
    .A(_00646_));
 sg13g2_buf_8 fanout1771 (.A(_00645_),
    .X(net1771));
 sg13g2_buf_4 fanout1772 (.X(net1772),
    .A(_00645_));
 sg13g2_buf_4 fanout1773 (.X(net1773),
    .A(_00643_));
 sg13g2_buf_4 fanout1774 (.X(net1774),
    .A(_00643_));
 sg13g2_buf_4 fanout1775 (.X(net1775),
    .A(_00642_));
 sg13g2_buf_2 fanout1776 (.A(_00642_),
    .X(net1776));
 sg13g2_buf_4 fanout1777 (.X(net1777),
    .A(_00641_));
 sg13g2_buf_4 fanout1778 (.X(net1778),
    .A(_00641_));
 sg13g2_buf_8 fanout1779 (.A(_00640_),
    .X(net1779));
 sg13g2_buf_4 fanout1780 (.X(net1780),
    .A(_00640_));
 sg13g2_buf_4 fanout1781 (.X(net1781),
    .A(net1782));
 sg13g2_buf_4 fanout1782 (.X(net1782),
    .A(_00639_));
 sg13g2_buf_4 fanout1783 (.X(net1783),
    .A(_00638_));
 sg13g2_buf_4 fanout1784 (.X(net1784),
    .A(_00638_));
 sg13g2_buf_4 fanout1785 (.X(net1785),
    .A(net1056));
 sg13g2_buf_2 fanout1786 (.A(net1110),
    .X(net1786));
 sg13g2_buf_4 fanout1787 (.X(net1787),
    .A(net1051));
 sg13g2_buf_2 fanout1788 (.A(\u_tiny_nn_top.state_q[13] ),
    .X(net1788));
 sg13g2_buf_2 fanout1789 (.A(\u_tiny_nn_top.core_mul_add_op_b_en ),
    .X(net1789));
 sg13g2_buf_2 fanout1790 (.A(\u_tiny_nn_top.core_mul_add_op_b_en ),
    .X(net1790));
 sg13g2_buf_4 fanout1791 (.X(net1791),
    .A(\u_tiny_nn_top.state_q[1] ));
 sg13g2_buf_2 fanout1792 (.A(\u_tiny_nn_top.state_q[1] ),
    .X(net1792));
 sg13g2_buf_2 fanout1793 (.A(net1098),
    .X(net1793));
 sg13g2_buf_2 fanout1794 (.A(net1796),
    .X(net1794));
 sg13g2_buf_2 fanout1795 (.A(net1796),
    .X(net1795));
 sg13g2_buf_2 fanout1796 (.A(net1797),
    .X(net1796));
 sg13g2_buf_2 fanout1797 (.A(\u_tiny_nn_top.param_write_q[7] ),
    .X(net1797));
 sg13g2_buf_2 fanout1798 (.A(net1799),
    .X(net1798));
 sg13g2_buf_2 fanout1799 (.A(net1800),
    .X(net1799));
 sg13g2_buf_4 fanout1800 (.X(net1800),
    .A(net1801));
 sg13g2_buf_4 fanout1801 (.X(net1801),
    .A(net1061));
 sg13g2_buf_4 fanout1802 (.X(net1802),
    .A(net1803));
 sg13g2_buf_2 fanout1803 (.A(net1805),
    .X(net1803));
 sg13g2_buf_4 fanout1804 (.X(net1804),
    .A(\u_tiny_nn_top.param_write_q[4] ));
 sg13g2_buf_1 fanout1805 (.A(\u_tiny_nn_top.param_write_q[4] ),
    .X(net1805));
 sg13g2_buf_4 fanout1806 (.X(net1806),
    .A(\u_tiny_nn_top.param_write_q[3] ));
 sg13g2_buf_2 fanout1807 (.A(net1809),
    .X(net1807));
 sg13g2_buf_2 fanout1808 (.A(net1809),
    .X(net1808));
 sg13g2_buf_2 fanout1809 (.A(net1113),
    .X(net1809));
 sg13g2_buf_4 fanout1810 (.X(net1810),
    .A(net1811));
 sg13g2_buf_2 fanout1811 (.A(\u_tiny_nn_top.param_write_q[2] ),
    .X(net1811));
 sg13g2_buf_4 fanout1812 (.X(net1812),
    .A(net1813));
 sg13g2_buf_2 fanout1813 (.A(net1091),
    .X(net1813));
 sg13g2_buf_4 fanout1814 (.X(net1814),
    .A(net1816));
 sg13g2_buf_2 fanout1815 (.A(net1816),
    .X(net1815));
 sg13g2_buf_2 fanout1816 (.A(\u_tiny_nn_top.param_write_q[1] ),
    .X(net1816));
 sg13g2_buf_4 fanout1817 (.X(net1817),
    .A(net1818));
 sg13g2_buf_2 fanout1818 (.A(\u_tiny_nn_top.param_write_q[1] ),
    .X(net1818));
 sg13g2_buf_4 fanout1819 (.X(net1819),
    .A(net1820));
 sg13g2_buf_2 fanout1820 (.A(net1821),
    .X(net1820));
 sg13g2_buf_2 fanout1821 (.A(net1822),
    .X(net1821));
 sg13g2_buf_4 fanout1822 (.X(net1822),
    .A(net1026));
 sg13g2_buf_4 fanout1823 (.X(net1823),
    .A(net1825));
 sg13g2_buf_2 fanout1824 (.A(net1825),
    .X(net1824));
 sg13g2_buf_4 fanout1825 (.X(net1825),
    .A(net1826));
 sg13g2_buf_4 fanout1826 (.X(net1826),
    .A(\u_tiny_nn_top.data_i_q[15] ));
 sg13g2_buf_4 fanout1827 (.X(net1827),
    .A(net750));
 sg13g2_buf_4 fanout1828 (.X(net1828),
    .A(net1088));
 sg13g2_buf_2 fanout1829 (.A(\u_tiny_nn_top.data_i_q[12] ),
    .X(net1829));
 sg13g2_buf_4 fanout1830 (.X(net1830),
    .A(net1831));
 sg13g2_buf_4 fanout1831 (.X(net1831),
    .A(net1832));
 sg13g2_buf_4 fanout1832 (.X(net1832),
    .A(net779));
 sg13g2_buf_2 fanout1833 (.A(net1834),
    .X(net1833));
 sg13g2_buf_2 fanout1834 (.A(net1835),
    .X(net1834));
 sg13g2_buf_4 fanout1835 (.X(net1835),
    .A(net1836));
 sg13g2_buf_8 fanout1836 (.A(\u_tiny_nn_top.data_i_q[7] ),
    .X(net1836));
 sg13g2_buf_4 fanout1837 (.X(net1837),
    .A(net1838));
 sg13g2_buf_4 fanout1838 (.X(net1838),
    .A(net1839));
 sg13g2_buf_8 fanout1839 (.A(\u_tiny_nn_top.data_i_q[6] ),
    .X(net1839));
 sg13g2_buf_4 fanout1840 (.X(net1840),
    .A(net1842));
 sg13g2_buf_2 fanout1841 (.A(net1842),
    .X(net1841));
 sg13g2_buf_8 fanout1842 (.A(\u_tiny_nn_top.data_i_q[5] ),
    .X(net1842));
 sg13g2_buf_4 fanout1843 (.X(net1843),
    .A(net1845));
 sg13g2_buf_2 fanout1844 (.A(net1845),
    .X(net1844));
 sg13g2_buf_8 fanout1845 (.A(\u_tiny_nn_top.data_i_q[4] ),
    .X(net1845));
 sg13g2_buf_8 fanout1846 (.A(net1848),
    .X(net1846));
 sg13g2_buf_2 fanout1847 (.A(net1848),
    .X(net1847));
 sg13g2_buf_8 fanout1848 (.A(\u_tiny_nn_top.data_i_q[3] ),
    .X(net1848));
 sg13g2_buf_4 fanout1849 (.X(net1849),
    .A(net1850));
 sg13g2_buf_8 fanout1850 (.A(net1851),
    .X(net1850));
 sg13g2_buf_8 fanout1851 (.A(\u_tiny_nn_top.data_i_q[1] ),
    .X(net1851));
 sg13g2_buf_2 fanout1852 (.A(net1853),
    .X(net1852));
 sg13g2_buf_2 fanout1853 (.A(net1854),
    .X(net1853));
 sg13g2_buf_2 fanout1854 (.A(\u_tiny_nn_top.phase_q ),
    .X(net1854));
 sg13g2_buf_4 fanout1855 (.X(net1855),
    .A(\u_tiny_nn_top.counter_q[1] ));
 sg13g2_buf_2 fanout1856 (.A(net1080),
    .X(net1856));
 sg13g2_buf_2 fanout1857 (.A(net1861),
    .X(net1857));
 sg13g2_buf_2 fanout1858 (.A(net1860),
    .X(net1858));
 sg13g2_buf_1 fanout1859 (.A(net1860),
    .X(net1859));
 sg13g2_buf_2 fanout1860 (.A(net1861),
    .X(net1860));
 sg13g2_buf_2 fanout1861 (.A(\u_tiny_nn_top.counter_q[0] ),
    .X(net1861));
 sg13g2_buf_2 fanout1862 (.A(net1863),
    .X(net1862));
 sg13g2_buf_2 fanout1863 (.A(net1865),
    .X(net1863));
 sg13g2_buf_4 fanout1864 (.X(net1864),
    .A(net1865));
 sg13g2_buf_2 fanout1865 (.A(net1059),
    .X(net1865));
 sg13g2_buf_4 fanout1866 (.X(net1866),
    .A(net1868));
 sg13g2_buf_4 fanout1867 (.X(net1867),
    .A(net1868));
 sg13g2_buf_2 fanout1868 (.A(rst_n),
    .X(net1868));
 sg13g2_buf_4 fanout1869 (.X(net1869),
    .A(net1870));
 sg13g2_buf_4 fanout1870 (.X(net1870),
    .A(net1872));
 sg13g2_buf_4 fanout1871 (.X(net1871),
    .A(net1872));
 sg13g2_buf_2 fanout1872 (.A(rst_n),
    .X(net1872));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_tielo tt_um_gregac_tiny_nn_17 (.L_LO(net17));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_4_8_0_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_4_9_0_clk));
 sg13g2_buf_1 clkload9 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_11_0_clk));
 sg13g2_buf_1 clkload11 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_13_0_clk));
 sg13g2_buf_1 clkload13 (.A(clknet_4_14_0_clk));
 sg13g2_buf_2 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_inv_8 clkload15 (.A(clknet_leaf_1_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_3_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_66_clk));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_8_clk));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_6_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_15_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_18_clk));
 sg13g2_inv_8 clkload22 (.A(clknet_leaf_20_clk));
 sg13g2_inv_4 clkload23 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload25 (.A(clknet_leaf_21_clk));
 sg13g2_inv_4 clkload26 (.A(clknet_leaf_13_clk));
 sg13g2_inv_1 clkload27 (.A(clknet_leaf_30_clk));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_50_clk));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_53_clk));
 sg13g2_inv_2 clkload30 (.A(clknet_leaf_56_clk));
 sg13g2_inv_8 clkload31 (.A(clknet_leaf_57_clk));
 sg13g2_inv_1 clkload32 (.A(clknet_leaf_49_clk));
 sg13g2_inv_4 clkload33 (.A(clknet_leaf_31_clk));
 sg13g2_inv_8 clkload34 (.A(clknet_leaf_33_clk));
 sg13g2_inv_4 clkload35 (.A(clknet_leaf_42_clk));
 sg13g2_inv_4 clkload36 (.A(clknet_leaf_43_clk));
 sg13g2_inv_4 clkload37 (.A(clknet_leaf_46_clk));
 sg13g2_inv_4 clkload38 (.A(clknet_leaf_47_clk));
 sg13g2_inv_4 clkload39 (.A(clknet_leaf_37_clk));
 sg13g2_inv_4 clkload40 (.A(clknet_leaf_40_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][11] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold2 (.A(_00441_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold3 (.A(_00165_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold4 (.A(_00007_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold5 (.A(_00167_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold6 (.A(_00015_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold7 (.A(_00164_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold8 (.A(_00008_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold9 (.A(_00169_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold10 (.A(_00206_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold11 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][10] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold12 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][13] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold13 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][14] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold14 (.A(_00572_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold15 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][2] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold16 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][9] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold17 (.A(_00551_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold18 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][13] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold19 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][2] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold20 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][12] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold21 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][14] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold22 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][0] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold23 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][13] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold24 (.A(_05316_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold25 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][2] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold26 (.A(_05267_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold27 (.A(_00480_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold28 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][14] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold29 (.A(_05317_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold30 (.A(_00620_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold31 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][12] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold32 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][2] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][5] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold34 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][2] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold35 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][4] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold36 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][12] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold37 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][4] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold38 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][11] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold39 (.A(\u_tiny_nn_top.state_q[2] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold40 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][11] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold41 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][4] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold42 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][0] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold43 (.A(_05301_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold44 (.A(_00574_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold45 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][5] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold46 (.A(_00483_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold47 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][4] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold48 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][0] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold49 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][2] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold50 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][1] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold51 (.A(_00255_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold52 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][9] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold53 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][3] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold54 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][4] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold55 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][5] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold56 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][12] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold57 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][4] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold58 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][3] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold59 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][4] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold60 (.A(_00482_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold61 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][1] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold62 (.A(_00607_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold63 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][0] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold64 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][5] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold65 (.A(_00611_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold66 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][1] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold67 (.A(_00479_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold68 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][5] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold69 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][5] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold70 (.A(_00579_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold71 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][4] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold72 (.A(_00578_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold73 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][1] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold74 (.A(_00511_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold75 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][5] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold76 (.A(_00627_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold77 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][3] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold78 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[1][0] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold79 (.A(_00494_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold80 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][2] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold81 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][5] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold82 (.A(_00547_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold83 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][3] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold84 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][12] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold85 (.A(_00634_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold86 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][10] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold87 (.A(_00584_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold88 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][7] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold89 (.A(_00629_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold90 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][6] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold91 (.A(_00628_),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold92 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][6] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold93 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][15] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold94 (.A(_00621_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold95 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][12] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold96 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][9] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold97 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][13] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold98 (.A(_00635_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold99 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][6] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold100 (.A(_00580_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold101 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][8] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold102 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][3] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold103 (.A(_00609_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold104 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][14] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold105 (.A(_05308_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold106 (.A(_00588_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold107 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][14] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold108 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][11] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold109 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][1] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold110 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][3] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold111 (.A(_00625_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold112 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][6] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold113 (.A(_00260_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold114 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][9] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold115 (.A(_05312_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold116 (.A(_00615_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold117 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][14] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold118 (.A(_02866_),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold119 (.A(_00268_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold120 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][14] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold121 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][12] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold122 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][9] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold123 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][13] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold124 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][12] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold125 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][10] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold126 (.A(_00632_),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold127 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][2] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold128 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][3] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold129 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][11] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold130 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][11] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold131 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][8] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold132 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][15] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold133 (.A(_00637_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold134 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][9] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold135 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][10] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold136 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][9] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold137 (.A(_00631_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold138 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][5] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold139 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][6] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold140 (.A(_00612_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold141 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][8] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold142 (.A(_00614_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold143 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][2] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold144 (.A(_00624_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold145 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][13] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold146 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][10] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold147 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][9] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold148 (.A(_05268_),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold149 (.A(_00487_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold150 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][8] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold151 (.A(_00630_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold152 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][9] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold153 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][15] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold154 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][15] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold155 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][7] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold156 (.A(_00613_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold157 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][15] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold158 (.A(_00269_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold159 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][11] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold160 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][1] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold161 (.A(_00623_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold162 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][14] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold163 (.A(_00636_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold164 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][13] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold165 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][13] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold166 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][8] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold167 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][10] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold168 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][10] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold169 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][12] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold170 (.A(\u_tiny_nn_top.u_core.param_val_op_q[2][10] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold171 (.A(_05313_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold172 (.A(_00616_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold173 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][8] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold174 (.A(_02860_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold175 (.A(_00262_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold176 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][0] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold177 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][0] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold178 (.A(_05266_),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold179 (.A(_00478_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold180 (.A(\u_tiny_nn_top.u_core.param_val_op_q[6][7] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold181 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][11] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold182 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][3] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold183 (.A(_00257_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold184 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][13] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold185 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][12] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold186 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][0] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold187 (.A(_00622_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold188 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][0] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold189 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][14] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold190 (.A(_05256_),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold191 (.A(_00428_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold192 (.A(\u_tiny_nn_top.state_q[9] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold193 (.A(_00231_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold194 (.A(_00162_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold195 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[3][13] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold196 (.A(_00507_),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold197 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][9] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold198 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][10] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold199 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][6] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold200 (.A(_00516_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold201 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][11] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold202 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][0] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold203 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][15] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold204 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][11] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold205 (.A(_00633_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold206 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][0] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold207 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][6] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold208 (.A(_00484_),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold209 (.A(\u_tiny_nn_top.core_accumulate_result[2] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold210 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][3] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold211 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][8] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold212 (.A(_00566_),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold213 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][0] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold214 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][4] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold215 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][7] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold216 (.A(_00485_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold217 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][8] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold218 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][14] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold219 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][13] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold220 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][8] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold221 (.A(_00486_),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold222 (.A(\u_tiny_nn_top.max_val_skid_q[0] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold223 (.A(_00207_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold224 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[0][4] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold225 (.A(_00626_),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold226 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][7] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold227 (.A(_00421_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold228 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][8] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold229 (.A(_00518_),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold230 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][1] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold231 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][14] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold232 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][13] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold233 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][15] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold234 (.A(_00493_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold235 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][1] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold236 (.A(_00575_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold237 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][1] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold238 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][6] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold239 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][7] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold240 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][10] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold241 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][8] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold242 (.A(_00454_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold243 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][10] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold244 (.A(_05278_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold245 (.A(_00520_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold246 (.A(\u_tiny_nn_top.u_core.param_val_op_q[4][2] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold247 (.A(_05302_),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold248 (.A(_00576_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold249 (.A(\u_tiny_nn_top.u_core.param_val_op_q[3][3] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold250 (.A(_00481_),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold251 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][1] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold252 (.A(\u_tiny_nn_top.core_accumulate_result[14] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold253 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][6] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold254 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][14] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold255 (.A(_05282_),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold256 (.A(_00524_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold257 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][15] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold258 (.A(_00573_),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold259 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][5] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold260 (.A(_00595_),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold261 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][9] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold262 (.A(_00599_),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold263 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][12] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold264 (.A(_00602_),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold265 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][9] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold266 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][2] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold267 (.A(_00592_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold268 (.A(\u_tiny_nn_top.data_i_q[14] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold269 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][7] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold270 (.A(_00597_),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold271 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][9] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold272 (.A(_00567_),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold273 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][15] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold274 (.A(_00525_),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold275 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][10] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold276 (.A(_00568_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold277 (.A(\u_tiny_nn_top.start_count_q[4] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold278 (.A(\u_tiny_nn_top.start_count_q[2] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold279 (.A(\u_tiny_nn_top.start_count_q[5] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold280 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][12] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold281 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][6] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold282 (.A(\u_tiny_nn_top.u_core.param_val_op_q[7][15] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold283 (.A(_00429_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold284 (.A(\u_tiny_nn_top.u_core.param_val_op_q[0][7] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold285 (.A(_00261_),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold286 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][5] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold287 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][4] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold288 (.A(_00594_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold289 (.A(\u_tiny_nn_top.core_accumulate_result[12] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold290 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][12] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold291 (.A(\u_tiny_nn_top.max_val_skid_q[5] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold292 (.A(_00212_),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold293 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][3] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold294 (.A(_00561_),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold295 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][13] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold296 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][0] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold297 (.A(\u_tiny_nn_top.data_i_q[8] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold298 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][4] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold299 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][7] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold300 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][5] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold301 (.A(_00563_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold302 (.A(\u_tiny_nn_top.start_count_q[1] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold303 (.A(_00191_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold304 (.A(\u_tiny_nn_top.core_accumulate_result[8] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold305 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][14] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold306 (.A(_00604_),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold307 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][13] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold308 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][11] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold309 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][12] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold310 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][9] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold311 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][3] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold312 (.A(\u_tiny_nn_top.core_accumulate_result[5] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold313 (.A(\u_tiny_nn_top.core_accumulate_result[9] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold314 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][4] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold315 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][6] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold316 (.A(\u_tiny_nn_top.core_accumulate_result[7] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold317 (.A(\u_tiny_nn_top.start_count_q[6] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold318 (.A(_00196_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold319 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][6] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold320 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][3] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold321 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][3] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold322 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][10] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold323 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][4] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold324 (.A(_00166_),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold325 (.A(_00004_),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold326 (.A(\u_tiny_nn_top.start_count_q[7] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold327 (.A(_00197_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold328 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][5] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold329 (.A(\u_tiny_nn_top.core_accumulate_result[11] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold330 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][10] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold331 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][6] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold332 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][5] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold333 (.A(\u_tiny_nn_top.core_accumulate_result[3] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold334 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][15] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold335 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[1][8] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold336 (.A(_00502_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold337 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][2] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold338 (.A(\u_tiny_nn_top.core_accumulate_result[0] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold339 (.A(\u_tiny_nn_top.u_core.param_val_op_q[5][7] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold340 (.A(_00453_),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold341 (.A(\u_tiny_nn_top.core_accumulate_result[1] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold342 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][2] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold343 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[1][11] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold344 (.A(_00505_),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold345 (.A(\u_tiny_nn_top.start_count_q[3] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold346 (.A(_00193_),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold347 (.A(\u_tiny_nn_top.max_val_skid_q[4] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold348 (.A(_00211_),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold349 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][7] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold350 (.A(\u_tiny_nn_top.core_accumulate_result[10] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold351 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[1][2] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold352 (.A(_00496_),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold353 (.A(\u_tiny_nn_top.max_val_skid_q[3] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold354 (.A(_00210_),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold355 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[1][7] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold356 (.A(_00501_),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold357 (.A(\u_tiny_nn_top.start_count_q[0] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold358 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][1] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold359 (.A(\u_tiny_nn_top.core_accumulate_result[4] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold360 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][14] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold361 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][11] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold362 (.A(_00601_),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold363 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][6] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold364 (.A(_00436_),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold365 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[3][15] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold366 (.A(_00509_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold367 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][13] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold368 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[1][12] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold369 (.A(_00506_),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold370 (.A(\u_tiny_nn_top.max_val_skid_q[6] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold371 (.A(_00213_),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold372 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][0] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold373 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][2] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold374 (.A(\u_tiny_nn_top.u_core.param_val_op_q[1][7] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold375 (.A(_00517_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold376 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][2] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold377 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[3][10] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold378 (.A(_00504_),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold379 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][3] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold380 (.A(_00465_),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold381 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][8] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold382 (.A(_00598_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold383 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][15] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold384 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][4] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold385 (.A(_00466_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold386 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][3] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold387 (.A(_03332_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold388 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[1][1] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold389 (.A(_00495_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold390 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][1] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold391 (.A(_00431_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold392 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][4] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold393 (.A(_03338_),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold394 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][1] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold395 (.A(\u_tiny_nn_top.max_val_skid_q[1] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold396 (.A(_00208_),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold397 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][12] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold398 (.A(_00474_),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold399 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][10] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold400 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[1][4] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold401 (.A(_00498_),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold402 (.A(\u_tiny_nn_top.state_q[5] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold403 (.A(_00009_),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold404 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[6][11] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold405 (.A(\u_tiny_nn_top.core_accumulate_result[6] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold406 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[1][5] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold407 (.A(_00499_),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold408 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][2] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold409 (.A(_03326_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold410 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[3][0] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold411 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][1] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold412 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[1][14] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold413 (.A(_00508_),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold414 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][15] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold415 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[1][9] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold416 (.A(_00503_),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold417 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][3] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold418 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][4] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold419 (.A(\u_tiny_nn_top.max_val_skid_q[2] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold420 (.A(_00209_),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold421 (.A(\u_tiny_nn_top.relu_q ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold422 (.A(_00188_),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold423 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][1] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold424 (.A(_03320_),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold425 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[3][7] ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold426 (.A(_00469_),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold427 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][0] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold428 (.A(_00590_),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold429 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][9] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold430 (.A(_00471_),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold431 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[2][1] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold432 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][7] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold433 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[1][3] ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold434 (.A(_00497_),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold435 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[3][14] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold436 (.A(_00098_),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold437 (.A(_00186_),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold438 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][13] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold439 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][11] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold440 (.A(_00473_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold441 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[3][6] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold442 (.A(_00468_),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold443 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][5] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold444 (.A(_00435_),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold445 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[1][6] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold446 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[6] ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold447 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[4][2] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold448 (.A(\u_tiny_nn_top.core_accumulate_result[15] ),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold449 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[3][5] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold450 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[0] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold451 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[3][1] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold452 (.A(_00463_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold453 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[6] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold454 (.A(\u_tiny_nn_top.max_val_skid_q[7] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold455 (.A(_00214_),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold456 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][15] ),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold457 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[5] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold458 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[3][2] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold459 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][3] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold460 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[1] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold461 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[0] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold462 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][5] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold463 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[6] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold464 (.A(\u_tiny_nn_top.max_val_q[8] ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold465 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[12] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold466 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][7] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold467 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[1] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold468 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[7][8] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold469 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[5][8] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold470 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[5] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold471 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][4] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold472 (.A(\u_tiny_nn_top.max_val_q[9] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold473 (.A(_00247_),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold474 (.A(\u_tiny_nn_top.core_accumulate_result[13] ),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold475 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][6] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold476 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][5] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold477 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[2] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold478 (.A(\u_tiny_nn_top.max_val_q[12] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold479 (.A(_00250_),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold480 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[3] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold481 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[4] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold482 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[5] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold483 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[4] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold484 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[2] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold485 (.A(\u_tiny_nn_top.u_core.mul_val_op_q[3][8] ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold486 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[1] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold487 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[0] ),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold488 (.A(\u_tiny_nn_top.max_val_q[14] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold489 (.A(\u_tiny_nn_top.max_val_q[3] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold490 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][0] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold491 (.A(\u_tiny_nn_top.max_val_q[13] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold492 (.A(_00251_),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold493 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][1] ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold494 (.A(\u_tiny_nn_top.state_q[16] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold495 (.A(_00011_),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold496 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][15] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold497 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[4] ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold498 (.A(\u_tiny_nn_top.max_val_q[5] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold499 (.A(\u_tiny_nn_top.max_val_q[10] ),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold500 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][0] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold501 (.A(\u_tiny_nn_top.state_q[6] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold502 (.A(_01050_),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold503 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][2] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold504 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[3] ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold505 (.A(\u_tiny_nn_top.max_val_q[15] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold506 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[3] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold507 (.A(\u_tiny_nn_top.state_q[3] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold508 (.A(_00012_),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold509 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][8] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold510 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[2] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold511 (.A(\u_tiny_nn_top.state_q[4] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold512 (.A(_00013_),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold513 (.A(\u_tiny_nn_top.max_val_q[11] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold514 (.A(_00249_),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold515 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[9] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold516 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][15] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold517 (.A(\u_tiny_nn_top.max_val_q[2] ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold518 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][7] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold519 (.A(\u_tiny_nn_top.max_val_q[4] ),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold520 (.A(\u_tiny_nn_top.max_val_q[7] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold521 (.A(\u_tiny_nn_top.state_q[7] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold522 (.A(_00187_),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold523 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[14] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold524 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][6] ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold525 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][1] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold526 (.A(\u_tiny_nn_top.counter_q[7] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold527 (.A(_00205_),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold528 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][15] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold529 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][0] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold530 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[15] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold531 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[7] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold532 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][2] ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold533 (.A(\u_tiny_nn_top.max_val_q[1] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold534 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][6] ),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold535 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[13] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold536 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][0] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold537 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][3] ),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold538 (.A(\u_tiny_nn_top.max_val_q[6] ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold539 (.A(\u_tiny_nn_top.u_core.mul_add_op_a_q[1][5] ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold540 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][11] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold541 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][13] ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold542 (.A(\u_tiny_nn_top.counter_q[5] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold543 (.A(_00203_),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold544 (.A(\u_tiny_nn_top.param_write_q[0] ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold545 (.A(_00232_),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold546 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][11] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold547 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][13] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold548 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[15] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold549 (.A(\u_tiny_nn_top.counter_q[3] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold550 (.A(_00201_),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold551 (.A(\u_tiny_nn_top.max_val_q[0] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold552 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[15] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold553 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][12] ),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold554 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][13] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold555 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][14] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold556 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][8] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold557 (.A(\u_tiny_nn_top.counter_q[6] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold558 (.A(_00204_),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold559 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[7] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold560 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][4] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold561 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][12] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold562 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][12] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold563 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][9] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold564 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][15] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold565 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][9] ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold566 (.A(\u_tiny_nn_top.counter_q[2] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold567 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[8] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold568 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][7] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold569 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][13] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold570 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][12] ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold571 (.A(\u_tiny_nn_top.counter_q[4] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold572 (.A(_00202_),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold573 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[7] ),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold574 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][10] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold575 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][6] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold576 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][14] ),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold577 (.A(\u_tiny_nn_top.param_write_q[6] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold578 (.A(_00237_),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold579 (.A(\u_tiny_nn_top.param_write_q[5] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold580 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][7] ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold581 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[11] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold582 (.A(_00088_),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold583 (.A(_00989_),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold584 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[0][8] ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold585 (.A(_00094_),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold586 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][7] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold587 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[11] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold588 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][5] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold589 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[12] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold590 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][11] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold591 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[14] ),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold592 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][14] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold593 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[10] ),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold594 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][9] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold595 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][14] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold596 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][11] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold597 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[13] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold598 (.A(\u_tiny_nn_top.counter_q[1] ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold599 (.A(_00199_),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold600 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][9] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold601 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[8] ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold602 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[1].u_add.op_b_i[8] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold603 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[14] ),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold604 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[13] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold605 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][15] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold606 (.A(\u_tiny_nn_top.data_i_q[12] ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold607 (.A(_00000_),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold608 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[0][10] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold609 (.A(\u_tiny_nn_top.param_write_q[2] ),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold610 (.A(_00234_),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold611 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[11] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold612 (.A(_00090_),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold613 (.A(_00970_),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold614 (.A(_00096_),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold615 (.A(_00930_),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold616 (.A(\u_tiny_nn_top.state_q[0] ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold617 (.A(_00091_),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold618 (.A(_00086_),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold619 (.A(_00994_),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold620 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][7] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold621 (.A(\u_tiny_nn_top.state_q[12] ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold622 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[9] ),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold623 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][8] ),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold624 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[10] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold625 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[9] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold626 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_b_i[12] ),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold627 (.A(\u_tiny_nn_top.u_core.accumulate_level_1_q[1][10] ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold628 (.A(\u_tiny_nn_top.u_core.accumulate_level_0_q[1][10] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold629 (.A(\u_tiny_nn_top.u_core.g_accumulate_level_0_inner[0].u_add.op_a_i[10] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold630 (.A(_00100_),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold631 (.A(\u_tiny_nn_top.param_write_q[3] ),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold632 (.A(\u_tiny_nn_top.data_i_q[14] ),
    .X(net1114));
 sg13g2_antennanp ANTENNA_1 (.A(\u_tiny_nn_top.max_val_skid_q[1] ));
 sg13g2_antennanp ANTENNA_2 (.A(\u_tiny_nn_top.max_val_skid_q[1] ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_945 ();
 sg13g2_decap_8 FILLER_0_952 ();
 sg13g2_decap_8 FILLER_0_959 ();
 sg13g2_decap_8 FILLER_0_966 ();
 sg13g2_decap_8 FILLER_0_973 ();
 sg13g2_decap_8 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_987 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_decap_8 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1008 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1022 ();
 sg13g2_decap_8 FILLER_0_1029 ();
 sg13g2_decap_8 FILLER_0_1036 ();
 sg13g2_decap_8 FILLER_0_1043 ();
 sg13g2_decap_8 FILLER_0_1050 ();
 sg13g2_decap_8 FILLER_0_1057 ();
 sg13g2_decap_8 FILLER_0_1064 ();
 sg13g2_decap_8 FILLER_0_1071 ();
 sg13g2_decap_8 FILLER_0_1078 ();
 sg13g2_decap_8 FILLER_0_1085 ();
 sg13g2_decap_8 FILLER_0_1092 ();
 sg13g2_decap_8 FILLER_0_1099 ();
 sg13g2_decap_8 FILLER_0_1106 ();
 sg13g2_decap_8 FILLER_0_1113 ();
 sg13g2_decap_8 FILLER_0_1120 ();
 sg13g2_decap_8 FILLER_0_1127 ();
 sg13g2_decap_8 FILLER_0_1134 ();
 sg13g2_decap_8 FILLER_0_1141 ();
 sg13g2_decap_8 FILLER_0_1148 ();
 sg13g2_decap_8 FILLER_0_1155 ();
 sg13g2_decap_8 FILLER_0_1162 ();
 sg13g2_decap_8 FILLER_0_1169 ();
 sg13g2_decap_8 FILLER_0_1176 ();
 sg13g2_decap_8 FILLER_0_1183 ();
 sg13g2_decap_8 FILLER_0_1190 ();
 sg13g2_decap_8 FILLER_0_1197 ();
 sg13g2_decap_8 FILLER_0_1204 ();
 sg13g2_decap_8 FILLER_0_1211 ();
 sg13g2_decap_8 FILLER_0_1218 ();
 sg13g2_decap_8 FILLER_0_1225 ();
 sg13g2_decap_8 FILLER_0_1232 ();
 sg13g2_decap_8 FILLER_0_1239 ();
 sg13g2_decap_8 FILLER_0_1246 ();
 sg13g2_decap_8 FILLER_0_1253 ();
 sg13g2_decap_8 FILLER_0_1260 ();
 sg13g2_decap_8 FILLER_0_1267 ();
 sg13g2_decap_8 FILLER_0_1274 ();
 sg13g2_decap_8 FILLER_0_1281 ();
 sg13g2_decap_8 FILLER_0_1288 ();
 sg13g2_decap_8 FILLER_0_1295 ();
 sg13g2_decap_8 FILLER_0_1302 ();
 sg13g2_decap_8 FILLER_0_1309 ();
 sg13g2_decap_8 FILLER_0_1316 ();
 sg13g2_decap_8 FILLER_0_1323 ();
 sg13g2_decap_8 FILLER_0_1330 ();
 sg13g2_decap_8 FILLER_0_1337 ();
 sg13g2_decap_8 FILLER_0_1344 ();
 sg13g2_decap_8 FILLER_0_1351 ();
 sg13g2_decap_8 FILLER_0_1358 ();
 sg13g2_decap_8 FILLER_0_1365 ();
 sg13g2_decap_8 FILLER_0_1372 ();
 sg13g2_decap_8 FILLER_0_1379 ();
 sg13g2_decap_8 FILLER_0_1386 ();
 sg13g2_decap_8 FILLER_0_1393 ();
 sg13g2_decap_8 FILLER_0_1400 ();
 sg13g2_decap_8 FILLER_0_1407 ();
 sg13g2_decap_8 FILLER_0_1414 ();
 sg13g2_decap_8 FILLER_0_1421 ();
 sg13g2_decap_8 FILLER_0_1428 ();
 sg13g2_decap_8 FILLER_0_1435 ();
 sg13g2_decap_8 FILLER_0_1442 ();
 sg13g2_decap_8 FILLER_0_1449 ();
 sg13g2_decap_8 FILLER_0_1456 ();
 sg13g2_decap_8 FILLER_0_1463 ();
 sg13g2_decap_8 FILLER_0_1470 ();
 sg13g2_decap_8 FILLER_0_1477 ();
 sg13g2_decap_8 FILLER_0_1484 ();
 sg13g2_decap_8 FILLER_0_1491 ();
 sg13g2_decap_8 FILLER_0_1498 ();
 sg13g2_decap_8 FILLER_0_1505 ();
 sg13g2_decap_8 FILLER_0_1512 ();
 sg13g2_decap_8 FILLER_0_1519 ();
 sg13g2_decap_8 FILLER_0_1526 ();
 sg13g2_decap_8 FILLER_0_1533 ();
 sg13g2_decap_8 FILLER_0_1540 ();
 sg13g2_decap_8 FILLER_0_1547 ();
 sg13g2_decap_8 FILLER_0_1554 ();
 sg13g2_decap_8 FILLER_0_1561 ();
 sg13g2_decap_8 FILLER_0_1568 ();
 sg13g2_decap_8 FILLER_0_1575 ();
 sg13g2_decap_8 FILLER_0_1582 ();
 sg13g2_decap_8 FILLER_0_1589 ();
 sg13g2_decap_8 FILLER_0_1596 ();
 sg13g2_decap_8 FILLER_0_1603 ();
 sg13g2_decap_8 FILLER_0_1610 ();
 sg13g2_decap_8 FILLER_0_1617 ();
 sg13g2_decap_8 FILLER_0_1624 ();
 sg13g2_decap_8 FILLER_0_1631 ();
 sg13g2_decap_8 FILLER_0_1638 ();
 sg13g2_decap_8 FILLER_0_1645 ();
 sg13g2_decap_8 FILLER_0_1652 ();
 sg13g2_decap_8 FILLER_0_1659 ();
 sg13g2_decap_8 FILLER_0_1666 ();
 sg13g2_decap_8 FILLER_0_1673 ();
 sg13g2_decap_8 FILLER_0_1680 ();
 sg13g2_decap_8 FILLER_0_1687 ();
 sg13g2_decap_8 FILLER_0_1694 ();
 sg13g2_decap_8 FILLER_0_1701 ();
 sg13g2_decap_8 FILLER_0_1708 ();
 sg13g2_decap_8 FILLER_0_1715 ();
 sg13g2_decap_8 FILLER_0_1722 ();
 sg13g2_decap_8 FILLER_0_1729 ();
 sg13g2_decap_8 FILLER_0_1736 ();
 sg13g2_decap_8 FILLER_0_1743 ();
 sg13g2_decap_8 FILLER_0_1750 ();
 sg13g2_decap_8 FILLER_0_1757 ();
 sg13g2_decap_4 FILLER_0_1764 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_decap_8 FILLER_1_875 ();
 sg13g2_decap_8 FILLER_1_882 ();
 sg13g2_decap_8 FILLER_1_889 ();
 sg13g2_decap_8 FILLER_1_896 ();
 sg13g2_decap_8 FILLER_1_903 ();
 sg13g2_decap_8 FILLER_1_910 ();
 sg13g2_decap_8 FILLER_1_917 ();
 sg13g2_decap_8 FILLER_1_924 ();
 sg13g2_decap_8 FILLER_1_931 ();
 sg13g2_decap_8 FILLER_1_938 ();
 sg13g2_decap_8 FILLER_1_945 ();
 sg13g2_decap_8 FILLER_1_952 ();
 sg13g2_decap_8 FILLER_1_959 ();
 sg13g2_decap_8 FILLER_1_966 ();
 sg13g2_decap_8 FILLER_1_973 ();
 sg13g2_decap_8 FILLER_1_980 ();
 sg13g2_decap_8 FILLER_1_987 ();
 sg13g2_decap_8 FILLER_1_994 ();
 sg13g2_decap_8 FILLER_1_1001 ();
 sg13g2_decap_8 FILLER_1_1008 ();
 sg13g2_decap_8 FILLER_1_1015 ();
 sg13g2_decap_8 FILLER_1_1022 ();
 sg13g2_decap_8 FILLER_1_1029 ();
 sg13g2_decap_8 FILLER_1_1036 ();
 sg13g2_decap_8 FILLER_1_1043 ();
 sg13g2_decap_8 FILLER_1_1050 ();
 sg13g2_decap_8 FILLER_1_1057 ();
 sg13g2_decap_8 FILLER_1_1064 ();
 sg13g2_decap_8 FILLER_1_1071 ();
 sg13g2_decap_8 FILLER_1_1078 ();
 sg13g2_decap_8 FILLER_1_1085 ();
 sg13g2_decap_8 FILLER_1_1092 ();
 sg13g2_decap_8 FILLER_1_1099 ();
 sg13g2_decap_8 FILLER_1_1106 ();
 sg13g2_decap_8 FILLER_1_1113 ();
 sg13g2_decap_8 FILLER_1_1120 ();
 sg13g2_decap_8 FILLER_1_1127 ();
 sg13g2_decap_8 FILLER_1_1134 ();
 sg13g2_decap_8 FILLER_1_1141 ();
 sg13g2_decap_8 FILLER_1_1148 ();
 sg13g2_decap_8 FILLER_1_1155 ();
 sg13g2_decap_8 FILLER_1_1162 ();
 sg13g2_decap_8 FILLER_1_1169 ();
 sg13g2_decap_8 FILLER_1_1176 ();
 sg13g2_decap_8 FILLER_1_1183 ();
 sg13g2_decap_8 FILLER_1_1190 ();
 sg13g2_decap_8 FILLER_1_1197 ();
 sg13g2_decap_8 FILLER_1_1204 ();
 sg13g2_decap_8 FILLER_1_1211 ();
 sg13g2_decap_8 FILLER_1_1218 ();
 sg13g2_decap_8 FILLER_1_1225 ();
 sg13g2_decap_8 FILLER_1_1232 ();
 sg13g2_decap_8 FILLER_1_1239 ();
 sg13g2_decap_8 FILLER_1_1246 ();
 sg13g2_decap_8 FILLER_1_1253 ();
 sg13g2_decap_8 FILLER_1_1260 ();
 sg13g2_decap_8 FILLER_1_1267 ();
 sg13g2_decap_8 FILLER_1_1274 ();
 sg13g2_decap_8 FILLER_1_1281 ();
 sg13g2_decap_8 FILLER_1_1288 ();
 sg13g2_decap_8 FILLER_1_1295 ();
 sg13g2_decap_8 FILLER_1_1302 ();
 sg13g2_decap_8 FILLER_1_1309 ();
 sg13g2_decap_8 FILLER_1_1316 ();
 sg13g2_decap_8 FILLER_1_1323 ();
 sg13g2_decap_8 FILLER_1_1330 ();
 sg13g2_decap_8 FILLER_1_1337 ();
 sg13g2_decap_8 FILLER_1_1344 ();
 sg13g2_decap_8 FILLER_1_1351 ();
 sg13g2_decap_8 FILLER_1_1358 ();
 sg13g2_decap_8 FILLER_1_1365 ();
 sg13g2_decap_8 FILLER_1_1372 ();
 sg13g2_decap_8 FILLER_1_1379 ();
 sg13g2_decap_8 FILLER_1_1386 ();
 sg13g2_decap_8 FILLER_1_1393 ();
 sg13g2_decap_8 FILLER_1_1400 ();
 sg13g2_decap_8 FILLER_1_1407 ();
 sg13g2_decap_8 FILLER_1_1414 ();
 sg13g2_decap_8 FILLER_1_1421 ();
 sg13g2_decap_8 FILLER_1_1428 ();
 sg13g2_decap_8 FILLER_1_1435 ();
 sg13g2_decap_8 FILLER_1_1442 ();
 sg13g2_decap_8 FILLER_1_1449 ();
 sg13g2_decap_8 FILLER_1_1456 ();
 sg13g2_decap_8 FILLER_1_1463 ();
 sg13g2_decap_8 FILLER_1_1470 ();
 sg13g2_decap_8 FILLER_1_1477 ();
 sg13g2_decap_8 FILLER_1_1484 ();
 sg13g2_decap_8 FILLER_1_1491 ();
 sg13g2_decap_8 FILLER_1_1498 ();
 sg13g2_decap_8 FILLER_1_1505 ();
 sg13g2_decap_8 FILLER_1_1512 ();
 sg13g2_decap_8 FILLER_1_1519 ();
 sg13g2_decap_8 FILLER_1_1526 ();
 sg13g2_decap_8 FILLER_1_1533 ();
 sg13g2_decap_8 FILLER_1_1540 ();
 sg13g2_decap_8 FILLER_1_1547 ();
 sg13g2_decap_8 FILLER_1_1554 ();
 sg13g2_decap_8 FILLER_1_1561 ();
 sg13g2_decap_8 FILLER_1_1568 ();
 sg13g2_decap_8 FILLER_1_1575 ();
 sg13g2_decap_8 FILLER_1_1582 ();
 sg13g2_decap_8 FILLER_1_1589 ();
 sg13g2_decap_8 FILLER_1_1596 ();
 sg13g2_decap_8 FILLER_1_1603 ();
 sg13g2_decap_8 FILLER_1_1610 ();
 sg13g2_decap_8 FILLER_1_1617 ();
 sg13g2_decap_8 FILLER_1_1624 ();
 sg13g2_decap_8 FILLER_1_1631 ();
 sg13g2_decap_8 FILLER_1_1638 ();
 sg13g2_decap_8 FILLER_1_1645 ();
 sg13g2_decap_8 FILLER_1_1652 ();
 sg13g2_decap_8 FILLER_1_1659 ();
 sg13g2_decap_8 FILLER_1_1666 ();
 sg13g2_decap_8 FILLER_1_1673 ();
 sg13g2_decap_8 FILLER_1_1680 ();
 sg13g2_decap_8 FILLER_1_1687 ();
 sg13g2_decap_8 FILLER_1_1694 ();
 sg13g2_decap_8 FILLER_1_1701 ();
 sg13g2_decap_8 FILLER_1_1708 ();
 sg13g2_decap_8 FILLER_1_1715 ();
 sg13g2_decap_8 FILLER_1_1722 ();
 sg13g2_decap_8 FILLER_1_1729 ();
 sg13g2_decap_8 FILLER_1_1736 ();
 sg13g2_decap_8 FILLER_1_1743 ();
 sg13g2_decap_8 FILLER_1_1750 ();
 sg13g2_decap_8 FILLER_1_1757 ();
 sg13g2_decap_4 FILLER_1_1764 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_4 FILLER_2_441 ();
 sg13g2_fill_1 FILLER_2_445 ();
 sg13g2_fill_1 FILLER_2_451 ();
 sg13g2_fill_1 FILLER_2_455 ();
 sg13g2_decap_4 FILLER_2_460 ();
 sg13g2_decap_8 FILLER_2_468 ();
 sg13g2_decap_8 FILLER_2_475 ();
 sg13g2_fill_1 FILLER_2_482 ();
 sg13g2_decap_8 FILLER_2_487 ();
 sg13g2_decap_8 FILLER_2_494 ();
 sg13g2_decap_8 FILLER_2_501 ();
 sg13g2_decap_8 FILLER_2_508 ();
 sg13g2_decap_8 FILLER_2_515 ();
 sg13g2_decap_8 FILLER_2_522 ();
 sg13g2_decap_8 FILLER_2_529 ();
 sg13g2_decap_8 FILLER_2_536 ();
 sg13g2_decap_8 FILLER_2_543 ();
 sg13g2_decap_8 FILLER_2_550 ();
 sg13g2_decap_8 FILLER_2_557 ();
 sg13g2_decap_8 FILLER_2_564 ();
 sg13g2_decap_8 FILLER_2_571 ();
 sg13g2_decap_8 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_585 ();
 sg13g2_decap_8 FILLER_2_592 ();
 sg13g2_decap_8 FILLER_2_599 ();
 sg13g2_decap_8 FILLER_2_606 ();
 sg13g2_decap_8 FILLER_2_613 ();
 sg13g2_decap_8 FILLER_2_620 ();
 sg13g2_decap_8 FILLER_2_627 ();
 sg13g2_decap_8 FILLER_2_634 ();
 sg13g2_decap_8 FILLER_2_641 ();
 sg13g2_decap_8 FILLER_2_648 ();
 sg13g2_decap_8 FILLER_2_655 ();
 sg13g2_decap_8 FILLER_2_662 ();
 sg13g2_decap_8 FILLER_2_669 ();
 sg13g2_decap_8 FILLER_2_676 ();
 sg13g2_decap_8 FILLER_2_683 ();
 sg13g2_decap_8 FILLER_2_690 ();
 sg13g2_decap_8 FILLER_2_697 ();
 sg13g2_decap_8 FILLER_2_704 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_decap_8 FILLER_2_718 ();
 sg13g2_decap_8 FILLER_2_725 ();
 sg13g2_decap_8 FILLER_2_732 ();
 sg13g2_decap_8 FILLER_2_739 ();
 sg13g2_decap_8 FILLER_2_746 ();
 sg13g2_decap_8 FILLER_2_753 ();
 sg13g2_decap_8 FILLER_2_760 ();
 sg13g2_decap_8 FILLER_2_767 ();
 sg13g2_decap_8 FILLER_2_774 ();
 sg13g2_decap_8 FILLER_2_781 ();
 sg13g2_decap_8 FILLER_2_788 ();
 sg13g2_decap_8 FILLER_2_795 ();
 sg13g2_decap_8 FILLER_2_802 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_8 FILLER_2_858 ();
 sg13g2_decap_8 FILLER_2_865 ();
 sg13g2_decap_8 FILLER_2_872 ();
 sg13g2_decap_8 FILLER_2_879 ();
 sg13g2_decap_8 FILLER_2_886 ();
 sg13g2_decap_8 FILLER_2_893 ();
 sg13g2_decap_8 FILLER_2_900 ();
 sg13g2_decap_8 FILLER_2_907 ();
 sg13g2_decap_8 FILLER_2_914 ();
 sg13g2_decap_8 FILLER_2_921 ();
 sg13g2_decap_8 FILLER_2_928 ();
 sg13g2_decap_8 FILLER_2_935 ();
 sg13g2_decap_8 FILLER_2_942 ();
 sg13g2_decap_8 FILLER_2_949 ();
 sg13g2_decap_8 FILLER_2_956 ();
 sg13g2_decap_8 FILLER_2_963 ();
 sg13g2_decap_8 FILLER_2_970 ();
 sg13g2_decap_8 FILLER_2_977 ();
 sg13g2_decap_8 FILLER_2_984 ();
 sg13g2_decap_8 FILLER_2_991 ();
 sg13g2_decap_8 FILLER_2_998 ();
 sg13g2_decap_8 FILLER_2_1005 ();
 sg13g2_decap_8 FILLER_2_1012 ();
 sg13g2_decap_8 FILLER_2_1019 ();
 sg13g2_decap_8 FILLER_2_1026 ();
 sg13g2_decap_8 FILLER_2_1033 ();
 sg13g2_decap_8 FILLER_2_1040 ();
 sg13g2_decap_8 FILLER_2_1047 ();
 sg13g2_decap_8 FILLER_2_1054 ();
 sg13g2_decap_8 FILLER_2_1061 ();
 sg13g2_decap_8 FILLER_2_1068 ();
 sg13g2_decap_8 FILLER_2_1075 ();
 sg13g2_decap_8 FILLER_2_1082 ();
 sg13g2_decap_8 FILLER_2_1089 ();
 sg13g2_decap_8 FILLER_2_1096 ();
 sg13g2_decap_8 FILLER_2_1103 ();
 sg13g2_decap_8 FILLER_2_1110 ();
 sg13g2_decap_8 FILLER_2_1117 ();
 sg13g2_decap_8 FILLER_2_1124 ();
 sg13g2_decap_8 FILLER_2_1131 ();
 sg13g2_decap_8 FILLER_2_1138 ();
 sg13g2_decap_8 FILLER_2_1145 ();
 sg13g2_decap_8 FILLER_2_1152 ();
 sg13g2_decap_8 FILLER_2_1159 ();
 sg13g2_decap_8 FILLER_2_1166 ();
 sg13g2_decap_8 FILLER_2_1173 ();
 sg13g2_decap_8 FILLER_2_1180 ();
 sg13g2_decap_8 FILLER_2_1187 ();
 sg13g2_decap_8 FILLER_2_1194 ();
 sg13g2_decap_8 FILLER_2_1201 ();
 sg13g2_decap_8 FILLER_2_1208 ();
 sg13g2_decap_8 FILLER_2_1215 ();
 sg13g2_decap_8 FILLER_2_1222 ();
 sg13g2_decap_8 FILLER_2_1229 ();
 sg13g2_decap_8 FILLER_2_1236 ();
 sg13g2_decap_8 FILLER_2_1243 ();
 sg13g2_decap_8 FILLER_2_1250 ();
 sg13g2_decap_8 FILLER_2_1257 ();
 sg13g2_decap_8 FILLER_2_1264 ();
 sg13g2_decap_8 FILLER_2_1271 ();
 sg13g2_decap_8 FILLER_2_1278 ();
 sg13g2_decap_8 FILLER_2_1285 ();
 sg13g2_decap_8 FILLER_2_1292 ();
 sg13g2_decap_8 FILLER_2_1299 ();
 sg13g2_decap_8 FILLER_2_1306 ();
 sg13g2_decap_8 FILLER_2_1313 ();
 sg13g2_decap_8 FILLER_2_1320 ();
 sg13g2_decap_8 FILLER_2_1327 ();
 sg13g2_decap_8 FILLER_2_1334 ();
 sg13g2_decap_8 FILLER_2_1341 ();
 sg13g2_decap_8 FILLER_2_1348 ();
 sg13g2_decap_8 FILLER_2_1355 ();
 sg13g2_decap_8 FILLER_2_1362 ();
 sg13g2_decap_8 FILLER_2_1369 ();
 sg13g2_decap_8 FILLER_2_1376 ();
 sg13g2_decap_8 FILLER_2_1383 ();
 sg13g2_decap_8 FILLER_2_1390 ();
 sg13g2_decap_8 FILLER_2_1397 ();
 sg13g2_decap_8 FILLER_2_1404 ();
 sg13g2_decap_8 FILLER_2_1411 ();
 sg13g2_decap_8 FILLER_2_1418 ();
 sg13g2_decap_8 FILLER_2_1425 ();
 sg13g2_decap_8 FILLER_2_1432 ();
 sg13g2_decap_8 FILLER_2_1439 ();
 sg13g2_decap_8 FILLER_2_1446 ();
 sg13g2_decap_8 FILLER_2_1453 ();
 sg13g2_decap_8 FILLER_2_1460 ();
 sg13g2_decap_8 FILLER_2_1467 ();
 sg13g2_decap_8 FILLER_2_1474 ();
 sg13g2_decap_8 FILLER_2_1481 ();
 sg13g2_decap_8 FILLER_2_1488 ();
 sg13g2_decap_8 FILLER_2_1495 ();
 sg13g2_decap_8 FILLER_2_1502 ();
 sg13g2_decap_8 FILLER_2_1509 ();
 sg13g2_decap_8 FILLER_2_1516 ();
 sg13g2_decap_8 FILLER_2_1523 ();
 sg13g2_decap_8 FILLER_2_1530 ();
 sg13g2_decap_8 FILLER_2_1537 ();
 sg13g2_decap_8 FILLER_2_1544 ();
 sg13g2_decap_8 FILLER_2_1551 ();
 sg13g2_decap_8 FILLER_2_1558 ();
 sg13g2_decap_8 FILLER_2_1565 ();
 sg13g2_decap_8 FILLER_2_1572 ();
 sg13g2_decap_8 FILLER_2_1579 ();
 sg13g2_decap_8 FILLER_2_1586 ();
 sg13g2_decap_8 FILLER_2_1593 ();
 sg13g2_decap_8 FILLER_2_1600 ();
 sg13g2_decap_8 FILLER_2_1607 ();
 sg13g2_decap_8 FILLER_2_1614 ();
 sg13g2_decap_8 FILLER_2_1621 ();
 sg13g2_decap_8 FILLER_2_1628 ();
 sg13g2_decap_8 FILLER_2_1635 ();
 sg13g2_decap_8 FILLER_2_1642 ();
 sg13g2_decap_8 FILLER_2_1649 ();
 sg13g2_decap_8 FILLER_2_1656 ();
 sg13g2_decap_8 FILLER_2_1663 ();
 sg13g2_decap_8 FILLER_2_1670 ();
 sg13g2_decap_8 FILLER_2_1677 ();
 sg13g2_decap_8 FILLER_2_1684 ();
 sg13g2_decap_8 FILLER_2_1691 ();
 sg13g2_decap_8 FILLER_2_1698 ();
 sg13g2_decap_8 FILLER_2_1705 ();
 sg13g2_decap_8 FILLER_2_1712 ();
 sg13g2_decap_8 FILLER_2_1719 ();
 sg13g2_decap_8 FILLER_2_1726 ();
 sg13g2_decap_8 FILLER_2_1733 ();
 sg13g2_decap_8 FILLER_2_1740 ();
 sg13g2_decap_8 FILLER_2_1747 ();
 sg13g2_decap_8 FILLER_2_1754 ();
 sg13g2_decap_8 FILLER_2_1761 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_fill_2 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_499 ();
 sg13g2_decap_8 FILLER_3_506 ();
 sg13g2_fill_2 FILLER_3_513 ();
 sg13g2_fill_1 FILLER_3_515 ();
 sg13g2_decap_8 FILLER_3_531 ();
 sg13g2_decap_8 FILLER_3_538 ();
 sg13g2_decap_8 FILLER_3_545 ();
 sg13g2_decap_8 FILLER_3_552 ();
 sg13g2_decap_8 FILLER_3_559 ();
 sg13g2_decap_8 FILLER_3_566 ();
 sg13g2_decap_8 FILLER_3_573 ();
 sg13g2_decap_8 FILLER_3_580 ();
 sg13g2_decap_8 FILLER_3_587 ();
 sg13g2_decap_8 FILLER_3_594 ();
 sg13g2_decap_8 FILLER_3_601 ();
 sg13g2_decap_8 FILLER_3_608 ();
 sg13g2_decap_8 FILLER_3_615 ();
 sg13g2_decap_8 FILLER_3_622 ();
 sg13g2_decap_8 FILLER_3_629 ();
 sg13g2_decap_8 FILLER_3_636 ();
 sg13g2_decap_8 FILLER_3_643 ();
 sg13g2_decap_8 FILLER_3_650 ();
 sg13g2_decap_8 FILLER_3_657 ();
 sg13g2_decap_8 FILLER_3_664 ();
 sg13g2_decap_8 FILLER_3_671 ();
 sg13g2_decap_8 FILLER_3_678 ();
 sg13g2_decap_8 FILLER_3_685 ();
 sg13g2_decap_8 FILLER_3_692 ();
 sg13g2_decap_8 FILLER_3_699 ();
 sg13g2_decap_8 FILLER_3_706 ();
 sg13g2_decap_8 FILLER_3_713 ();
 sg13g2_decap_8 FILLER_3_720 ();
 sg13g2_decap_8 FILLER_3_727 ();
 sg13g2_decap_8 FILLER_3_734 ();
 sg13g2_decap_8 FILLER_3_741 ();
 sg13g2_decap_8 FILLER_3_748 ();
 sg13g2_decap_8 FILLER_3_755 ();
 sg13g2_decap_8 FILLER_3_762 ();
 sg13g2_decap_8 FILLER_3_769 ();
 sg13g2_decap_8 FILLER_3_776 ();
 sg13g2_decap_8 FILLER_3_783 ();
 sg13g2_decap_8 FILLER_3_790 ();
 sg13g2_decap_8 FILLER_3_797 ();
 sg13g2_decap_8 FILLER_3_804 ();
 sg13g2_decap_8 FILLER_3_811 ();
 sg13g2_decap_8 FILLER_3_818 ();
 sg13g2_decap_8 FILLER_3_825 ();
 sg13g2_decap_8 FILLER_3_832 ();
 sg13g2_decap_8 FILLER_3_839 ();
 sg13g2_decap_8 FILLER_3_846 ();
 sg13g2_decap_8 FILLER_3_853 ();
 sg13g2_decap_8 FILLER_3_860 ();
 sg13g2_decap_8 FILLER_3_867 ();
 sg13g2_decap_8 FILLER_3_874 ();
 sg13g2_decap_8 FILLER_3_881 ();
 sg13g2_decap_8 FILLER_3_888 ();
 sg13g2_decap_8 FILLER_3_895 ();
 sg13g2_decap_8 FILLER_3_902 ();
 sg13g2_decap_8 FILLER_3_909 ();
 sg13g2_decap_8 FILLER_3_916 ();
 sg13g2_decap_8 FILLER_3_923 ();
 sg13g2_decap_8 FILLER_3_930 ();
 sg13g2_decap_8 FILLER_3_937 ();
 sg13g2_decap_8 FILLER_3_944 ();
 sg13g2_decap_8 FILLER_3_951 ();
 sg13g2_decap_8 FILLER_3_958 ();
 sg13g2_decap_8 FILLER_3_965 ();
 sg13g2_decap_8 FILLER_3_972 ();
 sg13g2_decap_8 FILLER_3_979 ();
 sg13g2_decap_8 FILLER_3_986 ();
 sg13g2_decap_8 FILLER_3_993 ();
 sg13g2_decap_8 FILLER_3_1000 ();
 sg13g2_decap_8 FILLER_3_1007 ();
 sg13g2_decap_8 FILLER_3_1014 ();
 sg13g2_decap_8 FILLER_3_1021 ();
 sg13g2_decap_8 FILLER_3_1028 ();
 sg13g2_decap_8 FILLER_3_1035 ();
 sg13g2_decap_8 FILLER_3_1042 ();
 sg13g2_decap_8 FILLER_3_1049 ();
 sg13g2_decap_8 FILLER_3_1056 ();
 sg13g2_decap_8 FILLER_3_1063 ();
 sg13g2_decap_8 FILLER_3_1070 ();
 sg13g2_decap_8 FILLER_3_1077 ();
 sg13g2_decap_8 FILLER_3_1084 ();
 sg13g2_decap_8 FILLER_3_1091 ();
 sg13g2_decap_8 FILLER_3_1098 ();
 sg13g2_decap_8 FILLER_3_1105 ();
 sg13g2_decap_8 FILLER_3_1112 ();
 sg13g2_decap_8 FILLER_3_1119 ();
 sg13g2_decap_8 FILLER_3_1126 ();
 sg13g2_decap_8 FILLER_3_1133 ();
 sg13g2_decap_8 FILLER_3_1140 ();
 sg13g2_decap_8 FILLER_3_1147 ();
 sg13g2_decap_8 FILLER_3_1154 ();
 sg13g2_decap_8 FILLER_3_1161 ();
 sg13g2_decap_8 FILLER_3_1168 ();
 sg13g2_decap_8 FILLER_3_1175 ();
 sg13g2_decap_8 FILLER_3_1182 ();
 sg13g2_decap_8 FILLER_3_1189 ();
 sg13g2_decap_8 FILLER_3_1196 ();
 sg13g2_decap_8 FILLER_3_1203 ();
 sg13g2_decap_8 FILLER_3_1210 ();
 sg13g2_decap_8 FILLER_3_1217 ();
 sg13g2_decap_8 FILLER_3_1224 ();
 sg13g2_decap_8 FILLER_3_1231 ();
 sg13g2_decap_8 FILLER_3_1238 ();
 sg13g2_decap_8 FILLER_3_1245 ();
 sg13g2_decap_8 FILLER_3_1252 ();
 sg13g2_decap_8 FILLER_3_1259 ();
 sg13g2_decap_8 FILLER_3_1266 ();
 sg13g2_decap_8 FILLER_3_1273 ();
 sg13g2_decap_8 FILLER_3_1280 ();
 sg13g2_decap_8 FILLER_3_1287 ();
 sg13g2_decap_8 FILLER_3_1294 ();
 sg13g2_decap_8 FILLER_3_1301 ();
 sg13g2_decap_8 FILLER_3_1308 ();
 sg13g2_decap_8 FILLER_3_1315 ();
 sg13g2_decap_8 FILLER_3_1322 ();
 sg13g2_decap_8 FILLER_3_1329 ();
 sg13g2_decap_8 FILLER_3_1336 ();
 sg13g2_decap_8 FILLER_3_1343 ();
 sg13g2_decap_8 FILLER_3_1350 ();
 sg13g2_decap_8 FILLER_3_1357 ();
 sg13g2_decap_8 FILLER_3_1364 ();
 sg13g2_decap_8 FILLER_3_1371 ();
 sg13g2_decap_8 FILLER_3_1378 ();
 sg13g2_decap_8 FILLER_3_1385 ();
 sg13g2_decap_8 FILLER_3_1392 ();
 sg13g2_decap_8 FILLER_3_1399 ();
 sg13g2_decap_8 FILLER_3_1406 ();
 sg13g2_decap_8 FILLER_3_1413 ();
 sg13g2_decap_8 FILLER_3_1420 ();
 sg13g2_decap_8 FILLER_3_1427 ();
 sg13g2_decap_8 FILLER_3_1434 ();
 sg13g2_decap_8 FILLER_3_1441 ();
 sg13g2_decap_8 FILLER_3_1448 ();
 sg13g2_decap_8 FILLER_3_1455 ();
 sg13g2_decap_8 FILLER_3_1462 ();
 sg13g2_decap_8 FILLER_3_1469 ();
 sg13g2_decap_8 FILLER_3_1476 ();
 sg13g2_decap_8 FILLER_3_1483 ();
 sg13g2_decap_8 FILLER_3_1490 ();
 sg13g2_decap_8 FILLER_3_1497 ();
 sg13g2_decap_8 FILLER_3_1504 ();
 sg13g2_decap_8 FILLER_3_1511 ();
 sg13g2_decap_8 FILLER_3_1518 ();
 sg13g2_decap_8 FILLER_3_1525 ();
 sg13g2_decap_8 FILLER_3_1532 ();
 sg13g2_decap_8 FILLER_3_1539 ();
 sg13g2_decap_8 FILLER_3_1546 ();
 sg13g2_decap_8 FILLER_3_1553 ();
 sg13g2_decap_8 FILLER_3_1560 ();
 sg13g2_decap_8 FILLER_3_1567 ();
 sg13g2_decap_8 FILLER_3_1574 ();
 sg13g2_decap_8 FILLER_3_1581 ();
 sg13g2_decap_8 FILLER_3_1588 ();
 sg13g2_decap_8 FILLER_3_1595 ();
 sg13g2_decap_8 FILLER_3_1602 ();
 sg13g2_decap_8 FILLER_3_1609 ();
 sg13g2_decap_8 FILLER_3_1616 ();
 sg13g2_decap_8 FILLER_3_1623 ();
 sg13g2_decap_8 FILLER_3_1630 ();
 sg13g2_decap_8 FILLER_3_1637 ();
 sg13g2_decap_8 FILLER_3_1644 ();
 sg13g2_decap_8 FILLER_3_1651 ();
 sg13g2_decap_8 FILLER_3_1658 ();
 sg13g2_decap_8 FILLER_3_1665 ();
 sg13g2_decap_8 FILLER_3_1672 ();
 sg13g2_decap_8 FILLER_3_1679 ();
 sg13g2_decap_8 FILLER_3_1686 ();
 sg13g2_decap_8 FILLER_3_1693 ();
 sg13g2_decap_8 FILLER_3_1700 ();
 sg13g2_decap_8 FILLER_3_1707 ();
 sg13g2_decap_8 FILLER_3_1714 ();
 sg13g2_decap_8 FILLER_3_1721 ();
 sg13g2_decap_8 FILLER_3_1728 ();
 sg13g2_decap_8 FILLER_3_1735 ();
 sg13g2_decap_8 FILLER_3_1742 ();
 sg13g2_decap_8 FILLER_3_1749 ();
 sg13g2_decap_8 FILLER_3_1756 ();
 sg13g2_decap_4 FILLER_3_1763 ();
 sg13g2_fill_1 FILLER_3_1767 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_fill_2 FILLER_4_413 ();
 sg13g2_fill_1 FILLER_4_415 ();
 sg13g2_fill_1 FILLER_4_441 ();
 sg13g2_fill_1 FILLER_4_447 ();
 sg13g2_decap_8 FILLER_4_452 ();
 sg13g2_fill_2 FILLER_4_459 ();
 sg13g2_fill_1 FILLER_4_465 ();
 sg13g2_decap_8 FILLER_4_475 ();
 sg13g2_decap_8 FILLER_4_482 ();
 sg13g2_fill_1 FILLER_4_489 ();
 sg13g2_fill_1 FILLER_4_506 ();
 sg13g2_decap_4 FILLER_4_542 ();
 sg13g2_fill_2 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_559 ();
 sg13g2_decap_8 FILLER_4_566 ();
 sg13g2_decap_8 FILLER_4_573 ();
 sg13g2_decap_8 FILLER_4_580 ();
 sg13g2_decap_8 FILLER_4_587 ();
 sg13g2_decap_8 FILLER_4_594 ();
 sg13g2_decap_8 FILLER_4_601 ();
 sg13g2_decap_8 FILLER_4_608 ();
 sg13g2_decap_8 FILLER_4_615 ();
 sg13g2_decap_8 FILLER_4_622 ();
 sg13g2_decap_8 FILLER_4_629 ();
 sg13g2_decap_8 FILLER_4_636 ();
 sg13g2_decap_8 FILLER_4_643 ();
 sg13g2_decap_8 FILLER_4_650 ();
 sg13g2_decap_8 FILLER_4_657 ();
 sg13g2_decap_8 FILLER_4_664 ();
 sg13g2_decap_8 FILLER_4_671 ();
 sg13g2_decap_8 FILLER_4_678 ();
 sg13g2_decap_8 FILLER_4_685 ();
 sg13g2_decap_8 FILLER_4_692 ();
 sg13g2_decap_8 FILLER_4_699 ();
 sg13g2_decap_8 FILLER_4_706 ();
 sg13g2_decap_8 FILLER_4_713 ();
 sg13g2_decap_8 FILLER_4_720 ();
 sg13g2_decap_8 FILLER_4_727 ();
 sg13g2_decap_8 FILLER_4_734 ();
 sg13g2_decap_8 FILLER_4_741 ();
 sg13g2_decap_8 FILLER_4_748 ();
 sg13g2_decap_8 FILLER_4_755 ();
 sg13g2_decap_8 FILLER_4_762 ();
 sg13g2_decap_8 FILLER_4_769 ();
 sg13g2_decap_8 FILLER_4_776 ();
 sg13g2_decap_8 FILLER_4_783 ();
 sg13g2_decap_8 FILLER_4_790 ();
 sg13g2_decap_8 FILLER_4_797 ();
 sg13g2_decap_8 FILLER_4_804 ();
 sg13g2_decap_8 FILLER_4_811 ();
 sg13g2_decap_8 FILLER_4_818 ();
 sg13g2_decap_8 FILLER_4_825 ();
 sg13g2_decap_8 FILLER_4_832 ();
 sg13g2_decap_8 FILLER_4_839 ();
 sg13g2_decap_8 FILLER_4_846 ();
 sg13g2_decap_8 FILLER_4_853 ();
 sg13g2_decap_8 FILLER_4_860 ();
 sg13g2_decap_8 FILLER_4_867 ();
 sg13g2_decap_8 FILLER_4_874 ();
 sg13g2_decap_8 FILLER_4_881 ();
 sg13g2_decap_8 FILLER_4_888 ();
 sg13g2_decap_8 FILLER_4_895 ();
 sg13g2_decap_8 FILLER_4_902 ();
 sg13g2_decap_8 FILLER_4_909 ();
 sg13g2_decap_8 FILLER_4_916 ();
 sg13g2_decap_8 FILLER_4_923 ();
 sg13g2_decap_8 FILLER_4_930 ();
 sg13g2_decap_8 FILLER_4_937 ();
 sg13g2_decap_8 FILLER_4_944 ();
 sg13g2_decap_8 FILLER_4_951 ();
 sg13g2_decap_8 FILLER_4_958 ();
 sg13g2_decap_8 FILLER_4_965 ();
 sg13g2_decap_8 FILLER_4_972 ();
 sg13g2_decap_8 FILLER_4_979 ();
 sg13g2_decap_8 FILLER_4_986 ();
 sg13g2_decap_8 FILLER_4_993 ();
 sg13g2_decap_8 FILLER_4_1000 ();
 sg13g2_decap_8 FILLER_4_1007 ();
 sg13g2_decap_8 FILLER_4_1014 ();
 sg13g2_decap_8 FILLER_4_1021 ();
 sg13g2_decap_8 FILLER_4_1028 ();
 sg13g2_decap_8 FILLER_4_1035 ();
 sg13g2_decap_8 FILLER_4_1042 ();
 sg13g2_decap_8 FILLER_4_1049 ();
 sg13g2_decap_8 FILLER_4_1056 ();
 sg13g2_decap_8 FILLER_4_1063 ();
 sg13g2_decap_8 FILLER_4_1070 ();
 sg13g2_decap_8 FILLER_4_1077 ();
 sg13g2_decap_8 FILLER_4_1084 ();
 sg13g2_decap_8 FILLER_4_1091 ();
 sg13g2_decap_8 FILLER_4_1098 ();
 sg13g2_decap_8 FILLER_4_1105 ();
 sg13g2_decap_8 FILLER_4_1112 ();
 sg13g2_decap_8 FILLER_4_1119 ();
 sg13g2_decap_8 FILLER_4_1126 ();
 sg13g2_decap_8 FILLER_4_1133 ();
 sg13g2_decap_8 FILLER_4_1140 ();
 sg13g2_decap_8 FILLER_4_1147 ();
 sg13g2_decap_8 FILLER_4_1154 ();
 sg13g2_decap_8 FILLER_4_1161 ();
 sg13g2_decap_8 FILLER_4_1168 ();
 sg13g2_decap_8 FILLER_4_1175 ();
 sg13g2_decap_8 FILLER_4_1182 ();
 sg13g2_decap_8 FILLER_4_1189 ();
 sg13g2_decap_8 FILLER_4_1196 ();
 sg13g2_decap_8 FILLER_4_1203 ();
 sg13g2_decap_8 FILLER_4_1210 ();
 sg13g2_decap_8 FILLER_4_1217 ();
 sg13g2_decap_8 FILLER_4_1224 ();
 sg13g2_decap_8 FILLER_4_1231 ();
 sg13g2_decap_8 FILLER_4_1238 ();
 sg13g2_decap_8 FILLER_4_1245 ();
 sg13g2_decap_8 FILLER_4_1252 ();
 sg13g2_decap_8 FILLER_4_1259 ();
 sg13g2_decap_8 FILLER_4_1266 ();
 sg13g2_decap_8 FILLER_4_1273 ();
 sg13g2_decap_8 FILLER_4_1280 ();
 sg13g2_decap_8 FILLER_4_1287 ();
 sg13g2_decap_8 FILLER_4_1294 ();
 sg13g2_decap_8 FILLER_4_1301 ();
 sg13g2_decap_8 FILLER_4_1308 ();
 sg13g2_decap_8 FILLER_4_1315 ();
 sg13g2_decap_8 FILLER_4_1322 ();
 sg13g2_decap_8 FILLER_4_1329 ();
 sg13g2_decap_8 FILLER_4_1336 ();
 sg13g2_decap_8 FILLER_4_1343 ();
 sg13g2_decap_8 FILLER_4_1350 ();
 sg13g2_decap_8 FILLER_4_1357 ();
 sg13g2_decap_8 FILLER_4_1364 ();
 sg13g2_decap_8 FILLER_4_1371 ();
 sg13g2_decap_8 FILLER_4_1378 ();
 sg13g2_decap_8 FILLER_4_1385 ();
 sg13g2_decap_8 FILLER_4_1392 ();
 sg13g2_decap_8 FILLER_4_1399 ();
 sg13g2_decap_8 FILLER_4_1406 ();
 sg13g2_decap_8 FILLER_4_1413 ();
 sg13g2_decap_8 FILLER_4_1420 ();
 sg13g2_decap_8 FILLER_4_1427 ();
 sg13g2_decap_8 FILLER_4_1434 ();
 sg13g2_decap_8 FILLER_4_1441 ();
 sg13g2_decap_8 FILLER_4_1448 ();
 sg13g2_decap_8 FILLER_4_1455 ();
 sg13g2_decap_8 FILLER_4_1462 ();
 sg13g2_decap_8 FILLER_4_1469 ();
 sg13g2_decap_8 FILLER_4_1476 ();
 sg13g2_decap_8 FILLER_4_1483 ();
 sg13g2_decap_8 FILLER_4_1490 ();
 sg13g2_decap_8 FILLER_4_1497 ();
 sg13g2_decap_8 FILLER_4_1504 ();
 sg13g2_decap_8 FILLER_4_1511 ();
 sg13g2_decap_8 FILLER_4_1518 ();
 sg13g2_decap_8 FILLER_4_1525 ();
 sg13g2_decap_8 FILLER_4_1532 ();
 sg13g2_decap_8 FILLER_4_1539 ();
 sg13g2_decap_8 FILLER_4_1546 ();
 sg13g2_decap_8 FILLER_4_1553 ();
 sg13g2_decap_8 FILLER_4_1560 ();
 sg13g2_decap_8 FILLER_4_1567 ();
 sg13g2_decap_8 FILLER_4_1574 ();
 sg13g2_decap_8 FILLER_4_1581 ();
 sg13g2_decap_8 FILLER_4_1588 ();
 sg13g2_decap_8 FILLER_4_1595 ();
 sg13g2_decap_8 FILLER_4_1602 ();
 sg13g2_decap_8 FILLER_4_1609 ();
 sg13g2_decap_8 FILLER_4_1616 ();
 sg13g2_decap_8 FILLER_4_1623 ();
 sg13g2_decap_8 FILLER_4_1630 ();
 sg13g2_decap_8 FILLER_4_1637 ();
 sg13g2_decap_8 FILLER_4_1644 ();
 sg13g2_decap_8 FILLER_4_1651 ();
 sg13g2_decap_8 FILLER_4_1658 ();
 sg13g2_decap_8 FILLER_4_1665 ();
 sg13g2_decap_8 FILLER_4_1672 ();
 sg13g2_decap_8 FILLER_4_1679 ();
 sg13g2_decap_8 FILLER_4_1686 ();
 sg13g2_decap_8 FILLER_4_1693 ();
 sg13g2_decap_8 FILLER_4_1700 ();
 sg13g2_decap_8 FILLER_4_1707 ();
 sg13g2_decap_8 FILLER_4_1714 ();
 sg13g2_decap_8 FILLER_4_1721 ();
 sg13g2_decap_8 FILLER_4_1728 ();
 sg13g2_decap_8 FILLER_4_1735 ();
 sg13g2_decap_8 FILLER_4_1742 ();
 sg13g2_decap_8 FILLER_4_1749 ();
 sg13g2_decap_8 FILLER_4_1756 ();
 sg13g2_decap_4 FILLER_4_1763 ();
 sg13g2_fill_1 FILLER_4_1767 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_1 FILLER_5_439 ();
 sg13g2_fill_2 FILLER_5_445 ();
 sg13g2_fill_1 FILLER_5_456 ();
 sg13g2_decap_4 FILLER_5_471 ();
 sg13g2_fill_2 FILLER_5_475 ();
 sg13g2_decap_4 FILLER_5_503 ();
 sg13g2_fill_1 FILLER_5_507 ();
 sg13g2_fill_2 FILLER_5_518 ();
 sg13g2_decap_4 FILLER_5_532 ();
 sg13g2_fill_2 FILLER_5_536 ();
 sg13g2_fill_2 FILLER_5_543 ();
 sg13g2_decap_4 FILLER_5_558 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_fill_1 FILLER_5_651 ();
 sg13g2_decap_4 FILLER_5_655 ();
 sg13g2_fill_1 FILLER_5_659 ();
 sg13g2_decap_8 FILLER_5_670 ();
 sg13g2_decap_8 FILLER_5_677 ();
 sg13g2_decap_8 FILLER_5_684 ();
 sg13g2_decap_8 FILLER_5_691 ();
 sg13g2_decap_8 FILLER_5_698 ();
 sg13g2_decap_8 FILLER_5_705 ();
 sg13g2_decap_8 FILLER_5_712 ();
 sg13g2_decap_8 FILLER_5_724 ();
 sg13g2_decap_8 FILLER_5_731 ();
 sg13g2_decap_8 FILLER_5_738 ();
 sg13g2_decap_8 FILLER_5_745 ();
 sg13g2_decap_8 FILLER_5_752 ();
 sg13g2_decap_8 FILLER_5_759 ();
 sg13g2_decap_8 FILLER_5_766 ();
 sg13g2_decap_8 FILLER_5_773 ();
 sg13g2_decap_8 FILLER_5_780 ();
 sg13g2_decap_8 FILLER_5_787 ();
 sg13g2_decap_8 FILLER_5_794 ();
 sg13g2_decap_8 FILLER_5_801 ();
 sg13g2_decap_8 FILLER_5_808 ();
 sg13g2_decap_8 FILLER_5_815 ();
 sg13g2_decap_8 FILLER_5_822 ();
 sg13g2_decap_8 FILLER_5_829 ();
 sg13g2_decap_8 FILLER_5_836 ();
 sg13g2_decap_8 FILLER_5_843 ();
 sg13g2_decap_8 FILLER_5_850 ();
 sg13g2_decap_8 FILLER_5_857 ();
 sg13g2_decap_8 FILLER_5_864 ();
 sg13g2_decap_8 FILLER_5_871 ();
 sg13g2_decap_8 FILLER_5_878 ();
 sg13g2_decap_8 FILLER_5_885 ();
 sg13g2_decap_8 FILLER_5_892 ();
 sg13g2_decap_8 FILLER_5_899 ();
 sg13g2_decap_8 FILLER_5_906 ();
 sg13g2_decap_8 FILLER_5_913 ();
 sg13g2_decap_8 FILLER_5_920 ();
 sg13g2_decap_8 FILLER_5_927 ();
 sg13g2_decap_8 FILLER_5_934 ();
 sg13g2_decap_8 FILLER_5_941 ();
 sg13g2_decap_8 FILLER_5_948 ();
 sg13g2_decap_8 FILLER_5_955 ();
 sg13g2_decap_8 FILLER_5_962 ();
 sg13g2_decap_8 FILLER_5_969 ();
 sg13g2_decap_8 FILLER_5_976 ();
 sg13g2_decap_8 FILLER_5_983 ();
 sg13g2_decap_8 FILLER_5_990 ();
 sg13g2_decap_8 FILLER_5_997 ();
 sg13g2_decap_8 FILLER_5_1004 ();
 sg13g2_decap_8 FILLER_5_1011 ();
 sg13g2_decap_8 FILLER_5_1018 ();
 sg13g2_decap_8 FILLER_5_1025 ();
 sg13g2_decap_8 FILLER_5_1032 ();
 sg13g2_decap_8 FILLER_5_1039 ();
 sg13g2_decap_8 FILLER_5_1046 ();
 sg13g2_decap_8 FILLER_5_1053 ();
 sg13g2_decap_8 FILLER_5_1060 ();
 sg13g2_decap_8 FILLER_5_1067 ();
 sg13g2_decap_8 FILLER_5_1074 ();
 sg13g2_decap_8 FILLER_5_1081 ();
 sg13g2_decap_8 FILLER_5_1088 ();
 sg13g2_decap_8 FILLER_5_1095 ();
 sg13g2_decap_8 FILLER_5_1102 ();
 sg13g2_decap_8 FILLER_5_1109 ();
 sg13g2_decap_8 FILLER_5_1116 ();
 sg13g2_decap_8 FILLER_5_1123 ();
 sg13g2_decap_8 FILLER_5_1130 ();
 sg13g2_decap_8 FILLER_5_1137 ();
 sg13g2_decap_8 FILLER_5_1144 ();
 sg13g2_decap_8 FILLER_5_1151 ();
 sg13g2_decap_8 FILLER_5_1158 ();
 sg13g2_decap_8 FILLER_5_1165 ();
 sg13g2_decap_8 FILLER_5_1172 ();
 sg13g2_decap_8 FILLER_5_1179 ();
 sg13g2_decap_8 FILLER_5_1186 ();
 sg13g2_decap_8 FILLER_5_1193 ();
 sg13g2_decap_8 FILLER_5_1200 ();
 sg13g2_decap_8 FILLER_5_1207 ();
 sg13g2_decap_8 FILLER_5_1214 ();
 sg13g2_decap_8 FILLER_5_1221 ();
 sg13g2_decap_8 FILLER_5_1228 ();
 sg13g2_decap_8 FILLER_5_1235 ();
 sg13g2_decap_8 FILLER_5_1242 ();
 sg13g2_decap_8 FILLER_5_1249 ();
 sg13g2_decap_8 FILLER_5_1256 ();
 sg13g2_decap_8 FILLER_5_1263 ();
 sg13g2_decap_8 FILLER_5_1270 ();
 sg13g2_decap_8 FILLER_5_1277 ();
 sg13g2_decap_8 FILLER_5_1284 ();
 sg13g2_decap_8 FILLER_5_1291 ();
 sg13g2_decap_8 FILLER_5_1298 ();
 sg13g2_decap_8 FILLER_5_1305 ();
 sg13g2_decap_8 FILLER_5_1312 ();
 sg13g2_decap_8 FILLER_5_1319 ();
 sg13g2_decap_8 FILLER_5_1326 ();
 sg13g2_decap_8 FILLER_5_1333 ();
 sg13g2_decap_8 FILLER_5_1340 ();
 sg13g2_decap_8 FILLER_5_1347 ();
 sg13g2_decap_8 FILLER_5_1354 ();
 sg13g2_decap_8 FILLER_5_1361 ();
 sg13g2_decap_8 FILLER_5_1368 ();
 sg13g2_decap_8 FILLER_5_1375 ();
 sg13g2_decap_8 FILLER_5_1382 ();
 sg13g2_decap_8 FILLER_5_1389 ();
 sg13g2_decap_8 FILLER_5_1396 ();
 sg13g2_decap_8 FILLER_5_1403 ();
 sg13g2_decap_8 FILLER_5_1410 ();
 sg13g2_decap_8 FILLER_5_1417 ();
 sg13g2_decap_8 FILLER_5_1424 ();
 sg13g2_decap_8 FILLER_5_1431 ();
 sg13g2_decap_8 FILLER_5_1438 ();
 sg13g2_decap_8 FILLER_5_1445 ();
 sg13g2_decap_8 FILLER_5_1452 ();
 sg13g2_decap_8 FILLER_5_1459 ();
 sg13g2_decap_8 FILLER_5_1466 ();
 sg13g2_decap_8 FILLER_5_1473 ();
 sg13g2_decap_8 FILLER_5_1480 ();
 sg13g2_decap_8 FILLER_5_1487 ();
 sg13g2_decap_8 FILLER_5_1494 ();
 sg13g2_decap_8 FILLER_5_1501 ();
 sg13g2_decap_8 FILLER_5_1508 ();
 sg13g2_decap_8 FILLER_5_1515 ();
 sg13g2_decap_8 FILLER_5_1522 ();
 sg13g2_decap_8 FILLER_5_1529 ();
 sg13g2_decap_8 FILLER_5_1536 ();
 sg13g2_decap_8 FILLER_5_1543 ();
 sg13g2_decap_8 FILLER_5_1550 ();
 sg13g2_decap_8 FILLER_5_1557 ();
 sg13g2_decap_8 FILLER_5_1564 ();
 sg13g2_decap_8 FILLER_5_1571 ();
 sg13g2_decap_8 FILLER_5_1578 ();
 sg13g2_decap_8 FILLER_5_1585 ();
 sg13g2_decap_8 FILLER_5_1592 ();
 sg13g2_decap_8 FILLER_5_1599 ();
 sg13g2_decap_8 FILLER_5_1606 ();
 sg13g2_decap_8 FILLER_5_1613 ();
 sg13g2_decap_8 FILLER_5_1620 ();
 sg13g2_decap_8 FILLER_5_1627 ();
 sg13g2_decap_8 FILLER_5_1634 ();
 sg13g2_decap_8 FILLER_5_1641 ();
 sg13g2_decap_8 FILLER_5_1648 ();
 sg13g2_decap_8 FILLER_5_1655 ();
 sg13g2_decap_8 FILLER_5_1662 ();
 sg13g2_decap_8 FILLER_5_1669 ();
 sg13g2_decap_8 FILLER_5_1676 ();
 sg13g2_decap_8 FILLER_5_1683 ();
 sg13g2_decap_8 FILLER_5_1690 ();
 sg13g2_decap_8 FILLER_5_1697 ();
 sg13g2_decap_8 FILLER_5_1704 ();
 sg13g2_decap_8 FILLER_5_1711 ();
 sg13g2_decap_8 FILLER_5_1718 ();
 sg13g2_decap_8 FILLER_5_1725 ();
 sg13g2_decap_8 FILLER_5_1732 ();
 sg13g2_decap_8 FILLER_5_1739 ();
 sg13g2_decap_8 FILLER_5_1746 ();
 sg13g2_decap_8 FILLER_5_1753 ();
 sg13g2_decap_8 FILLER_5_1760 ();
 sg13g2_fill_1 FILLER_5_1767 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_4 FILLER_6_413 ();
 sg13g2_decap_4 FILLER_6_440 ();
 sg13g2_fill_2 FILLER_6_444 ();
 sg13g2_decap_8 FILLER_6_492 ();
 sg13g2_decap_4 FILLER_6_499 ();
 sg13g2_fill_2 FILLER_6_503 ();
 sg13g2_decap_8 FILLER_6_521 ();
 sg13g2_decap_4 FILLER_6_528 ();
 sg13g2_fill_1 FILLER_6_532 ();
 sg13g2_fill_1 FILLER_6_561 ();
 sg13g2_decap_8 FILLER_6_579 ();
 sg13g2_decap_8 FILLER_6_586 ();
 sg13g2_decap_8 FILLER_6_593 ();
 sg13g2_decap_4 FILLER_6_600 ();
 sg13g2_fill_2 FILLER_6_604 ();
 sg13g2_decap_8 FILLER_6_615 ();
 sg13g2_decap_8 FILLER_6_622 ();
 sg13g2_decap_8 FILLER_6_629 ();
 sg13g2_decap_8 FILLER_6_636 ();
 sg13g2_fill_2 FILLER_6_643 ();
 sg13g2_fill_2 FILLER_6_664 ();
 sg13g2_fill_1 FILLER_6_666 ();
 sg13g2_decap_8 FILLER_6_684 ();
 sg13g2_fill_2 FILLER_6_691 ();
 sg13g2_fill_1 FILLER_6_693 ();
 sg13g2_fill_2 FILLER_6_700 ();
 sg13g2_decap_4 FILLER_6_707 ();
 sg13g2_fill_1 FILLER_6_711 ();
 sg13g2_decap_4 FILLER_6_736 ();
 sg13g2_decap_8 FILLER_6_764 ();
 sg13g2_decap_8 FILLER_6_771 ();
 sg13g2_decap_8 FILLER_6_778 ();
 sg13g2_decap_8 FILLER_6_785 ();
 sg13g2_decap_8 FILLER_6_792 ();
 sg13g2_decap_8 FILLER_6_799 ();
 sg13g2_decap_8 FILLER_6_806 ();
 sg13g2_decap_8 FILLER_6_813 ();
 sg13g2_decap_8 FILLER_6_820 ();
 sg13g2_decap_8 FILLER_6_827 ();
 sg13g2_decap_8 FILLER_6_834 ();
 sg13g2_decap_8 FILLER_6_841 ();
 sg13g2_decap_8 FILLER_6_848 ();
 sg13g2_decap_8 FILLER_6_855 ();
 sg13g2_decap_8 FILLER_6_862 ();
 sg13g2_decap_8 FILLER_6_869 ();
 sg13g2_decap_8 FILLER_6_876 ();
 sg13g2_decap_8 FILLER_6_883 ();
 sg13g2_decap_8 FILLER_6_890 ();
 sg13g2_decap_8 FILLER_6_897 ();
 sg13g2_decap_8 FILLER_6_904 ();
 sg13g2_decap_8 FILLER_6_911 ();
 sg13g2_decap_8 FILLER_6_918 ();
 sg13g2_decap_8 FILLER_6_925 ();
 sg13g2_decap_8 FILLER_6_932 ();
 sg13g2_decap_8 FILLER_6_939 ();
 sg13g2_decap_8 FILLER_6_946 ();
 sg13g2_decap_8 FILLER_6_953 ();
 sg13g2_decap_8 FILLER_6_960 ();
 sg13g2_decap_8 FILLER_6_967 ();
 sg13g2_decap_8 FILLER_6_974 ();
 sg13g2_decap_8 FILLER_6_981 ();
 sg13g2_decap_8 FILLER_6_988 ();
 sg13g2_decap_8 FILLER_6_995 ();
 sg13g2_decap_8 FILLER_6_1002 ();
 sg13g2_decap_8 FILLER_6_1009 ();
 sg13g2_decap_8 FILLER_6_1016 ();
 sg13g2_decap_8 FILLER_6_1023 ();
 sg13g2_decap_8 FILLER_6_1030 ();
 sg13g2_decap_8 FILLER_6_1037 ();
 sg13g2_decap_8 FILLER_6_1044 ();
 sg13g2_decap_8 FILLER_6_1051 ();
 sg13g2_decap_8 FILLER_6_1058 ();
 sg13g2_decap_8 FILLER_6_1065 ();
 sg13g2_decap_8 FILLER_6_1072 ();
 sg13g2_decap_8 FILLER_6_1079 ();
 sg13g2_decap_8 FILLER_6_1086 ();
 sg13g2_decap_8 FILLER_6_1093 ();
 sg13g2_decap_8 FILLER_6_1100 ();
 sg13g2_decap_8 FILLER_6_1107 ();
 sg13g2_decap_8 FILLER_6_1114 ();
 sg13g2_decap_8 FILLER_6_1121 ();
 sg13g2_decap_8 FILLER_6_1128 ();
 sg13g2_decap_8 FILLER_6_1135 ();
 sg13g2_decap_8 FILLER_6_1142 ();
 sg13g2_decap_8 FILLER_6_1149 ();
 sg13g2_decap_8 FILLER_6_1156 ();
 sg13g2_decap_8 FILLER_6_1163 ();
 sg13g2_decap_8 FILLER_6_1170 ();
 sg13g2_decap_8 FILLER_6_1177 ();
 sg13g2_decap_8 FILLER_6_1184 ();
 sg13g2_decap_8 FILLER_6_1191 ();
 sg13g2_decap_8 FILLER_6_1198 ();
 sg13g2_decap_8 FILLER_6_1205 ();
 sg13g2_decap_8 FILLER_6_1212 ();
 sg13g2_decap_8 FILLER_6_1219 ();
 sg13g2_decap_8 FILLER_6_1226 ();
 sg13g2_decap_8 FILLER_6_1233 ();
 sg13g2_decap_8 FILLER_6_1240 ();
 sg13g2_decap_8 FILLER_6_1247 ();
 sg13g2_decap_8 FILLER_6_1254 ();
 sg13g2_decap_8 FILLER_6_1261 ();
 sg13g2_decap_8 FILLER_6_1268 ();
 sg13g2_decap_8 FILLER_6_1275 ();
 sg13g2_decap_8 FILLER_6_1282 ();
 sg13g2_decap_8 FILLER_6_1289 ();
 sg13g2_decap_8 FILLER_6_1296 ();
 sg13g2_decap_8 FILLER_6_1303 ();
 sg13g2_decap_8 FILLER_6_1310 ();
 sg13g2_decap_8 FILLER_6_1317 ();
 sg13g2_decap_8 FILLER_6_1324 ();
 sg13g2_decap_8 FILLER_6_1331 ();
 sg13g2_decap_8 FILLER_6_1338 ();
 sg13g2_decap_8 FILLER_6_1345 ();
 sg13g2_decap_8 FILLER_6_1352 ();
 sg13g2_decap_8 FILLER_6_1359 ();
 sg13g2_decap_8 FILLER_6_1366 ();
 sg13g2_decap_8 FILLER_6_1373 ();
 sg13g2_decap_8 FILLER_6_1380 ();
 sg13g2_decap_8 FILLER_6_1387 ();
 sg13g2_decap_8 FILLER_6_1394 ();
 sg13g2_decap_8 FILLER_6_1401 ();
 sg13g2_decap_8 FILLER_6_1408 ();
 sg13g2_decap_8 FILLER_6_1415 ();
 sg13g2_decap_8 FILLER_6_1422 ();
 sg13g2_decap_8 FILLER_6_1429 ();
 sg13g2_decap_8 FILLER_6_1436 ();
 sg13g2_decap_8 FILLER_6_1443 ();
 sg13g2_decap_8 FILLER_6_1450 ();
 sg13g2_decap_8 FILLER_6_1457 ();
 sg13g2_decap_8 FILLER_6_1464 ();
 sg13g2_decap_8 FILLER_6_1471 ();
 sg13g2_decap_8 FILLER_6_1478 ();
 sg13g2_decap_8 FILLER_6_1485 ();
 sg13g2_decap_8 FILLER_6_1492 ();
 sg13g2_decap_8 FILLER_6_1499 ();
 sg13g2_decap_8 FILLER_6_1506 ();
 sg13g2_decap_8 FILLER_6_1513 ();
 sg13g2_decap_8 FILLER_6_1520 ();
 sg13g2_decap_8 FILLER_6_1527 ();
 sg13g2_decap_8 FILLER_6_1534 ();
 sg13g2_decap_8 FILLER_6_1541 ();
 sg13g2_decap_8 FILLER_6_1548 ();
 sg13g2_decap_8 FILLER_6_1555 ();
 sg13g2_decap_8 FILLER_6_1562 ();
 sg13g2_decap_8 FILLER_6_1569 ();
 sg13g2_decap_8 FILLER_6_1576 ();
 sg13g2_decap_8 FILLER_6_1583 ();
 sg13g2_decap_8 FILLER_6_1590 ();
 sg13g2_decap_8 FILLER_6_1597 ();
 sg13g2_decap_8 FILLER_6_1604 ();
 sg13g2_decap_8 FILLER_6_1611 ();
 sg13g2_decap_8 FILLER_6_1618 ();
 sg13g2_decap_8 FILLER_6_1625 ();
 sg13g2_decap_8 FILLER_6_1632 ();
 sg13g2_decap_8 FILLER_6_1639 ();
 sg13g2_decap_8 FILLER_6_1646 ();
 sg13g2_decap_8 FILLER_6_1653 ();
 sg13g2_decap_8 FILLER_6_1660 ();
 sg13g2_decap_8 FILLER_6_1667 ();
 sg13g2_decap_8 FILLER_6_1674 ();
 sg13g2_decap_8 FILLER_6_1681 ();
 sg13g2_decap_8 FILLER_6_1688 ();
 sg13g2_decap_8 FILLER_6_1695 ();
 sg13g2_decap_8 FILLER_6_1702 ();
 sg13g2_decap_8 FILLER_6_1709 ();
 sg13g2_decap_8 FILLER_6_1716 ();
 sg13g2_decap_8 FILLER_6_1723 ();
 sg13g2_decap_8 FILLER_6_1730 ();
 sg13g2_decap_8 FILLER_6_1737 ();
 sg13g2_decap_8 FILLER_6_1744 ();
 sg13g2_decap_8 FILLER_6_1751 ();
 sg13g2_decap_8 FILLER_6_1758 ();
 sg13g2_fill_2 FILLER_6_1765 ();
 sg13g2_fill_1 FILLER_6_1767 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_fill_2 FILLER_7_343 ();
 sg13g2_fill_1 FILLER_7_345 ();
 sg13g2_decap_8 FILLER_7_359 ();
 sg13g2_decap_8 FILLER_7_366 ();
 sg13g2_decap_8 FILLER_7_373 ();
 sg13g2_fill_2 FILLER_7_380 ();
 sg13g2_decap_4 FILLER_7_408 ();
 sg13g2_fill_1 FILLER_7_412 ();
 sg13g2_fill_1 FILLER_7_443 ();
 sg13g2_fill_2 FILLER_7_454 ();
 sg13g2_decap_8 FILLER_7_466 ();
 sg13g2_decap_4 FILLER_7_473 ();
 sg13g2_fill_1 FILLER_7_477 ();
 sg13g2_fill_2 FILLER_7_493 ();
 sg13g2_fill_1 FILLER_7_507 ();
 sg13g2_decap_4 FILLER_7_526 ();
 sg13g2_fill_2 FILLER_7_530 ();
 sg13g2_fill_2 FILLER_7_549 ();
 sg13g2_fill_1 FILLER_7_551 ();
 sg13g2_fill_2 FILLER_7_556 ();
 sg13g2_decap_8 FILLER_7_576 ();
 sg13g2_decap_8 FILLER_7_583 ();
 sg13g2_decap_8 FILLER_7_590 ();
 sg13g2_fill_2 FILLER_7_597 ();
 sg13g2_decap_8 FILLER_7_625 ();
 sg13g2_decap_8 FILLER_7_632 ();
 sg13g2_fill_2 FILLER_7_639 ();
 sg13g2_fill_1 FILLER_7_641 ();
 sg13g2_fill_2 FILLER_7_664 ();
 sg13g2_fill_1 FILLER_7_666 ();
 sg13g2_fill_2 FILLER_7_733 ();
 sg13g2_decap_4 FILLER_7_740 ();
 sg13g2_decap_4 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_785 ();
 sg13g2_decap_8 FILLER_7_792 ();
 sg13g2_decap_8 FILLER_7_799 ();
 sg13g2_decap_8 FILLER_7_806 ();
 sg13g2_decap_8 FILLER_7_813 ();
 sg13g2_decap_8 FILLER_7_820 ();
 sg13g2_decap_8 FILLER_7_827 ();
 sg13g2_decap_8 FILLER_7_834 ();
 sg13g2_decap_8 FILLER_7_841 ();
 sg13g2_decap_8 FILLER_7_848 ();
 sg13g2_decap_8 FILLER_7_855 ();
 sg13g2_decap_8 FILLER_7_862 ();
 sg13g2_decap_8 FILLER_7_869 ();
 sg13g2_decap_8 FILLER_7_876 ();
 sg13g2_decap_8 FILLER_7_883 ();
 sg13g2_decap_8 FILLER_7_890 ();
 sg13g2_decap_8 FILLER_7_897 ();
 sg13g2_decap_8 FILLER_7_904 ();
 sg13g2_decap_8 FILLER_7_911 ();
 sg13g2_decap_8 FILLER_7_918 ();
 sg13g2_decap_8 FILLER_7_925 ();
 sg13g2_decap_8 FILLER_7_932 ();
 sg13g2_decap_8 FILLER_7_939 ();
 sg13g2_decap_8 FILLER_7_946 ();
 sg13g2_decap_8 FILLER_7_953 ();
 sg13g2_decap_8 FILLER_7_960 ();
 sg13g2_decap_8 FILLER_7_967 ();
 sg13g2_decap_8 FILLER_7_974 ();
 sg13g2_decap_8 FILLER_7_981 ();
 sg13g2_decap_8 FILLER_7_988 ();
 sg13g2_decap_8 FILLER_7_995 ();
 sg13g2_decap_8 FILLER_7_1002 ();
 sg13g2_decap_8 FILLER_7_1009 ();
 sg13g2_decap_8 FILLER_7_1016 ();
 sg13g2_decap_8 FILLER_7_1023 ();
 sg13g2_decap_8 FILLER_7_1030 ();
 sg13g2_decap_8 FILLER_7_1037 ();
 sg13g2_decap_8 FILLER_7_1044 ();
 sg13g2_decap_8 FILLER_7_1051 ();
 sg13g2_decap_8 FILLER_7_1058 ();
 sg13g2_decap_8 FILLER_7_1065 ();
 sg13g2_decap_8 FILLER_7_1072 ();
 sg13g2_decap_8 FILLER_7_1079 ();
 sg13g2_decap_8 FILLER_7_1086 ();
 sg13g2_decap_8 FILLER_7_1093 ();
 sg13g2_decap_8 FILLER_7_1100 ();
 sg13g2_decap_8 FILLER_7_1107 ();
 sg13g2_decap_8 FILLER_7_1114 ();
 sg13g2_decap_8 FILLER_7_1121 ();
 sg13g2_decap_8 FILLER_7_1128 ();
 sg13g2_decap_8 FILLER_7_1135 ();
 sg13g2_decap_8 FILLER_7_1142 ();
 sg13g2_decap_8 FILLER_7_1149 ();
 sg13g2_decap_8 FILLER_7_1156 ();
 sg13g2_decap_8 FILLER_7_1163 ();
 sg13g2_decap_8 FILLER_7_1170 ();
 sg13g2_decap_8 FILLER_7_1177 ();
 sg13g2_decap_8 FILLER_7_1184 ();
 sg13g2_decap_8 FILLER_7_1191 ();
 sg13g2_decap_8 FILLER_7_1198 ();
 sg13g2_decap_8 FILLER_7_1205 ();
 sg13g2_decap_8 FILLER_7_1212 ();
 sg13g2_decap_8 FILLER_7_1219 ();
 sg13g2_decap_8 FILLER_7_1226 ();
 sg13g2_decap_8 FILLER_7_1233 ();
 sg13g2_decap_8 FILLER_7_1240 ();
 sg13g2_decap_8 FILLER_7_1247 ();
 sg13g2_decap_8 FILLER_7_1254 ();
 sg13g2_decap_8 FILLER_7_1261 ();
 sg13g2_decap_8 FILLER_7_1268 ();
 sg13g2_decap_8 FILLER_7_1275 ();
 sg13g2_decap_8 FILLER_7_1282 ();
 sg13g2_decap_8 FILLER_7_1289 ();
 sg13g2_decap_8 FILLER_7_1296 ();
 sg13g2_decap_8 FILLER_7_1303 ();
 sg13g2_decap_8 FILLER_7_1310 ();
 sg13g2_decap_8 FILLER_7_1317 ();
 sg13g2_decap_8 FILLER_7_1324 ();
 sg13g2_decap_8 FILLER_7_1331 ();
 sg13g2_decap_8 FILLER_7_1338 ();
 sg13g2_decap_8 FILLER_7_1345 ();
 sg13g2_decap_8 FILLER_7_1352 ();
 sg13g2_decap_8 FILLER_7_1359 ();
 sg13g2_decap_8 FILLER_7_1366 ();
 sg13g2_decap_8 FILLER_7_1373 ();
 sg13g2_decap_8 FILLER_7_1380 ();
 sg13g2_decap_8 FILLER_7_1387 ();
 sg13g2_decap_8 FILLER_7_1394 ();
 sg13g2_decap_8 FILLER_7_1401 ();
 sg13g2_decap_8 FILLER_7_1408 ();
 sg13g2_decap_8 FILLER_7_1415 ();
 sg13g2_decap_8 FILLER_7_1422 ();
 sg13g2_decap_8 FILLER_7_1429 ();
 sg13g2_decap_8 FILLER_7_1436 ();
 sg13g2_decap_8 FILLER_7_1443 ();
 sg13g2_decap_8 FILLER_7_1450 ();
 sg13g2_decap_8 FILLER_7_1457 ();
 sg13g2_decap_8 FILLER_7_1464 ();
 sg13g2_decap_8 FILLER_7_1471 ();
 sg13g2_decap_8 FILLER_7_1478 ();
 sg13g2_decap_8 FILLER_7_1485 ();
 sg13g2_decap_8 FILLER_7_1492 ();
 sg13g2_decap_8 FILLER_7_1499 ();
 sg13g2_decap_8 FILLER_7_1506 ();
 sg13g2_decap_8 FILLER_7_1513 ();
 sg13g2_decap_8 FILLER_7_1520 ();
 sg13g2_decap_8 FILLER_7_1527 ();
 sg13g2_decap_8 FILLER_7_1534 ();
 sg13g2_decap_8 FILLER_7_1541 ();
 sg13g2_decap_8 FILLER_7_1548 ();
 sg13g2_decap_8 FILLER_7_1555 ();
 sg13g2_decap_8 FILLER_7_1562 ();
 sg13g2_decap_8 FILLER_7_1569 ();
 sg13g2_decap_8 FILLER_7_1576 ();
 sg13g2_decap_8 FILLER_7_1583 ();
 sg13g2_decap_8 FILLER_7_1590 ();
 sg13g2_decap_8 FILLER_7_1597 ();
 sg13g2_decap_8 FILLER_7_1604 ();
 sg13g2_decap_8 FILLER_7_1611 ();
 sg13g2_decap_8 FILLER_7_1618 ();
 sg13g2_decap_8 FILLER_7_1625 ();
 sg13g2_decap_8 FILLER_7_1632 ();
 sg13g2_decap_8 FILLER_7_1639 ();
 sg13g2_decap_8 FILLER_7_1646 ();
 sg13g2_decap_8 FILLER_7_1653 ();
 sg13g2_decap_8 FILLER_7_1660 ();
 sg13g2_decap_8 FILLER_7_1667 ();
 sg13g2_decap_8 FILLER_7_1674 ();
 sg13g2_decap_8 FILLER_7_1681 ();
 sg13g2_decap_8 FILLER_7_1688 ();
 sg13g2_decap_8 FILLER_7_1695 ();
 sg13g2_decap_8 FILLER_7_1702 ();
 sg13g2_decap_8 FILLER_7_1709 ();
 sg13g2_decap_8 FILLER_7_1716 ();
 sg13g2_decap_8 FILLER_7_1723 ();
 sg13g2_decap_8 FILLER_7_1730 ();
 sg13g2_decap_8 FILLER_7_1737 ();
 sg13g2_decap_8 FILLER_7_1744 ();
 sg13g2_decap_8 FILLER_7_1751 ();
 sg13g2_decap_8 FILLER_7_1758 ();
 sg13g2_fill_2 FILLER_7_1765 ();
 sg13g2_fill_1 FILLER_7_1767 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_fill_2 FILLER_8_273 ();
 sg13g2_fill_1 FILLER_8_275 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_4 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_316 ();
 sg13g2_decap_4 FILLER_8_323 ();
 sg13g2_fill_2 FILLER_8_361 ();
 sg13g2_fill_2 FILLER_8_371 ();
 sg13g2_fill_1 FILLER_8_373 ();
 sg13g2_fill_1 FILLER_8_378 ();
 sg13g2_fill_1 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_438 ();
 sg13g2_decap_8 FILLER_8_445 ();
 sg13g2_fill_1 FILLER_8_452 ();
 sg13g2_fill_1 FILLER_8_466 ();
 sg13g2_decap_4 FILLER_8_499 ();
 sg13g2_fill_2 FILLER_8_503 ();
 sg13g2_fill_1 FILLER_8_525 ();
 sg13g2_fill_2 FILLER_8_548 ();
 sg13g2_fill_1 FILLER_8_550 ();
 sg13g2_fill_2 FILLER_8_567 ();
 sg13g2_fill_1 FILLER_8_569 ();
 sg13g2_decap_8 FILLER_8_583 ();
 sg13g2_decap_8 FILLER_8_590 ();
 sg13g2_fill_2 FILLER_8_606 ();
 sg13g2_fill_2 FILLER_8_634 ();
 sg13g2_fill_1 FILLER_8_636 ();
 sg13g2_decap_8 FILLER_8_690 ();
 sg13g2_decap_4 FILLER_8_697 ();
 sg13g2_fill_2 FILLER_8_711 ();
 sg13g2_decap_8 FILLER_8_718 ();
 sg13g2_fill_2 FILLER_8_760 ();
 sg13g2_fill_1 FILLER_8_762 ();
 sg13g2_decap_8 FILLER_8_789 ();
 sg13g2_decap_8 FILLER_8_796 ();
 sg13g2_decap_8 FILLER_8_803 ();
 sg13g2_decap_8 FILLER_8_810 ();
 sg13g2_decap_8 FILLER_8_817 ();
 sg13g2_decap_8 FILLER_8_824 ();
 sg13g2_decap_8 FILLER_8_831 ();
 sg13g2_decap_8 FILLER_8_838 ();
 sg13g2_decap_8 FILLER_8_845 ();
 sg13g2_decap_8 FILLER_8_852 ();
 sg13g2_decap_8 FILLER_8_859 ();
 sg13g2_decap_8 FILLER_8_866 ();
 sg13g2_decap_8 FILLER_8_873 ();
 sg13g2_decap_8 FILLER_8_880 ();
 sg13g2_decap_8 FILLER_8_887 ();
 sg13g2_decap_8 FILLER_8_894 ();
 sg13g2_decap_8 FILLER_8_901 ();
 sg13g2_decap_8 FILLER_8_908 ();
 sg13g2_decap_8 FILLER_8_915 ();
 sg13g2_decap_8 FILLER_8_922 ();
 sg13g2_decap_8 FILLER_8_929 ();
 sg13g2_decap_8 FILLER_8_936 ();
 sg13g2_decap_8 FILLER_8_943 ();
 sg13g2_decap_8 FILLER_8_950 ();
 sg13g2_decap_8 FILLER_8_957 ();
 sg13g2_decap_8 FILLER_8_964 ();
 sg13g2_decap_8 FILLER_8_971 ();
 sg13g2_decap_8 FILLER_8_978 ();
 sg13g2_decap_8 FILLER_8_985 ();
 sg13g2_decap_8 FILLER_8_992 ();
 sg13g2_decap_8 FILLER_8_999 ();
 sg13g2_decap_8 FILLER_8_1006 ();
 sg13g2_decap_8 FILLER_8_1013 ();
 sg13g2_decap_8 FILLER_8_1020 ();
 sg13g2_decap_8 FILLER_8_1027 ();
 sg13g2_decap_8 FILLER_8_1034 ();
 sg13g2_decap_8 FILLER_8_1041 ();
 sg13g2_decap_8 FILLER_8_1048 ();
 sg13g2_decap_8 FILLER_8_1055 ();
 sg13g2_decap_8 FILLER_8_1062 ();
 sg13g2_decap_8 FILLER_8_1069 ();
 sg13g2_decap_8 FILLER_8_1076 ();
 sg13g2_decap_8 FILLER_8_1083 ();
 sg13g2_decap_8 FILLER_8_1090 ();
 sg13g2_decap_8 FILLER_8_1097 ();
 sg13g2_decap_8 FILLER_8_1104 ();
 sg13g2_decap_8 FILLER_8_1111 ();
 sg13g2_decap_8 FILLER_8_1118 ();
 sg13g2_decap_8 FILLER_8_1125 ();
 sg13g2_decap_8 FILLER_8_1132 ();
 sg13g2_decap_8 FILLER_8_1139 ();
 sg13g2_decap_8 FILLER_8_1146 ();
 sg13g2_decap_8 FILLER_8_1153 ();
 sg13g2_decap_8 FILLER_8_1160 ();
 sg13g2_decap_8 FILLER_8_1167 ();
 sg13g2_decap_8 FILLER_8_1174 ();
 sg13g2_decap_8 FILLER_8_1181 ();
 sg13g2_decap_8 FILLER_8_1188 ();
 sg13g2_decap_8 FILLER_8_1195 ();
 sg13g2_decap_8 FILLER_8_1202 ();
 sg13g2_decap_8 FILLER_8_1209 ();
 sg13g2_decap_8 FILLER_8_1216 ();
 sg13g2_decap_8 FILLER_8_1223 ();
 sg13g2_decap_8 FILLER_8_1230 ();
 sg13g2_decap_8 FILLER_8_1237 ();
 sg13g2_decap_8 FILLER_8_1244 ();
 sg13g2_decap_8 FILLER_8_1251 ();
 sg13g2_decap_8 FILLER_8_1258 ();
 sg13g2_decap_8 FILLER_8_1265 ();
 sg13g2_decap_8 FILLER_8_1272 ();
 sg13g2_decap_8 FILLER_8_1279 ();
 sg13g2_decap_8 FILLER_8_1286 ();
 sg13g2_decap_8 FILLER_8_1293 ();
 sg13g2_decap_8 FILLER_8_1300 ();
 sg13g2_decap_8 FILLER_8_1307 ();
 sg13g2_decap_8 FILLER_8_1314 ();
 sg13g2_decap_8 FILLER_8_1321 ();
 sg13g2_decap_8 FILLER_8_1328 ();
 sg13g2_decap_8 FILLER_8_1335 ();
 sg13g2_decap_8 FILLER_8_1342 ();
 sg13g2_decap_8 FILLER_8_1349 ();
 sg13g2_decap_8 FILLER_8_1356 ();
 sg13g2_decap_8 FILLER_8_1363 ();
 sg13g2_decap_8 FILLER_8_1370 ();
 sg13g2_decap_8 FILLER_8_1377 ();
 sg13g2_decap_8 FILLER_8_1384 ();
 sg13g2_decap_8 FILLER_8_1391 ();
 sg13g2_decap_8 FILLER_8_1398 ();
 sg13g2_decap_8 FILLER_8_1405 ();
 sg13g2_decap_8 FILLER_8_1412 ();
 sg13g2_decap_8 FILLER_8_1419 ();
 sg13g2_decap_8 FILLER_8_1426 ();
 sg13g2_decap_8 FILLER_8_1433 ();
 sg13g2_decap_8 FILLER_8_1440 ();
 sg13g2_decap_8 FILLER_8_1447 ();
 sg13g2_decap_8 FILLER_8_1454 ();
 sg13g2_decap_8 FILLER_8_1461 ();
 sg13g2_decap_8 FILLER_8_1468 ();
 sg13g2_decap_8 FILLER_8_1475 ();
 sg13g2_decap_8 FILLER_8_1482 ();
 sg13g2_decap_8 FILLER_8_1489 ();
 sg13g2_decap_8 FILLER_8_1496 ();
 sg13g2_decap_8 FILLER_8_1503 ();
 sg13g2_decap_8 FILLER_8_1510 ();
 sg13g2_decap_8 FILLER_8_1517 ();
 sg13g2_decap_8 FILLER_8_1524 ();
 sg13g2_decap_8 FILLER_8_1531 ();
 sg13g2_decap_8 FILLER_8_1538 ();
 sg13g2_decap_8 FILLER_8_1545 ();
 sg13g2_decap_8 FILLER_8_1552 ();
 sg13g2_decap_8 FILLER_8_1559 ();
 sg13g2_decap_8 FILLER_8_1566 ();
 sg13g2_decap_8 FILLER_8_1573 ();
 sg13g2_decap_8 FILLER_8_1580 ();
 sg13g2_decap_8 FILLER_8_1587 ();
 sg13g2_decap_8 FILLER_8_1594 ();
 sg13g2_decap_8 FILLER_8_1601 ();
 sg13g2_decap_8 FILLER_8_1608 ();
 sg13g2_decap_8 FILLER_8_1615 ();
 sg13g2_decap_8 FILLER_8_1622 ();
 sg13g2_decap_8 FILLER_8_1629 ();
 sg13g2_decap_8 FILLER_8_1636 ();
 sg13g2_decap_8 FILLER_8_1643 ();
 sg13g2_decap_8 FILLER_8_1650 ();
 sg13g2_decap_8 FILLER_8_1657 ();
 sg13g2_decap_8 FILLER_8_1664 ();
 sg13g2_decap_8 FILLER_8_1671 ();
 sg13g2_decap_8 FILLER_8_1678 ();
 sg13g2_decap_8 FILLER_8_1685 ();
 sg13g2_decap_8 FILLER_8_1692 ();
 sg13g2_decap_8 FILLER_8_1699 ();
 sg13g2_decap_8 FILLER_8_1706 ();
 sg13g2_decap_8 FILLER_8_1713 ();
 sg13g2_decap_8 FILLER_8_1720 ();
 sg13g2_decap_8 FILLER_8_1727 ();
 sg13g2_decap_8 FILLER_8_1734 ();
 sg13g2_decap_8 FILLER_8_1741 ();
 sg13g2_decap_8 FILLER_8_1748 ();
 sg13g2_decap_8 FILLER_8_1755 ();
 sg13g2_decap_4 FILLER_8_1762 ();
 sg13g2_fill_2 FILLER_8_1766 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_4 FILLER_9_91 ();
 sg13g2_fill_1 FILLER_9_95 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_4 FILLER_9_126 ();
 sg13g2_fill_2 FILLER_9_130 ();
 sg13g2_fill_2 FILLER_9_141 ();
 sg13g2_fill_1 FILLER_9_143 ();
 sg13g2_decap_8 FILLER_9_148 ();
 sg13g2_decap_8 FILLER_9_155 ();
 sg13g2_decap_8 FILLER_9_162 ();
 sg13g2_decap_8 FILLER_9_169 ();
 sg13g2_decap_8 FILLER_9_176 ();
 sg13g2_decap_8 FILLER_9_183 ();
 sg13g2_decap_8 FILLER_9_190 ();
 sg13g2_decap_8 FILLER_9_197 ();
 sg13g2_decap_4 FILLER_9_204 ();
 sg13g2_fill_2 FILLER_9_208 ();
 sg13g2_fill_2 FILLER_9_236 ();
 sg13g2_fill_1 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_248 ();
 sg13g2_decap_4 FILLER_9_255 ();
 sg13g2_fill_2 FILLER_9_259 ();
 sg13g2_fill_1 FILLER_9_274 ();
 sg13g2_fill_1 FILLER_9_343 ();
 sg13g2_fill_1 FILLER_9_371 ();
 sg13g2_fill_2 FILLER_9_418 ();
 sg13g2_fill_1 FILLER_9_430 ();
 sg13g2_fill_2 FILLER_9_435 ();
 sg13g2_fill_1 FILLER_9_437 ();
 sg13g2_fill_1 FILLER_9_465 ();
 sg13g2_fill_1 FILLER_9_471 ();
 sg13g2_decap_8 FILLER_9_486 ();
 sg13g2_decap_4 FILLER_9_493 ();
 sg13g2_fill_2 FILLER_9_497 ();
 sg13g2_fill_1 FILLER_9_504 ();
 sg13g2_decap_4 FILLER_9_518 ();
 sg13g2_fill_1 FILLER_9_522 ();
 sg13g2_decap_8 FILLER_9_535 ();
 sg13g2_decap_8 FILLER_9_550 ();
 sg13g2_decap_4 FILLER_9_557 ();
 sg13g2_fill_2 FILLER_9_561 ();
 sg13g2_fill_1 FILLER_9_571 ();
 sg13g2_fill_2 FILLER_9_577 ();
 sg13g2_fill_2 FILLER_9_605 ();
 sg13g2_fill_2 FILLER_9_616 ();
 sg13g2_fill_2 FILLER_9_628 ();
 sg13g2_fill_2 FILLER_9_639 ();
 sg13g2_fill_1 FILLER_9_641 ();
 sg13g2_fill_2 FILLER_9_651 ();
 sg13g2_fill_2 FILLER_9_657 ();
 sg13g2_decap_4 FILLER_9_671 ();
 sg13g2_fill_2 FILLER_9_675 ();
 sg13g2_fill_2 FILLER_9_706 ();
 sg13g2_fill_2 FILLER_9_720 ();
 sg13g2_decap_4 FILLER_9_734 ();
 sg13g2_fill_2 FILLER_9_738 ();
 sg13g2_fill_1 FILLER_9_743 ();
 sg13g2_decap_4 FILLER_9_757 ();
 sg13g2_decap_8 FILLER_9_765 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_decap_8 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_9_868 ();
 sg13g2_decap_8 FILLER_9_875 ();
 sg13g2_decap_8 FILLER_9_882 ();
 sg13g2_decap_8 FILLER_9_889 ();
 sg13g2_decap_8 FILLER_9_896 ();
 sg13g2_decap_8 FILLER_9_903 ();
 sg13g2_decap_8 FILLER_9_910 ();
 sg13g2_decap_8 FILLER_9_917 ();
 sg13g2_decap_8 FILLER_9_924 ();
 sg13g2_decap_8 FILLER_9_931 ();
 sg13g2_decap_8 FILLER_9_938 ();
 sg13g2_decap_8 FILLER_9_945 ();
 sg13g2_decap_8 FILLER_9_952 ();
 sg13g2_decap_8 FILLER_9_959 ();
 sg13g2_decap_8 FILLER_9_966 ();
 sg13g2_decap_8 FILLER_9_973 ();
 sg13g2_decap_8 FILLER_9_980 ();
 sg13g2_decap_8 FILLER_9_987 ();
 sg13g2_decap_8 FILLER_9_994 ();
 sg13g2_decap_8 FILLER_9_1001 ();
 sg13g2_decap_8 FILLER_9_1008 ();
 sg13g2_decap_8 FILLER_9_1015 ();
 sg13g2_decap_8 FILLER_9_1022 ();
 sg13g2_decap_8 FILLER_9_1029 ();
 sg13g2_decap_8 FILLER_9_1036 ();
 sg13g2_decap_8 FILLER_9_1043 ();
 sg13g2_decap_8 FILLER_9_1050 ();
 sg13g2_decap_8 FILLER_9_1057 ();
 sg13g2_decap_8 FILLER_9_1064 ();
 sg13g2_decap_8 FILLER_9_1071 ();
 sg13g2_decap_8 FILLER_9_1078 ();
 sg13g2_decap_8 FILLER_9_1085 ();
 sg13g2_decap_8 FILLER_9_1092 ();
 sg13g2_decap_8 FILLER_9_1099 ();
 sg13g2_decap_8 FILLER_9_1106 ();
 sg13g2_decap_8 FILLER_9_1113 ();
 sg13g2_decap_8 FILLER_9_1120 ();
 sg13g2_decap_8 FILLER_9_1127 ();
 sg13g2_decap_8 FILLER_9_1134 ();
 sg13g2_decap_8 FILLER_9_1141 ();
 sg13g2_decap_8 FILLER_9_1148 ();
 sg13g2_decap_8 FILLER_9_1155 ();
 sg13g2_decap_8 FILLER_9_1162 ();
 sg13g2_decap_8 FILLER_9_1169 ();
 sg13g2_decap_8 FILLER_9_1176 ();
 sg13g2_decap_8 FILLER_9_1183 ();
 sg13g2_decap_8 FILLER_9_1190 ();
 sg13g2_decap_8 FILLER_9_1197 ();
 sg13g2_decap_8 FILLER_9_1204 ();
 sg13g2_decap_8 FILLER_9_1211 ();
 sg13g2_decap_8 FILLER_9_1218 ();
 sg13g2_decap_8 FILLER_9_1225 ();
 sg13g2_decap_8 FILLER_9_1232 ();
 sg13g2_decap_8 FILLER_9_1239 ();
 sg13g2_decap_8 FILLER_9_1246 ();
 sg13g2_decap_8 FILLER_9_1253 ();
 sg13g2_decap_8 FILLER_9_1260 ();
 sg13g2_decap_8 FILLER_9_1267 ();
 sg13g2_decap_8 FILLER_9_1274 ();
 sg13g2_decap_8 FILLER_9_1281 ();
 sg13g2_decap_8 FILLER_9_1288 ();
 sg13g2_decap_8 FILLER_9_1295 ();
 sg13g2_decap_8 FILLER_9_1302 ();
 sg13g2_decap_8 FILLER_9_1309 ();
 sg13g2_decap_8 FILLER_9_1316 ();
 sg13g2_decap_8 FILLER_9_1323 ();
 sg13g2_decap_8 FILLER_9_1330 ();
 sg13g2_decap_8 FILLER_9_1337 ();
 sg13g2_decap_8 FILLER_9_1344 ();
 sg13g2_decap_8 FILLER_9_1351 ();
 sg13g2_decap_8 FILLER_9_1358 ();
 sg13g2_decap_8 FILLER_9_1365 ();
 sg13g2_decap_8 FILLER_9_1372 ();
 sg13g2_decap_8 FILLER_9_1379 ();
 sg13g2_decap_8 FILLER_9_1386 ();
 sg13g2_decap_8 FILLER_9_1393 ();
 sg13g2_decap_8 FILLER_9_1400 ();
 sg13g2_decap_8 FILLER_9_1407 ();
 sg13g2_decap_8 FILLER_9_1414 ();
 sg13g2_decap_8 FILLER_9_1421 ();
 sg13g2_decap_8 FILLER_9_1428 ();
 sg13g2_decap_8 FILLER_9_1435 ();
 sg13g2_decap_8 FILLER_9_1442 ();
 sg13g2_decap_8 FILLER_9_1449 ();
 sg13g2_decap_8 FILLER_9_1456 ();
 sg13g2_decap_8 FILLER_9_1463 ();
 sg13g2_decap_8 FILLER_9_1470 ();
 sg13g2_decap_8 FILLER_9_1477 ();
 sg13g2_decap_8 FILLER_9_1484 ();
 sg13g2_decap_8 FILLER_9_1491 ();
 sg13g2_decap_8 FILLER_9_1498 ();
 sg13g2_decap_8 FILLER_9_1505 ();
 sg13g2_decap_8 FILLER_9_1512 ();
 sg13g2_decap_8 FILLER_9_1519 ();
 sg13g2_decap_8 FILLER_9_1526 ();
 sg13g2_decap_8 FILLER_9_1533 ();
 sg13g2_decap_8 FILLER_9_1540 ();
 sg13g2_decap_8 FILLER_9_1547 ();
 sg13g2_decap_8 FILLER_9_1554 ();
 sg13g2_decap_8 FILLER_9_1561 ();
 sg13g2_decap_8 FILLER_9_1568 ();
 sg13g2_decap_8 FILLER_9_1575 ();
 sg13g2_decap_8 FILLER_9_1582 ();
 sg13g2_decap_8 FILLER_9_1589 ();
 sg13g2_decap_8 FILLER_9_1596 ();
 sg13g2_decap_8 FILLER_9_1603 ();
 sg13g2_decap_8 FILLER_9_1610 ();
 sg13g2_decap_8 FILLER_9_1617 ();
 sg13g2_decap_8 FILLER_9_1624 ();
 sg13g2_decap_8 FILLER_9_1631 ();
 sg13g2_decap_8 FILLER_9_1638 ();
 sg13g2_decap_8 FILLER_9_1645 ();
 sg13g2_decap_8 FILLER_9_1652 ();
 sg13g2_decap_8 FILLER_9_1659 ();
 sg13g2_decap_8 FILLER_9_1666 ();
 sg13g2_decap_8 FILLER_9_1673 ();
 sg13g2_decap_8 FILLER_9_1680 ();
 sg13g2_decap_8 FILLER_9_1687 ();
 sg13g2_decap_8 FILLER_9_1694 ();
 sg13g2_decap_8 FILLER_9_1701 ();
 sg13g2_decap_8 FILLER_9_1708 ();
 sg13g2_decap_8 FILLER_9_1715 ();
 sg13g2_decap_8 FILLER_9_1722 ();
 sg13g2_decap_8 FILLER_9_1729 ();
 sg13g2_decap_8 FILLER_9_1736 ();
 sg13g2_decap_8 FILLER_9_1743 ();
 sg13g2_decap_8 FILLER_9_1750 ();
 sg13g2_decap_8 FILLER_9_1757 ();
 sg13g2_decap_4 FILLER_9_1764 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_fill_2 FILLER_10_63 ();
 sg13g2_fill_2 FILLER_10_74 ();
 sg13g2_fill_1 FILLER_10_76 ();
 sg13g2_decap_8 FILLER_10_81 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_fill_2 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_fill_2 FILLER_10_130 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_decap_8 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_172 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_fill_1 FILLER_10_200 ();
 sg13g2_fill_1 FILLER_10_211 ();
 sg13g2_fill_2 FILLER_10_229 ();
 sg13g2_decap_4 FILLER_10_241 ();
 sg13g2_fill_1 FILLER_10_245 ();
 sg13g2_fill_2 FILLER_10_345 ();
 sg13g2_fill_2 FILLER_10_394 ();
 sg13g2_fill_1 FILLER_10_396 ();
 sg13g2_fill_2 FILLER_10_449 ();
 sg13g2_fill_2 FILLER_10_473 ();
 sg13g2_decap_8 FILLER_10_487 ();
 sg13g2_fill_1 FILLER_10_494 ();
 sg13g2_fill_1 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_517 ();
 sg13g2_fill_2 FILLER_10_524 ();
 sg13g2_fill_1 FILLER_10_526 ();
 sg13g2_decap_8 FILLER_10_548 ();
 sg13g2_decap_8 FILLER_10_568 ();
 sg13g2_decap_8 FILLER_10_575 ();
 sg13g2_fill_1 FILLER_10_582 ();
 sg13g2_decap_4 FILLER_10_626 ();
 sg13g2_fill_1 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_655 ();
 sg13g2_fill_2 FILLER_10_676 ();
 sg13g2_fill_1 FILLER_10_678 ();
 sg13g2_decap_4 FILLER_10_684 ();
 sg13g2_fill_1 FILLER_10_688 ();
 sg13g2_decap_8 FILLER_10_708 ();
 sg13g2_decap_4 FILLER_10_715 ();
 sg13g2_fill_2 FILLER_10_719 ();
 sg13g2_decap_8 FILLER_10_726 ();
 sg13g2_decap_4 FILLER_10_750 ();
 sg13g2_fill_1 FILLER_10_754 ();
 sg13g2_decap_4 FILLER_10_767 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_decap_8 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_10_868 ();
 sg13g2_decap_8 FILLER_10_875 ();
 sg13g2_decap_8 FILLER_10_882 ();
 sg13g2_decap_8 FILLER_10_889 ();
 sg13g2_decap_8 FILLER_10_896 ();
 sg13g2_decap_8 FILLER_10_903 ();
 sg13g2_decap_8 FILLER_10_910 ();
 sg13g2_decap_8 FILLER_10_917 ();
 sg13g2_decap_8 FILLER_10_924 ();
 sg13g2_decap_8 FILLER_10_931 ();
 sg13g2_decap_8 FILLER_10_938 ();
 sg13g2_decap_8 FILLER_10_945 ();
 sg13g2_decap_8 FILLER_10_952 ();
 sg13g2_decap_8 FILLER_10_959 ();
 sg13g2_decap_8 FILLER_10_966 ();
 sg13g2_decap_8 FILLER_10_973 ();
 sg13g2_decap_8 FILLER_10_980 ();
 sg13g2_decap_8 FILLER_10_987 ();
 sg13g2_decap_8 FILLER_10_994 ();
 sg13g2_decap_8 FILLER_10_1001 ();
 sg13g2_decap_8 FILLER_10_1008 ();
 sg13g2_decap_8 FILLER_10_1015 ();
 sg13g2_decap_8 FILLER_10_1022 ();
 sg13g2_decap_8 FILLER_10_1029 ();
 sg13g2_decap_8 FILLER_10_1036 ();
 sg13g2_decap_8 FILLER_10_1043 ();
 sg13g2_decap_8 FILLER_10_1050 ();
 sg13g2_decap_8 FILLER_10_1057 ();
 sg13g2_decap_8 FILLER_10_1064 ();
 sg13g2_decap_8 FILLER_10_1071 ();
 sg13g2_decap_8 FILLER_10_1078 ();
 sg13g2_decap_8 FILLER_10_1085 ();
 sg13g2_decap_8 FILLER_10_1092 ();
 sg13g2_decap_8 FILLER_10_1099 ();
 sg13g2_decap_8 FILLER_10_1106 ();
 sg13g2_decap_8 FILLER_10_1113 ();
 sg13g2_decap_8 FILLER_10_1120 ();
 sg13g2_decap_8 FILLER_10_1127 ();
 sg13g2_decap_8 FILLER_10_1134 ();
 sg13g2_decap_8 FILLER_10_1141 ();
 sg13g2_decap_8 FILLER_10_1148 ();
 sg13g2_decap_8 FILLER_10_1155 ();
 sg13g2_decap_8 FILLER_10_1162 ();
 sg13g2_decap_8 FILLER_10_1169 ();
 sg13g2_decap_8 FILLER_10_1176 ();
 sg13g2_decap_8 FILLER_10_1183 ();
 sg13g2_decap_8 FILLER_10_1190 ();
 sg13g2_decap_8 FILLER_10_1197 ();
 sg13g2_decap_8 FILLER_10_1204 ();
 sg13g2_decap_8 FILLER_10_1211 ();
 sg13g2_decap_8 FILLER_10_1218 ();
 sg13g2_decap_8 FILLER_10_1225 ();
 sg13g2_decap_8 FILLER_10_1232 ();
 sg13g2_decap_8 FILLER_10_1239 ();
 sg13g2_decap_8 FILLER_10_1246 ();
 sg13g2_decap_8 FILLER_10_1253 ();
 sg13g2_decap_8 FILLER_10_1260 ();
 sg13g2_decap_8 FILLER_10_1267 ();
 sg13g2_decap_8 FILLER_10_1274 ();
 sg13g2_decap_8 FILLER_10_1281 ();
 sg13g2_decap_8 FILLER_10_1288 ();
 sg13g2_decap_8 FILLER_10_1295 ();
 sg13g2_decap_8 FILLER_10_1302 ();
 sg13g2_decap_8 FILLER_10_1309 ();
 sg13g2_decap_8 FILLER_10_1316 ();
 sg13g2_decap_8 FILLER_10_1323 ();
 sg13g2_decap_8 FILLER_10_1330 ();
 sg13g2_decap_8 FILLER_10_1337 ();
 sg13g2_decap_8 FILLER_10_1344 ();
 sg13g2_decap_8 FILLER_10_1351 ();
 sg13g2_decap_8 FILLER_10_1358 ();
 sg13g2_decap_8 FILLER_10_1365 ();
 sg13g2_decap_8 FILLER_10_1372 ();
 sg13g2_decap_8 FILLER_10_1379 ();
 sg13g2_decap_8 FILLER_10_1386 ();
 sg13g2_decap_8 FILLER_10_1393 ();
 sg13g2_decap_8 FILLER_10_1400 ();
 sg13g2_decap_8 FILLER_10_1407 ();
 sg13g2_decap_8 FILLER_10_1414 ();
 sg13g2_decap_8 FILLER_10_1421 ();
 sg13g2_decap_8 FILLER_10_1428 ();
 sg13g2_decap_8 FILLER_10_1435 ();
 sg13g2_decap_8 FILLER_10_1442 ();
 sg13g2_decap_8 FILLER_10_1449 ();
 sg13g2_decap_8 FILLER_10_1456 ();
 sg13g2_decap_8 FILLER_10_1463 ();
 sg13g2_decap_8 FILLER_10_1470 ();
 sg13g2_decap_8 FILLER_10_1477 ();
 sg13g2_decap_8 FILLER_10_1484 ();
 sg13g2_decap_8 FILLER_10_1491 ();
 sg13g2_decap_8 FILLER_10_1498 ();
 sg13g2_decap_8 FILLER_10_1505 ();
 sg13g2_decap_8 FILLER_10_1512 ();
 sg13g2_decap_8 FILLER_10_1519 ();
 sg13g2_decap_8 FILLER_10_1526 ();
 sg13g2_decap_8 FILLER_10_1533 ();
 sg13g2_decap_8 FILLER_10_1540 ();
 sg13g2_decap_8 FILLER_10_1547 ();
 sg13g2_decap_8 FILLER_10_1554 ();
 sg13g2_decap_8 FILLER_10_1561 ();
 sg13g2_decap_8 FILLER_10_1568 ();
 sg13g2_decap_8 FILLER_10_1575 ();
 sg13g2_decap_8 FILLER_10_1582 ();
 sg13g2_decap_8 FILLER_10_1589 ();
 sg13g2_decap_8 FILLER_10_1596 ();
 sg13g2_decap_8 FILLER_10_1603 ();
 sg13g2_decap_8 FILLER_10_1610 ();
 sg13g2_decap_8 FILLER_10_1617 ();
 sg13g2_decap_8 FILLER_10_1624 ();
 sg13g2_decap_8 FILLER_10_1631 ();
 sg13g2_decap_8 FILLER_10_1638 ();
 sg13g2_decap_8 FILLER_10_1645 ();
 sg13g2_decap_8 FILLER_10_1652 ();
 sg13g2_decap_8 FILLER_10_1659 ();
 sg13g2_decap_8 FILLER_10_1666 ();
 sg13g2_decap_8 FILLER_10_1673 ();
 sg13g2_decap_8 FILLER_10_1680 ();
 sg13g2_decap_8 FILLER_10_1687 ();
 sg13g2_decap_8 FILLER_10_1694 ();
 sg13g2_decap_8 FILLER_10_1701 ();
 sg13g2_decap_8 FILLER_10_1708 ();
 sg13g2_decap_8 FILLER_10_1715 ();
 sg13g2_decap_8 FILLER_10_1722 ();
 sg13g2_decap_8 FILLER_10_1729 ();
 sg13g2_decap_8 FILLER_10_1736 ();
 sg13g2_decap_8 FILLER_10_1743 ();
 sg13g2_decap_8 FILLER_10_1750 ();
 sg13g2_decap_8 FILLER_10_1757 ();
 sg13g2_decap_4 FILLER_10_1764 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_fill_2 FILLER_11_49 ();
 sg13g2_fill_1 FILLER_11_51 ();
 sg13g2_decap_4 FILLER_11_62 ();
 sg13g2_fill_1 FILLER_11_92 ();
 sg13g2_fill_1 FILLER_11_136 ();
 sg13g2_fill_2 FILLER_11_190 ();
 sg13g2_fill_1 FILLER_11_192 ();
 sg13g2_fill_1 FILLER_11_229 ();
 sg13g2_fill_2 FILLER_11_351 ();
 sg13g2_fill_2 FILLER_11_367 ();
 sg13g2_fill_2 FILLER_11_383 ();
 sg13g2_fill_1 FILLER_11_385 ();
 sg13g2_decap_4 FILLER_11_436 ();
 sg13g2_fill_2 FILLER_11_440 ();
 sg13g2_decap_8 FILLER_11_447 ();
 sg13g2_fill_2 FILLER_11_454 ();
 sg13g2_fill_2 FILLER_11_461 ();
 sg13g2_fill_1 FILLER_11_463 ();
 sg13g2_fill_1 FILLER_11_473 ();
 sg13g2_decap_8 FILLER_11_486 ();
 sg13g2_fill_2 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_512 ();
 sg13g2_decap_4 FILLER_11_540 ();
 sg13g2_fill_2 FILLER_11_544 ();
 sg13g2_fill_2 FILLER_11_563 ();
 sg13g2_fill_1 FILLER_11_565 ();
 sg13g2_decap_4 FILLER_11_570 ();
 sg13g2_fill_1 FILLER_11_574 ();
 sg13g2_fill_1 FILLER_11_585 ();
 sg13g2_fill_2 FILLER_11_596 ();
 sg13g2_fill_1 FILLER_11_598 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_fill_2 FILLER_11_630 ();
 sg13g2_fill_2 FILLER_11_640 ();
 sg13g2_decap_8 FILLER_11_650 ();
 sg13g2_fill_1 FILLER_11_657 ();
 sg13g2_fill_2 FILLER_11_678 ();
 sg13g2_fill_1 FILLER_11_680 ();
 sg13g2_decap_4 FILLER_11_691 ();
 sg13g2_decap_4 FILLER_11_700 ();
 sg13g2_fill_2 FILLER_11_708 ();
 sg13g2_decap_8 FILLER_11_733 ();
 sg13g2_fill_1 FILLER_11_740 ();
 sg13g2_decap_8 FILLER_11_769 ();
 sg13g2_fill_2 FILLER_11_776 ();
 sg13g2_fill_1 FILLER_11_778 ();
 sg13g2_decap_8 FILLER_11_789 ();
 sg13g2_decap_8 FILLER_11_796 ();
 sg13g2_decap_8 FILLER_11_803 ();
 sg13g2_decap_8 FILLER_11_810 ();
 sg13g2_decap_8 FILLER_11_817 ();
 sg13g2_decap_8 FILLER_11_824 ();
 sg13g2_decap_8 FILLER_11_831 ();
 sg13g2_decap_8 FILLER_11_838 ();
 sg13g2_decap_8 FILLER_11_845 ();
 sg13g2_decap_8 FILLER_11_852 ();
 sg13g2_decap_8 FILLER_11_859 ();
 sg13g2_decap_8 FILLER_11_866 ();
 sg13g2_decap_8 FILLER_11_873 ();
 sg13g2_decap_8 FILLER_11_880 ();
 sg13g2_decap_8 FILLER_11_887 ();
 sg13g2_decap_8 FILLER_11_894 ();
 sg13g2_decap_8 FILLER_11_901 ();
 sg13g2_decap_8 FILLER_11_908 ();
 sg13g2_decap_8 FILLER_11_915 ();
 sg13g2_decap_8 FILLER_11_922 ();
 sg13g2_decap_8 FILLER_11_929 ();
 sg13g2_decap_8 FILLER_11_936 ();
 sg13g2_decap_8 FILLER_11_943 ();
 sg13g2_decap_8 FILLER_11_950 ();
 sg13g2_decap_8 FILLER_11_957 ();
 sg13g2_decap_8 FILLER_11_964 ();
 sg13g2_decap_8 FILLER_11_971 ();
 sg13g2_decap_8 FILLER_11_978 ();
 sg13g2_decap_8 FILLER_11_985 ();
 sg13g2_decap_8 FILLER_11_992 ();
 sg13g2_decap_8 FILLER_11_999 ();
 sg13g2_decap_8 FILLER_11_1006 ();
 sg13g2_decap_8 FILLER_11_1013 ();
 sg13g2_decap_8 FILLER_11_1020 ();
 sg13g2_decap_8 FILLER_11_1027 ();
 sg13g2_decap_8 FILLER_11_1034 ();
 sg13g2_decap_8 FILLER_11_1041 ();
 sg13g2_decap_8 FILLER_11_1048 ();
 sg13g2_decap_8 FILLER_11_1055 ();
 sg13g2_decap_8 FILLER_11_1062 ();
 sg13g2_decap_8 FILLER_11_1069 ();
 sg13g2_decap_8 FILLER_11_1076 ();
 sg13g2_decap_8 FILLER_11_1083 ();
 sg13g2_decap_8 FILLER_11_1090 ();
 sg13g2_decap_8 FILLER_11_1097 ();
 sg13g2_decap_8 FILLER_11_1104 ();
 sg13g2_decap_8 FILLER_11_1111 ();
 sg13g2_decap_8 FILLER_11_1118 ();
 sg13g2_decap_8 FILLER_11_1125 ();
 sg13g2_decap_8 FILLER_11_1132 ();
 sg13g2_decap_8 FILLER_11_1139 ();
 sg13g2_decap_8 FILLER_11_1146 ();
 sg13g2_decap_8 FILLER_11_1153 ();
 sg13g2_decap_8 FILLER_11_1160 ();
 sg13g2_decap_8 FILLER_11_1167 ();
 sg13g2_decap_8 FILLER_11_1174 ();
 sg13g2_decap_8 FILLER_11_1181 ();
 sg13g2_decap_8 FILLER_11_1188 ();
 sg13g2_decap_8 FILLER_11_1195 ();
 sg13g2_decap_8 FILLER_11_1202 ();
 sg13g2_decap_8 FILLER_11_1209 ();
 sg13g2_decap_8 FILLER_11_1216 ();
 sg13g2_decap_8 FILLER_11_1223 ();
 sg13g2_decap_8 FILLER_11_1230 ();
 sg13g2_decap_8 FILLER_11_1237 ();
 sg13g2_decap_8 FILLER_11_1244 ();
 sg13g2_decap_8 FILLER_11_1251 ();
 sg13g2_decap_8 FILLER_11_1258 ();
 sg13g2_decap_8 FILLER_11_1265 ();
 sg13g2_decap_8 FILLER_11_1272 ();
 sg13g2_decap_8 FILLER_11_1279 ();
 sg13g2_decap_8 FILLER_11_1286 ();
 sg13g2_decap_8 FILLER_11_1293 ();
 sg13g2_decap_8 FILLER_11_1300 ();
 sg13g2_decap_8 FILLER_11_1307 ();
 sg13g2_decap_8 FILLER_11_1314 ();
 sg13g2_decap_8 FILLER_11_1321 ();
 sg13g2_decap_8 FILLER_11_1328 ();
 sg13g2_decap_8 FILLER_11_1335 ();
 sg13g2_decap_8 FILLER_11_1342 ();
 sg13g2_decap_8 FILLER_11_1349 ();
 sg13g2_decap_8 FILLER_11_1356 ();
 sg13g2_decap_8 FILLER_11_1363 ();
 sg13g2_decap_8 FILLER_11_1370 ();
 sg13g2_decap_8 FILLER_11_1377 ();
 sg13g2_decap_8 FILLER_11_1384 ();
 sg13g2_decap_8 FILLER_11_1391 ();
 sg13g2_decap_8 FILLER_11_1398 ();
 sg13g2_decap_8 FILLER_11_1405 ();
 sg13g2_decap_8 FILLER_11_1412 ();
 sg13g2_decap_8 FILLER_11_1419 ();
 sg13g2_decap_8 FILLER_11_1426 ();
 sg13g2_decap_8 FILLER_11_1433 ();
 sg13g2_decap_8 FILLER_11_1440 ();
 sg13g2_decap_8 FILLER_11_1447 ();
 sg13g2_decap_8 FILLER_11_1454 ();
 sg13g2_decap_8 FILLER_11_1461 ();
 sg13g2_decap_8 FILLER_11_1468 ();
 sg13g2_decap_8 FILLER_11_1475 ();
 sg13g2_decap_8 FILLER_11_1482 ();
 sg13g2_decap_8 FILLER_11_1489 ();
 sg13g2_decap_8 FILLER_11_1496 ();
 sg13g2_decap_8 FILLER_11_1503 ();
 sg13g2_decap_8 FILLER_11_1510 ();
 sg13g2_decap_8 FILLER_11_1517 ();
 sg13g2_decap_8 FILLER_11_1524 ();
 sg13g2_decap_8 FILLER_11_1531 ();
 sg13g2_decap_8 FILLER_11_1538 ();
 sg13g2_decap_8 FILLER_11_1545 ();
 sg13g2_decap_8 FILLER_11_1552 ();
 sg13g2_decap_8 FILLER_11_1559 ();
 sg13g2_decap_8 FILLER_11_1566 ();
 sg13g2_decap_8 FILLER_11_1573 ();
 sg13g2_decap_8 FILLER_11_1580 ();
 sg13g2_decap_8 FILLER_11_1587 ();
 sg13g2_decap_8 FILLER_11_1594 ();
 sg13g2_decap_8 FILLER_11_1601 ();
 sg13g2_decap_8 FILLER_11_1608 ();
 sg13g2_decap_8 FILLER_11_1615 ();
 sg13g2_decap_8 FILLER_11_1622 ();
 sg13g2_decap_8 FILLER_11_1629 ();
 sg13g2_decap_8 FILLER_11_1636 ();
 sg13g2_decap_8 FILLER_11_1643 ();
 sg13g2_decap_8 FILLER_11_1650 ();
 sg13g2_decap_8 FILLER_11_1657 ();
 sg13g2_decap_8 FILLER_11_1664 ();
 sg13g2_decap_8 FILLER_11_1671 ();
 sg13g2_decap_8 FILLER_11_1678 ();
 sg13g2_decap_8 FILLER_11_1685 ();
 sg13g2_decap_8 FILLER_11_1692 ();
 sg13g2_decap_8 FILLER_11_1699 ();
 sg13g2_decap_8 FILLER_11_1706 ();
 sg13g2_decap_8 FILLER_11_1713 ();
 sg13g2_decap_8 FILLER_11_1720 ();
 sg13g2_decap_8 FILLER_11_1727 ();
 sg13g2_decap_8 FILLER_11_1734 ();
 sg13g2_decap_8 FILLER_11_1741 ();
 sg13g2_decap_8 FILLER_11_1748 ();
 sg13g2_decap_8 FILLER_11_1755 ();
 sg13g2_decap_4 FILLER_11_1762 ();
 sg13g2_fill_2 FILLER_11_1766 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_4 FILLER_12_42 ();
 sg13g2_fill_2 FILLER_12_46 ();
 sg13g2_decap_8 FILLER_12_74 ();
 sg13g2_fill_1 FILLER_12_81 ();
 sg13g2_fill_1 FILLER_12_159 ();
 sg13g2_fill_2 FILLER_12_195 ();
 sg13g2_decap_4 FILLER_12_231 ();
 sg13g2_fill_1 FILLER_12_294 ();
 sg13g2_fill_1 FILLER_12_321 ();
 sg13g2_fill_1 FILLER_12_353 ();
 sg13g2_fill_2 FILLER_12_433 ();
 sg13g2_fill_1 FILLER_12_451 ();
 sg13g2_fill_2 FILLER_12_459 ();
 sg13g2_fill_1 FILLER_12_461 ();
 sg13g2_fill_1 FILLER_12_476 ();
 sg13g2_fill_2 FILLER_12_488 ();
 sg13g2_fill_1 FILLER_12_490 ();
 sg13g2_fill_2 FILLER_12_522 ();
 sg13g2_fill_1 FILLER_12_524 ();
 sg13g2_fill_2 FILLER_12_532 ();
 sg13g2_fill_1 FILLER_12_534 ();
 sg13g2_fill_2 FILLER_12_556 ();
 sg13g2_fill_1 FILLER_12_566 ();
 sg13g2_fill_2 FILLER_12_575 ();
 sg13g2_fill_2 FILLER_12_636 ();
 sg13g2_fill_1 FILLER_12_653 ();
 sg13g2_decap_4 FILLER_12_675 ();
 sg13g2_fill_1 FILLER_12_679 ();
 sg13g2_fill_1 FILLER_12_688 ();
 sg13g2_fill_2 FILLER_12_694 ();
 sg13g2_fill_1 FILLER_12_696 ();
 sg13g2_fill_1 FILLER_12_734 ();
 sg13g2_fill_1 FILLER_12_747 ();
 sg13g2_decap_8 FILLER_12_758 ();
 sg13g2_decap_4 FILLER_12_765 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_794 ();
 sg13g2_decap_8 FILLER_12_801 ();
 sg13g2_decap_8 FILLER_12_808 ();
 sg13g2_decap_8 FILLER_12_815 ();
 sg13g2_decap_8 FILLER_12_822 ();
 sg13g2_decap_8 FILLER_12_829 ();
 sg13g2_decap_8 FILLER_12_836 ();
 sg13g2_decap_8 FILLER_12_843 ();
 sg13g2_decap_8 FILLER_12_850 ();
 sg13g2_decap_8 FILLER_12_857 ();
 sg13g2_decap_8 FILLER_12_864 ();
 sg13g2_decap_8 FILLER_12_871 ();
 sg13g2_decap_8 FILLER_12_878 ();
 sg13g2_decap_8 FILLER_12_885 ();
 sg13g2_decap_8 FILLER_12_892 ();
 sg13g2_decap_8 FILLER_12_899 ();
 sg13g2_decap_8 FILLER_12_906 ();
 sg13g2_decap_8 FILLER_12_913 ();
 sg13g2_decap_8 FILLER_12_920 ();
 sg13g2_decap_8 FILLER_12_927 ();
 sg13g2_decap_8 FILLER_12_934 ();
 sg13g2_decap_8 FILLER_12_941 ();
 sg13g2_decap_8 FILLER_12_948 ();
 sg13g2_decap_8 FILLER_12_955 ();
 sg13g2_decap_8 FILLER_12_962 ();
 sg13g2_decap_8 FILLER_12_969 ();
 sg13g2_decap_8 FILLER_12_976 ();
 sg13g2_decap_8 FILLER_12_983 ();
 sg13g2_decap_8 FILLER_12_990 ();
 sg13g2_decap_8 FILLER_12_997 ();
 sg13g2_decap_8 FILLER_12_1004 ();
 sg13g2_decap_8 FILLER_12_1011 ();
 sg13g2_decap_8 FILLER_12_1018 ();
 sg13g2_decap_8 FILLER_12_1025 ();
 sg13g2_decap_8 FILLER_12_1032 ();
 sg13g2_decap_8 FILLER_12_1039 ();
 sg13g2_decap_8 FILLER_12_1046 ();
 sg13g2_decap_8 FILLER_12_1053 ();
 sg13g2_decap_8 FILLER_12_1060 ();
 sg13g2_decap_8 FILLER_12_1067 ();
 sg13g2_decap_8 FILLER_12_1074 ();
 sg13g2_decap_8 FILLER_12_1081 ();
 sg13g2_decap_8 FILLER_12_1088 ();
 sg13g2_decap_8 FILLER_12_1095 ();
 sg13g2_decap_8 FILLER_12_1102 ();
 sg13g2_decap_8 FILLER_12_1109 ();
 sg13g2_decap_8 FILLER_12_1116 ();
 sg13g2_decap_8 FILLER_12_1123 ();
 sg13g2_decap_8 FILLER_12_1130 ();
 sg13g2_decap_8 FILLER_12_1137 ();
 sg13g2_decap_8 FILLER_12_1144 ();
 sg13g2_decap_8 FILLER_12_1151 ();
 sg13g2_decap_8 FILLER_12_1158 ();
 sg13g2_decap_8 FILLER_12_1165 ();
 sg13g2_decap_8 FILLER_12_1172 ();
 sg13g2_decap_8 FILLER_12_1179 ();
 sg13g2_decap_8 FILLER_12_1186 ();
 sg13g2_decap_8 FILLER_12_1193 ();
 sg13g2_decap_8 FILLER_12_1200 ();
 sg13g2_decap_8 FILLER_12_1207 ();
 sg13g2_decap_8 FILLER_12_1214 ();
 sg13g2_decap_8 FILLER_12_1221 ();
 sg13g2_decap_8 FILLER_12_1228 ();
 sg13g2_decap_8 FILLER_12_1235 ();
 sg13g2_decap_8 FILLER_12_1242 ();
 sg13g2_decap_8 FILLER_12_1249 ();
 sg13g2_decap_8 FILLER_12_1256 ();
 sg13g2_decap_8 FILLER_12_1263 ();
 sg13g2_decap_8 FILLER_12_1270 ();
 sg13g2_decap_8 FILLER_12_1277 ();
 sg13g2_decap_8 FILLER_12_1284 ();
 sg13g2_decap_8 FILLER_12_1291 ();
 sg13g2_decap_8 FILLER_12_1298 ();
 sg13g2_decap_8 FILLER_12_1305 ();
 sg13g2_decap_8 FILLER_12_1312 ();
 sg13g2_decap_8 FILLER_12_1319 ();
 sg13g2_decap_8 FILLER_12_1326 ();
 sg13g2_decap_8 FILLER_12_1333 ();
 sg13g2_decap_8 FILLER_12_1340 ();
 sg13g2_decap_8 FILLER_12_1347 ();
 sg13g2_decap_8 FILLER_12_1354 ();
 sg13g2_decap_8 FILLER_12_1361 ();
 sg13g2_decap_8 FILLER_12_1368 ();
 sg13g2_decap_8 FILLER_12_1375 ();
 sg13g2_decap_8 FILLER_12_1382 ();
 sg13g2_decap_8 FILLER_12_1389 ();
 sg13g2_decap_8 FILLER_12_1396 ();
 sg13g2_decap_8 FILLER_12_1403 ();
 sg13g2_decap_8 FILLER_12_1410 ();
 sg13g2_decap_8 FILLER_12_1417 ();
 sg13g2_decap_8 FILLER_12_1424 ();
 sg13g2_decap_8 FILLER_12_1431 ();
 sg13g2_decap_8 FILLER_12_1438 ();
 sg13g2_decap_8 FILLER_12_1445 ();
 sg13g2_decap_8 FILLER_12_1452 ();
 sg13g2_decap_8 FILLER_12_1459 ();
 sg13g2_decap_8 FILLER_12_1466 ();
 sg13g2_decap_8 FILLER_12_1473 ();
 sg13g2_decap_8 FILLER_12_1480 ();
 sg13g2_decap_8 FILLER_12_1487 ();
 sg13g2_decap_8 FILLER_12_1494 ();
 sg13g2_decap_8 FILLER_12_1501 ();
 sg13g2_decap_8 FILLER_12_1508 ();
 sg13g2_decap_8 FILLER_12_1515 ();
 sg13g2_decap_8 FILLER_12_1522 ();
 sg13g2_decap_8 FILLER_12_1529 ();
 sg13g2_decap_8 FILLER_12_1536 ();
 sg13g2_decap_8 FILLER_12_1543 ();
 sg13g2_decap_8 FILLER_12_1550 ();
 sg13g2_decap_8 FILLER_12_1557 ();
 sg13g2_decap_8 FILLER_12_1564 ();
 sg13g2_decap_8 FILLER_12_1571 ();
 sg13g2_decap_8 FILLER_12_1578 ();
 sg13g2_decap_8 FILLER_12_1585 ();
 sg13g2_decap_8 FILLER_12_1592 ();
 sg13g2_decap_8 FILLER_12_1599 ();
 sg13g2_decap_8 FILLER_12_1606 ();
 sg13g2_decap_8 FILLER_12_1613 ();
 sg13g2_decap_8 FILLER_12_1620 ();
 sg13g2_decap_8 FILLER_12_1627 ();
 sg13g2_decap_8 FILLER_12_1634 ();
 sg13g2_decap_8 FILLER_12_1641 ();
 sg13g2_decap_8 FILLER_12_1648 ();
 sg13g2_decap_8 FILLER_12_1655 ();
 sg13g2_decap_8 FILLER_12_1662 ();
 sg13g2_decap_8 FILLER_12_1669 ();
 sg13g2_decap_8 FILLER_12_1676 ();
 sg13g2_decap_8 FILLER_12_1683 ();
 sg13g2_decap_8 FILLER_12_1690 ();
 sg13g2_decap_8 FILLER_12_1697 ();
 sg13g2_decap_8 FILLER_12_1704 ();
 sg13g2_decap_8 FILLER_12_1711 ();
 sg13g2_decap_8 FILLER_12_1718 ();
 sg13g2_decap_8 FILLER_12_1725 ();
 sg13g2_decap_8 FILLER_12_1732 ();
 sg13g2_decap_8 FILLER_12_1739 ();
 sg13g2_decap_8 FILLER_12_1746 ();
 sg13g2_decap_8 FILLER_12_1753 ();
 sg13g2_decap_8 FILLER_12_1760 ();
 sg13g2_fill_1 FILLER_12_1767 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_fill_2 FILLER_13_49 ();
 sg13g2_fill_1 FILLER_13_51 ();
 sg13g2_fill_2 FILLER_13_92 ();
 sg13g2_decap_4 FILLER_13_116 ();
 sg13g2_fill_2 FILLER_13_120 ();
 sg13g2_fill_2 FILLER_13_154 ();
 sg13g2_fill_2 FILLER_13_166 ();
 sg13g2_decap_8 FILLER_13_194 ();
 sg13g2_fill_1 FILLER_13_201 ();
 sg13g2_fill_2 FILLER_13_251 ();
 sg13g2_fill_1 FILLER_13_253 ();
 sg13g2_fill_2 FILLER_13_280 ();
 sg13g2_fill_1 FILLER_13_282 ();
 sg13g2_fill_2 FILLER_13_297 ();
 sg13g2_fill_2 FILLER_13_318 ();
 sg13g2_fill_1 FILLER_13_320 ();
 sg13g2_fill_1 FILLER_13_329 ();
 sg13g2_fill_2 FILLER_13_379 ();
 sg13g2_fill_2 FILLER_13_404 ();
 sg13g2_decap_4 FILLER_13_443 ();
 sg13g2_fill_2 FILLER_13_447 ();
 sg13g2_decap_8 FILLER_13_457 ();
 sg13g2_decap_4 FILLER_13_473 ();
 sg13g2_fill_2 FILLER_13_489 ();
 sg13g2_fill_1 FILLER_13_519 ();
 sg13g2_fill_2 FILLER_13_523 ();
 sg13g2_fill_1 FILLER_13_525 ();
 sg13g2_decap_4 FILLER_13_534 ();
 sg13g2_fill_2 FILLER_13_547 ();
 sg13g2_fill_1 FILLER_13_549 ();
 sg13g2_fill_1 FILLER_13_558 ();
 sg13g2_fill_2 FILLER_13_563 ();
 sg13g2_fill_1 FILLER_13_569 ();
 sg13g2_decap_8 FILLER_13_621 ();
 sg13g2_fill_1 FILLER_13_628 ();
 sg13g2_decap_4 FILLER_13_652 ();
 sg13g2_fill_2 FILLER_13_665 ();
 sg13g2_fill_1 FILLER_13_667 ();
 sg13g2_fill_2 FILLER_13_673 ();
 sg13g2_fill_1 FILLER_13_696 ();
 sg13g2_decap_8 FILLER_13_702 ();
 sg13g2_fill_2 FILLER_13_709 ();
 sg13g2_decap_8 FILLER_13_723 ();
 sg13g2_decap_4 FILLER_13_746 ();
 sg13g2_fill_2 FILLER_13_783 ();
 sg13g2_fill_1 FILLER_13_785 ();
 sg13g2_decap_8 FILLER_13_799 ();
 sg13g2_decap_8 FILLER_13_806 ();
 sg13g2_decap_8 FILLER_13_813 ();
 sg13g2_decap_8 FILLER_13_820 ();
 sg13g2_decap_8 FILLER_13_827 ();
 sg13g2_decap_8 FILLER_13_834 ();
 sg13g2_decap_8 FILLER_13_841 ();
 sg13g2_decap_8 FILLER_13_848 ();
 sg13g2_decap_8 FILLER_13_855 ();
 sg13g2_decap_8 FILLER_13_862 ();
 sg13g2_decap_8 FILLER_13_869 ();
 sg13g2_decap_8 FILLER_13_876 ();
 sg13g2_decap_8 FILLER_13_883 ();
 sg13g2_decap_8 FILLER_13_890 ();
 sg13g2_decap_8 FILLER_13_897 ();
 sg13g2_decap_8 FILLER_13_904 ();
 sg13g2_decap_8 FILLER_13_911 ();
 sg13g2_decap_8 FILLER_13_918 ();
 sg13g2_decap_8 FILLER_13_925 ();
 sg13g2_decap_8 FILLER_13_932 ();
 sg13g2_decap_8 FILLER_13_939 ();
 sg13g2_decap_8 FILLER_13_946 ();
 sg13g2_decap_8 FILLER_13_953 ();
 sg13g2_decap_8 FILLER_13_960 ();
 sg13g2_decap_8 FILLER_13_967 ();
 sg13g2_decap_8 FILLER_13_974 ();
 sg13g2_decap_8 FILLER_13_981 ();
 sg13g2_decap_8 FILLER_13_988 ();
 sg13g2_decap_8 FILLER_13_995 ();
 sg13g2_decap_8 FILLER_13_1002 ();
 sg13g2_decap_8 FILLER_13_1009 ();
 sg13g2_decap_8 FILLER_13_1016 ();
 sg13g2_decap_8 FILLER_13_1023 ();
 sg13g2_decap_8 FILLER_13_1030 ();
 sg13g2_decap_8 FILLER_13_1037 ();
 sg13g2_decap_8 FILLER_13_1044 ();
 sg13g2_decap_8 FILLER_13_1051 ();
 sg13g2_decap_8 FILLER_13_1058 ();
 sg13g2_decap_8 FILLER_13_1065 ();
 sg13g2_decap_8 FILLER_13_1072 ();
 sg13g2_decap_8 FILLER_13_1079 ();
 sg13g2_decap_8 FILLER_13_1086 ();
 sg13g2_decap_8 FILLER_13_1093 ();
 sg13g2_decap_8 FILLER_13_1100 ();
 sg13g2_decap_8 FILLER_13_1107 ();
 sg13g2_decap_8 FILLER_13_1114 ();
 sg13g2_decap_8 FILLER_13_1121 ();
 sg13g2_decap_8 FILLER_13_1128 ();
 sg13g2_decap_8 FILLER_13_1135 ();
 sg13g2_decap_8 FILLER_13_1142 ();
 sg13g2_decap_8 FILLER_13_1149 ();
 sg13g2_decap_8 FILLER_13_1156 ();
 sg13g2_decap_8 FILLER_13_1163 ();
 sg13g2_decap_8 FILLER_13_1170 ();
 sg13g2_decap_8 FILLER_13_1177 ();
 sg13g2_decap_8 FILLER_13_1184 ();
 sg13g2_decap_8 FILLER_13_1191 ();
 sg13g2_decap_8 FILLER_13_1198 ();
 sg13g2_decap_8 FILLER_13_1205 ();
 sg13g2_decap_8 FILLER_13_1212 ();
 sg13g2_decap_8 FILLER_13_1219 ();
 sg13g2_decap_8 FILLER_13_1226 ();
 sg13g2_decap_8 FILLER_13_1233 ();
 sg13g2_decap_8 FILLER_13_1240 ();
 sg13g2_decap_8 FILLER_13_1247 ();
 sg13g2_decap_8 FILLER_13_1254 ();
 sg13g2_decap_8 FILLER_13_1261 ();
 sg13g2_decap_8 FILLER_13_1268 ();
 sg13g2_decap_8 FILLER_13_1275 ();
 sg13g2_decap_8 FILLER_13_1282 ();
 sg13g2_decap_8 FILLER_13_1289 ();
 sg13g2_decap_8 FILLER_13_1296 ();
 sg13g2_decap_8 FILLER_13_1303 ();
 sg13g2_decap_8 FILLER_13_1310 ();
 sg13g2_decap_8 FILLER_13_1317 ();
 sg13g2_decap_8 FILLER_13_1324 ();
 sg13g2_decap_8 FILLER_13_1331 ();
 sg13g2_decap_8 FILLER_13_1338 ();
 sg13g2_decap_8 FILLER_13_1345 ();
 sg13g2_decap_8 FILLER_13_1352 ();
 sg13g2_decap_8 FILLER_13_1359 ();
 sg13g2_decap_8 FILLER_13_1366 ();
 sg13g2_decap_8 FILLER_13_1373 ();
 sg13g2_decap_8 FILLER_13_1380 ();
 sg13g2_decap_8 FILLER_13_1387 ();
 sg13g2_decap_8 FILLER_13_1394 ();
 sg13g2_decap_8 FILLER_13_1401 ();
 sg13g2_decap_8 FILLER_13_1408 ();
 sg13g2_decap_8 FILLER_13_1415 ();
 sg13g2_decap_8 FILLER_13_1422 ();
 sg13g2_decap_8 FILLER_13_1429 ();
 sg13g2_decap_8 FILLER_13_1436 ();
 sg13g2_decap_8 FILLER_13_1443 ();
 sg13g2_decap_8 FILLER_13_1450 ();
 sg13g2_decap_8 FILLER_13_1457 ();
 sg13g2_decap_8 FILLER_13_1464 ();
 sg13g2_decap_8 FILLER_13_1471 ();
 sg13g2_decap_8 FILLER_13_1478 ();
 sg13g2_decap_8 FILLER_13_1485 ();
 sg13g2_decap_8 FILLER_13_1492 ();
 sg13g2_decap_8 FILLER_13_1499 ();
 sg13g2_decap_8 FILLER_13_1506 ();
 sg13g2_decap_8 FILLER_13_1513 ();
 sg13g2_decap_8 FILLER_13_1520 ();
 sg13g2_decap_8 FILLER_13_1527 ();
 sg13g2_decap_8 FILLER_13_1534 ();
 sg13g2_decap_8 FILLER_13_1541 ();
 sg13g2_decap_8 FILLER_13_1548 ();
 sg13g2_decap_8 FILLER_13_1555 ();
 sg13g2_decap_8 FILLER_13_1562 ();
 sg13g2_decap_8 FILLER_13_1569 ();
 sg13g2_decap_8 FILLER_13_1576 ();
 sg13g2_decap_8 FILLER_13_1583 ();
 sg13g2_decap_8 FILLER_13_1590 ();
 sg13g2_decap_8 FILLER_13_1597 ();
 sg13g2_decap_8 FILLER_13_1604 ();
 sg13g2_decap_8 FILLER_13_1611 ();
 sg13g2_decap_8 FILLER_13_1618 ();
 sg13g2_decap_8 FILLER_13_1625 ();
 sg13g2_decap_8 FILLER_13_1632 ();
 sg13g2_decap_8 FILLER_13_1639 ();
 sg13g2_decap_8 FILLER_13_1646 ();
 sg13g2_decap_8 FILLER_13_1653 ();
 sg13g2_decap_8 FILLER_13_1660 ();
 sg13g2_decap_8 FILLER_13_1667 ();
 sg13g2_decap_8 FILLER_13_1674 ();
 sg13g2_decap_8 FILLER_13_1681 ();
 sg13g2_decap_8 FILLER_13_1688 ();
 sg13g2_decap_8 FILLER_13_1695 ();
 sg13g2_decap_8 FILLER_13_1702 ();
 sg13g2_decap_8 FILLER_13_1709 ();
 sg13g2_decap_8 FILLER_13_1716 ();
 sg13g2_decap_8 FILLER_13_1723 ();
 sg13g2_decap_8 FILLER_13_1730 ();
 sg13g2_decap_8 FILLER_13_1737 ();
 sg13g2_decap_8 FILLER_13_1744 ();
 sg13g2_decap_8 FILLER_13_1751 ();
 sg13g2_decap_8 FILLER_13_1758 ();
 sg13g2_fill_2 FILLER_13_1765 ();
 sg13g2_fill_1 FILLER_13_1767 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_4 FILLER_14_21 ();
 sg13g2_fill_2 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_113 ();
 sg13g2_fill_2 FILLER_14_120 ();
 sg13g2_decap_4 FILLER_14_158 ();
 sg13g2_fill_2 FILLER_14_162 ();
 sg13g2_fill_2 FILLER_14_190 ();
 sg13g2_fill_1 FILLER_14_212 ();
 sg13g2_fill_1 FILLER_14_229 ();
 sg13g2_decap_4 FILLER_14_239 ();
 sg13g2_fill_2 FILLER_14_253 ();
 sg13g2_fill_2 FILLER_14_296 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_2 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_4 FILLER_14_440 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_fill_1 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_481 ();
 sg13g2_decap_4 FILLER_14_488 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_fill_1 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_510 ();
 sg13g2_fill_2 FILLER_14_547 ();
 sg13g2_fill_1 FILLER_14_549 ();
 sg13g2_fill_2 FILLER_14_554 ();
 sg13g2_decap_8 FILLER_14_622 ();
 sg13g2_fill_1 FILLER_14_629 ();
 sg13g2_decap_8 FILLER_14_668 ();
 sg13g2_fill_1 FILLER_14_675 ();
 sg13g2_fill_1 FILLER_14_682 ();
 sg13g2_fill_2 FILLER_14_691 ();
 sg13g2_fill_2 FILLER_14_710 ();
 sg13g2_decap_4 FILLER_14_725 ();
 sg13g2_fill_1 FILLER_14_729 ();
 sg13g2_decap_8 FILLER_14_737 ();
 sg13g2_decap_4 FILLER_14_744 ();
 sg13g2_fill_2 FILLER_14_760 ();
 sg13g2_fill_1 FILLER_14_762 ();
 sg13g2_decap_8 FILLER_14_768 ();
 sg13g2_decap_4 FILLER_14_775 ();
 sg13g2_decap_8 FILLER_14_789 ();
 sg13g2_decap_8 FILLER_14_796 ();
 sg13g2_decap_8 FILLER_14_803 ();
 sg13g2_decap_8 FILLER_14_810 ();
 sg13g2_decap_8 FILLER_14_817 ();
 sg13g2_decap_8 FILLER_14_824 ();
 sg13g2_decap_8 FILLER_14_831 ();
 sg13g2_decap_8 FILLER_14_838 ();
 sg13g2_decap_8 FILLER_14_845 ();
 sg13g2_decap_8 FILLER_14_852 ();
 sg13g2_decap_8 FILLER_14_859 ();
 sg13g2_decap_8 FILLER_14_866 ();
 sg13g2_decap_8 FILLER_14_873 ();
 sg13g2_decap_8 FILLER_14_880 ();
 sg13g2_decap_8 FILLER_14_887 ();
 sg13g2_decap_8 FILLER_14_894 ();
 sg13g2_decap_8 FILLER_14_901 ();
 sg13g2_decap_8 FILLER_14_908 ();
 sg13g2_decap_8 FILLER_14_915 ();
 sg13g2_decap_8 FILLER_14_922 ();
 sg13g2_decap_8 FILLER_14_929 ();
 sg13g2_decap_8 FILLER_14_936 ();
 sg13g2_decap_8 FILLER_14_943 ();
 sg13g2_decap_8 FILLER_14_950 ();
 sg13g2_decap_8 FILLER_14_957 ();
 sg13g2_decap_8 FILLER_14_964 ();
 sg13g2_decap_8 FILLER_14_971 ();
 sg13g2_decap_8 FILLER_14_978 ();
 sg13g2_decap_8 FILLER_14_985 ();
 sg13g2_decap_8 FILLER_14_992 ();
 sg13g2_decap_8 FILLER_14_999 ();
 sg13g2_decap_8 FILLER_14_1006 ();
 sg13g2_decap_8 FILLER_14_1013 ();
 sg13g2_decap_8 FILLER_14_1020 ();
 sg13g2_decap_8 FILLER_14_1027 ();
 sg13g2_decap_8 FILLER_14_1034 ();
 sg13g2_decap_8 FILLER_14_1041 ();
 sg13g2_decap_8 FILLER_14_1048 ();
 sg13g2_decap_8 FILLER_14_1055 ();
 sg13g2_decap_8 FILLER_14_1062 ();
 sg13g2_decap_8 FILLER_14_1069 ();
 sg13g2_decap_8 FILLER_14_1076 ();
 sg13g2_decap_8 FILLER_14_1083 ();
 sg13g2_decap_8 FILLER_14_1090 ();
 sg13g2_decap_8 FILLER_14_1097 ();
 sg13g2_decap_8 FILLER_14_1104 ();
 sg13g2_decap_8 FILLER_14_1111 ();
 sg13g2_decap_8 FILLER_14_1118 ();
 sg13g2_decap_8 FILLER_14_1125 ();
 sg13g2_decap_8 FILLER_14_1132 ();
 sg13g2_decap_8 FILLER_14_1139 ();
 sg13g2_decap_8 FILLER_14_1146 ();
 sg13g2_decap_8 FILLER_14_1153 ();
 sg13g2_decap_8 FILLER_14_1160 ();
 sg13g2_decap_8 FILLER_14_1167 ();
 sg13g2_decap_8 FILLER_14_1174 ();
 sg13g2_decap_8 FILLER_14_1181 ();
 sg13g2_decap_8 FILLER_14_1188 ();
 sg13g2_decap_8 FILLER_14_1195 ();
 sg13g2_decap_8 FILLER_14_1202 ();
 sg13g2_decap_8 FILLER_14_1209 ();
 sg13g2_decap_8 FILLER_14_1216 ();
 sg13g2_decap_8 FILLER_14_1223 ();
 sg13g2_decap_8 FILLER_14_1230 ();
 sg13g2_decap_8 FILLER_14_1237 ();
 sg13g2_decap_8 FILLER_14_1244 ();
 sg13g2_decap_8 FILLER_14_1251 ();
 sg13g2_decap_8 FILLER_14_1258 ();
 sg13g2_decap_8 FILLER_14_1265 ();
 sg13g2_decap_8 FILLER_14_1272 ();
 sg13g2_decap_8 FILLER_14_1279 ();
 sg13g2_decap_8 FILLER_14_1286 ();
 sg13g2_decap_8 FILLER_14_1293 ();
 sg13g2_decap_8 FILLER_14_1300 ();
 sg13g2_decap_8 FILLER_14_1307 ();
 sg13g2_decap_8 FILLER_14_1314 ();
 sg13g2_decap_8 FILLER_14_1321 ();
 sg13g2_decap_8 FILLER_14_1328 ();
 sg13g2_decap_8 FILLER_14_1335 ();
 sg13g2_decap_8 FILLER_14_1342 ();
 sg13g2_decap_8 FILLER_14_1349 ();
 sg13g2_decap_8 FILLER_14_1356 ();
 sg13g2_decap_8 FILLER_14_1363 ();
 sg13g2_decap_8 FILLER_14_1370 ();
 sg13g2_decap_8 FILLER_14_1377 ();
 sg13g2_decap_8 FILLER_14_1384 ();
 sg13g2_decap_8 FILLER_14_1391 ();
 sg13g2_decap_8 FILLER_14_1398 ();
 sg13g2_decap_8 FILLER_14_1405 ();
 sg13g2_decap_8 FILLER_14_1412 ();
 sg13g2_decap_8 FILLER_14_1419 ();
 sg13g2_decap_8 FILLER_14_1426 ();
 sg13g2_decap_8 FILLER_14_1433 ();
 sg13g2_decap_8 FILLER_14_1440 ();
 sg13g2_decap_8 FILLER_14_1447 ();
 sg13g2_decap_8 FILLER_14_1454 ();
 sg13g2_decap_8 FILLER_14_1461 ();
 sg13g2_decap_8 FILLER_14_1468 ();
 sg13g2_decap_8 FILLER_14_1475 ();
 sg13g2_decap_8 FILLER_14_1482 ();
 sg13g2_decap_8 FILLER_14_1489 ();
 sg13g2_decap_8 FILLER_14_1496 ();
 sg13g2_decap_8 FILLER_14_1503 ();
 sg13g2_decap_8 FILLER_14_1510 ();
 sg13g2_decap_8 FILLER_14_1517 ();
 sg13g2_decap_8 FILLER_14_1524 ();
 sg13g2_decap_8 FILLER_14_1531 ();
 sg13g2_decap_8 FILLER_14_1538 ();
 sg13g2_decap_8 FILLER_14_1545 ();
 sg13g2_decap_8 FILLER_14_1552 ();
 sg13g2_decap_8 FILLER_14_1559 ();
 sg13g2_decap_8 FILLER_14_1566 ();
 sg13g2_decap_8 FILLER_14_1573 ();
 sg13g2_decap_8 FILLER_14_1580 ();
 sg13g2_decap_8 FILLER_14_1587 ();
 sg13g2_decap_8 FILLER_14_1594 ();
 sg13g2_decap_8 FILLER_14_1601 ();
 sg13g2_decap_8 FILLER_14_1608 ();
 sg13g2_decap_8 FILLER_14_1615 ();
 sg13g2_decap_8 FILLER_14_1622 ();
 sg13g2_decap_8 FILLER_14_1629 ();
 sg13g2_decap_8 FILLER_14_1636 ();
 sg13g2_decap_8 FILLER_14_1643 ();
 sg13g2_decap_8 FILLER_14_1650 ();
 sg13g2_decap_8 FILLER_14_1657 ();
 sg13g2_decap_8 FILLER_14_1664 ();
 sg13g2_decap_8 FILLER_14_1671 ();
 sg13g2_decap_8 FILLER_14_1678 ();
 sg13g2_decap_8 FILLER_14_1685 ();
 sg13g2_decap_8 FILLER_14_1692 ();
 sg13g2_decap_8 FILLER_14_1699 ();
 sg13g2_decap_8 FILLER_14_1706 ();
 sg13g2_decap_8 FILLER_14_1713 ();
 sg13g2_decap_8 FILLER_14_1720 ();
 sg13g2_decap_8 FILLER_14_1727 ();
 sg13g2_decap_8 FILLER_14_1734 ();
 sg13g2_decap_8 FILLER_14_1741 ();
 sg13g2_decap_8 FILLER_14_1748 ();
 sg13g2_decap_8 FILLER_14_1755 ();
 sg13g2_decap_4 FILLER_14_1762 ();
 sg13g2_fill_2 FILLER_14_1766 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_4 FILLER_15_60 ();
 sg13g2_fill_1 FILLER_15_64 ();
 sg13g2_decap_4 FILLER_15_78 ();
 sg13g2_fill_1 FILLER_15_82 ();
 sg13g2_fill_2 FILLER_15_119 ();
 sg13g2_fill_1 FILLER_15_121 ();
 sg13g2_fill_2 FILLER_15_148 ();
 sg13g2_fill_2 FILLER_15_170 ();
 sg13g2_fill_2 FILLER_15_323 ();
 sg13g2_fill_1 FILLER_15_325 ();
 sg13g2_fill_2 FILLER_15_335 ();
 sg13g2_fill_1 FILLER_15_346 ();
 sg13g2_decap_4 FILLER_15_372 ();
 sg13g2_fill_2 FILLER_15_376 ();
 sg13g2_fill_2 FILLER_15_395 ();
 sg13g2_fill_1 FILLER_15_397 ();
 sg13g2_fill_2 FILLER_15_402 ();
 sg13g2_fill_2 FILLER_15_422 ();
 sg13g2_fill_1 FILLER_15_424 ();
 sg13g2_fill_1 FILLER_15_436 ();
 sg13g2_fill_2 FILLER_15_451 ();
 sg13g2_fill_1 FILLER_15_453 ();
 sg13g2_fill_2 FILLER_15_505 ();
 sg13g2_fill_1 FILLER_15_514 ();
 sg13g2_decap_8 FILLER_15_531 ();
 sg13g2_decap_4 FILLER_15_543 ();
 sg13g2_fill_2 FILLER_15_547 ();
 sg13g2_fill_1 FILLER_15_552 ();
 sg13g2_fill_1 FILLER_15_557 ();
 sg13g2_fill_2 FILLER_15_563 ();
 sg13g2_fill_2 FILLER_15_574 ();
 sg13g2_fill_1 FILLER_15_576 ();
 sg13g2_fill_1 FILLER_15_581 ();
 sg13g2_fill_2 FILLER_15_632 ();
 sg13g2_fill_1 FILLER_15_634 ();
 sg13g2_fill_2 FILLER_15_647 ();
 sg13g2_fill_1 FILLER_15_662 ();
 sg13g2_decap_8 FILLER_15_675 ();
 sg13g2_fill_1 FILLER_15_686 ();
 sg13g2_decap_4 FILLER_15_704 ();
 sg13g2_fill_2 FILLER_15_708 ();
 sg13g2_fill_2 FILLER_15_723 ();
 sg13g2_fill_1 FILLER_15_751 ();
 sg13g2_fill_2 FILLER_15_773 ();
 sg13g2_fill_1 FILLER_15_775 ();
 sg13g2_decap_8 FILLER_15_797 ();
 sg13g2_decap_8 FILLER_15_804 ();
 sg13g2_decap_8 FILLER_15_811 ();
 sg13g2_decap_8 FILLER_15_818 ();
 sg13g2_decap_8 FILLER_15_825 ();
 sg13g2_decap_8 FILLER_15_832 ();
 sg13g2_decap_8 FILLER_15_839 ();
 sg13g2_decap_8 FILLER_15_846 ();
 sg13g2_decap_8 FILLER_15_853 ();
 sg13g2_decap_8 FILLER_15_860 ();
 sg13g2_decap_8 FILLER_15_867 ();
 sg13g2_decap_8 FILLER_15_874 ();
 sg13g2_decap_8 FILLER_15_881 ();
 sg13g2_decap_8 FILLER_15_888 ();
 sg13g2_decap_8 FILLER_15_895 ();
 sg13g2_decap_8 FILLER_15_902 ();
 sg13g2_decap_8 FILLER_15_909 ();
 sg13g2_decap_8 FILLER_15_916 ();
 sg13g2_decap_8 FILLER_15_923 ();
 sg13g2_decap_8 FILLER_15_930 ();
 sg13g2_decap_8 FILLER_15_937 ();
 sg13g2_decap_8 FILLER_15_944 ();
 sg13g2_decap_8 FILLER_15_951 ();
 sg13g2_decap_8 FILLER_15_958 ();
 sg13g2_decap_8 FILLER_15_965 ();
 sg13g2_decap_8 FILLER_15_972 ();
 sg13g2_decap_8 FILLER_15_979 ();
 sg13g2_decap_8 FILLER_15_986 ();
 sg13g2_decap_8 FILLER_15_993 ();
 sg13g2_decap_8 FILLER_15_1000 ();
 sg13g2_decap_8 FILLER_15_1007 ();
 sg13g2_decap_8 FILLER_15_1014 ();
 sg13g2_decap_8 FILLER_15_1021 ();
 sg13g2_decap_8 FILLER_15_1028 ();
 sg13g2_decap_8 FILLER_15_1035 ();
 sg13g2_decap_8 FILLER_15_1042 ();
 sg13g2_decap_8 FILLER_15_1049 ();
 sg13g2_decap_8 FILLER_15_1056 ();
 sg13g2_decap_8 FILLER_15_1063 ();
 sg13g2_decap_8 FILLER_15_1070 ();
 sg13g2_decap_8 FILLER_15_1077 ();
 sg13g2_decap_8 FILLER_15_1084 ();
 sg13g2_decap_8 FILLER_15_1091 ();
 sg13g2_decap_8 FILLER_15_1098 ();
 sg13g2_decap_8 FILLER_15_1105 ();
 sg13g2_decap_8 FILLER_15_1112 ();
 sg13g2_decap_8 FILLER_15_1119 ();
 sg13g2_decap_8 FILLER_15_1126 ();
 sg13g2_decap_8 FILLER_15_1133 ();
 sg13g2_decap_8 FILLER_15_1140 ();
 sg13g2_decap_8 FILLER_15_1147 ();
 sg13g2_decap_8 FILLER_15_1154 ();
 sg13g2_decap_8 FILLER_15_1161 ();
 sg13g2_decap_8 FILLER_15_1168 ();
 sg13g2_decap_8 FILLER_15_1175 ();
 sg13g2_decap_8 FILLER_15_1182 ();
 sg13g2_decap_8 FILLER_15_1189 ();
 sg13g2_decap_8 FILLER_15_1196 ();
 sg13g2_decap_8 FILLER_15_1203 ();
 sg13g2_decap_8 FILLER_15_1210 ();
 sg13g2_decap_8 FILLER_15_1217 ();
 sg13g2_decap_8 FILLER_15_1224 ();
 sg13g2_decap_8 FILLER_15_1231 ();
 sg13g2_decap_8 FILLER_15_1238 ();
 sg13g2_decap_8 FILLER_15_1245 ();
 sg13g2_decap_8 FILLER_15_1252 ();
 sg13g2_decap_8 FILLER_15_1259 ();
 sg13g2_decap_8 FILLER_15_1266 ();
 sg13g2_decap_8 FILLER_15_1273 ();
 sg13g2_decap_8 FILLER_15_1280 ();
 sg13g2_decap_8 FILLER_15_1287 ();
 sg13g2_decap_8 FILLER_15_1294 ();
 sg13g2_decap_8 FILLER_15_1301 ();
 sg13g2_decap_8 FILLER_15_1308 ();
 sg13g2_decap_8 FILLER_15_1315 ();
 sg13g2_decap_8 FILLER_15_1322 ();
 sg13g2_decap_8 FILLER_15_1329 ();
 sg13g2_decap_8 FILLER_15_1336 ();
 sg13g2_decap_8 FILLER_15_1343 ();
 sg13g2_decap_8 FILLER_15_1350 ();
 sg13g2_decap_8 FILLER_15_1357 ();
 sg13g2_decap_8 FILLER_15_1364 ();
 sg13g2_decap_8 FILLER_15_1371 ();
 sg13g2_decap_8 FILLER_15_1378 ();
 sg13g2_decap_8 FILLER_15_1385 ();
 sg13g2_decap_8 FILLER_15_1392 ();
 sg13g2_decap_8 FILLER_15_1399 ();
 sg13g2_decap_8 FILLER_15_1406 ();
 sg13g2_decap_8 FILLER_15_1413 ();
 sg13g2_decap_8 FILLER_15_1420 ();
 sg13g2_decap_8 FILLER_15_1427 ();
 sg13g2_decap_8 FILLER_15_1434 ();
 sg13g2_decap_8 FILLER_15_1441 ();
 sg13g2_decap_8 FILLER_15_1448 ();
 sg13g2_decap_8 FILLER_15_1455 ();
 sg13g2_decap_8 FILLER_15_1462 ();
 sg13g2_decap_8 FILLER_15_1469 ();
 sg13g2_decap_8 FILLER_15_1476 ();
 sg13g2_decap_8 FILLER_15_1483 ();
 sg13g2_decap_8 FILLER_15_1490 ();
 sg13g2_decap_8 FILLER_15_1497 ();
 sg13g2_decap_8 FILLER_15_1504 ();
 sg13g2_decap_8 FILLER_15_1511 ();
 sg13g2_decap_8 FILLER_15_1518 ();
 sg13g2_decap_8 FILLER_15_1525 ();
 sg13g2_decap_8 FILLER_15_1532 ();
 sg13g2_decap_8 FILLER_15_1539 ();
 sg13g2_decap_8 FILLER_15_1546 ();
 sg13g2_decap_8 FILLER_15_1553 ();
 sg13g2_decap_8 FILLER_15_1560 ();
 sg13g2_decap_8 FILLER_15_1567 ();
 sg13g2_decap_8 FILLER_15_1574 ();
 sg13g2_decap_8 FILLER_15_1581 ();
 sg13g2_decap_8 FILLER_15_1588 ();
 sg13g2_decap_8 FILLER_15_1595 ();
 sg13g2_decap_8 FILLER_15_1602 ();
 sg13g2_decap_8 FILLER_15_1609 ();
 sg13g2_decap_8 FILLER_15_1616 ();
 sg13g2_decap_8 FILLER_15_1623 ();
 sg13g2_decap_8 FILLER_15_1630 ();
 sg13g2_decap_8 FILLER_15_1637 ();
 sg13g2_decap_8 FILLER_15_1644 ();
 sg13g2_decap_8 FILLER_15_1651 ();
 sg13g2_decap_8 FILLER_15_1658 ();
 sg13g2_decap_8 FILLER_15_1665 ();
 sg13g2_decap_8 FILLER_15_1672 ();
 sg13g2_decap_8 FILLER_15_1679 ();
 sg13g2_decap_8 FILLER_15_1686 ();
 sg13g2_decap_8 FILLER_15_1693 ();
 sg13g2_decap_8 FILLER_15_1700 ();
 sg13g2_decap_8 FILLER_15_1707 ();
 sg13g2_decap_8 FILLER_15_1714 ();
 sg13g2_decap_8 FILLER_15_1721 ();
 sg13g2_decap_8 FILLER_15_1728 ();
 sg13g2_decap_8 FILLER_15_1735 ();
 sg13g2_decap_8 FILLER_15_1742 ();
 sg13g2_decap_8 FILLER_15_1749 ();
 sg13g2_decap_8 FILLER_15_1756 ();
 sg13g2_decap_4 FILLER_15_1763 ();
 sg13g2_fill_1 FILLER_15_1767 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_14 ();
 sg13g2_fill_1 FILLER_16_42 ();
 sg13g2_decap_4 FILLER_16_80 ();
 sg13g2_decap_8 FILLER_16_95 ();
 sg13g2_decap_8 FILLER_16_102 ();
 sg13g2_decap_8 FILLER_16_109 ();
 sg13g2_fill_2 FILLER_16_147 ();
 sg13g2_fill_1 FILLER_16_149 ();
 sg13g2_fill_2 FILLER_16_161 ();
 sg13g2_fill_1 FILLER_16_163 ();
 sg13g2_fill_2 FILLER_16_181 ();
 sg13g2_fill_1 FILLER_16_183 ();
 sg13g2_fill_2 FILLER_16_206 ();
 sg13g2_fill_1 FILLER_16_217 ();
 sg13g2_fill_1 FILLER_16_227 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_fill_1 FILLER_16_259 ();
 sg13g2_fill_1 FILLER_16_269 ();
 sg13g2_fill_2 FILLER_16_280 ();
 sg13g2_fill_2 FILLER_16_305 ();
 sg13g2_fill_1 FILLER_16_307 ();
 sg13g2_fill_2 FILLER_16_381 ();
 sg13g2_fill_2 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_405 ();
 sg13g2_fill_1 FILLER_16_412 ();
 sg13g2_fill_2 FILLER_16_426 ();
 sg13g2_fill_2 FILLER_16_475 ();
 sg13g2_decap_8 FILLER_16_487 ();
 sg13g2_fill_2 FILLER_16_494 ();
 sg13g2_fill_2 FILLER_16_506 ();
 sg13g2_fill_1 FILLER_16_508 ();
 sg13g2_fill_1 FILLER_16_514 ();
 sg13g2_decap_8 FILLER_16_519 ();
 sg13g2_fill_1 FILLER_16_526 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_fill_2 FILLER_16_539 ();
 sg13g2_fill_2 FILLER_16_549 ();
 sg13g2_fill_1 FILLER_16_559 ();
 sg13g2_fill_1 FILLER_16_565 ();
 sg13g2_decap_8 FILLER_16_597 ();
 sg13g2_fill_2 FILLER_16_604 ();
 sg13g2_decap_8 FILLER_16_610 ();
 sg13g2_decap_8 FILLER_16_617 ();
 sg13g2_decap_4 FILLER_16_624 ();
 sg13g2_fill_2 FILLER_16_628 ();
 sg13g2_fill_2 FILLER_16_635 ();
 sg13g2_decap_4 FILLER_16_649 ();
 sg13g2_fill_1 FILLER_16_653 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_fill_2 FILLER_16_679 ();
 sg13g2_fill_1 FILLER_16_681 ();
 sg13g2_decap_8 FILLER_16_694 ();
 sg13g2_decap_8 FILLER_16_701 ();
 sg13g2_decap_8 FILLER_16_716 ();
 sg13g2_decap_4 FILLER_16_723 ();
 sg13g2_fill_1 FILLER_16_727 ();
 sg13g2_fill_2 FILLER_16_731 ();
 sg13g2_fill_1 FILLER_16_733 ();
 sg13g2_decap_4 FILLER_16_755 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_fill_2 FILLER_16_784 ();
 sg13g2_fill_1 FILLER_16_786 ();
 sg13g2_decap_8 FILLER_16_797 ();
 sg13g2_decap_8 FILLER_16_804 ();
 sg13g2_decap_8 FILLER_16_811 ();
 sg13g2_decap_8 FILLER_16_818 ();
 sg13g2_decap_8 FILLER_16_825 ();
 sg13g2_decap_8 FILLER_16_832 ();
 sg13g2_decap_8 FILLER_16_839 ();
 sg13g2_decap_8 FILLER_16_846 ();
 sg13g2_decap_8 FILLER_16_853 ();
 sg13g2_decap_8 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_16_867 ();
 sg13g2_decap_8 FILLER_16_874 ();
 sg13g2_decap_8 FILLER_16_881 ();
 sg13g2_decap_8 FILLER_16_888 ();
 sg13g2_decap_8 FILLER_16_895 ();
 sg13g2_decap_8 FILLER_16_902 ();
 sg13g2_decap_8 FILLER_16_909 ();
 sg13g2_decap_8 FILLER_16_916 ();
 sg13g2_decap_8 FILLER_16_923 ();
 sg13g2_decap_8 FILLER_16_930 ();
 sg13g2_decap_8 FILLER_16_937 ();
 sg13g2_decap_8 FILLER_16_944 ();
 sg13g2_decap_8 FILLER_16_951 ();
 sg13g2_decap_8 FILLER_16_958 ();
 sg13g2_decap_8 FILLER_16_965 ();
 sg13g2_decap_8 FILLER_16_972 ();
 sg13g2_decap_8 FILLER_16_979 ();
 sg13g2_decap_8 FILLER_16_986 ();
 sg13g2_decap_8 FILLER_16_993 ();
 sg13g2_decap_8 FILLER_16_1000 ();
 sg13g2_decap_8 FILLER_16_1007 ();
 sg13g2_decap_8 FILLER_16_1014 ();
 sg13g2_decap_8 FILLER_16_1021 ();
 sg13g2_decap_8 FILLER_16_1028 ();
 sg13g2_decap_8 FILLER_16_1035 ();
 sg13g2_decap_8 FILLER_16_1042 ();
 sg13g2_decap_8 FILLER_16_1049 ();
 sg13g2_decap_8 FILLER_16_1056 ();
 sg13g2_decap_8 FILLER_16_1063 ();
 sg13g2_decap_8 FILLER_16_1070 ();
 sg13g2_decap_8 FILLER_16_1077 ();
 sg13g2_decap_8 FILLER_16_1084 ();
 sg13g2_decap_8 FILLER_16_1091 ();
 sg13g2_decap_8 FILLER_16_1098 ();
 sg13g2_decap_8 FILLER_16_1105 ();
 sg13g2_decap_8 FILLER_16_1112 ();
 sg13g2_decap_8 FILLER_16_1119 ();
 sg13g2_decap_8 FILLER_16_1126 ();
 sg13g2_decap_8 FILLER_16_1133 ();
 sg13g2_decap_8 FILLER_16_1140 ();
 sg13g2_decap_8 FILLER_16_1147 ();
 sg13g2_decap_8 FILLER_16_1154 ();
 sg13g2_decap_8 FILLER_16_1161 ();
 sg13g2_decap_8 FILLER_16_1168 ();
 sg13g2_decap_8 FILLER_16_1175 ();
 sg13g2_decap_8 FILLER_16_1182 ();
 sg13g2_decap_8 FILLER_16_1189 ();
 sg13g2_decap_8 FILLER_16_1196 ();
 sg13g2_decap_8 FILLER_16_1203 ();
 sg13g2_decap_8 FILLER_16_1210 ();
 sg13g2_decap_8 FILLER_16_1217 ();
 sg13g2_decap_8 FILLER_16_1224 ();
 sg13g2_decap_8 FILLER_16_1231 ();
 sg13g2_decap_8 FILLER_16_1238 ();
 sg13g2_decap_8 FILLER_16_1245 ();
 sg13g2_decap_8 FILLER_16_1252 ();
 sg13g2_decap_8 FILLER_16_1259 ();
 sg13g2_decap_8 FILLER_16_1266 ();
 sg13g2_decap_8 FILLER_16_1273 ();
 sg13g2_decap_8 FILLER_16_1280 ();
 sg13g2_decap_8 FILLER_16_1287 ();
 sg13g2_decap_8 FILLER_16_1294 ();
 sg13g2_decap_8 FILLER_16_1301 ();
 sg13g2_decap_8 FILLER_16_1308 ();
 sg13g2_decap_8 FILLER_16_1315 ();
 sg13g2_decap_8 FILLER_16_1322 ();
 sg13g2_decap_8 FILLER_16_1329 ();
 sg13g2_decap_8 FILLER_16_1336 ();
 sg13g2_decap_8 FILLER_16_1343 ();
 sg13g2_decap_8 FILLER_16_1350 ();
 sg13g2_decap_8 FILLER_16_1357 ();
 sg13g2_decap_8 FILLER_16_1364 ();
 sg13g2_decap_8 FILLER_16_1371 ();
 sg13g2_decap_8 FILLER_16_1378 ();
 sg13g2_decap_8 FILLER_16_1385 ();
 sg13g2_decap_8 FILLER_16_1392 ();
 sg13g2_decap_8 FILLER_16_1399 ();
 sg13g2_decap_8 FILLER_16_1406 ();
 sg13g2_decap_8 FILLER_16_1413 ();
 sg13g2_decap_8 FILLER_16_1420 ();
 sg13g2_decap_8 FILLER_16_1427 ();
 sg13g2_decap_8 FILLER_16_1434 ();
 sg13g2_decap_8 FILLER_16_1441 ();
 sg13g2_decap_8 FILLER_16_1448 ();
 sg13g2_decap_8 FILLER_16_1455 ();
 sg13g2_decap_8 FILLER_16_1462 ();
 sg13g2_decap_8 FILLER_16_1469 ();
 sg13g2_decap_8 FILLER_16_1476 ();
 sg13g2_decap_8 FILLER_16_1483 ();
 sg13g2_decap_8 FILLER_16_1490 ();
 sg13g2_decap_8 FILLER_16_1497 ();
 sg13g2_decap_8 FILLER_16_1504 ();
 sg13g2_decap_8 FILLER_16_1511 ();
 sg13g2_decap_8 FILLER_16_1518 ();
 sg13g2_decap_8 FILLER_16_1525 ();
 sg13g2_decap_8 FILLER_16_1532 ();
 sg13g2_decap_8 FILLER_16_1539 ();
 sg13g2_decap_8 FILLER_16_1546 ();
 sg13g2_decap_8 FILLER_16_1553 ();
 sg13g2_decap_8 FILLER_16_1560 ();
 sg13g2_decap_8 FILLER_16_1567 ();
 sg13g2_decap_8 FILLER_16_1574 ();
 sg13g2_decap_8 FILLER_16_1581 ();
 sg13g2_decap_8 FILLER_16_1588 ();
 sg13g2_decap_8 FILLER_16_1595 ();
 sg13g2_decap_8 FILLER_16_1602 ();
 sg13g2_decap_8 FILLER_16_1609 ();
 sg13g2_decap_8 FILLER_16_1616 ();
 sg13g2_decap_8 FILLER_16_1623 ();
 sg13g2_decap_8 FILLER_16_1630 ();
 sg13g2_decap_8 FILLER_16_1637 ();
 sg13g2_decap_8 FILLER_16_1644 ();
 sg13g2_decap_8 FILLER_16_1651 ();
 sg13g2_decap_8 FILLER_16_1658 ();
 sg13g2_decap_8 FILLER_16_1665 ();
 sg13g2_decap_8 FILLER_16_1672 ();
 sg13g2_decap_8 FILLER_16_1679 ();
 sg13g2_decap_8 FILLER_16_1686 ();
 sg13g2_decap_8 FILLER_16_1693 ();
 sg13g2_decap_8 FILLER_16_1700 ();
 sg13g2_decap_8 FILLER_16_1707 ();
 sg13g2_decap_8 FILLER_16_1714 ();
 sg13g2_decap_8 FILLER_16_1721 ();
 sg13g2_decap_8 FILLER_16_1728 ();
 sg13g2_decap_8 FILLER_16_1735 ();
 sg13g2_decap_8 FILLER_16_1742 ();
 sg13g2_decap_8 FILLER_16_1749 ();
 sg13g2_decap_8 FILLER_16_1756 ();
 sg13g2_decap_4 FILLER_16_1763 ();
 sg13g2_fill_1 FILLER_16_1767 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_21 ();
 sg13g2_fill_2 FILLER_17_36 ();
 sg13g2_decap_8 FILLER_17_46 ();
 sg13g2_decap_4 FILLER_17_53 ();
 sg13g2_fill_1 FILLER_17_57 ();
 sg13g2_fill_2 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_69 ();
 sg13g2_fill_2 FILLER_17_76 ();
 sg13g2_fill_1 FILLER_17_78 ();
 sg13g2_fill_2 FILLER_17_127 ();
 sg13g2_fill_1 FILLER_17_129 ();
 sg13g2_fill_2 FILLER_17_145 ();
 sg13g2_fill_1 FILLER_17_147 ();
 sg13g2_fill_2 FILLER_17_183 ();
 sg13g2_fill_2 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_228 ();
 sg13g2_fill_2 FILLER_17_429 ();
 sg13g2_fill_1 FILLER_17_431 ();
 sg13g2_decap_4 FILLER_17_449 ();
 sg13g2_fill_2 FILLER_17_480 ();
 sg13g2_fill_2 FILLER_17_508 ();
 sg13g2_fill_2 FILLER_17_518 ();
 sg13g2_fill_1 FILLER_17_520 ();
 sg13g2_decap_8 FILLER_17_537 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_fill_2 FILLER_17_560 ();
 sg13g2_fill_1 FILLER_17_562 ();
 sg13g2_decap_8 FILLER_17_568 ();
 sg13g2_fill_1 FILLER_17_575 ();
 sg13g2_fill_1 FILLER_17_643 ();
 sg13g2_fill_2 FILLER_17_667 ();
 sg13g2_fill_1 FILLER_17_673 ();
 sg13g2_fill_2 FILLER_17_694 ();
 sg13g2_fill_2 FILLER_17_725 ();
 sg13g2_decap_8 FILLER_17_732 ();
 sg13g2_decap_4 FILLER_17_742 ();
 sg13g2_decap_4 FILLER_17_751 ();
 sg13g2_decap_8 FILLER_17_760 ();
 sg13g2_fill_1 FILLER_17_767 ();
 sg13g2_fill_1 FILLER_17_775 ();
 sg13g2_decap_4 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_decap_8 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_17_868 ();
 sg13g2_decap_8 FILLER_17_875 ();
 sg13g2_decap_8 FILLER_17_882 ();
 sg13g2_decap_8 FILLER_17_889 ();
 sg13g2_decap_8 FILLER_17_896 ();
 sg13g2_decap_8 FILLER_17_903 ();
 sg13g2_decap_8 FILLER_17_910 ();
 sg13g2_decap_8 FILLER_17_917 ();
 sg13g2_decap_8 FILLER_17_924 ();
 sg13g2_decap_8 FILLER_17_931 ();
 sg13g2_decap_8 FILLER_17_938 ();
 sg13g2_decap_8 FILLER_17_945 ();
 sg13g2_decap_8 FILLER_17_952 ();
 sg13g2_decap_8 FILLER_17_959 ();
 sg13g2_decap_8 FILLER_17_966 ();
 sg13g2_decap_8 FILLER_17_973 ();
 sg13g2_decap_8 FILLER_17_980 ();
 sg13g2_decap_8 FILLER_17_987 ();
 sg13g2_decap_8 FILLER_17_994 ();
 sg13g2_decap_8 FILLER_17_1001 ();
 sg13g2_decap_8 FILLER_17_1008 ();
 sg13g2_decap_8 FILLER_17_1015 ();
 sg13g2_decap_8 FILLER_17_1022 ();
 sg13g2_decap_8 FILLER_17_1029 ();
 sg13g2_decap_8 FILLER_17_1036 ();
 sg13g2_decap_8 FILLER_17_1043 ();
 sg13g2_decap_8 FILLER_17_1050 ();
 sg13g2_decap_8 FILLER_17_1057 ();
 sg13g2_decap_8 FILLER_17_1064 ();
 sg13g2_decap_8 FILLER_17_1071 ();
 sg13g2_decap_8 FILLER_17_1078 ();
 sg13g2_decap_8 FILLER_17_1085 ();
 sg13g2_decap_8 FILLER_17_1092 ();
 sg13g2_decap_8 FILLER_17_1099 ();
 sg13g2_decap_8 FILLER_17_1106 ();
 sg13g2_decap_8 FILLER_17_1113 ();
 sg13g2_decap_8 FILLER_17_1120 ();
 sg13g2_decap_8 FILLER_17_1127 ();
 sg13g2_decap_8 FILLER_17_1134 ();
 sg13g2_decap_8 FILLER_17_1141 ();
 sg13g2_decap_8 FILLER_17_1148 ();
 sg13g2_decap_8 FILLER_17_1155 ();
 sg13g2_decap_8 FILLER_17_1162 ();
 sg13g2_decap_8 FILLER_17_1169 ();
 sg13g2_decap_8 FILLER_17_1176 ();
 sg13g2_decap_8 FILLER_17_1183 ();
 sg13g2_decap_8 FILLER_17_1190 ();
 sg13g2_decap_8 FILLER_17_1197 ();
 sg13g2_decap_8 FILLER_17_1204 ();
 sg13g2_decap_8 FILLER_17_1211 ();
 sg13g2_decap_8 FILLER_17_1218 ();
 sg13g2_decap_8 FILLER_17_1225 ();
 sg13g2_decap_8 FILLER_17_1232 ();
 sg13g2_decap_8 FILLER_17_1239 ();
 sg13g2_decap_8 FILLER_17_1246 ();
 sg13g2_decap_8 FILLER_17_1253 ();
 sg13g2_decap_8 FILLER_17_1260 ();
 sg13g2_decap_8 FILLER_17_1267 ();
 sg13g2_decap_8 FILLER_17_1274 ();
 sg13g2_decap_8 FILLER_17_1281 ();
 sg13g2_decap_8 FILLER_17_1288 ();
 sg13g2_decap_8 FILLER_17_1295 ();
 sg13g2_decap_8 FILLER_17_1302 ();
 sg13g2_decap_8 FILLER_17_1309 ();
 sg13g2_decap_8 FILLER_17_1316 ();
 sg13g2_decap_8 FILLER_17_1323 ();
 sg13g2_decap_8 FILLER_17_1330 ();
 sg13g2_decap_8 FILLER_17_1337 ();
 sg13g2_decap_8 FILLER_17_1344 ();
 sg13g2_decap_8 FILLER_17_1351 ();
 sg13g2_decap_8 FILLER_17_1358 ();
 sg13g2_decap_8 FILLER_17_1365 ();
 sg13g2_decap_8 FILLER_17_1372 ();
 sg13g2_decap_8 FILLER_17_1379 ();
 sg13g2_decap_8 FILLER_17_1386 ();
 sg13g2_decap_8 FILLER_17_1393 ();
 sg13g2_decap_8 FILLER_17_1400 ();
 sg13g2_decap_8 FILLER_17_1407 ();
 sg13g2_decap_8 FILLER_17_1414 ();
 sg13g2_decap_8 FILLER_17_1421 ();
 sg13g2_decap_8 FILLER_17_1428 ();
 sg13g2_decap_8 FILLER_17_1435 ();
 sg13g2_decap_8 FILLER_17_1442 ();
 sg13g2_decap_8 FILLER_17_1449 ();
 sg13g2_decap_8 FILLER_17_1456 ();
 sg13g2_decap_8 FILLER_17_1463 ();
 sg13g2_decap_8 FILLER_17_1470 ();
 sg13g2_decap_8 FILLER_17_1477 ();
 sg13g2_decap_8 FILLER_17_1484 ();
 sg13g2_decap_8 FILLER_17_1491 ();
 sg13g2_decap_8 FILLER_17_1498 ();
 sg13g2_decap_8 FILLER_17_1505 ();
 sg13g2_decap_8 FILLER_17_1512 ();
 sg13g2_decap_8 FILLER_17_1519 ();
 sg13g2_decap_8 FILLER_17_1526 ();
 sg13g2_decap_8 FILLER_17_1533 ();
 sg13g2_decap_8 FILLER_17_1540 ();
 sg13g2_decap_8 FILLER_17_1547 ();
 sg13g2_decap_8 FILLER_17_1554 ();
 sg13g2_decap_8 FILLER_17_1561 ();
 sg13g2_decap_8 FILLER_17_1568 ();
 sg13g2_decap_8 FILLER_17_1575 ();
 sg13g2_decap_8 FILLER_17_1582 ();
 sg13g2_decap_8 FILLER_17_1589 ();
 sg13g2_decap_8 FILLER_17_1596 ();
 sg13g2_decap_8 FILLER_17_1603 ();
 sg13g2_decap_8 FILLER_17_1610 ();
 sg13g2_decap_8 FILLER_17_1617 ();
 sg13g2_decap_8 FILLER_17_1624 ();
 sg13g2_decap_8 FILLER_17_1631 ();
 sg13g2_decap_8 FILLER_17_1638 ();
 sg13g2_decap_8 FILLER_17_1645 ();
 sg13g2_decap_8 FILLER_17_1652 ();
 sg13g2_decap_8 FILLER_17_1659 ();
 sg13g2_decap_8 FILLER_17_1666 ();
 sg13g2_decap_8 FILLER_17_1673 ();
 sg13g2_decap_8 FILLER_17_1680 ();
 sg13g2_decap_8 FILLER_17_1687 ();
 sg13g2_decap_8 FILLER_17_1694 ();
 sg13g2_decap_8 FILLER_17_1701 ();
 sg13g2_decap_8 FILLER_17_1708 ();
 sg13g2_decap_8 FILLER_17_1715 ();
 sg13g2_decap_8 FILLER_17_1722 ();
 sg13g2_decap_8 FILLER_17_1729 ();
 sg13g2_decap_8 FILLER_17_1736 ();
 sg13g2_decap_8 FILLER_17_1743 ();
 sg13g2_decap_8 FILLER_17_1750 ();
 sg13g2_decap_8 FILLER_17_1757 ();
 sg13g2_decap_4 FILLER_17_1764 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_4 ();
 sg13g2_decap_8 FILLER_18_57 ();
 sg13g2_decap_4 FILLER_18_64 ();
 sg13g2_fill_2 FILLER_18_68 ();
 sg13g2_fill_2 FILLER_18_93 ();
 sg13g2_decap_8 FILLER_18_100 ();
 sg13g2_fill_2 FILLER_18_107 ();
 sg13g2_fill_2 FILLER_18_122 ();
 sg13g2_fill_1 FILLER_18_124 ();
 sg13g2_fill_1 FILLER_18_157 ();
 sg13g2_fill_1 FILLER_18_167 ();
 sg13g2_decap_8 FILLER_18_194 ();
 sg13g2_fill_2 FILLER_18_201 ();
 sg13g2_fill_1 FILLER_18_203 ();
 sg13g2_fill_1 FILLER_18_249 ();
 sg13g2_fill_2 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_282 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_fill_2 FILLER_18_309 ();
 sg13g2_fill_2 FILLER_18_324 ();
 sg13g2_fill_1 FILLER_18_326 ();
 sg13g2_fill_2 FILLER_18_363 ();
 sg13g2_fill_1 FILLER_18_365 ();
 sg13g2_fill_1 FILLER_18_411 ();
 sg13g2_fill_1 FILLER_18_422 ();
 sg13g2_decap_4 FILLER_18_469 ();
 sg13g2_fill_2 FILLER_18_489 ();
 sg13g2_fill_2 FILLER_18_499 ();
 sg13g2_fill_2 FILLER_18_522 ();
 sg13g2_fill_1 FILLER_18_524 ();
 sg13g2_fill_2 FILLER_18_541 ();
 sg13g2_fill_1 FILLER_18_543 ();
 sg13g2_fill_2 FILLER_18_552 ();
 sg13g2_decap_4 FILLER_18_566 ();
 sg13g2_fill_1 FILLER_18_570 ();
 sg13g2_fill_2 FILLER_18_581 ();
 sg13g2_fill_1 FILLER_18_583 ();
 sg13g2_decap_8 FILLER_18_598 ();
 sg13g2_fill_1 FILLER_18_628 ();
 sg13g2_decap_4 FILLER_18_645 ();
 sg13g2_decap_8 FILLER_18_667 ();
 sg13g2_decap_8 FILLER_18_674 ();
 sg13g2_fill_1 FILLER_18_681 ();
 sg13g2_fill_1 FILLER_18_700 ();
 sg13g2_fill_2 FILLER_18_719 ();
 sg13g2_fill_2 FILLER_18_742 ();
 sg13g2_fill_1 FILLER_18_744 ();
 sg13g2_fill_2 FILLER_18_758 ();
 sg13g2_fill_1 FILLER_18_760 ();
 sg13g2_decap_4 FILLER_18_769 ();
 sg13g2_fill_2 FILLER_18_773 ();
 sg13g2_decap_8 FILLER_18_795 ();
 sg13g2_decap_8 FILLER_18_802 ();
 sg13g2_fill_1 FILLER_18_809 ();
 sg13g2_decap_8 FILLER_18_860 ();
 sg13g2_decap_8 FILLER_18_867 ();
 sg13g2_fill_1 FILLER_18_874 ();
 sg13g2_decap_8 FILLER_18_880 ();
 sg13g2_decap_8 FILLER_18_887 ();
 sg13g2_decap_8 FILLER_18_894 ();
 sg13g2_decap_8 FILLER_18_905 ();
 sg13g2_decap_8 FILLER_18_912 ();
 sg13g2_decap_8 FILLER_18_919 ();
 sg13g2_decap_8 FILLER_18_926 ();
 sg13g2_decap_4 FILLER_18_933 ();
 sg13g2_fill_2 FILLER_18_937 ();
 sg13g2_decap_8 FILLER_18_960 ();
 sg13g2_decap_8 FILLER_18_967 ();
 sg13g2_decap_8 FILLER_18_974 ();
 sg13g2_decap_8 FILLER_18_981 ();
 sg13g2_decap_8 FILLER_18_988 ();
 sg13g2_decap_8 FILLER_18_995 ();
 sg13g2_decap_8 FILLER_18_1002 ();
 sg13g2_decap_8 FILLER_18_1009 ();
 sg13g2_decap_8 FILLER_18_1016 ();
 sg13g2_decap_8 FILLER_18_1023 ();
 sg13g2_decap_8 FILLER_18_1030 ();
 sg13g2_decap_8 FILLER_18_1037 ();
 sg13g2_decap_8 FILLER_18_1044 ();
 sg13g2_decap_8 FILLER_18_1051 ();
 sg13g2_decap_8 FILLER_18_1058 ();
 sg13g2_decap_8 FILLER_18_1065 ();
 sg13g2_decap_8 FILLER_18_1072 ();
 sg13g2_decap_8 FILLER_18_1079 ();
 sg13g2_decap_8 FILLER_18_1086 ();
 sg13g2_decap_8 FILLER_18_1093 ();
 sg13g2_decap_8 FILLER_18_1100 ();
 sg13g2_decap_8 FILLER_18_1107 ();
 sg13g2_decap_8 FILLER_18_1114 ();
 sg13g2_decap_8 FILLER_18_1121 ();
 sg13g2_decap_8 FILLER_18_1128 ();
 sg13g2_decap_8 FILLER_18_1135 ();
 sg13g2_decap_8 FILLER_18_1142 ();
 sg13g2_decap_8 FILLER_18_1149 ();
 sg13g2_decap_8 FILLER_18_1156 ();
 sg13g2_decap_8 FILLER_18_1163 ();
 sg13g2_decap_8 FILLER_18_1170 ();
 sg13g2_decap_8 FILLER_18_1177 ();
 sg13g2_decap_8 FILLER_18_1184 ();
 sg13g2_decap_8 FILLER_18_1191 ();
 sg13g2_decap_8 FILLER_18_1198 ();
 sg13g2_decap_8 FILLER_18_1205 ();
 sg13g2_decap_8 FILLER_18_1212 ();
 sg13g2_decap_8 FILLER_18_1219 ();
 sg13g2_decap_8 FILLER_18_1226 ();
 sg13g2_decap_8 FILLER_18_1233 ();
 sg13g2_decap_8 FILLER_18_1240 ();
 sg13g2_decap_8 FILLER_18_1247 ();
 sg13g2_decap_8 FILLER_18_1254 ();
 sg13g2_decap_8 FILLER_18_1261 ();
 sg13g2_decap_8 FILLER_18_1268 ();
 sg13g2_decap_8 FILLER_18_1275 ();
 sg13g2_decap_8 FILLER_18_1282 ();
 sg13g2_decap_8 FILLER_18_1289 ();
 sg13g2_decap_8 FILLER_18_1296 ();
 sg13g2_decap_8 FILLER_18_1303 ();
 sg13g2_decap_8 FILLER_18_1310 ();
 sg13g2_decap_8 FILLER_18_1317 ();
 sg13g2_decap_8 FILLER_18_1324 ();
 sg13g2_decap_8 FILLER_18_1331 ();
 sg13g2_decap_8 FILLER_18_1338 ();
 sg13g2_decap_8 FILLER_18_1345 ();
 sg13g2_decap_8 FILLER_18_1352 ();
 sg13g2_decap_8 FILLER_18_1359 ();
 sg13g2_decap_8 FILLER_18_1366 ();
 sg13g2_decap_8 FILLER_18_1373 ();
 sg13g2_decap_8 FILLER_18_1380 ();
 sg13g2_decap_8 FILLER_18_1387 ();
 sg13g2_decap_8 FILLER_18_1394 ();
 sg13g2_decap_8 FILLER_18_1401 ();
 sg13g2_decap_8 FILLER_18_1408 ();
 sg13g2_decap_8 FILLER_18_1415 ();
 sg13g2_decap_8 FILLER_18_1422 ();
 sg13g2_decap_8 FILLER_18_1429 ();
 sg13g2_decap_8 FILLER_18_1436 ();
 sg13g2_decap_8 FILLER_18_1443 ();
 sg13g2_decap_8 FILLER_18_1450 ();
 sg13g2_decap_8 FILLER_18_1457 ();
 sg13g2_decap_8 FILLER_18_1464 ();
 sg13g2_decap_8 FILLER_18_1471 ();
 sg13g2_decap_8 FILLER_18_1478 ();
 sg13g2_decap_8 FILLER_18_1485 ();
 sg13g2_decap_8 FILLER_18_1492 ();
 sg13g2_decap_8 FILLER_18_1499 ();
 sg13g2_decap_8 FILLER_18_1506 ();
 sg13g2_decap_8 FILLER_18_1513 ();
 sg13g2_decap_8 FILLER_18_1520 ();
 sg13g2_decap_8 FILLER_18_1527 ();
 sg13g2_decap_8 FILLER_18_1534 ();
 sg13g2_decap_8 FILLER_18_1541 ();
 sg13g2_decap_8 FILLER_18_1548 ();
 sg13g2_decap_8 FILLER_18_1555 ();
 sg13g2_decap_8 FILLER_18_1562 ();
 sg13g2_decap_8 FILLER_18_1569 ();
 sg13g2_decap_8 FILLER_18_1576 ();
 sg13g2_decap_8 FILLER_18_1583 ();
 sg13g2_decap_8 FILLER_18_1590 ();
 sg13g2_decap_8 FILLER_18_1597 ();
 sg13g2_decap_8 FILLER_18_1604 ();
 sg13g2_decap_8 FILLER_18_1611 ();
 sg13g2_decap_8 FILLER_18_1618 ();
 sg13g2_decap_8 FILLER_18_1625 ();
 sg13g2_decap_8 FILLER_18_1632 ();
 sg13g2_decap_8 FILLER_18_1639 ();
 sg13g2_decap_8 FILLER_18_1646 ();
 sg13g2_decap_8 FILLER_18_1653 ();
 sg13g2_decap_8 FILLER_18_1660 ();
 sg13g2_decap_8 FILLER_18_1667 ();
 sg13g2_decap_8 FILLER_18_1674 ();
 sg13g2_decap_8 FILLER_18_1681 ();
 sg13g2_decap_8 FILLER_18_1688 ();
 sg13g2_decap_8 FILLER_18_1695 ();
 sg13g2_decap_8 FILLER_18_1702 ();
 sg13g2_decap_8 FILLER_18_1709 ();
 sg13g2_decap_8 FILLER_18_1716 ();
 sg13g2_decap_8 FILLER_18_1723 ();
 sg13g2_decap_8 FILLER_18_1730 ();
 sg13g2_decap_8 FILLER_18_1737 ();
 sg13g2_decap_8 FILLER_18_1744 ();
 sg13g2_decap_8 FILLER_18_1751 ();
 sg13g2_decap_8 FILLER_18_1758 ();
 sg13g2_fill_2 FILLER_18_1765 ();
 sg13g2_fill_1 FILLER_18_1767 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_4 FILLER_19_14 ();
 sg13g2_fill_2 FILLER_19_18 ();
 sg13g2_fill_2 FILLER_19_71 ();
 sg13g2_fill_1 FILLER_19_73 ();
 sg13g2_fill_1 FILLER_19_78 ();
 sg13g2_fill_2 FILLER_19_105 ();
 sg13g2_fill_2 FILLER_19_117 ();
 sg13g2_fill_2 FILLER_19_139 ();
 sg13g2_fill_1 FILLER_19_141 ();
 sg13g2_fill_2 FILLER_19_172 ();
 sg13g2_fill_1 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_179 ();
 sg13g2_fill_2 FILLER_19_226 ();
 sg13g2_fill_2 FILLER_19_238 ();
 sg13g2_fill_1 FILLER_19_240 ();
 sg13g2_fill_2 FILLER_19_294 ();
 sg13g2_fill_1 FILLER_19_300 ();
 sg13g2_fill_2 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_317 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_fill_2 FILLER_19_480 ();
 sg13g2_fill_1 FILLER_19_482 ();
 sg13g2_fill_2 FILLER_19_496 ();
 sg13g2_fill_1 FILLER_19_498 ();
 sg13g2_fill_2 FILLER_19_512 ();
 sg13g2_fill_2 FILLER_19_540 ();
 sg13g2_fill_2 FILLER_19_554 ();
 sg13g2_fill_1 FILLER_19_556 ();
 sg13g2_fill_1 FILLER_19_582 ();
 sg13g2_decap_4 FILLER_19_592 ();
 sg13g2_fill_1 FILLER_19_596 ();
 sg13g2_decap_8 FILLER_19_610 ();
 sg13g2_decap_4 FILLER_19_617 ();
 sg13g2_fill_1 FILLER_19_621 ();
 sg13g2_decap_4 FILLER_19_653 ();
 sg13g2_decap_4 FILLER_19_668 ();
 sg13g2_fill_2 FILLER_19_672 ();
 sg13g2_fill_2 FILLER_19_681 ();
 sg13g2_fill_1 FILLER_19_683 ();
 sg13g2_decap_4 FILLER_19_690 ();
 sg13g2_decap_4 FILLER_19_727 ();
 sg13g2_fill_2 FILLER_19_748 ();
 sg13g2_decap_8 FILLER_19_758 ();
 sg13g2_fill_2 FILLER_19_775 ();
 sg13g2_fill_1 FILLER_19_777 ();
 sg13g2_fill_2 FILLER_19_782 ();
 sg13g2_fill_1 FILLER_19_784 ();
 sg13g2_fill_1 FILLER_19_835 ();
 sg13g2_fill_1 FILLER_19_847 ();
 sg13g2_decap_4 FILLER_19_863 ();
 sg13g2_fill_1 FILLER_19_867 ();
 sg13g2_decap_4 FILLER_19_887 ();
 sg13g2_decap_8 FILLER_19_911 ();
 sg13g2_decap_8 FILLER_19_968 ();
 sg13g2_decap_8 FILLER_19_975 ();
 sg13g2_decap_8 FILLER_19_982 ();
 sg13g2_decap_8 FILLER_19_989 ();
 sg13g2_decap_8 FILLER_19_996 ();
 sg13g2_decap_8 FILLER_19_1003 ();
 sg13g2_decap_8 FILLER_19_1010 ();
 sg13g2_decap_8 FILLER_19_1017 ();
 sg13g2_decap_8 FILLER_19_1024 ();
 sg13g2_decap_8 FILLER_19_1031 ();
 sg13g2_decap_8 FILLER_19_1038 ();
 sg13g2_decap_8 FILLER_19_1045 ();
 sg13g2_decap_8 FILLER_19_1052 ();
 sg13g2_decap_8 FILLER_19_1059 ();
 sg13g2_decap_8 FILLER_19_1066 ();
 sg13g2_decap_8 FILLER_19_1073 ();
 sg13g2_decap_8 FILLER_19_1080 ();
 sg13g2_decap_8 FILLER_19_1087 ();
 sg13g2_decap_8 FILLER_19_1094 ();
 sg13g2_decap_8 FILLER_19_1101 ();
 sg13g2_decap_8 FILLER_19_1108 ();
 sg13g2_decap_8 FILLER_19_1115 ();
 sg13g2_decap_8 FILLER_19_1122 ();
 sg13g2_decap_8 FILLER_19_1129 ();
 sg13g2_decap_8 FILLER_19_1136 ();
 sg13g2_decap_8 FILLER_19_1143 ();
 sg13g2_decap_8 FILLER_19_1150 ();
 sg13g2_decap_8 FILLER_19_1157 ();
 sg13g2_decap_8 FILLER_19_1164 ();
 sg13g2_decap_8 FILLER_19_1171 ();
 sg13g2_decap_8 FILLER_19_1178 ();
 sg13g2_decap_8 FILLER_19_1185 ();
 sg13g2_decap_8 FILLER_19_1192 ();
 sg13g2_decap_8 FILLER_19_1199 ();
 sg13g2_decap_8 FILLER_19_1206 ();
 sg13g2_decap_8 FILLER_19_1213 ();
 sg13g2_decap_8 FILLER_19_1220 ();
 sg13g2_decap_8 FILLER_19_1227 ();
 sg13g2_decap_8 FILLER_19_1234 ();
 sg13g2_decap_8 FILLER_19_1241 ();
 sg13g2_decap_8 FILLER_19_1248 ();
 sg13g2_decap_8 FILLER_19_1255 ();
 sg13g2_decap_8 FILLER_19_1262 ();
 sg13g2_decap_8 FILLER_19_1269 ();
 sg13g2_decap_8 FILLER_19_1276 ();
 sg13g2_decap_8 FILLER_19_1283 ();
 sg13g2_decap_8 FILLER_19_1290 ();
 sg13g2_decap_8 FILLER_19_1297 ();
 sg13g2_decap_8 FILLER_19_1304 ();
 sg13g2_decap_8 FILLER_19_1311 ();
 sg13g2_decap_8 FILLER_19_1318 ();
 sg13g2_decap_8 FILLER_19_1325 ();
 sg13g2_decap_8 FILLER_19_1332 ();
 sg13g2_decap_8 FILLER_19_1339 ();
 sg13g2_decap_8 FILLER_19_1346 ();
 sg13g2_decap_8 FILLER_19_1353 ();
 sg13g2_decap_8 FILLER_19_1360 ();
 sg13g2_decap_8 FILLER_19_1367 ();
 sg13g2_decap_8 FILLER_19_1374 ();
 sg13g2_decap_8 FILLER_19_1381 ();
 sg13g2_decap_8 FILLER_19_1388 ();
 sg13g2_decap_8 FILLER_19_1395 ();
 sg13g2_decap_8 FILLER_19_1402 ();
 sg13g2_decap_8 FILLER_19_1409 ();
 sg13g2_decap_8 FILLER_19_1416 ();
 sg13g2_decap_8 FILLER_19_1423 ();
 sg13g2_decap_8 FILLER_19_1430 ();
 sg13g2_decap_8 FILLER_19_1437 ();
 sg13g2_decap_8 FILLER_19_1444 ();
 sg13g2_decap_8 FILLER_19_1451 ();
 sg13g2_decap_8 FILLER_19_1458 ();
 sg13g2_decap_8 FILLER_19_1465 ();
 sg13g2_decap_8 FILLER_19_1472 ();
 sg13g2_decap_8 FILLER_19_1479 ();
 sg13g2_decap_8 FILLER_19_1486 ();
 sg13g2_decap_8 FILLER_19_1493 ();
 sg13g2_decap_8 FILLER_19_1500 ();
 sg13g2_decap_8 FILLER_19_1507 ();
 sg13g2_decap_8 FILLER_19_1514 ();
 sg13g2_decap_8 FILLER_19_1521 ();
 sg13g2_decap_8 FILLER_19_1528 ();
 sg13g2_decap_8 FILLER_19_1535 ();
 sg13g2_decap_8 FILLER_19_1542 ();
 sg13g2_decap_8 FILLER_19_1549 ();
 sg13g2_decap_8 FILLER_19_1556 ();
 sg13g2_decap_8 FILLER_19_1563 ();
 sg13g2_decap_8 FILLER_19_1570 ();
 sg13g2_decap_8 FILLER_19_1577 ();
 sg13g2_decap_8 FILLER_19_1584 ();
 sg13g2_decap_8 FILLER_19_1591 ();
 sg13g2_decap_8 FILLER_19_1598 ();
 sg13g2_decap_8 FILLER_19_1605 ();
 sg13g2_decap_8 FILLER_19_1612 ();
 sg13g2_decap_8 FILLER_19_1619 ();
 sg13g2_decap_8 FILLER_19_1626 ();
 sg13g2_decap_8 FILLER_19_1633 ();
 sg13g2_decap_8 FILLER_19_1640 ();
 sg13g2_decap_8 FILLER_19_1647 ();
 sg13g2_decap_8 FILLER_19_1654 ();
 sg13g2_decap_8 FILLER_19_1661 ();
 sg13g2_decap_8 FILLER_19_1668 ();
 sg13g2_decap_8 FILLER_19_1675 ();
 sg13g2_decap_8 FILLER_19_1682 ();
 sg13g2_decap_8 FILLER_19_1689 ();
 sg13g2_decap_8 FILLER_19_1696 ();
 sg13g2_decap_8 FILLER_19_1703 ();
 sg13g2_decap_8 FILLER_19_1710 ();
 sg13g2_decap_8 FILLER_19_1717 ();
 sg13g2_decap_8 FILLER_19_1724 ();
 sg13g2_decap_8 FILLER_19_1731 ();
 sg13g2_decap_8 FILLER_19_1738 ();
 sg13g2_decap_8 FILLER_19_1745 ();
 sg13g2_decap_8 FILLER_19_1752 ();
 sg13g2_decap_8 FILLER_19_1759 ();
 sg13g2_fill_2 FILLER_19_1766 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_73 ();
 sg13g2_fill_2 FILLER_20_88 ();
 sg13g2_fill_1 FILLER_20_99 ();
 sg13g2_fill_2 FILLER_20_108 ();
 sg13g2_fill_2 FILLER_20_114 ();
 sg13g2_decap_4 FILLER_20_129 ();
 sg13g2_fill_2 FILLER_20_133 ();
 sg13g2_fill_2 FILLER_20_140 ();
 sg13g2_fill_1 FILLER_20_142 ();
 sg13g2_fill_2 FILLER_20_155 ();
 sg13g2_fill_1 FILLER_20_174 ();
 sg13g2_fill_2 FILLER_20_182 ();
 sg13g2_fill_1 FILLER_20_184 ();
 sg13g2_fill_2 FILLER_20_194 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_fill_1 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_262 ();
 sg13g2_fill_1 FILLER_20_264 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_fill_2 FILLER_20_342 ();
 sg13g2_fill_1 FILLER_20_344 ();
 sg13g2_fill_2 FILLER_20_359 ();
 sg13g2_fill_2 FILLER_20_463 ();
 sg13g2_fill_2 FILLER_20_501 ();
 sg13g2_decap_8 FILLER_20_519 ();
 sg13g2_fill_2 FILLER_20_526 ();
 sg13g2_fill_1 FILLER_20_528 ();
 sg13g2_decap_8 FILLER_20_551 ();
 sg13g2_decap_8 FILLER_20_558 ();
 sg13g2_fill_1 FILLER_20_579 ();
 sg13g2_decap_8 FILLER_20_584 ();
 sg13g2_decap_4 FILLER_20_617 ();
 sg13g2_fill_1 FILLER_20_621 ();
 sg13g2_fill_1 FILLER_20_626 ();
 sg13g2_fill_1 FILLER_20_644 ();
 sg13g2_fill_2 FILLER_20_666 ();
 sg13g2_fill_1 FILLER_20_684 ();
 sg13g2_decap_4 FILLER_20_710 ();
 sg13g2_decap_8 FILLER_20_746 ();
 sg13g2_decap_4 FILLER_20_753 ();
 sg13g2_fill_1 FILLER_20_757 ();
 sg13g2_fill_1 FILLER_20_810 ();
 sg13g2_fill_1 FILLER_20_823 ();
 sg13g2_fill_1 FILLER_20_846 ();
 sg13g2_fill_2 FILLER_20_856 ();
 sg13g2_fill_1 FILLER_20_864 ();
 sg13g2_decap_4 FILLER_20_872 ();
 sg13g2_decap_8 FILLER_20_881 ();
 sg13g2_decap_4 FILLER_20_888 ();
 sg13g2_decap_8 FILLER_20_896 ();
 sg13g2_decap_8 FILLER_20_903 ();
 sg13g2_decap_4 FILLER_20_910 ();
 sg13g2_fill_2 FILLER_20_914 ();
 sg13g2_decap_8 FILLER_20_935 ();
 sg13g2_decap_4 FILLER_20_942 ();
 sg13g2_decap_4 FILLER_20_949 ();
 sg13g2_fill_1 FILLER_20_953 ();
 sg13g2_decap_8 FILLER_20_962 ();
 sg13g2_decap_8 FILLER_20_969 ();
 sg13g2_decap_8 FILLER_20_976 ();
 sg13g2_decap_8 FILLER_20_983 ();
 sg13g2_decap_8 FILLER_20_990 ();
 sg13g2_decap_8 FILLER_20_997 ();
 sg13g2_decap_8 FILLER_20_1004 ();
 sg13g2_decap_8 FILLER_20_1011 ();
 sg13g2_decap_8 FILLER_20_1018 ();
 sg13g2_decap_8 FILLER_20_1025 ();
 sg13g2_decap_8 FILLER_20_1032 ();
 sg13g2_decap_8 FILLER_20_1039 ();
 sg13g2_decap_8 FILLER_20_1046 ();
 sg13g2_decap_8 FILLER_20_1053 ();
 sg13g2_decap_8 FILLER_20_1060 ();
 sg13g2_decap_8 FILLER_20_1067 ();
 sg13g2_decap_8 FILLER_20_1074 ();
 sg13g2_decap_8 FILLER_20_1081 ();
 sg13g2_decap_8 FILLER_20_1088 ();
 sg13g2_decap_8 FILLER_20_1095 ();
 sg13g2_decap_8 FILLER_20_1102 ();
 sg13g2_decap_8 FILLER_20_1109 ();
 sg13g2_decap_8 FILLER_20_1116 ();
 sg13g2_decap_8 FILLER_20_1123 ();
 sg13g2_decap_8 FILLER_20_1130 ();
 sg13g2_decap_8 FILLER_20_1137 ();
 sg13g2_decap_8 FILLER_20_1144 ();
 sg13g2_decap_8 FILLER_20_1151 ();
 sg13g2_decap_8 FILLER_20_1158 ();
 sg13g2_decap_8 FILLER_20_1165 ();
 sg13g2_decap_8 FILLER_20_1172 ();
 sg13g2_decap_8 FILLER_20_1179 ();
 sg13g2_decap_8 FILLER_20_1186 ();
 sg13g2_decap_8 FILLER_20_1193 ();
 sg13g2_decap_8 FILLER_20_1200 ();
 sg13g2_decap_8 FILLER_20_1207 ();
 sg13g2_decap_8 FILLER_20_1214 ();
 sg13g2_decap_8 FILLER_20_1221 ();
 sg13g2_decap_8 FILLER_20_1228 ();
 sg13g2_decap_8 FILLER_20_1235 ();
 sg13g2_decap_8 FILLER_20_1242 ();
 sg13g2_decap_8 FILLER_20_1249 ();
 sg13g2_decap_8 FILLER_20_1256 ();
 sg13g2_decap_8 FILLER_20_1263 ();
 sg13g2_decap_8 FILLER_20_1270 ();
 sg13g2_decap_8 FILLER_20_1277 ();
 sg13g2_decap_8 FILLER_20_1284 ();
 sg13g2_decap_8 FILLER_20_1291 ();
 sg13g2_decap_8 FILLER_20_1298 ();
 sg13g2_decap_8 FILLER_20_1305 ();
 sg13g2_decap_8 FILLER_20_1312 ();
 sg13g2_decap_8 FILLER_20_1319 ();
 sg13g2_decap_8 FILLER_20_1326 ();
 sg13g2_decap_8 FILLER_20_1333 ();
 sg13g2_decap_8 FILLER_20_1340 ();
 sg13g2_decap_8 FILLER_20_1347 ();
 sg13g2_decap_8 FILLER_20_1354 ();
 sg13g2_decap_8 FILLER_20_1361 ();
 sg13g2_decap_8 FILLER_20_1368 ();
 sg13g2_decap_8 FILLER_20_1375 ();
 sg13g2_decap_8 FILLER_20_1382 ();
 sg13g2_decap_8 FILLER_20_1389 ();
 sg13g2_decap_8 FILLER_20_1396 ();
 sg13g2_decap_8 FILLER_20_1403 ();
 sg13g2_decap_8 FILLER_20_1410 ();
 sg13g2_decap_8 FILLER_20_1417 ();
 sg13g2_decap_8 FILLER_20_1424 ();
 sg13g2_decap_8 FILLER_20_1431 ();
 sg13g2_decap_8 FILLER_20_1438 ();
 sg13g2_decap_8 FILLER_20_1445 ();
 sg13g2_decap_8 FILLER_20_1452 ();
 sg13g2_decap_8 FILLER_20_1459 ();
 sg13g2_decap_8 FILLER_20_1466 ();
 sg13g2_decap_8 FILLER_20_1473 ();
 sg13g2_decap_8 FILLER_20_1480 ();
 sg13g2_decap_8 FILLER_20_1487 ();
 sg13g2_decap_8 FILLER_20_1494 ();
 sg13g2_decap_8 FILLER_20_1501 ();
 sg13g2_decap_8 FILLER_20_1508 ();
 sg13g2_decap_8 FILLER_20_1515 ();
 sg13g2_decap_8 FILLER_20_1522 ();
 sg13g2_decap_8 FILLER_20_1529 ();
 sg13g2_decap_8 FILLER_20_1536 ();
 sg13g2_decap_8 FILLER_20_1543 ();
 sg13g2_decap_8 FILLER_20_1550 ();
 sg13g2_decap_8 FILLER_20_1557 ();
 sg13g2_decap_8 FILLER_20_1564 ();
 sg13g2_decap_8 FILLER_20_1571 ();
 sg13g2_decap_8 FILLER_20_1578 ();
 sg13g2_decap_8 FILLER_20_1585 ();
 sg13g2_decap_8 FILLER_20_1592 ();
 sg13g2_decap_8 FILLER_20_1599 ();
 sg13g2_decap_8 FILLER_20_1606 ();
 sg13g2_decap_8 FILLER_20_1613 ();
 sg13g2_decap_8 FILLER_20_1620 ();
 sg13g2_decap_8 FILLER_20_1627 ();
 sg13g2_decap_8 FILLER_20_1634 ();
 sg13g2_decap_8 FILLER_20_1641 ();
 sg13g2_decap_8 FILLER_20_1648 ();
 sg13g2_decap_8 FILLER_20_1655 ();
 sg13g2_decap_8 FILLER_20_1662 ();
 sg13g2_decap_8 FILLER_20_1669 ();
 sg13g2_decap_8 FILLER_20_1676 ();
 sg13g2_decap_8 FILLER_20_1683 ();
 sg13g2_decap_8 FILLER_20_1690 ();
 sg13g2_decap_8 FILLER_20_1697 ();
 sg13g2_decap_8 FILLER_20_1704 ();
 sg13g2_decap_8 FILLER_20_1711 ();
 sg13g2_decap_8 FILLER_20_1718 ();
 sg13g2_decap_8 FILLER_20_1725 ();
 sg13g2_decap_8 FILLER_20_1732 ();
 sg13g2_decap_8 FILLER_20_1739 ();
 sg13g2_decap_8 FILLER_20_1746 ();
 sg13g2_decap_8 FILLER_20_1753 ();
 sg13g2_decap_8 FILLER_20_1760 ();
 sg13g2_fill_1 FILLER_20_1767 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_11 ();
 sg13g2_fill_2 FILLER_21_75 ();
 sg13g2_fill_1 FILLER_21_77 ();
 sg13g2_fill_2 FILLER_21_87 ();
 sg13g2_fill_1 FILLER_21_89 ();
 sg13g2_fill_2 FILLER_21_94 ();
 sg13g2_fill_1 FILLER_21_107 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_4 FILLER_21_153 ();
 sg13g2_decap_8 FILLER_21_193 ();
 sg13g2_decap_4 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_fill_2 FILLER_21_215 ();
 sg13g2_fill_2 FILLER_21_226 ();
 sg13g2_fill_1 FILLER_21_242 ();
 sg13g2_fill_2 FILLER_21_262 ();
 sg13g2_fill_1 FILLER_21_264 ();
 sg13g2_fill_1 FILLER_21_433 ();
 sg13g2_fill_2 FILLER_21_458 ();
 sg13g2_fill_1 FILLER_21_460 ();
 sg13g2_fill_1 FILLER_21_471 ();
 sg13g2_fill_1 FILLER_21_498 ();
 sg13g2_decap_4 FILLER_21_503 ();
 sg13g2_fill_1 FILLER_21_507 ();
 sg13g2_decap_8 FILLER_21_517 ();
 sg13g2_fill_2 FILLER_21_524 ();
 sg13g2_decap_8 FILLER_21_530 ();
 sg13g2_decap_4 FILLER_21_537 ();
 sg13g2_fill_2 FILLER_21_581 ();
 sg13g2_fill_1 FILLER_21_597 ();
 sg13g2_fill_1 FILLER_21_670 ();
 sg13g2_fill_2 FILLER_21_686 ();
 sg13g2_fill_2 FILLER_21_702 ();
 sg13g2_fill_1 FILLER_21_704 ();
 sg13g2_decap_8 FILLER_21_711 ();
 sg13g2_decap_4 FILLER_21_718 ();
 sg13g2_fill_2 FILLER_21_727 ();
 sg13g2_fill_1 FILLER_21_729 ();
 sg13g2_fill_1 FILLER_21_736 ();
 sg13g2_fill_1 FILLER_21_741 ();
 sg13g2_decap_4 FILLER_21_791 ();
 sg13g2_fill_1 FILLER_21_799 ();
 sg13g2_fill_1 FILLER_21_806 ();
 sg13g2_fill_2 FILLER_21_833 ();
 sg13g2_fill_2 FILLER_21_854 ();
 sg13g2_decap_8 FILLER_21_970 ();
 sg13g2_decap_8 FILLER_21_977 ();
 sg13g2_decap_8 FILLER_21_984 ();
 sg13g2_decap_8 FILLER_21_991 ();
 sg13g2_decap_8 FILLER_21_998 ();
 sg13g2_decap_8 FILLER_21_1005 ();
 sg13g2_decap_8 FILLER_21_1012 ();
 sg13g2_decap_8 FILLER_21_1019 ();
 sg13g2_decap_8 FILLER_21_1026 ();
 sg13g2_decap_8 FILLER_21_1033 ();
 sg13g2_decap_8 FILLER_21_1040 ();
 sg13g2_decap_8 FILLER_21_1047 ();
 sg13g2_decap_8 FILLER_21_1054 ();
 sg13g2_decap_8 FILLER_21_1061 ();
 sg13g2_decap_8 FILLER_21_1068 ();
 sg13g2_decap_8 FILLER_21_1075 ();
 sg13g2_decap_8 FILLER_21_1082 ();
 sg13g2_decap_8 FILLER_21_1089 ();
 sg13g2_decap_8 FILLER_21_1096 ();
 sg13g2_decap_8 FILLER_21_1103 ();
 sg13g2_decap_8 FILLER_21_1110 ();
 sg13g2_decap_8 FILLER_21_1117 ();
 sg13g2_decap_8 FILLER_21_1124 ();
 sg13g2_decap_8 FILLER_21_1131 ();
 sg13g2_decap_8 FILLER_21_1138 ();
 sg13g2_decap_8 FILLER_21_1145 ();
 sg13g2_decap_8 FILLER_21_1152 ();
 sg13g2_decap_8 FILLER_21_1159 ();
 sg13g2_decap_8 FILLER_21_1166 ();
 sg13g2_decap_8 FILLER_21_1173 ();
 sg13g2_decap_8 FILLER_21_1180 ();
 sg13g2_decap_8 FILLER_21_1187 ();
 sg13g2_decap_8 FILLER_21_1194 ();
 sg13g2_decap_8 FILLER_21_1201 ();
 sg13g2_decap_8 FILLER_21_1208 ();
 sg13g2_decap_8 FILLER_21_1215 ();
 sg13g2_decap_8 FILLER_21_1222 ();
 sg13g2_decap_8 FILLER_21_1229 ();
 sg13g2_decap_8 FILLER_21_1236 ();
 sg13g2_decap_8 FILLER_21_1243 ();
 sg13g2_decap_8 FILLER_21_1250 ();
 sg13g2_decap_8 FILLER_21_1257 ();
 sg13g2_decap_8 FILLER_21_1264 ();
 sg13g2_decap_8 FILLER_21_1271 ();
 sg13g2_decap_8 FILLER_21_1278 ();
 sg13g2_decap_8 FILLER_21_1285 ();
 sg13g2_decap_8 FILLER_21_1292 ();
 sg13g2_decap_8 FILLER_21_1299 ();
 sg13g2_decap_8 FILLER_21_1306 ();
 sg13g2_decap_8 FILLER_21_1313 ();
 sg13g2_decap_8 FILLER_21_1320 ();
 sg13g2_decap_8 FILLER_21_1327 ();
 sg13g2_decap_8 FILLER_21_1334 ();
 sg13g2_decap_8 FILLER_21_1341 ();
 sg13g2_decap_8 FILLER_21_1348 ();
 sg13g2_decap_8 FILLER_21_1355 ();
 sg13g2_decap_8 FILLER_21_1362 ();
 sg13g2_decap_8 FILLER_21_1369 ();
 sg13g2_decap_8 FILLER_21_1376 ();
 sg13g2_decap_8 FILLER_21_1383 ();
 sg13g2_decap_8 FILLER_21_1390 ();
 sg13g2_decap_8 FILLER_21_1397 ();
 sg13g2_decap_8 FILLER_21_1404 ();
 sg13g2_decap_8 FILLER_21_1411 ();
 sg13g2_decap_8 FILLER_21_1418 ();
 sg13g2_decap_8 FILLER_21_1425 ();
 sg13g2_decap_8 FILLER_21_1432 ();
 sg13g2_decap_8 FILLER_21_1439 ();
 sg13g2_decap_8 FILLER_21_1446 ();
 sg13g2_decap_8 FILLER_21_1453 ();
 sg13g2_decap_8 FILLER_21_1460 ();
 sg13g2_decap_8 FILLER_21_1467 ();
 sg13g2_decap_8 FILLER_21_1474 ();
 sg13g2_decap_8 FILLER_21_1481 ();
 sg13g2_decap_8 FILLER_21_1488 ();
 sg13g2_decap_8 FILLER_21_1495 ();
 sg13g2_decap_8 FILLER_21_1502 ();
 sg13g2_decap_8 FILLER_21_1509 ();
 sg13g2_decap_8 FILLER_21_1516 ();
 sg13g2_decap_8 FILLER_21_1523 ();
 sg13g2_decap_8 FILLER_21_1530 ();
 sg13g2_decap_8 FILLER_21_1537 ();
 sg13g2_decap_8 FILLER_21_1544 ();
 sg13g2_decap_8 FILLER_21_1551 ();
 sg13g2_decap_8 FILLER_21_1558 ();
 sg13g2_decap_8 FILLER_21_1565 ();
 sg13g2_decap_8 FILLER_21_1572 ();
 sg13g2_decap_8 FILLER_21_1579 ();
 sg13g2_decap_8 FILLER_21_1586 ();
 sg13g2_decap_8 FILLER_21_1593 ();
 sg13g2_decap_8 FILLER_21_1600 ();
 sg13g2_decap_8 FILLER_21_1607 ();
 sg13g2_decap_8 FILLER_21_1614 ();
 sg13g2_decap_8 FILLER_21_1621 ();
 sg13g2_decap_8 FILLER_21_1628 ();
 sg13g2_decap_8 FILLER_21_1635 ();
 sg13g2_decap_8 FILLER_21_1642 ();
 sg13g2_decap_8 FILLER_21_1649 ();
 sg13g2_decap_8 FILLER_21_1656 ();
 sg13g2_decap_8 FILLER_21_1663 ();
 sg13g2_decap_8 FILLER_21_1670 ();
 sg13g2_decap_8 FILLER_21_1677 ();
 sg13g2_decap_8 FILLER_21_1684 ();
 sg13g2_decap_8 FILLER_21_1691 ();
 sg13g2_decap_8 FILLER_21_1698 ();
 sg13g2_decap_8 FILLER_21_1705 ();
 sg13g2_decap_8 FILLER_21_1712 ();
 sg13g2_decap_8 FILLER_21_1719 ();
 sg13g2_decap_8 FILLER_21_1726 ();
 sg13g2_decap_8 FILLER_21_1733 ();
 sg13g2_decap_8 FILLER_21_1740 ();
 sg13g2_decap_8 FILLER_21_1747 ();
 sg13g2_decap_8 FILLER_21_1754 ();
 sg13g2_decap_8 FILLER_21_1761 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_11 ();
 sg13g2_fill_2 FILLER_22_33 ();
 sg13g2_fill_1 FILLER_22_54 ();
 sg13g2_fill_2 FILLER_22_69 ();
 sg13g2_fill_1 FILLER_22_80 ();
 sg13g2_fill_2 FILLER_22_86 ();
 sg13g2_decap_8 FILLER_22_118 ();
 sg13g2_fill_2 FILLER_22_125 ();
 sg13g2_fill_1 FILLER_22_127 ();
 sg13g2_fill_1 FILLER_22_137 ();
 sg13g2_decap_8 FILLER_22_151 ();
 sg13g2_decap_4 FILLER_22_158 ();
 sg13g2_fill_1 FILLER_22_169 ();
 sg13g2_fill_2 FILLER_22_191 ();
 sg13g2_fill_2 FILLER_22_205 ();
 sg13g2_fill_2 FILLER_22_223 ();
 sg13g2_fill_2 FILLER_22_251 ();
 sg13g2_fill_1 FILLER_22_253 ();
 sg13g2_fill_2 FILLER_22_310 ();
 sg13g2_fill_1 FILLER_22_312 ();
 sg13g2_fill_2 FILLER_22_361 ();
 sg13g2_fill_2 FILLER_22_367 ();
 sg13g2_fill_1 FILLER_22_416 ();
 sg13g2_fill_1 FILLER_22_465 ();
 sg13g2_fill_1 FILLER_22_546 ();
 sg13g2_fill_1 FILLER_22_564 ();
 sg13g2_fill_1 FILLER_22_570 ();
 sg13g2_fill_2 FILLER_22_601 ();
 sg13g2_fill_1 FILLER_22_603 ();
 sg13g2_fill_1 FILLER_22_636 ();
 sg13g2_fill_2 FILLER_22_692 ();
 sg13g2_fill_1 FILLER_22_694 ();
 sg13g2_fill_2 FILLER_22_703 ();
 sg13g2_fill_1 FILLER_22_705 ();
 sg13g2_fill_1 FILLER_22_732 ();
 sg13g2_decap_4 FILLER_22_793 ();
 sg13g2_fill_1 FILLER_22_797 ();
 sg13g2_decap_8 FILLER_22_808 ();
 sg13g2_fill_2 FILLER_22_815 ();
 sg13g2_fill_1 FILLER_22_817 ();
 sg13g2_fill_2 FILLER_22_828 ();
 sg13g2_fill_1 FILLER_22_830 ();
 sg13g2_decap_4 FILLER_22_854 ();
 sg13g2_fill_2 FILLER_22_858 ();
 sg13g2_decap_8 FILLER_22_872 ();
 sg13g2_fill_1 FILLER_22_879 ();
 sg13g2_fill_2 FILLER_22_890 ();
 sg13g2_fill_1 FILLER_22_892 ();
 sg13g2_decap_4 FILLER_22_913 ();
 sg13g2_fill_2 FILLER_22_926 ();
 sg13g2_decap_8 FILLER_22_939 ();
 sg13g2_fill_1 FILLER_22_946 ();
 sg13g2_decap_4 FILLER_22_970 ();
 sg13g2_decap_8 FILLER_22_978 ();
 sg13g2_decap_8 FILLER_22_985 ();
 sg13g2_decap_8 FILLER_22_992 ();
 sg13g2_decap_8 FILLER_22_999 ();
 sg13g2_decap_8 FILLER_22_1006 ();
 sg13g2_decap_8 FILLER_22_1013 ();
 sg13g2_decap_8 FILLER_22_1020 ();
 sg13g2_decap_8 FILLER_22_1027 ();
 sg13g2_decap_8 FILLER_22_1034 ();
 sg13g2_decap_8 FILLER_22_1041 ();
 sg13g2_decap_8 FILLER_22_1048 ();
 sg13g2_decap_8 FILLER_22_1055 ();
 sg13g2_decap_8 FILLER_22_1062 ();
 sg13g2_decap_8 FILLER_22_1069 ();
 sg13g2_decap_8 FILLER_22_1076 ();
 sg13g2_decap_8 FILLER_22_1083 ();
 sg13g2_decap_8 FILLER_22_1090 ();
 sg13g2_decap_8 FILLER_22_1097 ();
 sg13g2_decap_8 FILLER_22_1104 ();
 sg13g2_decap_8 FILLER_22_1111 ();
 sg13g2_decap_8 FILLER_22_1118 ();
 sg13g2_decap_8 FILLER_22_1125 ();
 sg13g2_decap_8 FILLER_22_1132 ();
 sg13g2_decap_8 FILLER_22_1139 ();
 sg13g2_decap_8 FILLER_22_1146 ();
 sg13g2_decap_8 FILLER_22_1153 ();
 sg13g2_decap_8 FILLER_22_1160 ();
 sg13g2_decap_8 FILLER_22_1167 ();
 sg13g2_decap_8 FILLER_22_1174 ();
 sg13g2_decap_8 FILLER_22_1181 ();
 sg13g2_decap_8 FILLER_22_1188 ();
 sg13g2_decap_8 FILLER_22_1195 ();
 sg13g2_decap_8 FILLER_22_1202 ();
 sg13g2_decap_8 FILLER_22_1209 ();
 sg13g2_decap_8 FILLER_22_1216 ();
 sg13g2_decap_8 FILLER_22_1223 ();
 sg13g2_decap_8 FILLER_22_1230 ();
 sg13g2_decap_8 FILLER_22_1237 ();
 sg13g2_decap_8 FILLER_22_1244 ();
 sg13g2_decap_8 FILLER_22_1251 ();
 sg13g2_decap_8 FILLER_22_1258 ();
 sg13g2_decap_8 FILLER_22_1265 ();
 sg13g2_decap_8 FILLER_22_1272 ();
 sg13g2_decap_8 FILLER_22_1279 ();
 sg13g2_decap_8 FILLER_22_1286 ();
 sg13g2_decap_8 FILLER_22_1293 ();
 sg13g2_decap_8 FILLER_22_1300 ();
 sg13g2_decap_8 FILLER_22_1307 ();
 sg13g2_decap_8 FILLER_22_1314 ();
 sg13g2_decap_8 FILLER_22_1321 ();
 sg13g2_decap_8 FILLER_22_1328 ();
 sg13g2_decap_8 FILLER_22_1335 ();
 sg13g2_decap_8 FILLER_22_1342 ();
 sg13g2_decap_8 FILLER_22_1349 ();
 sg13g2_decap_8 FILLER_22_1356 ();
 sg13g2_decap_8 FILLER_22_1363 ();
 sg13g2_decap_8 FILLER_22_1370 ();
 sg13g2_decap_8 FILLER_22_1377 ();
 sg13g2_decap_8 FILLER_22_1384 ();
 sg13g2_decap_8 FILLER_22_1391 ();
 sg13g2_decap_8 FILLER_22_1398 ();
 sg13g2_decap_8 FILLER_22_1405 ();
 sg13g2_decap_8 FILLER_22_1412 ();
 sg13g2_decap_8 FILLER_22_1419 ();
 sg13g2_decap_8 FILLER_22_1426 ();
 sg13g2_decap_8 FILLER_22_1433 ();
 sg13g2_decap_8 FILLER_22_1440 ();
 sg13g2_decap_8 FILLER_22_1447 ();
 sg13g2_decap_8 FILLER_22_1454 ();
 sg13g2_decap_8 FILLER_22_1461 ();
 sg13g2_decap_8 FILLER_22_1468 ();
 sg13g2_decap_8 FILLER_22_1475 ();
 sg13g2_decap_8 FILLER_22_1482 ();
 sg13g2_decap_8 FILLER_22_1489 ();
 sg13g2_decap_8 FILLER_22_1496 ();
 sg13g2_decap_8 FILLER_22_1503 ();
 sg13g2_decap_8 FILLER_22_1510 ();
 sg13g2_decap_8 FILLER_22_1517 ();
 sg13g2_decap_8 FILLER_22_1524 ();
 sg13g2_decap_8 FILLER_22_1531 ();
 sg13g2_decap_8 FILLER_22_1538 ();
 sg13g2_decap_8 FILLER_22_1545 ();
 sg13g2_decap_8 FILLER_22_1552 ();
 sg13g2_decap_8 FILLER_22_1559 ();
 sg13g2_decap_8 FILLER_22_1566 ();
 sg13g2_decap_8 FILLER_22_1573 ();
 sg13g2_decap_8 FILLER_22_1580 ();
 sg13g2_decap_8 FILLER_22_1587 ();
 sg13g2_decap_8 FILLER_22_1594 ();
 sg13g2_decap_8 FILLER_22_1601 ();
 sg13g2_decap_8 FILLER_22_1608 ();
 sg13g2_decap_8 FILLER_22_1615 ();
 sg13g2_decap_8 FILLER_22_1622 ();
 sg13g2_decap_8 FILLER_22_1629 ();
 sg13g2_decap_8 FILLER_22_1636 ();
 sg13g2_decap_8 FILLER_22_1643 ();
 sg13g2_decap_8 FILLER_22_1650 ();
 sg13g2_decap_8 FILLER_22_1657 ();
 sg13g2_decap_8 FILLER_22_1664 ();
 sg13g2_decap_8 FILLER_22_1671 ();
 sg13g2_decap_8 FILLER_22_1678 ();
 sg13g2_decap_8 FILLER_22_1685 ();
 sg13g2_decap_8 FILLER_22_1692 ();
 sg13g2_decap_8 FILLER_22_1699 ();
 sg13g2_decap_8 FILLER_22_1706 ();
 sg13g2_decap_8 FILLER_22_1713 ();
 sg13g2_decap_8 FILLER_22_1720 ();
 sg13g2_decap_8 FILLER_22_1727 ();
 sg13g2_decap_8 FILLER_22_1734 ();
 sg13g2_decap_8 FILLER_22_1741 ();
 sg13g2_decap_8 FILLER_22_1748 ();
 sg13g2_decap_8 FILLER_22_1755 ();
 sg13g2_decap_4 FILLER_22_1762 ();
 sg13g2_fill_2 FILLER_22_1766 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_43 ();
 sg13g2_fill_2 FILLER_23_77 ();
 sg13g2_fill_1 FILLER_23_79 ();
 sg13g2_fill_1 FILLER_23_90 ();
 sg13g2_decap_4 FILLER_23_96 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_4 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_fill_2 FILLER_23_127 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_fill_2 FILLER_23_148 ();
 sg13g2_fill_2 FILLER_23_162 ();
 sg13g2_fill_1 FILLER_23_164 ();
 sg13g2_fill_2 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_181 ();
 sg13g2_fill_2 FILLER_23_213 ();
 sg13g2_fill_1 FILLER_23_215 ();
 sg13g2_fill_2 FILLER_23_230 ();
 sg13g2_fill_1 FILLER_23_232 ();
 sg13g2_fill_2 FILLER_23_238 ();
 sg13g2_fill_1 FILLER_23_249 ();
 sg13g2_fill_1 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_409 ();
 sg13g2_fill_1 FILLER_23_411 ();
 sg13g2_fill_1 FILLER_23_459 ();
 sg13g2_fill_1 FILLER_23_481 ();
 sg13g2_decap_4 FILLER_23_513 ();
 sg13g2_fill_1 FILLER_23_517 ();
 sg13g2_fill_1 FILLER_23_523 ();
 sg13g2_decap_4 FILLER_23_528 ();
 sg13g2_fill_2 FILLER_23_572 ();
 sg13g2_fill_1 FILLER_23_583 ();
 sg13g2_fill_2 FILLER_23_620 ();
 sg13g2_fill_1 FILLER_23_622 ();
 sg13g2_fill_2 FILLER_23_653 ();
 sg13g2_fill_1 FILLER_23_655 ();
 sg13g2_fill_2 FILLER_23_670 ();
 sg13g2_decap_4 FILLER_23_681 ();
 sg13g2_decap_8 FILLER_23_695 ();
 sg13g2_decap_8 FILLER_23_702 ();
 sg13g2_decap_8 FILLER_23_709 ();
 sg13g2_fill_1 FILLER_23_716 ();
 sg13g2_fill_2 FILLER_23_721 ();
 sg13g2_fill_2 FILLER_23_741 ();
 sg13g2_fill_1 FILLER_23_755 ();
 sg13g2_decap_4 FILLER_23_786 ();
 sg13g2_fill_1 FILLER_23_790 ();
 sg13g2_fill_2 FILLER_23_828 ();
 sg13g2_decap_4 FILLER_23_848 ();
 sg13g2_fill_2 FILLER_23_852 ();
 sg13g2_fill_2 FILLER_23_872 ();
 sg13g2_fill_1 FILLER_23_874 ();
 sg13g2_decap_8 FILLER_23_883 ();
 sg13g2_fill_2 FILLER_23_890 ();
 sg13g2_fill_1 FILLER_23_892 ();
 sg13g2_decap_8 FILLER_23_897 ();
 sg13g2_decap_4 FILLER_23_904 ();
 sg13g2_fill_1 FILLER_23_908 ();
 sg13g2_fill_1 FILLER_23_935 ();
 sg13g2_fill_2 FILLER_23_948 ();
 sg13g2_decap_4 FILLER_23_963 ();
 sg13g2_decap_8 FILLER_23_989 ();
 sg13g2_decap_8 FILLER_23_996 ();
 sg13g2_decap_8 FILLER_23_1003 ();
 sg13g2_decap_8 FILLER_23_1010 ();
 sg13g2_decap_8 FILLER_23_1017 ();
 sg13g2_decap_8 FILLER_23_1024 ();
 sg13g2_decap_8 FILLER_23_1031 ();
 sg13g2_decap_8 FILLER_23_1038 ();
 sg13g2_decap_8 FILLER_23_1045 ();
 sg13g2_decap_8 FILLER_23_1052 ();
 sg13g2_decap_8 FILLER_23_1059 ();
 sg13g2_decap_8 FILLER_23_1066 ();
 sg13g2_decap_8 FILLER_23_1073 ();
 sg13g2_decap_8 FILLER_23_1080 ();
 sg13g2_decap_8 FILLER_23_1087 ();
 sg13g2_decap_8 FILLER_23_1094 ();
 sg13g2_decap_8 FILLER_23_1101 ();
 sg13g2_decap_8 FILLER_23_1108 ();
 sg13g2_decap_8 FILLER_23_1115 ();
 sg13g2_decap_8 FILLER_23_1122 ();
 sg13g2_decap_8 FILLER_23_1129 ();
 sg13g2_decap_8 FILLER_23_1136 ();
 sg13g2_decap_8 FILLER_23_1143 ();
 sg13g2_decap_8 FILLER_23_1150 ();
 sg13g2_decap_8 FILLER_23_1157 ();
 sg13g2_decap_8 FILLER_23_1164 ();
 sg13g2_decap_8 FILLER_23_1171 ();
 sg13g2_decap_8 FILLER_23_1178 ();
 sg13g2_decap_8 FILLER_23_1185 ();
 sg13g2_decap_8 FILLER_23_1192 ();
 sg13g2_decap_8 FILLER_23_1199 ();
 sg13g2_decap_8 FILLER_23_1206 ();
 sg13g2_decap_8 FILLER_23_1213 ();
 sg13g2_decap_8 FILLER_23_1220 ();
 sg13g2_decap_8 FILLER_23_1227 ();
 sg13g2_decap_8 FILLER_23_1234 ();
 sg13g2_decap_8 FILLER_23_1241 ();
 sg13g2_decap_8 FILLER_23_1248 ();
 sg13g2_decap_8 FILLER_23_1255 ();
 sg13g2_decap_8 FILLER_23_1262 ();
 sg13g2_decap_8 FILLER_23_1269 ();
 sg13g2_decap_8 FILLER_23_1276 ();
 sg13g2_decap_8 FILLER_23_1283 ();
 sg13g2_decap_8 FILLER_23_1290 ();
 sg13g2_decap_8 FILLER_23_1297 ();
 sg13g2_decap_8 FILLER_23_1304 ();
 sg13g2_decap_8 FILLER_23_1311 ();
 sg13g2_decap_8 FILLER_23_1318 ();
 sg13g2_decap_8 FILLER_23_1325 ();
 sg13g2_decap_8 FILLER_23_1332 ();
 sg13g2_decap_8 FILLER_23_1339 ();
 sg13g2_decap_8 FILLER_23_1346 ();
 sg13g2_decap_8 FILLER_23_1353 ();
 sg13g2_decap_8 FILLER_23_1360 ();
 sg13g2_decap_8 FILLER_23_1367 ();
 sg13g2_decap_8 FILLER_23_1374 ();
 sg13g2_decap_8 FILLER_23_1381 ();
 sg13g2_decap_8 FILLER_23_1388 ();
 sg13g2_decap_8 FILLER_23_1395 ();
 sg13g2_decap_8 FILLER_23_1402 ();
 sg13g2_decap_8 FILLER_23_1409 ();
 sg13g2_decap_8 FILLER_23_1416 ();
 sg13g2_decap_8 FILLER_23_1423 ();
 sg13g2_decap_8 FILLER_23_1430 ();
 sg13g2_decap_8 FILLER_23_1437 ();
 sg13g2_decap_8 FILLER_23_1444 ();
 sg13g2_decap_8 FILLER_23_1451 ();
 sg13g2_decap_8 FILLER_23_1458 ();
 sg13g2_decap_8 FILLER_23_1465 ();
 sg13g2_decap_8 FILLER_23_1472 ();
 sg13g2_decap_8 FILLER_23_1479 ();
 sg13g2_decap_8 FILLER_23_1486 ();
 sg13g2_decap_8 FILLER_23_1493 ();
 sg13g2_decap_8 FILLER_23_1500 ();
 sg13g2_decap_8 FILLER_23_1507 ();
 sg13g2_decap_8 FILLER_23_1514 ();
 sg13g2_decap_8 FILLER_23_1521 ();
 sg13g2_decap_8 FILLER_23_1528 ();
 sg13g2_decap_8 FILLER_23_1535 ();
 sg13g2_decap_8 FILLER_23_1542 ();
 sg13g2_decap_8 FILLER_23_1549 ();
 sg13g2_decap_8 FILLER_23_1556 ();
 sg13g2_decap_8 FILLER_23_1563 ();
 sg13g2_decap_8 FILLER_23_1570 ();
 sg13g2_decap_8 FILLER_23_1577 ();
 sg13g2_decap_8 FILLER_23_1584 ();
 sg13g2_decap_8 FILLER_23_1591 ();
 sg13g2_decap_8 FILLER_23_1598 ();
 sg13g2_decap_8 FILLER_23_1605 ();
 sg13g2_decap_8 FILLER_23_1612 ();
 sg13g2_decap_8 FILLER_23_1619 ();
 sg13g2_decap_8 FILLER_23_1626 ();
 sg13g2_decap_8 FILLER_23_1633 ();
 sg13g2_decap_8 FILLER_23_1640 ();
 sg13g2_decap_8 FILLER_23_1647 ();
 sg13g2_decap_8 FILLER_23_1654 ();
 sg13g2_decap_8 FILLER_23_1661 ();
 sg13g2_decap_8 FILLER_23_1668 ();
 sg13g2_decap_8 FILLER_23_1675 ();
 sg13g2_decap_8 FILLER_23_1682 ();
 sg13g2_decap_8 FILLER_23_1689 ();
 sg13g2_decap_8 FILLER_23_1696 ();
 sg13g2_decap_8 FILLER_23_1703 ();
 sg13g2_decap_8 FILLER_23_1710 ();
 sg13g2_decap_8 FILLER_23_1717 ();
 sg13g2_decap_8 FILLER_23_1724 ();
 sg13g2_decap_8 FILLER_23_1731 ();
 sg13g2_decap_8 FILLER_23_1738 ();
 sg13g2_decap_8 FILLER_23_1745 ();
 sg13g2_decap_8 FILLER_23_1752 ();
 sg13g2_decap_8 FILLER_23_1759 ();
 sg13g2_fill_2 FILLER_23_1766 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_18 ();
 sg13g2_decap_8 FILLER_24_64 ();
 sg13g2_fill_2 FILLER_24_97 ();
 sg13g2_decap_8 FILLER_24_110 ();
 sg13g2_decap_4 FILLER_24_141 ();
 sg13g2_fill_2 FILLER_24_145 ();
 sg13g2_decap_4 FILLER_24_152 ();
 sg13g2_fill_1 FILLER_24_156 ();
 sg13g2_fill_2 FILLER_24_167 ();
 sg13g2_decap_4 FILLER_24_173 ();
 sg13g2_fill_1 FILLER_24_177 ();
 sg13g2_decap_4 FILLER_24_187 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_fill_2 FILLER_24_235 ();
 sg13g2_fill_2 FILLER_24_277 ();
 sg13g2_fill_2 FILLER_24_318 ();
 sg13g2_fill_1 FILLER_24_320 ();
 sg13g2_fill_2 FILLER_24_330 ();
 sg13g2_fill_1 FILLER_24_332 ();
 sg13g2_fill_1 FILLER_24_343 ();
 sg13g2_fill_2 FILLER_24_358 ();
 sg13g2_fill_2 FILLER_24_416 ();
 sg13g2_fill_2 FILLER_24_481 ();
 sg13g2_fill_2 FILLER_24_488 ();
 sg13g2_fill_1 FILLER_24_495 ();
 sg13g2_fill_1 FILLER_24_512 ();
 sg13g2_fill_2 FILLER_24_585 ();
 sg13g2_fill_1 FILLER_24_587 ();
 sg13g2_decap_8 FILLER_24_625 ();
 sg13g2_fill_2 FILLER_24_636 ();
 sg13g2_decap_4 FILLER_24_642 ();
 sg13g2_fill_1 FILLER_24_646 ();
 sg13g2_fill_1 FILLER_24_652 ();
 sg13g2_decap_8 FILLER_24_661 ();
 sg13g2_decap_8 FILLER_24_676 ();
 sg13g2_decap_8 FILLER_24_693 ();
 sg13g2_fill_2 FILLER_24_700 ();
 sg13g2_fill_1 FILLER_24_711 ();
 sg13g2_decap_8 FILLER_24_716 ();
 sg13g2_fill_2 FILLER_24_755 ();
 sg13g2_fill_1 FILLER_24_757 ();
 sg13g2_fill_1 FILLER_24_761 ();
 sg13g2_fill_1 FILLER_24_766 ();
 sg13g2_decap_8 FILLER_24_780 ();
 sg13g2_fill_2 FILLER_24_787 ();
 sg13g2_fill_1 FILLER_24_789 ();
 sg13g2_decap_4 FILLER_24_808 ();
 sg13g2_fill_1 FILLER_24_812 ();
 sg13g2_decap_4 FILLER_24_826 ();
 sg13g2_fill_2 FILLER_24_830 ();
 sg13g2_decap_4 FILLER_24_860 ();
 sg13g2_decap_4 FILLER_24_891 ();
 sg13g2_fill_2 FILLER_24_895 ();
 sg13g2_decap_4 FILLER_24_918 ();
 sg13g2_fill_2 FILLER_24_930 ();
 sg13g2_fill_2 FILLER_24_940 ();
 sg13g2_fill_1 FILLER_24_942 ();
 sg13g2_fill_2 FILLER_24_951 ();
 sg13g2_fill_1 FILLER_24_953 ();
 sg13g2_fill_2 FILLER_24_965 ();
 sg13g2_fill_1 FILLER_24_967 ();
 sg13g2_decap_8 FILLER_24_997 ();
 sg13g2_decap_8 FILLER_24_1004 ();
 sg13g2_decap_8 FILLER_24_1011 ();
 sg13g2_decap_8 FILLER_24_1018 ();
 sg13g2_decap_8 FILLER_24_1025 ();
 sg13g2_decap_8 FILLER_24_1032 ();
 sg13g2_decap_8 FILLER_24_1039 ();
 sg13g2_decap_8 FILLER_24_1046 ();
 sg13g2_decap_8 FILLER_24_1053 ();
 sg13g2_decap_8 FILLER_24_1060 ();
 sg13g2_decap_8 FILLER_24_1067 ();
 sg13g2_decap_8 FILLER_24_1074 ();
 sg13g2_decap_8 FILLER_24_1081 ();
 sg13g2_decap_8 FILLER_24_1088 ();
 sg13g2_decap_8 FILLER_24_1095 ();
 sg13g2_decap_8 FILLER_24_1102 ();
 sg13g2_decap_8 FILLER_24_1109 ();
 sg13g2_decap_8 FILLER_24_1116 ();
 sg13g2_decap_8 FILLER_24_1123 ();
 sg13g2_decap_8 FILLER_24_1130 ();
 sg13g2_decap_8 FILLER_24_1137 ();
 sg13g2_decap_8 FILLER_24_1144 ();
 sg13g2_decap_8 FILLER_24_1151 ();
 sg13g2_decap_8 FILLER_24_1158 ();
 sg13g2_decap_8 FILLER_24_1165 ();
 sg13g2_decap_8 FILLER_24_1172 ();
 sg13g2_decap_8 FILLER_24_1179 ();
 sg13g2_decap_8 FILLER_24_1186 ();
 sg13g2_decap_8 FILLER_24_1193 ();
 sg13g2_decap_8 FILLER_24_1200 ();
 sg13g2_decap_8 FILLER_24_1207 ();
 sg13g2_decap_8 FILLER_24_1214 ();
 sg13g2_decap_8 FILLER_24_1221 ();
 sg13g2_decap_8 FILLER_24_1228 ();
 sg13g2_decap_8 FILLER_24_1235 ();
 sg13g2_decap_8 FILLER_24_1242 ();
 sg13g2_decap_8 FILLER_24_1249 ();
 sg13g2_decap_8 FILLER_24_1256 ();
 sg13g2_decap_8 FILLER_24_1263 ();
 sg13g2_decap_8 FILLER_24_1270 ();
 sg13g2_decap_8 FILLER_24_1277 ();
 sg13g2_decap_8 FILLER_24_1284 ();
 sg13g2_decap_8 FILLER_24_1291 ();
 sg13g2_decap_8 FILLER_24_1298 ();
 sg13g2_decap_8 FILLER_24_1305 ();
 sg13g2_decap_8 FILLER_24_1312 ();
 sg13g2_decap_8 FILLER_24_1319 ();
 sg13g2_decap_8 FILLER_24_1326 ();
 sg13g2_decap_8 FILLER_24_1333 ();
 sg13g2_decap_8 FILLER_24_1340 ();
 sg13g2_decap_8 FILLER_24_1347 ();
 sg13g2_decap_8 FILLER_24_1354 ();
 sg13g2_decap_8 FILLER_24_1361 ();
 sg13g2_decap_8 FILLER_24_1368 ();
 sg13g2_decap_8 FILLER_24_1375 ();
 sg13g2_decap_8 FILLER_24_1382 ();
 sg13g2_decap_8 FILLER_24_1389 ();
 sg13g2_decap_8 FILLER_24_1396 ();
 sg13g2_decap_8 FILLER_24_1403 ();
 sg13g2_decap_8 FILLER_24_1410 ();
 sg13g2_decap_8 FILLER_24_1417 ();
 sg13g2_decap_8 FILLER_24_1424 ();
 sg13g2_decap_8 FILLER_24_1431 ();
 sg13g2_decap_8 FILLER_24_1438 ();
 sg13g2_decap_8 FILLER_24_1445 ();
 sg13g2_decap_8 FILLER_24_1452 ();
 sg13g2_decap_8 FILLER_24_1459 ();
 sg13g2_decap_8 FILLER_24_1466 ();
 sg13g2_decap_8 FILLER_24_1473 ();
 sg13g2_decap_8 FILLER_24_1480 ();
 sg13g2_decap_8 FILLER_24_1487 ();
 sg13g2_decap_8 FILLER_24_1494 ();
 sg13g2_decap_8 FILLER_24_1501 ();
 sg13g2_decap_8 FILLER_24_1508 ();
 sg13g2_decap_8 FILLER_24_1515 ();
 sg13g2_decap_8 FILLER_24_1522 ();
 sg13g2_decap_8 FILLER_24_1529 ();
 sg13g2_decap_8 FILLER_24_1536 ();
 sg13g2_decap_8 FILLER_24_1543 ();
 sg13g2_decap_8 FILLER_24_1550 ();
 sg13g2_decap_8 FILLER_24_1557 ();
 sg13g2_decap_8 FILLER_24_1564 ();
 sg13g2_decap_8 FILLER_24_1571 ();
 sg13g2_decap_8 FILLER_24_1578 ();
 sg13g2_decap_8 FILLER_24_1585 ();
 sg13g2_decap_8 FILLER_24_1592 ();
 sg13g2_decap_8 FILLER_24_1599 ();
 sg13g2_decap_8 FILLER_24_1606 ();
 sg13g2_decap_8 FILLER_24_1613 ();
 sg13g2_decap_8 FILLER_24_1620 ();
 sg13g2_decap_8 FILLER_24_1627 ();
 sg13g2_decap_8 FILLER_24_1634 ();
 sg13g2_decap_8 FILLER_24_1641 ();
 sg13g2_decap_8 FILLER_24_1648 ();
 sg13g2_decap_8 FILLER_24_1655 ();
 sg13g2_decap_8 FILLER_24_1662 ();
 sg13g2_decap_8 FILLER_24_1669 ();
 sg13g2_decap_8 FILLER_24_1676 ();
 sg13g2_decap_8 FILLER_24_1683 ();
 sg13g2_decap_8 FILLER_24_1690 ();
 sg13g2_decap_8 FILLER_24_1697 ();
 sg13g2_decap_8 FILLER_24_1704 ();
 sg13g2_decap_8 FILLER_24_1711 ();
 sg13g2_decap_8 FILLER_24_1718 ();
 sg13g2_decap_8 FILLER_24_1725 ();
 sg13g2_decap_8 FILLER_24_1732 ();
 sg13g2_decap_8 FILLER_24_1739 ();
 sg13g2_decap_8 FILLER_24_1746 ();
 sg13g2_decap_8 FILLER_24_1753 ();
 sg13g2_decap_8 FILLER_24_1760 ();
 sg13g2_fill_1 FILLER_24_1767 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_fill_2 FILLER_25_131 ();
 sg13g2_fill_2 FILLER_25_166 ();
 sg13g2_fill_2 FILLER_25_189 ();
 sg13g2_fill_1 FILLER_25_191 ();
 sg13g2_decap_8 FILLER_25_207 ();
 sg13g2_decap_4 FILLER_25_214 ();
 sg13g2_fill_1 FILLER_25_218 ();
 sg13g2_decap_4 FILLER_25_223 ();
 sg13g2_fill_2 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_394 ();
 sg13g2_fill_1 FILLER_25_396 ();
 sg13g2_fill_2 FILLER_25_475 ();
 sg13g2_fill_1 FILLER_25_477 ();
 sg13g2_fill_2 FILLER_25_504 ();
 sg13g2_fill_2 FILLER_25_547 ();
 sg13g2_fill_1 FILLER_25_573 ();
 sg13g2_fill_2 FILLER_25_583 ();
 sg13g2_decap_4 FILLER_25_589 ();
 sg13g2_fill_1 FILLER_25_593 ();
 sg13g2_decap_4 FILLER_25_618 ();
 sg13g2_fill_2 FILLER_25_630 ();
 sg13g2_fill_1 FILLER_25_661 ();
 sg13g2_decap_8 FILLER_25_691 ();
 sg13g2_fill_2 FILLER_25_698 ();
 sg13g2_fill_1 FILLER_25_700 ();
 sg13g2_decap_4 FILLER_25_736 ();
 sg13g2_fill_2 FILLER_25_744 ();
 sg13g2_fill_1 FILLER_25_746 ();
 sg13g2_fill_2 FILLER_25_819 ();
 sg13g2_fill_1 FILLER_25_841 ();
 sg13g2_fill_2 FILLER_25_853 ();
 sg13g2_fill_1 FILLER_25_855 ();
 sg13g2_fill_1 FILLER_25_871 ();
 sg13g2_fill_2 FILLER_25_890 ();
 sg13g2_fill_1 FILLER_25_892 ();
 sg13g2_fill_1 FILLER_25_904 ();
 sg13g2_fill_2 FILLER_25_918 ();
 sg13g2_fill_1 FILLER_25_920 ();
 sg13g2_decap_8 FILLER_25_940 ();
 sg13g2_decap_4 FILLER_25_947 ();
 sg13g2_fill_2 FILLER_25_951 ();
 sg13g2_decap_8 FILLER_25_961 ();
 sg13g2_decap_8 FILLER_25_968 ();
 sg13g2_fill_2 FILLER_25_975 ();
 sg13g2_fill_1 FILLER_25_977 ();
 sg13g2_decap_8 FILLER_25_986 ();
 sg13g2_decap_8 FILLER_25_993 ();
 sg13g2_decap_8 FILLER_25_1000 ();
 sg13g2_decap_8 FILLER_25_1007 ();
 sg13g2_decap_8 FILLER_25_1014 ();
 sg13g2_decap_8 FILLER_25_1021 ();
 sg13g2_decap_8 FILLER_25_1028 ();
 sg13g2_decap_8 FILLER_25_1035 ();
 sg13g2_decap_8 FILLER_25_1042 ();
 sg13g2_decap_8 FILLER_25_1049 ();
 sg13g2_decap_8 FILLER_25_1056 ();
 sg13g2_decap_8 FILLER_25_1063 ();
 sg13g2_decap_8 FILLER_25_1070 ();
 sg13g2_decap_8 FILLER_25_1077 ();
 sg13g2_decap_8 FILLER_25_1084 ();
 sg13g2_decap_8 FILLER_25_1091 ();
 sg13g2_decap_8 FILLER_25_1098 ();
 sg13g2_decap_8 FILLER_25_1105 ();
 sg13g2_decap_8 FILLER_25_1112 ();
 sg13g2_decap_8 FILLER_25_1119 ();
 sg13g2_decap_8 FILLER_25_1126 ();
 sg13g2_decap_8 FILLER_25_1133 ();
 sg13g2_decap_8 FILLER_25_1140 ();
 sg13g2_decap_8 FILLER_25_1147 ();
 sg13g2_decap_8 FILLER_25_1154 ();
 sg13g2_decap_8 FILLER_25_1161 ();
 sg13g2_decap_8 FILLER_25_1168 ();
 sg13g2_decap_8 FILLER_25_1175 ();
 sg13g2_decap_8 FILLER_25_1182 ();
 sg13g2_decap_8 FILLER_25_1189 ();
 sg13g2_decap_8 FILLER_25_1196 ();
 sg13g2_decap_8 FILLER_25_1203 ();
 sg13g2_decap_8 FILLER_25_1210 ();
 sg13g2_decap_8 FILLER_25_1217 ();
 sg13g2_decap_8 FILLER_25_1224 ();
 sg13g2_decap_8 FILLER_25_1231 ();
 sg13g2_decap_8 FILLER_25_1238 ();
 sg13g2_decap_8 FILLER_25_1245 ();
 sg13g2_decap_8 FILLER_25_1252 ();
 sg13g2_decap_8 FILLER_25_1259 ();
 sg13g2_decap_8 FILLER_25_1266 ();
 sg13g2_decap_8 FILLER_25_1273 ();
 sg13g2_decap_8 FILLER_25_1280 ();
 sg13g2_decap_8 FILLER_25_1287 ();
 sg13g2_decap_8 FILLER_25_1294 ();
 sg13g2_decap_8 FILLER_25_1301 ();
 sg13g2_decap_8 FILLER_25_1308 ();
 sg13g2_decap_8 FILLER_25_1315 ();
 sg13g2_decap_8 FILLER_25_1322 ();
 sg13g2_decap_8 FILLER_25_1329 ();
 sg13g2_decap_8 FILLER_25_1336 ();
 sg13g2_decap_8 FILLER_25_1343 ();
 sg13g2_decap_8 FILLER_25_1350 ();
 sg13g2_decap_8 FILLER_25_1357 ();
 sg13g2_decap_8 FILLER_25_1364 ();
 sg13g2_decap_8 FILLER_25_1371 ();
 sg13g2_decap_8 FILLER_25_1378 ();
 sg13g2_decap_8 FILLER_25_1385 ();
 sg13g2_decap_8 FILLER_25_1392 ();
 sg13g2_decap_8 FILLER_25_1399 ();
 sg13g2_decap_8 FILLER_25_1406 ();
 sg13g2_decap_8 FILLER_25_1413 ();
 sg13g2_decap_8 FILLER_25_1420 ();
 sg13g2_decap_8 FILLER_25_1427 ();
 sg13g2_decap_8 FILLER_25_1434 ();
 sg13g2_decap_8 FILLER_25_1441 ();
 sg13g2_decap_8 FILLER_25_1448 ();
 sg13g2_decap_8 FILLER_25_1455 ();
 sg13g2_decap_8 FILLER_25_1462 ();
 sg13g2_decap_8 FILLER_25_1469 ();
 sg13g2_decap_8 FILLER_25_1476 ();
 sg13g2_decap_8 FILLER_25_1483 ();
 sg13g2_decap_8 FILLER_25_1490 ();
 sg13g2_decap_8 FILLER_25_1497 ();
 sg13g2_decap_8 FILLER_25_1504 ();
 sg13g2_decap_8 FILLER_25_1511 ();
 sg13g2_decap_8 FILLER_25_1518 ();
 sg13g2_decap_8 FILLER_25_1525 ();
 sg13g2_decap_8 FILLER_25_1532 ();
 sg13g2_decap_8 FILLER_25_1539 ();
 sg13g2_decap_8 FILLER_25_1546 ();
 sg13g2_decap_8 FILLER_25_1553 ();
 sg13g2_decap_8 FILLER_25_1560 ();
 sg13g2_decap_8 FILLER_25_1567 ();
 sg13g2_decap_8 FILLER_25_1574 ();
 sg13g2_decap_8 FILLER_25_1581 ();
 sg13g2_decap_8 FILLER_25_1588 ();
 sg13g2_decap_8 FILLER_25_1595 ();
 sg13g2_decap_8 FILLER_25_1602 ();
 sg13g2_decap_8 FILLER_25_1609 ();
 sg13g2_decap_8 FILLER_25_1616 ();
 sg13g2_decap_8 FILLER_25_1623 ();
 sg13g2_decap_8 FILLER_25_1630 ();
 sg13g2_decap_8 FILLER_25_1637 ();
 sg13g2_decap_8 FILLER_25_1644 ();
 sg13g2_decap_8 FILLER_25_1651 ();
 sg13g2_decap_8 FILLER_25_1658 ();
 sg13g2_decap_8 FILLER_25_1665 ();
 sg13g2_decap_8 FILLER_25_1672 ();
 sg13g2_decap_8 FILLER_25_1679 ();
 sg13g2_decap_8 FILLER_25_1686 ();
 sg13g2_decap_8 FILLER_25_1693 ();
 sg13g2_decap_8 FILLER_25_1700 ();
 sg13g2_decap_8 FILLER_25_1707 ();
 sg13g2_decap_8 FILLER_25_1714 ();
 sg13g2_decap_8 FILLER_25_1721 ();
 sg13g2_decap_8 FILLER_25_1728 ();
 sg13g2_decap_8 FILLER_25_1735 ();
 sg13g2_decap_8 FILLER_25_1742 ();
 sg13g2_decap_8 FILLER_25_1749 ();
 sg13g2_decap_8 FILLER_25_1756 ();
 sg13g2_decap_4 FILLER_25_1763 ();
 sg13g2_fill_1 FILLER_25_1767 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_4 FILLER_26_35 ();
 sg13g2_fill_2 FILLER_26_43 ();
 sg13g2_fill_1 FILLER_26_55 ();
 sg13g2_decap_4 FILLER_26_68 ();
 sg13g2_fill_1 FILLER_26_82 ();
 sg13g2_decap_4 FILLER_26_95 ();
 sg13g2_fill_2 FILLER_26_99 ();
 sg13g2_fill_2 FILLER_26_114 ();
 sg13g2_fill_1 FILLER_26_116 ();
 sg13g2_fill_2 FILLER_26_122 ();
 sg13g2_decap_4 FILLER_26_141 ();
 sg13g2_fill_2 FILLER_26_145 ();
 sg13g2_decap_8 FILLER_26_152 ();
 sg13g2_decap_4 FILLER_26_159 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_fill_1 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_183 ();
 sg13g2_fill_2 FILLER_26_190 ();
 sg13g2_fill_2 FILLER_26_208 ();
 sg13g2_fill_1 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_265 ();
 sg13g2_fill_2 FILLER_26_272 ();
 sg13g2_fill_1 FILLER_26_274 ();
 sg13g2_fill_2 FILLER_26_288 ();
 sg13g2_fill_1 FILLER_26_290 ();
 sg13g2_fill_2 FILLER_26_385 ();
 sg13g2_fill_2 FILLER_26_415 ();
 sg13g2_fill_1 FILLER_26_417 ();
 sg13g2_fill_2 FILLER_26_435 ();
 sg13g2_fill_1 FILLER_26_441 ();
 sg13g2_fill_2 FILLER_26_485 ();
 sg13g2_fill_1 FILLER_26_487 ();
 sg13g2_decap_4 FILLER_26_525 ();
 sg13g2_fill_2 FILLER_26_565 ();
 sg13g2_fill_1 FILLER_26_567 ();
 sg13g2_decap_4 FILLER_26_626 ();
 sg13g2_fill_1 FILLER_26_640 ();
 sg13g2_fill_1 FILLER_26_685 ();
 sg13g2_decap_8 FILLER_26_695 ();
 sg13g2_decap_8 FILLER_26_702 ();
 sg13g2_decap_8 FILLER_26_709 ();
 sg13g2_fill_2 FILLER_26_716 ();
 sg13g2_fill_2 FILLER_26_766 ();
 sg13g2_fill_2 FILLER_26_799 ();
 sg13g2_fill_2 FILLER_26_806 ();
 sg13g2_fill_1 FILLER_26_820 ();
 sg13g2_decap_4 FILLER_26_836 ();
 sg13g2_fill_1 FILLER_26_840 ();
 sg13g2_decap_8 FILLER_26_872 ();
 sg13g2_fill_1 FILLER_26_879 ();
 sg13g2_decap_4 FILLER_26_886 ();
 sg13g2_fill_2 FILLER_26_890 ();
 sg13g2_decap_8 FILLER_26_923 ();
 sg13g2_decap_4 FILLER_26_930 ();
 sg13g2_fill_2 FILLER_26_934 ();
 sg13g2_decap_4 FILLER_26_941 ();
 sg13g2_fill_2 FILLER_26_945 ();
 sg13g2_fill_2 FILLER_26_951 ();
 sg13g2_decap_8 FILLER_26_997 ();
 sg13g2_decap_8 FILLER_26_1004 ();
 sg13g2_decap_8 FILLER_26_1011 ();
 sg13g2_decap_8 FILLER_26_1018 ();
 sg13g2_decap_8 FILLER_26_1025 ();
 sg13g2_decap_8 FILLER_26_1032 ();
 sg13g2_decap_8 FILLER_26_1039 ();
 sg13g2_decap_8 FILLER_26_1046 ();
 sg13g2_decap_8 FILLER_26_1053 ();
 sg13g2_decap_8 FILLER_26_1060 ();
 sg13g2_decap_8 FILLER_26_1067 ();
 sg13g2_decap_8 FILLER_26_1074 ();
 sg13g2_decap_8 FILLER_26_1081 ();
 sg13g2_decap_8 FILLER_26_1088 ();
 sg13g2_decap_8 FILLER_26_1095 ();
 sg13g2_decap_8 FILLER_26_1102 ();
 sg13g2_decap_8 FILLER_26_1109 ();
 sg13g2_decap_8 FILLER_26_1116 ();
 sg13g2_decap_8 FILLER_26_1123 ();
 sg13g2_decap_8 FILLER_26_1130 ();
 sg13g2_decap_8 FILLER_26_1137 ();
 sg13g2_decap_8 FILLER_26_1144 ();
 sg13g2_decap_8 FILLER_26_1151 ();
 sg13g2_decap_8 FILLER_26_1158 ();
 sg13g2_decap_8 FILLER_26_1165 ();
 sg13g2_decap_8 FILLER_26_1172 ();
 sg13g2_decap_8 FILLER_26_1179 ();
 sg13g2_decap_8 FILLER_26_1186 ();
 sg13g2_decap_8 FILLER_26_1193 ();
 sg13g2_decap_8 FILLER_26_1200 ();
 sg13g2_decap_8 FILLER_26_1207 ();
 sg13g2_decap_8 FILLER_26_1214 ();
 sg13g2_decap_8 FILLER_26_1221 ();
 sg13g2_decap_8 FILLER_26_1228 ();
 sg13g2_decap_8 FILLER_26_1235 ();
 sg13g2_decap_8 FILLER_26_1242 ();
 sg13g2_decap_8 FILLER_26_1249 ();
 sg13g2_decap_8 FILLER_26_1256 ();
 sg13g2_decap_8 FILLER_26_1263 ();
 sg13g2_decap_8 FILLER_26_1270 ();
 sg13g2_decap_8 FILLER_26_1277 ();
 sg13g2_decap_8 FILLER_26_1284 ();
 sg13g2_decap_8 FILLER_26_1291 ();
 sg13g2_decap_8 FILLER_26_1298 ();
 sg13g2_decap_8 FILLER_26_1305 ();
 sg13g2_decap_8 FILLER_26_1312 ();
 sg13g2_decap_8 FILLER_26_1319 ();
 sg13g2_decap_8 FILLER_26_1326 ();
 sg13g2_decap_8 FILLER_26_1333 ();
 sg13g2_decap_8 FILLER_26_1340 ();
 sg13g2_decap_8 FILLER_26_1347 ();
 sg13g2_decap_8 FILLER_26_1354 ();
 sg13g2_decap_8 FILLER_26_1361 ();
 sg13g2_decap_8 FILLER_26_1368 ();
 sg13g2_decap_8 FILLER_26_1375 ();
 sg13g2_decap_8 FILLER_26_1382 ();
 sg13g2_decap_8 FILLER_26_1389 ();
 sg13g2_decap_8 FILLER_26_1396 ();
 sg13g2_decap_8 FILLER_26_1403 ();
 sg13g2_decap_8 FILLER_26_1410 ();
 sg13g2_decap_8 FILLER_26_1417 ();
 sg13g2_decap_8 FILLER_26_1424 ();
 sg13g2_decap_8 FILLER_26_1431 ();
 sg13g2_decap_8 FILLER_26_1438 ();
 sg13g2_decap_8 FILLER_26_1445 ();
 sg13g2_decap_8 FILLER_26_1452 ();
 sg13g2_decap_8 FILLER_26_1459 ();
 sg13g2_decap_8 FILLER_26_1466 ();
 sg13g2_decap_8 FILLER_26_1473 ();
 sg13g2_decap_8 FILLER_26_1480 ();
 sg13g2_decap_8 FILLER_26_1487 ();
 sg13g2_decap_8 FILLER_26_1494 ();
 sg13g2_decap_8 FILLER_26_1501 ();
 sg13g2_decap_8 FILLER_26_1508 ();
 sg13g2_decap_8 FILLER_26_1515 ();
 sg13g2_decap_8 FILLER_26_1522 ();
 sg13g2_decap_8 FILLER_26_1529 ();
 sg13g2_decap_8 FILLER_26_1536 ();
 sg13g2_decap_8 FILLER_26_1543 ();
 sg13g2_decap_8 FILLER_26_1550 ();
 sg13g2_decap_8 FILLER_26_1557 ();
 sg13g2_decap_8 FILLER_26_1564 ();
 sg13g2_decap_8 FILLER_26_1571 ();
 sg13g2_decap_8 FILLER_26_1578 ();
 sg13g2_decap_8 FILLER_26_1585 ();
 sg13g2_decap_8 FILLER_26_1592 ();
 sg13g2_decap_8 FILLER_26_1599 ();
 sg13g2_decap_8 FILLER_26_1606 ();
 sg13g2_decap_8 FILLER_26_1613 ();
 sg13g2_decap_8 FILLER_26_1620 ();
 sg13g2_decap_8 FILLER_26_1627 ();
 sg13g2_decap_8 FILLER_26_1634 ();
 sg13g2_decap_8 FILLER_26_1641 ();
 sg13g2_decap_8 FILLER_26_1648 ();
 sg13g2_decap_8 FILLER_26_1655 ();
 sg13g2_decap_8 FILLER_26_1662 ();
 sg13g2_decap_8 FILLER_26_1669 ();
 sg13g2_decap_8 FILLER_26_1676 ();
 sg13g2_decap_8 FILLER_26_1683 ();
 sg13g2_decap_8 FILLER_26_1690 ();
 sg13g2_decap_8 FILLER_26_1697 ();
 sg13g2_decap_8 FILLER_26_1704 ();
 sg13g2_decap_8 FILLER_26_1711 ();
 sg13g2_decap_8 FILLER_26_1718 ();
 sg13g2_decap_8 FILLER_26_1725 ();
 sg13g2_decap_8 FILLER_26_1732 ();
 sg13g2_decap_8 FILLER_26_1739 ();
 sg13g2_decap_8 FILLER_26_1746 ();
 sg13g2_decap_8 FILLER_26_1753 ();
 sg13g2_decap_8 FILLER_26_1760 ();
 sg13g2_fill_1 FILLER_26_1767 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_25 ();
 sg13g2_decap_8 FILLER_27_68 ();
 sg13g2_decap_8 FILLER_27_96 ();
 sg13g2_fill_2 FILLER_27_150 ();
 sg13g2_fill_1 FILLER_27_152 ();
 sg13g2_fill_2 FILLER_27_163 ();
 sg13g2_fill_2 FILLER_27_178 ();
 sg13g2_decap_8 FILLER_27_188 ();
 sg13g2_fill_1 FILLER_27_195 ();
 sg13g2_fill_2 FILLER_27_200 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_fill_1 FILLER_27_231 ();
 sg13g2_fill_2 FILLER_27_263 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_297 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_1 FILLER_27_582 ();
 sg13g2_fill_2 FILLER_27_598 ();
 sg13g2_fill_1 FILLER_27_606 ();
 sg13g2_fill_2 FILLER_27_628 ();
 sg13g2_fill_1 FILLER_27_630 ();
 sg13g2_decap_4 FILLER_27_664 ();
 sg13g2_fill_2 FILLER_27_668 ();
 sg13g2_decap_8 FILLER_27_711 ();
 sg13g2_fill_1 FILLER_27_723 ();
 sg13g2_decap_8 FILLER_27_729 ();
 sg13g2_fill_1 FILLER_27_736 ();
 sg13g2_decap_4 FILLER_27_745 ();
 sg13g2_fill_1 FILLER_27_749 ();
 sg13g2_fill_1 FILLER_27_753 ();
 sg13g2_fill_1 FILLER_27_759 ();
 sg13g2_decap_8 FILLER_27_817 ();
 sg13g2_fill_2 FILLER_27_824 ();
 sg13g2_decap_8 FILLER_27_844 ();
 sg13g2_decap_4 FILLER_27_851 ();
 sg13g2_fill_2 FILLER_27_855 ();
 sg13g2_fill_2 FILLER_27_868 ();
 sg13g2_fill_1 FILLER_27_870 ();
 sg13g2_decap_8 FILLER_27_891 ();
 sg13g2_fill_1 FILLER_27_898 ();
 sg13g2_decap_4 FILLER_27_907 ();
 sg13g2_fill_2 FILLER_27_911 ();
 sg13g2_decap_4 FILLER_27_923 ();
 sg13g2_fill_1 FILLER_27_951 ();
 sg13g2_fill_2 FILLER_27_965 ();
 sg13g2_fill_1 FILLER_27_967 ();
 sg13g2_decap_8 FILLER_27_992 ();
 sg13g2_decap_8 FILLER_27_999 ();
 sg13g2_decap_8 FILLER_27_1006 ();
 sg13g2_decap_8 FILLER_27_1013 ();
 sg13g2_decap_8 FILLER_27_1020 ();
 sg13g2_decap_8 FILLER_27_1027 ();
 sg13g2_decap_8 FILLER_27_1034 ();
 sg13g2_decap_8 FILLER_27_1041 ();
 sg13g2_decap_8 FILLER_27_1048 ();
 sg13g2_decap_8 FILLER_27_1055 ();
 sg13g2_decap_8 FILLER_27_1062 ();
 sg13g2_decap_8 FILLER_27_1069 ();
 sg13g2_decap_8 FILLER_27_1076 ();
 sg13g2_decap_8 FILLER_27_1083 ();
 sg13g2_decap_8 FILLER_27_1090 ();
 sg13g2_decap_8 FILLER_27_1097 ();
 sg13g2_decap_8 FILLER_27_1104 ();
 sg13g2_decap_8 FILLER_27_1111 ();
 sg13g2_decap_8 FILLER_27_1118 ();
 sg13g2_decap_8 FILLER_27_1125 ();
 sg13g2_decap_8 FILLER_27_1132 ();
 sg13g2_decap_8 FILLER_27_1139 ();
 sg13g2_decap_8 FILLER_27_1146 ();
 sg13g2_decap_8 FILLER_27_1153 ();
 sg13g2_decap_8 FILLER_27_1160 ();
 sg13g2_decap_8 FILLER_27_1167 ();
 sg13g2_decap_8 FILLER_27_1174 ();
 sg13g2_decap_8 FILLER_27_1181 ();
 sg13g2_decap_8 FILLER_27_1188 ();
 sg13g2_decap_8 FILLER_27_1195 ();
 sg13g2_decap_8 FILLER_27_1202 ();
 sg13g2_decap_8 FILLER_27_1209 ();
 sg13g2_decap_8 FILLER_27_1216 ();
 sg13g2_decap_8 FILLER_27_1223 ();
 sg13g2_decap_8 FILLER_27_1230 ();
 sg13g2_decap_8 FILLER_27_1237 ();
 sg13g2_decap_8 FILLER_27_1244 ();
 sg13g2_decap_8 FILLER_27_1251 ();
 sg13g2_decap_8 FILLER_27_1258 ();
 sg13g2_decap_8 FILLER_27_1265 ();
 sg13g2_decap_8 FILLER_27_1272 ();
 sg13g2_decap_8 FILLER_27_1279 ();
 sg13g2_decap_8 FILLER_27_1286 ();
 sg13g2_decap_8 FILLER_27_1293 ();
 sg13g2_decap_8 FILLER_27_1300 ();
 sg13g2_decap_8 FILLER_27_1307 ();
 sg13g2_decap_8 FILLER_27_1314 ();
 sg13g2_decap_8 FILLER_27_1321 ();
 sg13g2_decap_8 FILLER_27_1328 ();
 sg13g2_decap_8 FILLER_27_1335 ();
 sg13g2_decap_8 FILLER_27_1342 ();
 sg13g2_decap_8 FILLER_27_1349 ();
 sg13g2_decap_8 FILLER_27_1356 ();
 sg13g2_decap_8 FILLER_27_1363 ();
 sg13g2_decap_8 FILLER_27_1370 ();
 sg13g2_decap_8 FILLER_27_1377 ();
 sg13g2_decap_8 FILLER_27_1384 ();
 sg13g2_decap_8 FILLER_27_1391 ();
 sg13g2_decap_8 FILLER_27_1398 ();
 sg13g2_decap_8 FILLER_27_1405 ();
 sg13g2_decap_8 FILLER_27_1412 ();
 sg13g2_decap_8 FILLER_27_1419 ();
 sg13g2_decap_8 FILLER_27_1426 ();
 sg13g2_decap_8 FILLER_27_1433 ();
 sg13g2_decap_8 FILLER_27_1440 ();
 sg13g2_decap_8 FILLER_27_1447 ();
 sg13g2_decap_8 FILLER_27_1454 ();
 sg13g2_decap_8 FILLER_27_1461 ();
 sg13g2_decap_8 FILLER_27_1468 ();
 sg13g2_decap_8 FILLER_27_1475 ();
 sg13g2_decap_8 FILLER_27_1482 ();
 sg13g2_decap_8 FILLER_27_1489 ();
 sg13g2_decap_8 FILLER_27_1496 ();
 sg13g2_decap_8 FILLER_27_1503 ();
 sg13g2_decap_8 FILLER_27_1510 ();
 sg13g2_decap_8 FILLER_27_1517 ();
 sg13g2_decap_8 FILLER_27_1524 ();
 sg13g2_decap_8 FILLER_27_1531 ();
 sg13g2_decap_8 FILLER_27_1538 ();
 sg13g2_decap_8 FILLER_27_1545 ();
 sg13g2_decap_8 FILLER_27_1552 ();
 sg13g2_decap_8 FILLER_27_1559 ();
 sg13g2_decap_8 FILLER_27_1566 ();
 sg13g2_decap_8 FILLER_27_1573 ();
 sg13g2_decap_8 FILLER_27_1580 ();
 sg13g2_decap_8 FILLER_27_1587 ();
 sg13g2_decap_8 FILLER_27_1594 ();
 sg13g2_decap_8 FILLER_27_1601 ();
 sg13g2_decap_8 FILLER_27_1608 ();
 sg13g2_decap_8 FILLER_27_1615 ();
 sg13g2_decap_8 FILLER_27_1622 ();
 sg13g2_decap_8 FILLER_27_1629 ();
 sg13g2_decap_8 FILLER_27_1636 ();
 sg13g2_decap_8 FILLER_27_1643 ();
 sg13g2_decap_8 FILLER_27_1650 ();
 sg13g2_decap_8 FILLER_27_1657 ();
 sg13g2_decap_8 FILLER_27_1664 ();
 sg13g2_decap_8 FILLER_27_1671 ();
 sg13g2_decap_8 FILLER_27_1678 ();
 sg13g2_decap_8 FILLER_27_1685 ();
 sg13g2_decap_8 FILLER_27_1692 ();
 sg13g2_decap_8 FILLER_27_1699 ();
 sg13g2_decap_8 FILLER_27_1706 ();
 sg13g2_decap_8 FILLER_27_1713 ();
 sg13g2_decap_8 FILLER_27_1720 ();
 sg13g2_decap_8 FILLER_27_1727 ();
 sg13g2_decap_8 FILLER_27_1734 ();
 sg13g2_decap_8 FILLER_27_1741 ();
 sg13g2_decap_8 FILLER_27_1748 ();
 sg13g2_decap_8 FILLER_27_1755 ();
 sg13g2_decap_4 FILLER_27_1762 ();
 sg13g2_fill_2 FILLER_27_1766 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_50 ();
 sg13g2_decap_4 FILLER_28_66 ();
 sg13g2_fill_2 FILLER_28_70 ();
 sg13g2_fill_1 FILLER_28_89 ();
 sg13g2_decap_8 FILLER_28_106 ();
 sg13g2_decap_4 FILLER_28_113 ();
 sg13g2_decap_8 FILLER_28_122 ();
 sg13g2_fill_2 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_131 ();
 sg13g2_fill_2 FILLER_28_141 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_decap_8 FILLER_28_148 ();
 sg13g2_fill_1 FILLER_28_163 ();
 sg13g2_fill_1 FILLER_28_181 ();
 sg13g2_fill_1 FILLER_28_190 ();
 sg13g2_decap_4 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_fill_1 FILLER_28_206 ();
 sg13g2_decap_8 FILLER_28_212 ();
 sg13g2_decap_4 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_254 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_450 ();
 sg13g2_fill_2 FILLER_28_463 ();
 sg13g2_fill_2 FILLER_28_474 ();
 sg13g2_fill_1 FILLER_28_495 ();
 sg13g2_fill_2 FILLER_28_522 ();
 sg13g2_fill_1 FILLER_28_524 ();
 sg13g2_fill_1 FILLER_28_543 ();
 sg13g2_decap_4 FILLER_28_596 ();
 sg13g2_fill_1 FILLER_28_600 ();
 sg13g2_decap_4 FILLER_28_611 ();
 sg13g2_fill_2 FILLER_28_615 ();
 sg13g2_decap_8 FILLER_28_622 ();
 sg13g2_decap_8 FILLER_28_629 ();
 sg13g2_decap_4 FILLER_28_636 ();
 sg13g2_decap_8 FILLER_28_658 ();
 sg13g2_fill_2 FILLER_28_665 ();
 sg13g2_fill_1 FILLER_28_667 ();
 sg13g2_fill_1 FILLER_28_693 ();
 sg13g2_fill_2 FILLER_28_699 ();
 sg13g2_fill_1 FILLER_28_701 ();
 sg13g2_decap_4 FILLER_28_716 ();
 sg13g2_fill_2 FILLER_28_772 ();
 sg13g2_fill_2 FILLER_28_789 ();
 sg13g2_fill_1 FILLER_28_796 ();
 sg13g2_decap_8 FILLER_28_807 ();
 sg13g2_decap_4 FILLER_28_814 ();
 sg13g2_fill_1 FILLER_28_818 ();
 sg13g2_fill_1 FILLER_28_828 ();
 sg13g2_decap_8 FILLER_28_855 ();
 sg13g2_decap_8 FILLER_28_862 ();
 sg13g2_decap_8 FILLER_28_869 ();
 sg13g2_decap_4 FILLER_28_876 ();
 sg13g2_fill_1 FILLER_28_880 ();
 sg13g2_fill_2 FILLER_28_885 ();
 sg13g2_fill_1 FILLER_28_887 ();
 sg13g2_decap_4 FILLER_28_893 ();
 sg13g2_fill_2 FILLER_28_907 ();
 sg13g2_fill_1 FILLER_28_909 ();
 sg13g2_decap_8 FILLER_28_921 ();
 sg13g2_decap_4 FILLER_28_928 ();
 sg13g2_fill_1 FILLER_28_932 ();
 sg13g2_decap_8 FILLER_28_942 ();
 sg13g2_fill_1 FILLER_28_949 ();
 sg13g2_fill_1 FILLER_28_962 ();
 sg13g2_decap_8 FILLER_28_967 ();
 sg13g2_fill_2 FILLER_28_974 ();
 sg13g2_fill_1 FILLER_28_980 ();
 sg13g2_decap_8 FILLER_28_994 ();
 sg13g2_decap_8 FILLER_28_1001 ();
 sg13g2_decap_8 FILLER_28_1008 ();
 sg13g2_decap_8 FILLER_28_1015 ();
 sg13g2_decap_8 FILLER_28_1022 ();
 sg13g2_decap_8 FILLER_28_1029 ();
 sg13g2_decap_8 FILLER_28_1036 ();
 sg13g2_decap_8 FILLER_28_1043 ();
 sg13g2_decap_8 FILLER_28_1050 ();
 sg13g2_decap_8 FILLER_28_1057 ();
 sg13g2_decap_8 FILLER_28_1064 ();
 sg13g2_decap_8 FILLER_28_1071 ();
 sg13g2_decap_8 FILLER_28_1078 ();
 sg13g2_decap_8 FILLER_28_1085 ();
 sg13g2_decap_8 FILLER_28_1092 ();
 sg13g2_decap_8 FILLER_28_1099 ();
 sg13g2_decap_8 FILLER_28_1106 ();
 sg13g2_decap_8 FILLER_28_1113 ();
 sg13g2_decap_8 FILLER_28_1120 ();
 sg13g2_decap_8 FILLER_28_1127 ();
 sg13g2_decap_8 FILLER_28_1134 ();
 sg13g2_decap_8 FILLER_28_1141 ();
 sg13g2_decap_8 FILLER_28_1148 ();
 sg13g2_decap_8 FILLER_28_1155 ();
 sg13g2_decap_8 FILLER_28_1162 ();
 sg13g2_decap_8 FILLER_28_1169 ();
 sg13g2_decap_8 FILLER_28_1176 ();
 sg13g2_decap_8 FILLER_28_1183 ();
 sg13g2_decap_8 FILLER_28_1190 ();
 sg13g2_decap_8 FILLER_28_1197 ();
 sg13g2_decap_8 FILLER_28_1204 ();
 sg13g2_decap_8 FILLER_28_1211 ();
 sg13g2_decap_8 FILLER_28_1218 ();
 sg13g2_decap_8 FILLER_28_1225 ();
 sg13g2_decap_8 FILLER_28_1232 ();
 sg13g2_decap_8 FILLER_28_1239 ();
 sg13g2_decap_8 FILLER_28_1246 ();
 sg13g2_decap_8 FILLER_28_1253 ();
 sg13g2_decap_8 FILLER_28_1260 ();
 sg13g2_decap_8 FILLER_28_1267 ();
 sg13g2_decap_8 FILLER_28_1274 ();
 sg13g2_decap_8 FILLER_28_1281 ();
 sg13g2_decap_8 FILLER_28_1288 ();
 sg13g2_decap_8 FILLER_28_1295 ();
 sg13g2_decap_8 FILLER_28_1302 ();
 sg13g2_decap_8 FILLER_28_1309 ();
 sg13g2_decap_8 FILLER_28_1316 ();
 sg13g2_decap_8 FILLER_28_1323 ();
 sg13g2_decap_8 FILLER_28_1330 ();
 sg13g2_decap_8 FILLER_28_1337 ();
 sg13g2_decap_8 FILLER_28_1344 ();
 sg13g2_decap_8 FILLER_28_1351 ();
 sg13g2_decap_8 FILLER_28_1358 ();
 sg13g2_decap_8 FILLER_28_1365 ();
 sg13g2_decap_8 FILLER_28_1372 ();
 sg13g2_decap_8 FILLER_28_1379 ();
 sg13g2_decap_8 FILLER_28_1386 ();
 sg13g2_decap_8 FILLER_28_1393 ();
 sg13g2_decap_8 FILLER_28_1400 ();
 sg13g2_decap_8 FILLER_28_1407 ();
 sg13g2_decap_8 FILLER_28_1414 ();
 sg13g2_decap_8 FILLER_28_1421 ();
 sg13g2_decap_8 FILLER_28_1428 ();
 sg13g2_decap_8 FILLER_28_1435 ();
 sg13g2_decap_8 FILLER_28_1442 ();
 sg13g2_decap_8 FILLER_28_1449 ();
 sg13g2_decap_8 FILLER_28_1456 ();
 sg13g2_decap_8 FILLER_28_1463 ();
 sg13g2_decap_8 FILLER_28_1470 ();
 sg13g2_decap_8 FILLER_28_1477 ();
 sg13g2_decap_8 FILLER_28_1484 ();
 sg13g2_decap_8 FILLER_28_1491 ();
 sg13g2_decap_8 FILLER_28_1498 ();
 sg13g2_decap_8 FILLER_28_1505 ();
 sg13g2_decap_8 FILLER_28_1512 ();
 sg13g2_decap_8 FILLER_28_1519 ();
 sg13g2_decap_8 FILLER_28_1526 ();
 sg13g2_decap_8 FILLER_28_1533 ();
 sg13g2_decap_8 FILLER_28_1540 ();
 sg13g2_decap_8 FILLER_28_1547 ();
 sg13g2_decap_8 FILLER_28_1554 ();
 sg13g2_decap_8 FILLER_28_1561 ();
 sg13g2_decap_8 FILLER_28_1568 ();
 sg13g2_decap_8 FILLER_28_1575 ();
 sg13g2_decap_8 FILLER_28_1582 ();
 sg13g2_decap_8 FILLER_28_1589 ();
 sg13g2_decap_8 FILLER_28_1596 ();
 sg13g2_decap_8 FILLER_28_1603 ();
 sg13g2_decap_8 FILLER_28_1610 ();
 sg13g2_decap_8 FILLER_28_1617 ();
 sg13g2_decap_8 FILLER_28_1624 ();
 sg13g2_decap_8 FILLER_28_1631 ();
 sg13g2_decap_8 FILLER_28_1638 ();
 sg13g2_decap_8 FILLER_28_1645 ();
 sg13g2_decap_8 FILLER_28_1652 ();
 sg13g2_decap_8 FILLER_28_1659 ();
 sg13g2_decap_8 FILLER_28_1666 ();
 sg13g2_decap_8 FILLER_28_1673 ();
 sg13g2_decap_8 FILLER_28_1680 ();
 sg13g2_decap_8 FILLER_28_1687 ();
 sg13g2_decap_8 FILLER_28_1694 ();
 sg13g2_decap_8 FILLER_28_1701 ();
 sg13g2_decap_8 FILLER_28_1708 ();
 sg13g2_decap_8 FILLER_28_1715 ();
 sg13g2_decap_8 FILLER_28_1722 ();
 sg13g2_decap_8 FILLER_28_1729 ();
 sg13g2_decap_8 FILLER_28_1736 ();
 sg13g2_decap_8 FILLER_28_1743 ();
 sg13g2_decap_8 FILLER_28_1750 ();
 sg13g2_decap_8 FILLER_28_1757 ();
 sg13g2_decap_4 FILLER_28_1764 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_fill_1 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_96 ();
 sg13g2_fill_1 FILLER_29_98 ();
 sg13g2_fill_2 FILLER_29_112 ();
 sg13g2_decap_4 FILLER_29_131 ();
 sg13g2_fill_1 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_169 ();
 sg13g2_fill_1 FILLER_29_171 ();
 sg13g2_fill_1 FILLER_29_180 ();
 sg13g2_decap_4 FILLER_29_213 ();
 sg13g2_fill_2 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_247 ();
 sg13g2_fill_2 FILLER_29_298 ();
 sg13g2_fill_1 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_338 ();
 sg13g2_fill_1 FILLER_29_390 ();
 sg13g2_fill_2 FILLER_29_405 ();
 sg13g2_fill_1 FILLER_29_407 ();
 sg13g2_fill_2 FILLER_29_457 ();
 sg13g2_fill_2 FILLER_29_557 ();
 sg13g2_fill_1 FILLER_29_559 ();
 sg13g2_decap_8 FILLER_29_574 ();
 sg13g2_fill_2 FILLER_29_581 ();
 sg13g2_decap_8 FILLER_29_592 ();
 sg13g2_fill_2 FILLER_29_599 ();
 sg13g2_fill_1 FILLER_29_601 ();
 sg13g2_decap_8 FILLER_29_630 ();
 sg13g2_fill_1 FILLER_29_637 ();
 sg13g2_decap_4 FILLER_29_643 ();
 sg13g2_fill_1 FILLER_29_660 ();
 sg13g2_decap_4 FILLER_29_681 ();
 sg13g2_fill_1 FILLER_29_692 ();
 sg13g2_decap_4 FILLER_29_707 ();
 sg13g2_fill_1 FILLER_29_711 ();
 sg13g2_fill_2 FILLER_29_751 ();
 sg13g2_fill_2 FILLER_29_769 ();
 sg13g2_fill_1 FILLER_29_777 ();
 sg13g2_decap_8 FILLER_29_790 ();
 sg13g2_fill_1 FILLER_29_801 ();
 sg13g2_decap_4 FILLER_29_841 ();
 sg13g2_fill_1 FILLER_29_881 ();
 sg13g2_fill_1 FILLER_29_898 ();
 sg13g2_fill_2 FILLER_29_920 ();
 sg13g2_fill_1 FILLER_29_949 ();
 sg13g2_fill_1 FILLER_29_976 ();
 sg13g2_decap_8 FILLER_29_993 ();
 sg13g2_decap_8 FILLER_29_1000 ();
 sg13g2_decap_8 FILLER_29_1007 ();
 sg13g2_decap_8 FILLER_29_1014 ();
 sg13g2_decap_8 FILLER_29_1021 ();
 sg13g2_decap_8 FILLER_29_1028 ();
 sg13g2_decap_8 FILLER_29_1035 ();
 sg13g2_decap_8 FILLER_29_1042 ();
 sg13g2_decap_8 FILLER_29_1049 ();
 sg13g2_decap_8 FILLER_29_1056 ();
 sg13g2_decap_8 FILLER_29_1063 ();
 sg13g2_decap_8 FILLER_29_1070 ();
 sg13g2_decap_8 FILLER_29_1077 ();
 sg13g2_decap_8 FILLER_29_1084 ();
 sg13g2_decap_8 FILLER_29_1091 ();
 sg13g2_decap_8 FILLER_29_1098 ();
 sg13g2_decap_8 FILLER_29_1105 ();
 sg13g2_decap_8 FILLER_29_1112 ();
 sg13g2_decap_8 FILLER_29_1119 ();
 sg13g2_decap_8 FILLER_29_1126 ();
 sg13g2_decap_8 FILLER_29_1133 ();
 sg13g2_decap_8 FILLER_29_1140 ();
 sg13g2_decap_8 FILLER_29_1147 ();
 sg13g2_decap_8 FILLER_29_1154 ();
 sg13g2_decap_8 FILLER_29_1161 ();
 sg13g2_decap_8 FILLER_29_1168 ();
 sg13g2_decap_8 FILLER_29_1175 ();
 sg13g2_decap_8 FILLER_29_1182 ();
 sg13g2_decap_8 FILLER_29_1189 ();
 sg13g2_decap_8 FILLER_29_1196 ();
 sg13g2_decap_8 FILLER_29_1203 ();
 sg13g2_decap_8 FILLER_29_1210 ();
 sg13g2_decap_8 FILLER_29_1217 ();
 sg13g2_decap_8 FILLER_29_1224 ();
 sg13g2_decap_8 FILLER_29_1231 ();
 sg13g2_decap_8 FILLER_29_1238 ();
 sg13g2_decap_8 FILLER_29_1245 ();
 sg13g2_decap_8 FILLER_29_1252 ();
 sg13g2_decap_8 FILLER_29_1259 ();
 sg13g2_decap_8 FILLER_29_1266 ();
 sg13g2_decap_8 FILLER_29_1273 ();
 sg13g2_decap_8 FILLER_29_1280 ();
 sg13g2_decap_8 FILLER_29_1287 ();
 sg13g2_decap_8 FILLER_29_1294 ();
 sg13g2_decap_8 FILLER_29_1301 ();
 sg13g2_decap_8 FILLER_29_1308 ();
 sg13g2_decap_8 FILLER_29_1315 ();
 sg13g2_decap_8 FILLER_29_1322 ();
 sg13g2_decap_8 FILLER_29_1329 ();
 sg13g2_decap_8 FILLER_29_1336 ();
 sg13g2_decap_8 FILLER_29_1343 ();
 sg13g2_decap_8 FILLER_29_1350 ();
 sg13g2_decap_8 FILLER_29_1357 ();
 sg13g2_decap_8 FILLER_29_1364 ();
 sg13g2_decap_8 FILLER_29_1371 ();
 sg13g2_decap_8 FILLER_29_1378 ();
 sg13g2_decap_8 FILLER_29_1385 ();
 sg13g2_decap_8 FILLER_29_1392 ();
 sg13g2_decap_8 FILLER_29_1399 ();
 sg13g2_decap_8 FILLER_29_1406 ();
 sg13g2_decap_8 FILLER_29_1413 ();
 sg13g2_decap_8 FILLER_29_1420 ();
 sg13g2_decap_8 FILLER_29_1427 ();
 sg13g2_decap_8 FILLER_29_1434 ();
 sg13g2_decap_8 FILLER_29_1441 ();
 sg13g2_decap_8 FILLER_29_1448 ();
 sg13g2_decap_8 FILLER_29_1455 ();
 sg13g2_decap_8 FILLER_29_1462 ();
 sg13g2_decap_8 FILLER_29_1469 ();
 sg13g2_decap_8 FILLER_29_1476 ();
 sg13g2_decap_8 FILLER_29_1483 ();
 sg13g2_decap_8 FILLER_29_1490 ();
 sg13g2_decap_8 FILLER_29_1497 ();
 sg13g2_decap_8 FILLER_29_1504 ();
 sg13g2_decap_8 FILLER_29_1511 ();
 sg13g2_decap_8 FILLER_29_1518 ();
 sg13g2_decap_8 FILLER_29_1525 ();
 sg13g2_decap_8 FILLER_29_1532 ();
 sg13g2_decap_8 FILLER_29_1539 ();
 sg13g2_decap_8 FILLER_29_1546 ();
 sg13g2_decap_8 FILLER_29_1553 ();
 sg13g2_decap_8 FILLER_29_1560 ();
 sg13g2_decap_8 FILLER_29_1567 ();
 sg13g2_decap_8 FILLER_29_1574 ();
 sg13g2_decap_8 FILLER_29_1581 ();
 sg13g2_decap_8 FILLER_29_1588 ();
 sg13g2_decap_8 FILLER_29_1595 ();
 sg13g2_decap_8 FILLER_29_1602 ();
 sg13g2_decap_8 FILLER_29_1609 ();
 sg13g2_decap_8 FILLER_29_1616 ();
 sg13g2_decap_8 FILLER_29_1623 ();
 sg13g2_decap_8 FILLER_29_1630 ();
 sg13g2_decap_8 FILLER_29_1637 ();
 sg13g2_decap_8 FILLER_29_1644 ();
 sg13g2_decap_8 FILLER_29_1651 ();
 sg13g2_decap_8 FILLER_29_1658 ();
 sg13g2_decap_8 FILLER_29_1665 ();
 sg13g2_decap_8 FILLER_29_1672 ();
 sg13g2_decap_8 FILLER_29_1679 ();
 sg13g2_decap_8 FILLER_29_1686 ();
 sg13g2_decap_8 FILLER_29_1693 ();
 sg13g2_decap_8 FILLER_29_1700 ();
 sg13g2_decap_8 FILLER_29_1707 ();
 sg13g2_decap_8 FILLER_29_1714 ();
 sg13g2_decap_8 FILLER_29_1721 ();
 sg13g2_decap_8 FILLER_29_1728 ();
 sg13g2_decap_8 FILLER_29_1735 ();
 sg13g2_decap_8 FILLER_29_1742 ();
 sg13g2_decap_8 FILLER_29_1749 ();
 sg13g2_decap_8 FILLER_29_1756 ();
 sg13g2_decap_4 FILLER_29_1763 ();
 sg13g2_fill_1 FILLER_29_1767 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_4 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_25 ();
 sg13g2_fill_1 FILLER_30_51 ();
 sg13g2_fill_2 FILLER_30_90 ();
 sg13g2_fill_1 FILLER_30_92 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_fill_2 FILLER_30_105 ();
 sg13g2_fill_1 FILLER_30_107 ();
 sg13g2_fill_2 FILLER_30_120 ();
 sg13g2_fill_1 FILLER_30_122 ();
 sg13g2_decap_8 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_143 ();
 sg13g2_decap_4 FILLER_30_150 ();
 sg13g2_fill_2 FILLER_30_154 ();
 sg13g2_fill_2 FILLER_30_160 ();
 sg13g2_fill_1 FILLER_30_162 ();
 sg13g2_decap_4 FILLER_30_167 ();
 sg13g2_decap_8 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_190 ();
 sg13g2_decap_4 FILLER_30_197 ();
 sg13g2_fill_1 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_206 ();
 sg13g2_fill_1 FILLER_30_213 ();
 sg13g2_decap_4 FILLER_30_249 ();
 sg13g2_fill_2 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_266 ();
 sg13g2_fill_2 FILLER_30_287 ();
 sg13g2_fill_1 FILLER_30_320 ();
 sg13g2_fill_2 FILLER_30_384 ();
 sg13g2_fill_2 FILLER_30_458 ();
 sg13g2_fill_1 FILLER_30_474 ();
 sg13g2_fill_1 FILLER_30_480 ();
 sg13g2_fill_2 FILLER_30_494 ();
 sg13g2_fill_2 FILLER_30_547 ();
 sg13g2_decap_8 FILLER_30_559 ();
 sg13g2_decap_8 FILLER_30_566 ();
 sg13g2_fill_1 FILLER_30_573 ();
 sg13g2_decap_8 FILLER_30_598 ();
 sg13g2_decap_8 FILLER_30_605 ();
 sg13g2_decap_4 FILLER_30_621 ();
 sg13g2_fill_1 FILLER_30_625 ();
 sg13g2_fill_2 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_664 ();
 sg13g2_fill_2 FILLER_30_671 ();
 sg13g2_decap_4 FILLER_30_681 ();
 sg13g2_fill_1 FILLER_30_713 ();
 sg13g2_fill_1 FILLER_30_779 ();
 sg13g2_fill_1 FILLER_30_815 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_4 FILLER_30_847 ();
 sg13g2_fill_2 FILLER_30_851 ();
 sg13g2_decap_8 FILLER_30_874 ();
 sg13g2_fill_1 FILLER_30_881 ();
 sg13g2_decap_4 FILLER_30_897 ();
 sg13g2_fill_2 FILLER_30_901 ();
 sg13g2_fill_1 FILLER_30_911 ();
 sg13g2_decap_4 FILLER_30_922 ();
 sg13g2_fill_1 FILLER_30_926 ();
 sg13g2_decap_4 FILLER_30_944 ();
 sg13g2_fill_2 FILLER_30_948 ();
 sg13g2_fill_2 FILLER_30_968 ();
 sg13g2_fill_1 FILLER_30_980 ();
 sg13g2_decap_8 FILLER_30_989 ();
 sg13g2_decap_8 FILLER_30_996 ();
 sg13g2_decap_8 FILLER_30_1003 ();
 sg13g2_decap_8 FILLER_30_1010 ();
 sg13g2_decap_8 FILLER_30_1017 ();
 sg13g2_decap_8 FILLER_30_1024 ();
 sg13g2_decap_8 FILLER_30_1031 ();
 sg13g2_decap_8 FILLER_30_1038 ();
 sg13g2_decap_8 FILLER_30_1045 ();
 sg13g2_decap_8 FILLER_30_1052 ();
 sg13g2_decap_8 FILLER_30_1059 ();
 sg13g2_decap_8 FILLER_30_1066 ();
 sg13g2_decap_8 FILLER_30_1073 ();
 sg13g2_decap_8 FILLER_30_1080 ();
 sg13g2_decap_8 FILLER_30_1087 ();
 sg13g2_decap_8 FILLER_30_1094 ();
 sg13g2_decap_8 FILLER_30_1101 ();
 sg13g2_decap_8 FILLER_30_1108 ();
 sg13g2_decap_8 FILLER_30_1115 ();
 sg13g2_decap_8 FILLER_30_1122 ();
 sg13g2_decap_8 FILLER_30_1129 ();
 sg13g2_decap_8 FILLER_30_1136 ();
 sg13g2_decap_8 FILLER_30_1143 ();
 sg13g2_decap_8 FILLER_30_1150 ();
 sg13g2_decap_8 FILLER_30_1157 ();
 sg13g2_decap_8 FILLER_30_1164 ();
 sg13g2_decap_8 FILLER_30_1171 ();
 sg13g2_decap_8 FILLER_30_1178 ();
 sg13g2_decap_8 FILLER_30_1185 ();
 sg13g2_decap_8 FILLER_30_1192 ();
 sg13g2_decap_8 FILLER_30_1199 ();
 sg13g2_decap_8 FILLER_30_1206 ();
 sg13g2_decap_8 FILLER_30_1213 ();
 sg13g2_decap_8 FILLER_30_1220 ();
 sg13g2_decap_8 FILLER_30_1227 ();
 sg13g2_decap_8 FILLER_30_1234 ();
 sg13g2_decap_8 FILLER_30_1241 ();
 sg13g2_decap_8 FILLER_30_1248 ();
 sg13g2_decap_8 FILLER_30_1255 ();
 sg13g2_decap_8 FILLER_30_1262 ();
 sg13g2_decap_8 FILLER_30_1269 ();
 sg13g2_decap_8 FILLER_30_1276 ();
 sg13g2_decap_8 FILLER_30_1283 ();
 sg13g2_decap_8 FILLER_30_1290 ();
 sg13g2_decap_8 FILLER_30_1297 ();
 sg13g2_decap_8 FILLER_30_1304 ();
 sg13g2_decap_8 FILLER_30_1311 ();
 sg13g2_decap_8 FILLER_30_1318 ();
 sg13g2_decap_8 FILLER_30_1325 ();
 sg13g2_decap_8 FILLER_30_1332 ();
 sg13g2_decap_8 FILLER_30_1339 ();
 sg13g2_decap_8 FILLER_30_1346 ();
 sg13g2_decap_8 FILLER_30_1353 ();
 sg13g2_decap_8 FILLER_30_1360 ();
 sg13g2_decap_8 FILLER_30_1367 ();
 sg13g2_decap_8 FILLER_30_1374 ();
 sg13g2_decap_8 FILLER_30_1381 ();
 sg13g2_decap_8 FILLER_30_1388 ();
 sg13g2_decap_8 FILLER_30_1395 ();
 sg13g2_decap_8 FILLER_30_1402 ();
 sg13g2_decap_8 FILLER_30_1409 ();
 sg13g2_decap_8 FILLER_30_1416 ();
 sg13g2_decap_8 FILLER_30_1423 ();
 sg13g2_decap_8 FILLER_30_1430 ();
 sg13g2_decap_8 FILLER_30_1437 ();
 sg13g2_decap_8 FILLER_30_1444 ();
 sg13g2_decap_8 FILLER_30_1451 ();
 sg13g2_decap_8 FILLER_30_1458 ();
 sg13g2_decap_8 FILLER_30_1465 ();
 sg13g2_decap_8 FILLER_30_1472 ();
 sg13g2_decap_8 FILLER_30_1479 ();
 sg13g2_decap_8 FILLER_30_1486 ();
 sg13g2_decap_8 FILLER_30_1493 ();
 sg13g2_decap_8 FILLER_30_1500 ();
 sg13g2_decap_8 FILLER_30_1507 ();
 sg13g2_decap_8 FILLER_30_1514 ();
 sg13g2_decap_8 FILLER_30_1521 ();
 sg13g2_decap_8 FILLER_30_1528 ();
 sg13g2_decap_8 FILLER_30_1535 ();
 sg13g2_decap_8 FILLER_30_1542 ();
 sg13g2_decap_8 FILLER_30_1549 ();
 sg13g2_decap_8 FILLER_30_1556 ();
 sg13g2_decap_8 FILLER_30_1563 ();
 sg13g2_decap_8 FILLER_30_1570 ();
 sg13g2_decap_8 FILLER_30_1577 ();
 sg13g2_decap_8 FILLER_30_1584 ();
 sg13g2_decap_8 FILLER_30_1591 ();
 sg13g2_decap_8 FILLER_30_1598 ();
 sg13g2_decap_8 FILLER_30_1605 ();
 sg13g2_decap_8 FILLER_30_1612 ();
 sg13g2_decap_8 FILLER_30_1619 ();
 sg13g2_decap_8 FILLER_30_1626 ();
 sg13g2_decap_8 FILLER_30_1633 ();
 sg13g2_decap_8 FILLER_30_1640 ();
 sg13g2_decap_8 FILLER_30_1647 ();
 sg13g2_decap_8 FILLER_30_1654 ();
 sg13g2_decap_8 FILLER_30_1661 ();
 sg13g2_decap_8 FILLER_30_1668 ();
 sg13g2_decap_8 FILLER_30_1675 ();
 sg13g2_decap_8 FILLER_30_1682 ();
 sg13g2_decap_8 FILLER_30_1689 ();
 sg13g2_decap_8 FILLER_30_1696 ();
 sg13g2_decap_8 FILLER_30_1703 ();
 sg13g2_decap_8 FILLER_30_1710 ();
 sg13g2_decap_8 FILLER_30_1717 ();
 sg13g2_decap_8 FILLER_30_1724 ();
 sg13g2_decap_8 FILLER_30_1731 ();
 sg13g2_decap_8 FILLER_30_1738 ();
 sg13g2_decap_8 FILLER_30_1745 ();
 sg13g2_decap_8 FILLER_30_1752 ();
 sg13g2_decap_8 FILLER_30_1759 ();
 sg13g2_fill_2 FILLER_30_1766 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_4 FILLER_31_28 ();
 sg13g2_fill_1 FILLER_31_72 ();
 sg13g2_fill_2 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_93 ();
 sg13g2_decap_4 FILLER_31_100 ();
 sg13g2_fill_2 FILLER_31_118 ();
 sg13g2_fill_2 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_fill_1 FILLER_31_153 ();
 sg13g2_fill_2 FILLER_31_162 ();
 sg13g2_decap_8 FILLER_31_206 ();
 sg13g2_decap_4 FILLER_31_213 ();
 sg13g2_fill_2 FILLER_31_217 ();
 sg13g2_decap_4 FILLER_31_265 ();
 sg13g2_fill_1 FILLER_31_269 ();
 sg13g2_fill_1 FILLER_31_281 ();
 sg13g2_fill_2 FILLER_31_381 ();
 sg13g2_fill_1 FILLER_31_383 ();
 sg13g2_fill_1 FILLER_31_394 ();
 sg13g2_fill_2 FILLER_31_455 ();
 sg13g2_fill_1 FILLER_31_499 ();
 sg13g2_fill_2 FILLER_31_510 ();
 sg13g2_fill_2 FILLER_31_516 ();
 sg13g2_fill_1 FILLER_31_518 ();
 sg13g2_fill_2 FILLER_31_523 ();
 sg13g2_fill_1 FILLER_31_525 ();
 sg13g2_decap_8 FILLER_31_547 ();
 sg13g2_decap_8 FILLER_31_554 ();
 sg13g2_fill_2 FILLER_31_561 ();
 sg13g2_fill_1 FILLER_31_563 ();
 sg13g2_fill_1 FILLER_31_605 ();
 sg13g2_decap_8 FILLER_31_628 ();
 sg13g2_decap_8 FILLER_31_635 ();
 sg13g2_fill_2 FILLER_31_642 ();
 sg13g2_decap_8 FILLER_31_649 ();
 sg13g2_fill_1 FILLER_31_656 ();
 sg13g2_decap_8 FILLER_31_661 ();
 sg13g2_decap_8 FILLER_31_668 ();
 sg13g2_decap_4 FILLER_31_675 ();
 sg13g2_fill_2 FILLER_31_687 ();
 sg13g2_fill_1 FILLER_31_715 ();
 sg13g2_decap_4 FILLER_31_719 ();
 sg13g2_decap_8 FILLER_31_730 ();
 sg13g2_decap_8 FILLER_31_742 ();
 sg13g2_decap_4 FILLER_31_749 ();
 sg13g2_fill_1 FILLER_31_753 ();
 sg13g2_fill_1 FILLER_31_761 ();
 sg13g2_decap_4 FILLER_31_767 ();
 sg13g2_fill_1 FILLER_31_771 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_4 FILLER_31_797 ();
 sg13g2_fill_1 FILLER_31_801 ();
 sg13g2_decap_8 FILLER_31_815 ();
 sg13g2_decap_4 FILLER_31_822 ();
 sg13g2_fill_1 FILLER_31_826 ();
 sg13g2_decap_4 FILLER_31_842 ();
 sg13g2_decap_8 FILLER_31_867 ();
 sg13g2_decap_4 FILLER_31_881 ();
 sg13g2_fill_2 FILLER_31_885 ();
 sg13g2_fill_2 FILLER_31_896 ();
 sg13g2_decap_8 FILLER_31_922 ();
 sg13g2_fill_1 FILLER_31_929 ();
 sg13g2_decap_8 FILLER_31_943 ();
 sg13g2_fill_2 FILLER_31_975 ();
 sg13g2_decap_8 FILLER_31_994 ();
 sg13g2_decap_8 FILLER_31_1001 ();
 sg13g2_decap_8 FILLER_31_1008 ();
 sg13g2_decap_8 FILLER_31_1015 ();
 sg13g2_decap_8 FILLER_31_1022 ();
 sg13g2_decap_8 FILLER_31_1029 ();
 sg13g2_decap_8 FILLER_31_1036 ();
 sg13g2_decap_8 FILLER_31_1043 ();
 sg13g2_decap_8 FILLER_31_1050 ();
 sg13g2_decap_8 FILLER_31_1057 ();
 sg13g2_decap_8 FILLER_31_1064 ();
 sg13g2_decap_8 FILLER_31_1071 ();
 sg13g2_decap_8 FILLER_31_1078 ();
 sg13g2_decap_8 FILLER_31_1085 ();
 sg13g2_decap_8 FILLER_31_1092 ();
 sg13g2_decap_8 FILLER_31_1099 ();
 sg13g2_decap_8 FILLER_31_1106 ();
 sg13g2_decap_8 FILLER_31_1113 ();
 sg13g2_decap_8 FILLER_31_1120 ();
 sg13g2_decap_8 FILLER_31_1127 ();
 sg13g2_decap_8 FILLER_31_1134 ();
 sg13g2_decap_8 FILLER_31_1141 ();
 sg13g2_decap_8 FILLER_31_1148 ();
 sg13g2_decap_8 FILLER_31_1155 ();
 sg13g2_decap_8 FILLER_31_1162 ();
 sg13g2_decap_8 FILLER_31_1169 ();
 sg13g2_decap_8 FILLER_31_1176 ();
 sg13g2_decap_8 FILLER_31_1183 ();
 sg13g2_decap_8 FILLER_31_1190 ();
 sg13g2_decap_8 FILLER_31_1197 ();
 sg13g2_decap_8 FILLER_31_1204 ();
 sg13g2_decap_8 FILLER_31_1211 ();
 sg13g2_decap_8 FILLER_31_1218 ();
 sg13g2_decap_8 FILLER_31_1225 ();
 sg13g2_decap_8 FILLER_31_1232 ();
 sg13g2_decap_8 FILLER_31_1239 ();
 sg13g2_decap_8 FILLER_31_1246 ();
 sg13g2_decap_8 FILLER_31_1253 ();
 sg13g2_decap_8 FILLER_31_1260 ();
 sg13g2_decap_8 FILLER_31_1267 ();
 sg13g2_decap_8 FILLER_31_1274 ();
 sg13g2_decap_8 FILLER_31_1281 ();
 sg13g2_decap_8 FILLER_31_1288 ();
 sg13g2_decap_8 FILLER_31_1295 ();
 sg13g2_decap_8 FILLER_31_1302 ();
 sg13g2_decap_8 FILLER_31_1309 ();
 sg13g2_decap_8 FILLER_31_1316 ();
 sg13g2_decap_8 FILLER_31_1323 ();
 sg13g2_decap_8 FILLER_31_1330 ();
 sg13g2_decap_8 FILLER_31_1337 ();
 sg13g2_decap_8 FILLER_31_1344 ();
 sg13g2_decap_8 FILLER_31_1351 ();
 sg13g2_decap_8 FILLER_31_1358 ();
 sg13g2_decap_8 FILLER_31_1365 ();
 sg13g2_decap_8 FILLER_31_1372 ();
 sg13g2_decap_8 FILLER_31_1379 ();
 sg13g2_decap_8 FILLER_31_1386 ();
 sg13g2_decap_8 FILLER_31_1393 ();
 sg13g2_decap_8 FILLER_31_1400 ();
 sg13g2_decap_8 FILLER_31_1407 ();
 sg13g2_decap_8 FILLER_31_1414 ();
 sg13g2_decap_8 FILLER_31_1421 ();
 sg13g2_decap_8 FILLER_31_1428 ();
 sg13g2_decap_8 FILLER_31_1435 ();
 sg13g2_decap_8 FILLER_31_1442 ();
 sg13g2_decap_8 FILLER_31_1449 ();
 sg13g2_decap_8 FILLER_31_1456 ();
 sg13g2_decap_8 FILLER_31_1463 ();
 sg13g2_decap_8 FILLER_31_1470 ();
 sg13g2_decap_8 FILLER_31_1477 ();
 sg13g2_decap_8 FILLER_31_1484 ();
 sg13g2_decap_8 FILLER_31_1491 ();
 sg13g2_decap_8 FILLER_31_1498 ();
 sg13g2_decap_8 FILLER_31_1505 ();
 sg13g2_decap_8 FILLER_31_1512 ();
 sg13g2_decap_8 FILLER_31_1519 ();
 sg13g2_decap_8 FILLER_31_1526 ();
 sg13g2_decap_8 FILLER_31_1533 ();
 sg13g2_decap_8 FILLER_31_1540 ();
 sg13g2_decap_8 FILLER_31_1547 ();
 sg13g2_decap_8 FILLER_31_1554 ();
 sg13g2_decap_8 FILLER_31_1561 ();
 sg13g2_decap_8 FILLER_31_1568 ();
 sg13g2_decap_8 FILLER_31_1575 ();
 sg13g2_decap_8 FILLER_31_1582 ();
 sg13g2_decap_8 FILLER_31_1589 ();
 sg13g2_decap_8 FILLER_31_1596 ();
 sg13g2_decap_8 FILLER_31_1603 ();
 sg13g2_decap_8 FILLER_31_1610 ();
 sg13g2_decap_8 FILLER_31_1617 ();
 sg13g2_decap_8 FILLER_31_1624 ();
 sg13g2_decap_8 FILLER_31_1631 ();
 sg13g2_decap_8 FILLER_31_1638 ();
 sg13g2_decap_8 FILLER_31_1645 ();
 sg13g2_decap_8 FILLER_31_1652 ();
 sg13g2_decap_8 FILLER_31_1659 ();
 sg13g2_decap_8 FILLER_31_1666 ();
 sg13g2_decap_8 FILLER_31_1673 ();
 sg13g2_decap_8 FILLER_31_1680 ();
 sg13g2_decap_8 FILLER_31_1687 ();
 sg13g2_decap_8 FILLER_31_1694 ();
 sg13g2_decap_8 FILLER_31_1701 ();
 sg13g2_decap_8 FILLER_31_1708 ();
 sg13g2_decap_8 FILLER_31_1715 ();
 sg13g2_decap_8 FILLER_31_1722 ();
 sg13g2_decap_8 FILLER_31_1729 ();
 sg13g2_decap_8 FILLER_31_1736 ();
 sg13g2_decap_8 FILLER_31_1743 ();
 sg13g2_decap_8 FILLER_31_1750 ();
 sg13g2_decap_8 FILLER_31_1757 ();
 sg13g2_decap_4 FILLER_31_1764 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_32 ();
 sg13g2_fill_1 FILLER_32_78 ();
 sg13g2_fill_2 FILLER_32_123 ();
 sg13g2_fill_1 FILLER_32_125 ();
 sg13g2_fill_2 FILLER_32_136 ();
 sg13g2_decap_8 FILLER_32_143 ();
 sg13g2_decap_8 FILLER_32_150 ();
 sg13g2_fill_2 FILLER_32_157 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_175 ();
 sg13g2_fill_1 FILLER_32_177 ();
 sg13g2_decap_8 FILLER_32_183 ();
 sg13g2_fill_2 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_240 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_decap_4 FILLER_32_298 ();
 sg13g2_fill_2 FILLER_32_302 ();
 sg13g2_fill_2 FILLER_32_314 ();
 sg13g2_decap_4 FILLER_32_331 ();
 sg13g2_fill_2 FILLER_32_361 ();
 sg13g2_fill_1 FILLER_32_363 ();
 sg13g2_fill_1 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_428 ();
 sg13g2_fill_1 FILLER_32_435 ();
 sg13g2_decap_4 FILLER_32_466 ();
 sg13g2_fill_2 FILLER_32_535 ();
 sg13g2_fill_1 FILLER_32_549 ();
 sg13g2_fill_1 FILLER_32_566 ();
 sg13g2_fill_1 FILLER_32_579 ();
 sg13g2_fill_2 FILLER_32_585 ();
 sg13g2_fill_1 FILLER_32_587 ();
 sg13g2_fill_1 FILLER_32_607 ();
 sg13g2_fill_1 FILLER_32_640 ();
 sg13g2_decap_8 FILLER_32_679 ();
 sg13g2_decap_8 FILLER_32_686 ();
 sg13g2_decap_8 FILLER_32_783 ();
 sg13g2_decap_4 FILLER_32_790 ();
 sg13g2_fill_2 FILLER_32_794 ();
 sg13g2_fill_1 FILLER_32_817 ();
 sg13g2_fill_2 FILLER_32_832 ();
 sg13g2_fill_1 FILLER_32_850 ();
 sg13g2_decap_8 FILLER_32_870 ();
 sg13g2_fill_2 FILLER_32_877 ();
 sg13g2_fill_2 FILLER_32_903 ();
 sg13g2_fill_1 FILLER_32_905 ();
 sg13g2_decap_4 FILLER_32_911 ();
 sg13g2_decap_4 FILLER_32_920 ();
 sg13g2_fill_2 FILLER_32_924 ();
 sg13g2_fill_1 FILLER_32_958 ();
 sg13g2_decap_8 FILLER_32_963 ();
 sg13g2_decap_8 FILLER_32_994 ();
 sg13g2_decap_8 FILLER_32_1001 ();
 sg13g2_decap_8 FILLER_32_1008 ();
 sg13g2_decap_8 FILLER_32_1015 ();
 sg13g2_decap_8 FILLER_32_1022 ();
 sg13g2_decap_8 FILLER_32_1029 ();
 sg13g2_decap_8 FILLER_32_1036 ();
 sg13g2_decap_8 FILLER_32_1043 ();
 sg13g2_decap_8 FILLER_32_1050 ();
 sg13g2_decap_8 FILLER_32_1057 ();
 sg13g2_decap_8 FILLER_32_1064 ();
 sg13g2_decap_8 FILLER_32_1071 ();
 sg13g2_decap_8 FILLER_32_1078 ();
 sg13g2_decap_8 FILLER_32_1085 ();
 sg13g2_decap_8 FILLER_32_1092 ();
 sg13g2_decap_8 FILLER_32_1099 ();
 sg13g2_decap_8 FILLER_32_1106 ();
 sg13g2_decap_8 FILLER_32_1113 ();
 sg13g2_decap_8 FILLER_32_1120 ();
 sg13g2_decap_8 FILLER_32_1127 ();
 sg13g2_decap_8 FILLER_32_1134 ();
 sg13g2_decap_8 FILLER_32_1141 ();
 sg13g2_decap_8 FILLER_32_1148 ();
 sg13g2_decap_8 FILLER_32_1155 ();
 sg13g2_decap_8 FILLER_32_1162 ();
 sg13g2_decap_8 FILLER_32_1169 ();
 sg13g2_decap_8 FILLER_32_1176 ();
 sg13g2_decap_8 FILLER_32_1183 ();
 sg13g2_decap_8 FILLER_32_1190 ();
 sg13g2_decap_8 FILLER_32_1197 ();
 sg13g2_decap_8 FILLER_32_1204 ();
 sg13g2_decap_8 FILLER_32_1211 ();
 sg13g2_decap_8 FILLER_32_1218 ();
 sg13g2_decap_8 FILLER_32_1225 ();
 sg13g2_decap_8 FILLER_32_1232 ();
 sg13g2_decap_8 FILLER_32_1239 ();
 sg13g2_decap_8 FILLER_32_1246 ();
 sg13g2_decap_8 FILLER_32_1253 ();
 sg13g2_decap_8 FILLER_32_1260 ();
 sg13g2_decap_8 FILLER_32_1267 ();
 sg13g2_decap_8 FILLER_32_1274 ();
 sg13g2_decap_8 FILLER_32_1281 ();
 sg13g2_decap_8 FILLER_32_1288 ();
 sg13g2_decap_8 FILLER_32_1295 ();
 sg13g2_decap_8 FILLER_32_1302 ();
 sg13g2_decap_8 FILLER_32_1309 ();
 sg13g2_decap_8 FILLER_32_1316 ();
 sg13g2_decap_8 FILLER_32_1323 ();
 sg13g2_decap_8 FILLER_32_1330 ();
 sg13g2_decap_8 FILLER_32_1337 ();
 sg13g2_decap_8 FILLER_32_1344 ();
 sg13g2_decap_8 FILLER_32_1351 ();
 sg13g2_decap_8 FILLER_32_1358 ();
 sg13g2_decap_8 FILLER_32_1365 ();
 sg13g2_decap_8 FILLER_32_1372 ();
 sg13g2_decap_8 FILLER_32_1379 ();
 sg13g2_decap_8 FILLER_32_1386 ();
 sg13g2_decap_8 FILLER_32_1393 ();
 sg13g2_decap_8 FILLER_32_1400 ();
 sg13g2_decap_8 FILLER_32_1407 ();
 sg13g2_decap_8 FILLER_32_1414 ();
 sg13g2_decap_8 FILLER_32_1421 ();
 sg13g2_decap_8 FILLER_32_1428 ();
 sg13g2_decap_8 FILLER_32_1435 ();
 sg13g2_decap_8 FILLER_32_1442 ();
 sg13g2_decap_8 FILLER_32_1449 ();
 sg13g2_decap_8 FILLER_32_1456 ();
 sg13g2_decap_8 FILLER_32_1463 ();
 sg13g2_decap_8 FILLER_32_1470 ();
 sg13g2_decap_8 FILLER_32_1477 ();
 sg13g2_decap_8 FILLER_32_1484 ();
 sg13g2_decap_8 FILLER_32_1491 ();
 sg13g2_decap_8 FILLER_32_1498 ();
 sg13g2_decap_8 FILLER_32_1505 ();
 sg13g2_decap_8 FILLER_32_1512 ();
 sg13g2_decap_8 FILLER_32_1519 ();
 sg13g2_decap_8 FILLER_32_1526 ();
 sg13g2_decap_8 FILLER_32_1533 ();
 sg13g2_decap_8 FILLER_32_1540 ();
 sg13g2_decap_8 FILLER_32_1547 ();
 sg13g2_decap_8 FILLER_32_1554 ();
 sg13g2_decap_8 FILLER_32_1561 ();
 sg13g2_decap_8 FILLER_32_1568 ();
 sg13g2_decap_8 FILLER_32_1575 ();
 sg13g2_decap_8 FILLER_32_1582 ();
 sg13g2_decap_8 FILLER_32_1589 ();
 sg13g2_decap_8 FILLER_32_1596 ();
 sg13g2_decap_8 FILLER_32_1603 ();
 sg13g2_decap_8 FILLER_32_1610 ();
 sg13g2_decap_8 FILLER_32_1617 ();
 sg13g2_decap_8 FILLER_32_1624 ();
 sg13g2_decap_8 FILLER_32_1631 ();
 sg13g2_decap_8 FILLER_32_1638 ();
 sg13g2_decap_8 FILLER_32_1645 ();
 sg13g2_decap_8 FILLER_32_1652 ();
 sg13g2_decap_8 FILLER_32_1659 ();
 sg13g2_decap_8 FILLER_32_1666 ();
 sg13g2_decap_8 FILLER_32_1673 ();
 sg13g2_decap_8 FILLER_32_1680 ();
 sg13g2_decap_8 FILLER_32_1687 ();
 sg13g2_decap_8 FILLER_32_1694 ();
 sg13g2_decap_8 FILLER_32_1701 ();
 sg13g2_decap_8 FILLER_32_1708 ();
 sg13g2_decap_8 FILLER_32_1715 ();
 sg13g2_decap_8 FILLER_32_1722 ();
 sg13g2_decap_8 FILLER_32_1729 ();
 sg13g2_decap_8 FILLER_32_1736 ();
 sg13g2_decap_8 FILLER_32_1743 ();
 sg13g2_decap_8 FILLER_32_1750 ();
 sg13g2_decap_8 FILLER_32_1757 ();
 sg13g2_decap_4 FILLER_32_1764 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_35 ();
 sg13g2_fill_1 FILLER_33_59 ();
 sg13g2_decap_4 FILLER_33_73 ();
 sg13g2_fill_2 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_83 ();
 sg13g2_decap_4 FILLER_33_94 ();
 sg13g2_fill_1 FILLER_33_98 ();
 sg13g2_decap_4 FILLER_33_130 ();
 sg13g2_fill_1 FILLER_33_149 ();
 sg13g2_fill_1 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_decap_4 FILLER_33_191 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_4 FILLER_33_210 ();
 sg13g2_fill_2 FILLER_33_214 ();
 sg13g2_fill_1 FILLER_33_228 ();
 sg13g2_fill_2 FILLER_33_234 ();
 sg13g2_decap_4 FILLER_33_244 ();
 sg13g2_fill_2 FILLER_33_262 ();
 sg13g2_fill_1 FILLER_33_278 ();
 sg13g2_decap_4 FILLER_33_324 ();
 sg13g2_fill_1 FILLER_33_328 ();
 sg13g2_fill_1 FILLER_33_348 ();
 sg13g2_fill_2 FILLER_33_358 ();
 sg13g2_fill_1 FILLER_33_360 ();
 sg13g2_fill_1 FILLER_33_370 ();
 sg13g2_fill_2 FILLER_33_411 ();
 sg13g2_fill_1 FILLER_33_469 ();
 sg13g2_fill_2 FILLER_33_488 ();
 sg13g2_fill_1 FILLER_33_490 ();
 sg13g2_fill_2 FILLER_33_502 ();
 sg13g2_fill_2 FILLER_33_509 ();
 sg13g2_fill_2 FILLER_33_515 ();
 sg13g2_decap_4 FILLER_33_578 ();
 sg13g2_fill_1 FILLER_33_582 ();
 sg13g2_fill_2 FILLER_33_596 ();
 sg13g2_decap_4 FILLER_33_606 ();
 sg13g2_fill_1 FILLER_33_610 ();
 sg13g2_fill_1 FILLER_33_616 ();
 sg13g2_fill_1 FILLER_33_620 ();
 sg13g2_decap_8 FILLER_33_626 ();
 sg13g2_fill_2 FILLER_33_633 ();
 sg13g2_decap_4 FILLER_33_655 ();
 sg13g2_fill_2 FILLER_33_659 ();
 sg13g2_fill_2 FILLER_33_675 ();
 sg13g2_fill_1 FILLER_33_677 ();
 sg13g2_fill_1 FILLER_33_694 ();
 sg13g2_fill_2 FILLER_33_707 ();
 sg13g2_fill_2 FILLER_33_724 ();
 sg13g2_decap_4 FILLER_33_754 ();
 sg13g2_fill_1 FILLER_33_794 ();
 sg13g2_fill_2 FILLER_33_812 ();
 sg13g2_decap_4 FILLER_33_834 ();
 sg13g2_fill_2 FILLER_33_838 ();
 sg13g2_decap_8 FILLER_33_845 ();
 sg13g2_decap_8 FILLER_33_852 ();
 sg13g2_decap_8 FILLER_33_859 ();
 sg13g2_decap_4 FILLER_33_866 ();
 sg13g2_fill_1 FILLER_33_870 ();
 sg13g2_fill_1 FILLER_33_882 ();
 sg13g2_fill_2 FILLER_33_891 ();
 sg13g2_decap_4 FILLER_33_900 ();
 sg13g2_fill_1 FILLER_33_904 ();
 sg13g2_decap_8 FILLER_33_925 ();
 sg13g2_fill_2 FILLER_33_937 ();
 sg13g2_fill_2 FILLER_33_943 ();
 sg13g2_fill_1 FILLER_33_945 ();
 sg13g2_fill_2 FILLER_33_964 ();
 sg13g2_fill_1 FILLER_33_966 ();
 sg13g2_decap_8 FILLER_33_993 ();
 sg13g2_decap_8 FILLER_33_1000 ();
 sg13g2_decap_8 FILLER_33_1007 ();
 sg13g2_decap_8 FILLER_33_1014 ();
 sg13g2_decap_8 FILLER_33_1021 ();
 sg13g2_decap_8 FILLER_33_1028 ();
 sg13g2_decap_8 FILLER_33_1035 ();
 sg13g2_decap_8 FILLER_33_1042 ();
 sg13g2_decap_8 FILLER_33_1049 ();
 sg13g2_decap_8 FILLER_33_1056 ();
 sg13g2_decap_8 FILLER_33_1063 ();
 sg13g2_decap_8 FILLER_33_1070 ();
 sg13g2_decap_8 FILLER_33_1077 ();
 sg13g2_decap_8 FILLER_33_1084 ();
 sg13g2_decap_8 FILLER_33_1091 ();
 sg13g2_decap_8 FILLER_33_1098 ();
 sg13g2_decap_8 FILLER_33_1105 ();
 sg13g2_decap_8 FILLER_33_1112 ();
 sg13g2_decap_8 FILLER_33_1119 ();
 sg13g2_decap_8 FILLER_33_1126 ();
 sg13g2_decap_8 FILLER_33_1133 ();
 sg13g2_decap_8 FILLER_33_1140 ();
 sg13g2_decap_8 FILLER_33_1147 ();
 sg13g2_decap_8 FILLER_33_1154 ();
 sg13g2_decap_8 FILLER_33_1161 ();
 sg13g2_decap_8 FILLER_33_1168 ();
 sg13g2_decap_8 FILLER_33_1175 ();
 sg13g2_decap_8 FILLER_33_1182 ();
 sg13g2_decap_8 FILLER_33_1189 ();
 sg13g2_decap_8 FILLER_33_1196 ();
 sg13g2_decap_8 FILLER_33_1203 ();
 sg13g2_decap_8 FILLER_33_1210 ();
 sg13g2_decap_8 FILLER_33_1217 ();
 sg13g2_decap_8 FILLER_33_1224 ();
 sg13g2_decap_8 FILLER_33_1231 ();
 sg13g2_decap_8 FILLER_33_1238 ();
 sg13g2_decap_8 FILLER_33_1245 ();
 sg13g2_decap_8 FILLER_33_1252 ();
 sg13g2_decap_8 FILLER_33_1259 ();
 sg13g2_decap_8 FILLER_33_1266 ();
 sg13g2_decap_8 FILLER_33_1273 ();
 sg13g2_decap_8 FILLER_33_1280 ();
 sg13g2_decap_8 FILLER_33_1287 ();
 sg13g2_decap_8 FILLER_33_1294 ();
 sg13g2_decap_8 FILLER_33_1301 ();
 sg13g2_decap_8 FILLER_33_1308 ();
 sg13g2_decap_8 FILLER_33_1315 ();
 sg13g2_decap_8 FILLER_33_1322 ();
 sg13g2_decap_8 FILLER_33_1329 ();
 sg13g2_decap_8 FILLER_33_1336 ();
 sg13g2_decap_8 FILLER_33_1343 ();
 sg13g2_decap_8 FILLER_33_1350 ();
 sg13g2_decap_8 FILLER_33_1357 ();
 sg13g2_decap_8 FILLER_33_1364 ();
 sg13g2_decap_8 FILLER_33_1371 ();
 sg13g2_decap_8 FILLER_33_1378 ();
 sg13g2_decap_8 FILLER_33_1385 ();
 sg13g2_decap_8 FILLER_33_1392 ();
 sg13g2_decap_8 FILLER_33_1399 ();
 sg13g2_decap_8 FILLER_33_1406 ();
 sg13g2_decap_8 FILLER_33_1413 ();
 sg13g2_decap_8 FILLER_33_1420 ();
 sg13g2_decap_8 FILLER_33_1427 ();
 sg13g2_decap_8 FILLER_33_1434 ();
 sg13g2_decap_8 FILLER_33_1441 ();
 sg13g2_decap_8 FILLER_33_1448 ();
 sg13g2_decap_8 FILLER_33_1455 ();
 sg13g2_decap_8 FILLER_33_1462 ();
 sg13g2_decap_8 FILLER_33_1469 ();
 sg13g2_decap_8 FILLER_33_1476 ();
 sg13g2_decap_8 FILLER_33_1483 ();
 sg13g2_decap_8 FILLER_33_1490 ();
 sg13g2_decap_8 FILLER_33_1497 ();
 sg13g2_decap_8 FILLER_33_1504 ();
 sg13g2_decap_8 FILLER_33_1511 ();
 sg13g2_decap_8 FILLER_33_1518 ();
 sg13g2_decap_8 FILLER_33_1525 ();
 sg13g2_decap_8 FILLER_33_1532 ();
 sg13g2_decap_8 FILLER_33_1539 ();
 sg13g2_decap_8 FILLER_33_1546 ();
 sg13g2_decap_8 FILLER_33_1553 ();
 sg13g2_decap_8 FILLER_33_1560 ();
 sg13g2_decap_8 FILLER_33_1567 ();
 sg13g2_decap_8 FILLER_33_1574 ();
 sg13g2_decap_8 FILLER_33_1581 ();
 sg13g2_decap_8 FILLER_33_1588 ();
 sg13g2_decap_8 FILLER_33_1595 ();
 sg13g2_decap_8 FILLER_33_1602 ();
 sg13g2_decap_8 FILLER_33_1609 ();
 sg13g2_decap_8 FILLER_33_1616 ();
 sg13g2_decap_8 FILLER_33_1623 ();
 sg13g2_decap_8 FILLER_33_1630 ();
 sg13g2_decap_8 FILLER_33_1637 ();
 sg13g2_decap_8 FILLER_33_1644 ();
 sg13g2_decap_8 FILLER_33_1651 ();
 sg13g2_decap_8 FILLER_33_1658 ();
 sg13g2_decap_8 FILLER_33_1665 ();
 sg13g2_decap_8 FILLER_33_1672 ();
 sg13g2_decap_8 FILLER_33_1679 ();
 sg13g2_decap_8 FILLER_33_1686 ();
 sg13g2_decap_8 FILLER_33_1693 ();
 sg13g2_decap_8 FILLER_33_1700 ();
 sg13g2_decap_8 FILLER_33_1707 ();
 sg13g2_decap_8 FILLER_33_1714 ();
 sg13g2_decap_8 FILLER_33_1721 ();
 sg13g2_decap_8 FILLER_33_1728 ();
 sg13g2_decap_8 FILLER_33_1735 ();
 sg13g2_decap_8 FILLER_33_1742 ();
 sg13g2_decap_8 FILLER_33_1749 ();
 sg13g2_decap_8 FILLER_33_1756 ();
 sg13g2_decap_4 FILLER_33_1763 ();
 sg13g2_fill_1 FILLER_33_1767 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_4 FILLER_34_103 ();
 sg13g2_fill_2 FILLER_34_107 ();
 sg13g2_fill_2 FILLER_34_127 ();
 sg13g2_fill_2 FILLER_34_133 ();
 sg13g2_fill_1 FILLER_34_135 ();
 sg13g2_decap_8 FILLER_34_148 ();
 sg13g2_fill_2 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_166 ();
 sg13g2_fill_1 FILLER_34_175 ();
 sg13g2_decap_4 FILLER_34_192 ();
 sg13g2_fill_2 FILLER_34_206 ();
 sg13g2_fill_2 FILLER_34_221 ();
 sg13g2_decap_4 FILLER_34_249 ();
 sg13g2_fill_1 FILLER_34_253 ();
 sg13g2_fill_2 FILLER_34_289 ();
 sg13g2_fill_1 FILLER_34_291 ();
 sg13g2_fill_2 FILLER_34_333 ();
 sg13g2_fill_2 FILLER_34_387 ();
 sg13g2_fill_2 FILLER_34_429 ();
 sg13g2_fill_1 FILLER_34_431 ();
 sg13g2_fill_1 FILLER_34_441 ();
 sg13g2_fill_2 FILLER_34_473 ();
 sg13g2_fill_2 FILLER_34_501 ();
 sg13g2_fill_2 FILLER_34_567 ();
 sg13g2_fill_1 FILLER_34_569 ();
 sg13g2_decap_4 FILLER_34_578 ();
 sg13g2_fill_2 FILLER_34_582 ();
 sg13g2_decap_4 FILLER_34_588 ();
 sg13g2_decap_8 FILLER_34_605 ();
 sg13g2_fill_2 FILLER_34_631 ();
 sg13g2_decap_4 FILLER_34_651 ();
 sg13g2_fill_2 FILLER_34_655 ();
 sg13g2_fill_1 FILLER_34_662 ();
 sg13g2_fill_1 FILLER_34_709 ();
 sg13g2_fill_1 FILLER_34_762 ();
 sg13g2_fill_1 FILLER_34_768 ();
 sg13g2_fill_2 FILLER_34_801 ();
 sg13g2_fill_1 FILLER_34_803 ();
 sg13g2_fill_2 FILLER_34_814 ();
 sg13g2_fill_1 FILLER_34_816 ();
 sg13g2_decap_4 FILLER_34_827 ();
 sg13g2_fill_2 FILLER_34_849 ();
 sg13g2_fill_1 FILLER_34_851 ();
 sg13g2_decap_4 FILLER_34_880 ();
 sg13g2_fill_2 FILLER_34_884 ();
 sg13g2_fill_2 FILLER_34_896 ();
 sg13g2_fill_2 FILLER_34_902 ();
 sg13g2_fill_1 FILLER_34_913 ();
 sg13g2_decap_8 FILLER_34_927 ();
 sg13g2_fill_1 FILLER_34_934 ();
 sg13g2_fill_2 FILLER_34_949 ();
 sg13g2_fill_1 FILLER_34_956 ();
 sg13g2_decap_8 FILLER_34_961 ();
 sg13g2_decap_8 FILLER_34_968 ();
 sg13g2_fill_1 FILLER_34_975 ();
 sg13g2_decap_8 FILLER_34_985 ();
 sg13g2_decap_8 FILLER_34_992 ();
 sg13g2_decap_8 FILLER_34_999 ();
 sg13g2_decap_8 FILLER_34_1006 ();
 sg13g2_decap_8 FILLER_34_1013 ();
 sg13g2_decap_8 FILLER_34_1020 ();
 sg13g2_decap_8 FILLER_34_1027 ();
 sg13g2_decap_8 FILLER_34_1034 ();
 sg13g2_decap_8 FILLER_34_1041 ();
 sg13g2_decap_8 FILLER_34_1048 ();
 sg13g2_decap_8 FILLER_34_1055 ();
 sg13g2_decap_8 FILLER_34_1062 ();
 sg13g2_decap_8 FILLER_34_1069 ();
 sg13g2_decap_8 FILLER_34_1076 ();
 sg13g2_decap_8 FILLER_34_1083 ();
 sg13g2_decap_8 FILLER_34_1090 ();
 sg13g2_decap_8 FILLER_34_1097 ();
 sg13g2_decap_8 FILLER_34_1104 ();
 sg13g2_decap_8 FILLER_34_1111 ();
 sg13g2_decap_8 FILLER_34_1118 ();
 sg13g2_decap_8 FILLER_34_1125 ();
 sg13g2_decap_8 FILLER_34_1132 ();
 sg13g2_decap_8 FILLER_34_1139 ();
 sg13g2_decap_8 FILLER_34_1146 ();
 sg13g2_decap_8 FILLER_34_1153 ();
 sg13g2_decap_8 FILLER_34_1160 ();
 sg13g2_decap_8 FILLER_34_1167 ();
 sg13g2_decap_8 FILLER_34_1174 ();
 sg13g2_decap_8 FILLER_34_1181 ();
 sg13g2_decap_8 FILLER_34_1188 ();
 sg13g2_decap_8 FILLER_34_1195 ();
 sg13g2_decap_8 FILLER_34_1202 ();
 sg13g2_decap_8 FILLER_34_1209 ();
 sg13g2_decap_8 FILLER_34_1216 ();
 sg13g2_decap_8 FILLER_34_1223 ();
 sg13g2_decap_8 FILLER_34_1230 ();
 sg13g2_decap_8 FILLER_34_1237 ();
 sg13g2_decap_8 FILLER_34_1244 ();
 sg13g2_decap_8 FILLER_34_1251 ();
 sg13g2_decap_8 FILLER_34_1258 ();
 sg13g2_decap_8 FILLER_34_1265 ();
 sg13g2_decap_8 FILLER_34_1272 ();
 sg13g2_decap_8 FILLER_34_1279 ();
 sg13g2_decap_8 FILLER_34_1286 ();
 sg13g2_decap_8 FILLER_34_1293 ();
 sg13g2_decap_8 FILLER_34_1300 ();
 sg13g2_decap_8 FILLER_34_1307 ();
 sg13g2_decap_8 FILLER_34_1314 ();
 sg13g2_decap_8 FILLER_34_1321 ();
 sg13g2_decap_8 FILLER_34_1328 ();
 sg13g2_decap_8 FILLER_34_1335 ();
 sg13g2_decap_8 FILLER_34_1342 ();
 sg13g2_decap_8 FILLER_34_1349 ();
 sg13g2_decap_8 FILLER_34_1356 ();
 sg13g2_decap_8 FILLER_34_1363 ();
 sg13g2_decap_8 FILLER_34_1370 ();
 sg13g2_decap_8 FILLER_34_1377 ();
 sg13g2_decap_8 FILLER_34_1384 ();
 sg13g2_decap_8 FILLER_34_1391 ();
 sg13g2_decap_8 FILLER_34_1398 ();
 sg13g2_decap_8 FILLER_34_1405 ();
 sg13g2_decap_8 FILLER_34_1412 ();
 sg13g2_decap_8 FILLER_34_1419 ();
 sg13g2_decap_8 FILLER_34_1426 ();
 sg13g2_decap_8 FILLER_34_1433 ();
 sg13g2_decap_8 FILLER_34_1440 ();
 sg13g2_decap_8 FILLER_34_1447 ();
 sg13g2_decap_8 FILLER_34_1454 ();
 sg13g2_decap_8 FILLER_34_1461 ();
 sg13g2_decap_8 FILLER_34_1468 ();
 sg13g2_decap_8 FILLER_34_1475 ();
 sg13g2_decap_8 FILLER_34_1482 ();
 sg13g2_decap_8 FILLER_34_1489 ();
 sg13g2_decap_8 FILLER_34_1496 ();
 sg13g2_decap_8 FILLER_34_1503 ();
 sg13g2_decap_8 FILLER_34_1510 ();
 sg13g2_decap_8 FILLER_34_1517 ();
 sg13g2_decap_8 FILLER_34_1524 ();
 sg13g2_decap_8 FILLER_34_1531 ();
 sg13g2_decap_8 FILLER_34_1538 ();
 sg13g2_decap_8 FILLER_34_1545 ();
 sg13g2_decap_8 FILLER_34_1552 ();
 sg13g2_decap_8 FILLER_34_1559 ();
 sg13g2_decap_8 FILLER_34_1566 ();
 sg13g2_decap_8 FILLER_34_1573 ();
 sg13g2_decap_8 FILLER_34_1580 ();
 sg13g2_decap_8 FILLER_34_1587 ();
 sg13g2_decap_8 FILLER_34_1594 ();
 sg13g2_decap_8 FILLER_34_1601 ();
 sg13g2_decap_8 FILLER_34_1608 ();
 sg13g2_decap_8 FILLER_34_1615 ();
 sg13g2_decap_8 FILLER_34_1622 ();
 sg13g2_decap_8 FILLER_34_1629 ();
 sg13g2_decap_8 FILLER_34_1636 ();
 sg13g2_decap_8 FILLER_34_1643 ();
 sg13g2_decap_8 FILLER_34_1650 ();
 sg13g2_decap_8 FILLER_34_1657 ();
 sg13g2_decap_8 FILLER_34_1664 ();
 sg13g2_decap_8 FILLER_34_1671 ();
 sg13g2_decap_8 FILLER_34_1678 ();
 sg13g2_decap_8 FILLER_34_1685 ();
 sg13g2_decap_8 FILLER_34_1692 ();
 sg13g2_decap_8 FILLER_34_1699 ();
 sg13g2_decap_8 FILLER_34_1706 ();
 sg13g2_decap_8 FILLER_34_1713 ();
 sg13g2_decap_8 FILLER_34_1720 ();
 sg13g2_decap_8 FILLER_34_1727 ();
 sg13g2_decap_8 FILLER_34_1734 ();
 sg13g2_decap_8 FILLER_34_1741 ();
 sg13g2_decap_8 FILLER_34_1748 ();
 sg13g2_decap_8 FILLER_34_1755 ();
 sg13g2_decap_4 FILLER_34_1762 ();
 sg13g2_fill_2 FILLER_34_1766 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_4 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_53 ();
 sg13g2_decap_8 FILLER_35_58 ();
 sg13g2_fill_2 FILLER_35_65 ();
 sg13g2_fill_1 FILLER_35_67 ();
 sg13g2_decap_4 FILLER_35_77 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_130 ();
 sg13g2_fill_1 FILLER_35_132 ();
 sg13g2_fill_1 FILLER_35_146 ();
 sg13g2_fill_2 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_fill_2 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_223 ();
 sg13g2_decap_4 FILLER_35_230 ();
 sg13g2_fill_2 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_fill_2 FILLER_35_265 ();
 sg13g2_fill_1 FILLER_35_277 ();
 sg13g2_fill_2 FILLER_35_304 ();
 sg13g2_fill_1 FILLER_35_306 ();
 sg13g2_fill_2 FILLER_35_333 ();
 sg13g2_fill_1 FILLER_35_335 ();
 sg13g2_fill_2 FILLER_35_377 ();
 sg13g2_decap_4 FILLER_35_389 ();
 sg13g2_fill_2 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_fill_1 FILLER_35_504 ();
 sg13g2_fill_1 FILLER_35_510 ();
 sg13g2_fill_2 FILLER_35_525 ();
 sg13g2_fill_1 FILLER_35_565 ();
 sg13g2_fill_2 FILLER_35_585 ();
 sg13g2_fill_2 FILLER_35_596 ();
 sg13g2_fill_2 FILLER_35_612 ();
 sg13g2_fill_1 FILLER_35_614 ();
 sg13g2_decap_4 FILLER_35_630 ();
 sg13g2_decap_8 FILLER_35_668 ();
 sg13g2_decap_4 FILLER_35_675 ();
 sg13g2_fill_1 FILLER_35_688 ();
 sg13g2_fill_2 FILLER_35_697 ();
 sg13g2_fill_1 FILLER_35_736 ();
 sg13g2_decap_4 FILLER_35_753 ();
 sg13g2_fill_2 FILLER_35_757 ();
 sg13g2_fill_2 FILLER_35_765 ();
 sg13g2_fill_1 FILLER_35_767 ();
 sg13g2_decap_8 FILLER_35_779 ();
 sg13g2_decap_8 FILLER_35_786 ();
 sg13g2_fill_2 FILLER_35_793 ();
 sg13g2_decap_8 FILLER_35_811 ();
 sg13g2_decap_4 FILLER_35_818 ();
 sg13g2_fill_1 FILLER_35_822 ();
 sg13g2_decap_8 FILLER_35_833 ();
 sg13g2_fill_1 FILLER_35_845 ();
 sg13g2_decap_4 FILLER_35_866 ();
 sg13g2_fill_2 FILLER_35_901 ();
 sg13g2_fill_1 FILLER_35_903 ();
 sg13g2_decap_8 FILLER_35_922 ();
 sg13g2_decap_8 FILLER_35_941 ();
 sg13g2_decap_8 FILLER_35_948 ();
 sg13g2_decap_8 FILLER_35_955 ();
 sg13g2_decap_8 FILLER_35_962 ();
 sg13g2_decap_8 FILLER_35_969 ();
 sg13g2_decap_8 FILLER_35_976 ();
 sg13g2_decap_8 FILLER_35_983 ();
 sg13g2_decap_8 FILLER_35_990 ();
 sg13g2_decap_8 FILLER_35_997 ();
 sg13g2_decap_8 FILLER_35_1004 ();
 sg13g2_decap_8 FILLER_35_1011 ();
 sg13g2_decap_8 FILLER_35_1018 ();
 sg13g2_decap_8 FILLER_35_1025 ();
 sg13g2_decap_8 FILLER_35_1032 ();
 sg13g2_decap_8 FILLER_35_1039 ();
 sg13g2_decap_8 FILLER_35_1046 ();
 sg13g2_decap_8 FILLER_35_1053 ();
 sg13g2_decap_8 FILLER_35_1060 ();
 sg13g2_decap_8 FILLER_35_1067 ();
 sg13g2_decap_8 FILLER_35_1074 ();
 sg13g2_decap_8 FILLER_35_1081 ();
 sg13g2_decap_8 FILLER_35_1088 ();
 sg13g2_decap_8 FILLER_35_1095 ();
 sg13g2_decap_8 FILLER_35_1102 ();
 sg13g2_decap_8 FILLER_35_1109 ();
 sg13g2_decap_8 FILLER_35_1116 ();
 sg13g2_decap_8 FILLER_35_1123 ();
 sg13g2_decap_8 FILLER_35_1130 ();
 sg13g2_decap_8 FILLER_35_1137 ();
 sg13g2_decap_8 FILLER_35_1144 ();
 sg13g2_decap_8 FILLER_35_1151 ();
 sg13g2_decap_8 FILLER_35_1158 ();
 sg13g2_decap_8 FILLER_35_1165 ();
 sg13g2_decap_8 FILLER_35_1172 ();
 sg13g2_decap_8 FILLER_35_1179 ();
 sg13g2_decap_8 FILLER_35_1186 ();
 sg13g2_decap_8 FILLER_35_1193 ();
 sg13g2_decap_8 FILLER_35_1200 ();
 sg13g2_decap_8 FILLER_35_1207 ();
 sg13g2_decap_8 FILLER_35_1214 ();
 sg13g2_decap_8 FILLER_35_1221 ();
 sg13g2_decap_8 FILLER_35_1228 ();
 sg13g2_decap_8 FILLER_35_1235 ();
 sg13g2_decap_8 FILLER_35_1242 ();
 sg13g2_decap_8 FILLER_35_1249 ();
 sg13g2_decap_8 FILLER_35_1256 ();
 sg13g2_decap_8 FILLER_35_1263 ();
 sg13g2_decap_8 FILLER_35_1270 ();
 sg13g2_decap_8 FILLER_35_1277 ();
 sg13g2_decap_8 FILLER_35_1284 ();
 sg13g2_decap_8 FILLER_35_1291 ();
 sg13g2_decap_8 FILLER_35_1298 ();
 sg13g2_decap_8 FILLER_35_1305 ();
 sg13g2_decap_8 FILLER_35_1312 ();
 sg13g2_decap_8 FILLER_35_1319 ();
 sg13g2_decap_8 FILLER_35_1326 ();
 sg13g2_decap_8 FILLER_35_1333 ();
 sg13g2_decap_8 FILLER_35_1340 ();
 sg13g2_decap_8 FILLER_35_1347 ();
 sg13g2_decap_8 FILLER_35_1354 ();
 sg13g2_decap_8 FILLER_35_1361 ();
 sg13g2_decap_8 FILLER_35_1368 ();
 sg13g2_decap_8 FILLER_35_1375 ();
 sg13g2_decap_8 FILLER_35_1382 ();
 sg13g2_decap_8 FILLER_35_1389 ();
 sg13g2_decap_8 FILLER_35_1396 ();
 sg13g2_decap_8 FILLER_35_1403 ();
 sg13g2_decap_8 FILLER_35_1410 ();
 sg13g2_decap_8 FILLER_35_1417 ();
 sg13g2_decap_8 FILLER_35_1424 ();
 sg13g2_decap_8 FILLER_35_1431 ();
 sg13g2_decap_8 FILLER_35_1438 ();
 sg13g2_decap_8 FILLER_35_1445 ();
 sg13g2_decap_8 FILLER_35_1452 ();
 sg13g2_decap_8 FILLER_35_1459 ();
 sg13g2_decap_8 FILLER_35_1466 ();
 sg13g2_decap_8 FILLER_35_1473 ();
 sg13g2_decap_8 FILLER_35_1480 ();
 sg13g2_decap_8 FILLER_35_1487 ();
 sg13g2_decap_8 FILLER_35_1494 ();
 sg13g2_decap_8 FILLER_35_1501 ();
 sg13g2_decap_8 FILLER_35_1508 ();
 sg13g2_decap_8 FILLER_35_1515 ();
 sg13g2_decap_8 FILLER_35_1522 ();
 sg13g2_decap_8 FILLER_35_1529 ();
 sg13g2_decap_8 FILLER_35_1536 ();
 sg13g2_decap_8 FILLER_35_1543 ();
 sg13g2_decap_8 FILLER_35_1550 ();
 sg13g2_decap_8 FILLER_35_1557 ();
 sg13g2_decap_8 FILLER_35_1564 ();
 sg13g2_decap_8 FILLER_35_1571 ();
 sg13g2_decap_8 FILLER_35_1578 ();
 sg13g2_decap_8 FILLER_35_1585 ();
 sg13g2_decap_8 FILLER_35_1592 ();
 sg13g2_decap_8 FILLER_35_1599 ();
 sg13g2_decap_8 FILLER_35_1606 ();
 sg13g2_decap_8 FILLER_35_1613 ();
 sg13g2_decap_8 FILLER_35_1620 ();
 sg13g2_decap_8 FILLER_35_1627 ();
 sg13g2_decap_8 FILLER_35_1634 ();
 sg13g2_decap_8 FILLER_35_1641 ();
 sg13g2_decap_8 FILLER_35_1648 ();
 sg13g2_decap_8 FILLER_35_1655 ();
 sg13g2_decap_8 FILLER_35_1662 ();
 sg13g2_decap_8 FILLER_35_1669 ();
 sg13g2_decap_8 FILLER_35_1676 ();
 sg13g2_decap_8 FILLER_35_1683 ();
 sg13g2_decap_8 FILLER_35_1690 ();
 sg13g2_decap_8 FILLER_35_1697 ();
 sg13g2_decap_8 FILLER_35_1704 ();
 sg13g2_decap_8 FILLER_35_1711 ();
 sg13g2_decap_8 FILLER_35_1718 ();
 sg13g2_decap_8 FILLER_35_1725 ();
 sg13g2_decap_8 FILLER_35_1732 ();
 sg13g2_decap_8 FILLER_35_1739 ();
 sg13g2_decap_8 FILLER_35_1746 ();
 sg13g2_decap_8 FILLER_35_1753 ();
 sg13g2_decap_8 FILLER_35_1760 ();
 sg13g2_fill_1 FILLER_35_1767 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_4 FILLER_36_49 ();
 sg13g2_decap_4 FILLER_36_87 ();
 sg13g2_fill_1 FILLER_36_91 ();
 sg13g2_fill_2 FILLER_36_118 ();
 sg13g2_fill_1 FILLER_36_120 ();
 sg13g2_fill_1 FILLER_36_135 ();
 sg13g2_fill_2 FILLER_36_141 ();
 sg13g2_fill_2 FILLER_36_174 ();
 sg13g2_fill_2 FILLER_36_189 ();
 sg13g2_fill_1 FILLER_36_191 ();
 sg13g2_decap_8 FILLER_36_202 ();
 sg13g2_fill_2 FILLER_36_209 ();
 sg13g2_decap_8 FILLER_36_236 ();
 sg13g2_fill_1 FILLER_36_243 ();
 sg13g2_fill_2 FILLER_36_253 ();
 sg13g2_decap_8 FILLER_36_271 ();
 sg13g2_fill_2 FILLER_36_278 ();
 sg13g2_decap_4 FILLER_36_284 ();
 sg13g2_decap_8 FILLER_36_292 ();
 sg13g2_decap_4 FILLER_36_299 ();
 sg13g2_fill_2 FILLER_36_303 ();
 sg13g2_fill_2 FILLER_36_318 ();
 sg13g2_fill_1 FILLER_36_320 ();
 sg13g2_fill_2 FILLER_36_330 ();
 sg13g2_fill_1 FILLER_36_332 ();
 sg13g2_fill_2 FILLER_36_344 ();
 sg13g2_decap_4 FILLER_36_377 ();
 sg13g2_decap_4 FILLER_36_428 ();
 sg13g2_fill_2 FILLER_36_441 ();
 sg13g2_fill_1 FILLER_36_443 ();
 sg13g2_fill_1 FILLER_36_454 ();
 sg13g2_fill_1 FILLER_36_501 ();
 sg13g2_fill_1 FILLER_36_573 ();
 sg13g2_fill_2 FILLER_36_600 ();
 sg13g2_fill_1 FILLER_36_602 ();
 sg13g2_decap_4 FILLER_36_607 ();
 sg13g2_fill_2 FILLER_36_611 ();
 sg13g2_decap_8 FILLER_36_634 ();
 sg13g2_decap_4 FILLER_36_641 ();
 sg13g2_decap_8 FILLER_36_649 ();
 sg13g2_decap_4 FILLER_36_666 ();
 sg13g2_fill_1 FILLER_36_670 ();
 sg13g2_fill_1 FILLER_36_677 ();
 sg13g2_fill_2 FILLER_36_684 ();
 sg13g2_fill_1 FILLER_36_686 ();
 sg13g2_decap_4 FILLER_36_748 ();
 sg13g2_fill_2 FILLER_36_809 ();
 sg13g2_fill_1 FILLER_36_811 ();
 sg13g2_fill_1 FILLER_36_832 ();
 sg13g2_fill_1 FILLER_36_838 ();
 sg13g2_fill_2 FILLER_36_849 ();
 sg13g2_decap_8 FILLER_36_862 ();
 sg13g2_decap_8 FILLER_36_869 ();
 sg13g2_decap_4 FILLER_36_881 ();
 sg13g2_decap_4 FILLER_36_891 ();
 sg13g2_fill_1 FILLER_36_895 ();
 sg13g2_fill_2 FILLER_36_901 ();
 sg13g2_decap_4 FILLER_36_912 ();
 sg13g2_fill_2 FILLER_36_916 ();
 sg13g2_decap_8 FILLER_36_933 ();
 sg13g2_decap_8 FILLER_36_940 ();
 sg13g2_decap_8 FILLER_36_947 ();
 sg13g2_decap_8 FILLER_36_954 ();
 sg13g2_decap_8 FILLER_36_961 ();
 sg13g2_decap_8 FILLER_36_968 ();
 sg13g2_decap_8 FILLER_36_975 ();
 sg13g2_decap_8 FILLER_36_982 ();
 sg13g2_decap_8 FILLER_36_989 ();
 sg13g2_decap_8 FILLER_36_996 ();
 sg13g2_decap_8 FILLER_36_1003 ();
 sg13g2_decap_8 FILLER_36_1010 ();
 sg13g2_decap_8 FILLER_36_1017 ();
 sg13g2_decap_8 FILLER_36_1024 ();
 sg13g2_decap_8 FILLER_36_1031 ();
 sg13g2_decap_8 FILLER_36_1038 ();
 sg13g2_decap_8 FILLER_36_1045 ();
 sg13g2_decap_8 FILLER_36_1052 ();
 sg13g2_decap_8 FILLER_36_1059 ();
 sg13g2_decap_8 FILLER_36_1066 ();
 sg13g2_decap_8 FILLER_36_1073 ();
 sg13g2_decap_8 FILLER_36_1080 ();
 sg13g2_decap_8 FILLER_36_1087 ();
 sg13g2_decap_8 FILLER_36_1094 ();
 sg13g2_decap_8 FILLER_36_1101 ();
 sg13g2_decap_8 FILLER_36_1108 ();
 sg13g2_decap_8 FILLER_36_1115 ();
 sg13g2_decap_8 FILLER_36_1122 ();
 sg13g2_decap_8 FILLER_36_1129 ();
 sg13g2_decap_8 FILLER_36_1136 ();
 sg13g2_decap_8 FILLER_36_1143 ();
 sg13g2_decap_8 FILLER_36_1150 ();
 sg13g2_decap_8 FILLER_36_1157 ();
 sg13g2_decap_8 FILLER_36_1164 ();
 sg13g2_decap_8 FILLER_36_1171 ();
 sg13g2_decap_8 FILLER_36_1178 ();
 sg13g2_decap_8 FILLER_36_1185 ();
 sg13g2_decap_8 FILLER_36_1192 ();
 sg13g2_decap_8 FILLER_36_1199 ();
 sg13g2_decap_8 FILLER_36_1206 ();
 sg13g2_decap_8 FILLER_36_1213 ();
 sg13g2_decap_8 FILLER_36_1220 ();
 sg13g2_decap_8 FILLER_36_1227 ();
 sg13g2_decap_8 FILLER_36_1234 ();
 sg13g2_decap_8 FILLER_36_1241 ();
 sg13g2_decap_8 FILLER_36_1248 ();
 sg13g2_decap_8 FILLER_36_1255 ();
 sg13g2_decap_8 FILLER_36_1262 ();
 sg13g2_decap_8 FILLER_36_1269 ();
 sg13g2_decap_8 FILLER_36_1276 ();
 sg13g2_decap_8 FILLER_36_1283 ();
 sg13g2_decap_8 FILLER_36_1290 ();
 sg13g2_decap_8 FILLER_36_1297 ();
 sg13g2_decap_8 FILLER_36_1304 ();
 sg13g2_decap_8 FILLER_36_1311 ();
 sg13g2_decap_8 FILLER_36_1318 ();
 sg13g2_decap_8 FILLER_36_1325 ();
 sg13g2_decap_8 FILLER_36_1332 ();
 sg13g2_decap_8 FILLER_36_1339 ();
 sg13g2_decap_8 FILLER_36_1346 ();
 sg13g2_decap_8 FILLER_36_1353 ();
 sg13g2_decap_8 FILLER_36_1360 ();
 sg13g2_decap_8 FILLER_36_1367 ();
 sg13g2_decap_8 FILLER_36_1374 ();
 sg13g2_decap_8 FILLER_36_1381 ();
 sg13g2_decap_8 FILLER_36_1388 ();
 sg13g2_decap_8 FILLER_36_1395 ();
 sg13g2_decap_8 FILLER_36_1402 ();
 sg13g2_decap_8 FILLER_36_1409 ();
 sg13g2_decap_8 FILLER_36_1416 ();
 sg13g2_decap_8 FILLER_36_1423 ();
 sg13g2_decap_8 FILLER_36_1430 ();
 sg13g2_decap_8 FILLER_36_1437 ();
 sg13g2_decap_8 FILLER_36_1444 ();
 sg13g2_decap_8 FILLER_36_1451 ();
 sg13g2_decap_8 FILLER_36_1458 ();
 sg13g2_decap_8 FILLER_36_1465 ();
 sg13g2_decap_8 FILLER_36_1472 ();
 sg13g2_decap_8 FILLER_36_1479 ();
 sg13g2_decap_8 FILLER_36_1486 ();
 sg13g2_decap_8 FILLER_36_1493 ();
 sg13g2_decap_8 FILLER_36_1500 ();
 sg13g2_decap_8 FILLER_36_1507 ();
 sg13g2_decap_8 FILLER_36_1514 ();
 sg13g2_decap_8 FILLER_36_1521 ();
 sg13g2_decap_8 FILLER_36_1528 ();
 sg13g2_decap_8 FILLER_36_1535 ();
 sg13g2_decap_8 FILLER_36_1542 ();
 sg13g2_decap_8 FILLER_36_1549 ();
 sg13g2_decap_8 FILLER_36_1556 ();
 sg13g2_decap_8 FILLER_36_1563 ();
 sg13g2_decap_8 FILLER_36_1570 ();
 sg13g2_decap_8 FILLER_36_1577 ();
 sg13g2_decap_8 FILLER_36_1584 ();
 sg13g2_decap_8 FILLER_36_1591 ();
 sg13g2_decap_8 FILLER_36_1598 ();
 sg13g2_decap_8 FILLER_36_1605 ();
 sg13g2_decap_8 FILLER_36_1612 ();
 sg13g2_decap_8 FILLER_36_1619 ();
 sg13g2_decap_8 FILLER_36_1626 ();
 sg13g2_decap_8 FILLER_36_1633 ();
 sg13g2_decap_8 FILLER_36_1640 ();
 sg13g2_decap_8 FILLER_36_1647 ();
 sg13g2_decap_8 FILLER_36_1654 ();
 sg13g2_decap_8 FILLER_36_1661 ();
 sg13g2_decap_8 FILLER_36_1668 ();
 sg13g2_decap_8 FILLER_36_1675 ();
 sg13g2_decap_8 FILLER_36_1682 ();
 sg13g2_decap_8 FILLER_36_1689 ();
 sg13g2_decap_8 FILLER_36_1696 ();
 sg13g2_decap_8 FILLER_36_1703 ();
 sg13g2_decap_8 FILLER_36_1710 ();
 sg13g2_decap_8 FILLER_36_1717 ();
 sg13g2_decap_8 FILLER_36_1724 ();
 sg13g2_decap_8 FILLER_36_1731 ();
 sg13g2_decap_8 FILLER_36_1738 ();
 sg13g2_decap_8 FILLER_36_1745 ();
 sg13g2_decap_8 FILLER_36_1752 ();
 sg13g2_decap_8 FILLER_36_1759 ();
 sg13g2_fill_2 FILLER_36_1766 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_fill_1 FILLER_37_70 ();
 sg13g2_decap_4 FILLER_37_80 ();
 sg13g2_fill_2 FILLER_37_84 ();
 sg13g2_fill_2 FILLER_37_107 ();
 sg13g2_fill_1 FILLER_37_139 ();
 sg13g2_fill_2 FILLER_37_148 ();
 sg13g2_fill_1 FILLER_37_150 ();
 sg13g2_decap_8 FILLER_37_177 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_220 ();
 sg13g2_fill_1 FILLER_37_226 ();
 sg13g2_fill_2 FILLER_37_243 ();
 sg13g2_fill_2 FILLER_37_264 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_fill_1 FILLER_37_279 ();
 sg13g2_fill_1 FILLER_37_288 ();
 sg13g2_decap_4 FILLER_37_307 ();
 sg13g2_fill_1 FILLER_37_337 ();
 sg13g2_decap_4 FILLER_37_347 ();
 sg13g2_fill_1 FILLER_37_351 ();
 sg13g2_fill_1 FILLER_37_421 ();
 sg13g2_fill_1 FILLER_37_463 ();
 sg13g2_fill_1 FILLER_37_474 ();
 sg13g2_fill_2 FILLER_37_488 ();
 sg13g2_fill_2 FILLER_37_503 ();
 sg13g2_fill_1 FILLER_37_505 ();
 sg13g2_fill_2 FILLER_37_515 ();
 sg13g2_fill_2 FILLER_37_554 ();
 sg13g2_decap_8 FILLER_37_628 ();
 sg13g2_fill_2 FILLER_37_661 ();
 sg13g2_fill_1 FILLER_37_699 ();
 sg13g2_fill_1 FILLER_37_713 ();
 sg13g2_fill_1 FILLER_37_739 ();
 sg13g2_fill_2 FILLER_37_746 ();
 sg13g2_decap_4 FILLER_37_761 ();
 sg13g2_fill_2 FILLER_37_811 ();
 sg13g2_decap_8 FILLER_37_831 ();
 sg13g2_fill_2 FILLER_37_863 ();
 sg13g2_fill_1 FILLER_37_865 ();
 sg13g2_fill_1 FILLER_37_873 ();
 sg13g2_fill_2 FILLER_37_884 ();
 sg13g2_fill_2 FILLER_37_898 ();
 sg13g2_fill_1 FILLER_37_900 ();
 sg13g2_decap_8 FILLER_37_922 ();
 sg13g2_decap_8 FILLER_37_929 ();
 sg13g2_decap_8 FILLER_37_936 ();
 sg13g2_decap_8 FILLER_37_943 ();
 sg13g2_decap_8 FILLER_37_950 ();
 sg13g2_decap_8 FILLER_37_957 ();
 sg13g2_decap_8 FILLER_37_964 ();
 sg13g2_decap_8 FILLER_37_971 ();
 sg13g2_decap_8 FILLER_37_978 ();
 sg13g2_decap_8 FILLER_37_985 ();
 sg13g2_decap_8 FILLER_37_992 ();
 sg13g2_decap_8 FILLER_37_999 ();
 sg13g2_decap_8 FILLER_37_1006 ();
 sg13g2_decap_8 FILLER_37_1013 ();
 sg13g2_decap_8 FILLER_37_1020 ();
 sg13g2_decap_8 FILLER_37_1027 ();
 sg13g2_decap_8 FILLER_37_1034 ();
 sg13g2_decap_8 FILLER_37_1041 ();
 sg13g2_decap_8 FILLER_37_1048 ();
 sg13g2_decap_8 FILLER_37_1055 ();
 sg13g2_decap_8 FILLER_37_1062 ();
 sg13g2_decap_8 FILLER_37_1069 ();
 sg13g2_decap_8 FILLER_37_1076 ();
 sg13g2_decap_8 FILLER_37_1083 ();
 sg13g2_decap_8 FILLER_37_1090 ();
 sg13g2_decap_8 FILLER_37_1097 ();
 sg13g2_decap_8 FILLER_37_1104 ();
 sg13g2_decap_8 FILLER_37_1111 ();
 sg13g2_decap_8 FILLER_37_1118 ();
 sg13g2_decap_8 FILLER_37_1125 ();
 sg13g2_decap_8 FILLER_37_1132 ();
 sg13g2_decap_8 FILLER_37_1139 ();
 sg13g2_decap_8 FILLER_37_1146 ();
 sg13g2_decap_8 FILLER_37_1153 ();
 sg13g2_decap_8 FILLER_37_1160 ();
 sg13g2_decap_8 FILLER_37_1167 ();
 sg13g2_decap_8 FILLER_37_1174 ();
 sg13g2_decap_8 FILLER_37_1181 ();
 sg13g2_decap_8 FILLER_37_1188 ();
 sg13g2_decap_8 FILLER_37_1195 ();
 sg13g2_decap_8 FILLER_37_1202 ();
 sg13g2_decap_8 FILLER_37_1209 ();
 sg13g2_decap_8 FILLER_37_1216 ();
 sg13g2_decap_8 FILLER_37_1223 ();
 sg13g2_decap_8 FILLER_37_1230 ();
 sg13g2_decap_8 FILLER_37_1237 ();
 sg13g2_decap_8 FILLER_37_1244 ();
 sg13g2_decap_8 FILLER_37_1251 ();
 sg13g2_decap_8 FILLER_37_1258 ();
 sg13g2_decap_8 FILLER_37_1265 ();
 sg13g2_decap_8 FILLER_37_1272 ();
 sg13g2_decap_8 FILLER_37_1279 ();
 sg13g2_decap_8 FILLER_37_1286 ();
 sg13g2_decap_8 FILLER_37_1293 ();
 sg13g2_decap_8 FILLER_37_1300 ();
 sg13g2_decap_8 FILLER_37_1307 ();
 sg13g2_decap_8 FILLER_37_1314 ();
 sg13g2_decap_8 FILLER_37_1321 ();
 sg13g2_decap_8 FILLER_37_1328 ();
 sg13g2_decap_8 FILLER_37_1335 ();
 sg13g2_decap_8 FILLER_37_1342 ();
 sg13g2_decap_8 FILLER_37_1349 ();
 sg13g2_decap_8 FILLER_37_1356 ();
 sg13g2_decap_8 FILLER_37_1363 ();
 sg13g2_decap_8 FILLER_37_1370 ();
 sg13g2_decap_8 FILLER_37_1377 ();
 sg13g2_decap_8 FILLER_37_1384 ();
 sg13g2_decap_8 FILLER_37_1391 ();
 sg13g2_decap_8 FILLER_37_1398 ();
 sg13g2_decap_8 FILLER_37_1405 ();
 sg13g2_decap_8 FILLER_37_1412 ();
 sg13g2_decap_8 FILLER_37_1419 ();
 sg13g2_decap_8 FILLER_37_1426 ();
 sg13g2_decap_8 FILLER_37_1433 ();
 sg13g2_decap_8 FILLER_37_1440 ();
 sg13g2_decap_8 FILLER_37_1447 ();
 sg13g2_decap_8 FILLER_37_1454 ();
 sg13g2_decap_8 FILLER_37_1461 ();
 sg13g2_decap_8 FILLER_37_1468 ();
 sg13g2_decap_8 FILLER_37_1475 ();
 sg13g2_decap_8 FILLER_37_1482 ();
 sg13g2_decap_8 FILLER_37_1489 ();
 sg13g2_decap_8 FILLER_37_1496 ();
 sg13g2_decap_8 FILLER_37_1503 ();
 sg13g2_decap_8 FILLER_37_1510 ();
 sg13g2_decap_8 FILLER_37_1517 ();
 sg13g2_decap_8 FILLER_37_1524 ();
 sg13g2_decap_8 FILLER_37_1531 ();
 sg13g2_decap_8 FILLER_37_1538 ();
 sg13g2_decap_8 FILLER_37_1545 ();
 sg13g2_decap_8 FILLER_37_1552 ();
 sg13g2_decap_8 FILLER_37_1559 ();
 sg13g2_decap_8 FILLER_37_1566 ();
 sg13g2_decap_8 FILLER_37_1573 ();
 sg13g2_decap_8 FILLER_37_1580 ();
 sg13g2_decap_8 FILLER_37_1587 ();
 sg13g2_decap_8 FILLER_37_1594 ();
 sg13g2_decap_8 FILLER_37_1601 ();
 sg13g2_decap_8 FILLER_37_1608 ();
 sg13g2_decap_8 FILLER_37_1615 ();
 sg13g2_decap_8 FILLER_37_1622 ();
 sg13g2_decap_8 FILLER_37_1629 ();
 sg13g2_decap_8 FILLER_37_1636 ();
 sg13g2_decap_8 FILLER_37_1643 ();
 sg13g2_decap_8 FILLER_37_1650 ();
 sg13g2_decap_8 FILLER_37_1657 ();
 sg13g2_decap_8 FILLER_37_1664 ();
 sg13g2_decap_8 FILLER_37_1671 ();
 sg13g2_decap_8 FILLER_37_1678 ();
 sg13g2_decap_8 FILLER_37_1685 ();
 sg13g2_decap_8 FILLER_37_1692 ();
 sg13g2_decap_8 FILLER_37_1699 ();
 sg13g2_decap_8 FILLER_37_1706 ();
 sg13g2_decap_8 FILLER_37_1713 ();
 sg13g2_decap_8 FILLER_37_1720 ();
 sg13g2_decap_8 FILLER_37_1727 ();
 sg13g2_decap_8 FILLER_37_1734 ();
 sg13g2_decap_8 FILLER_37_1741 ();
 sg13g2_decap_8 FILLER_37_1748 ();
 sg13g2_decap_8 FILLER_37_1755 ();
 sg13g2_decap_4 FILLER_37_1762 ();
 sg13g2_fill_2 FILLER_37_1766 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_56 ();
 sg13g2_fill_1 FILLER_38_86 ();
 sg13g2_fill_2 FILLER_38_113 ();
 sg13g2_fill_1 FILLER_38_115 ();
 sg13g2_decap_4 FILLER_38_195 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_fill_1 FILLER_38_227 ();
 sg13g2_decap_4 FILLER_38_244 ();
 sg13g2_decap_4 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_256 ();
 sg13g2_fill_2 FILLER_38_274 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_decap_4 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_321 ();
 sg13g2_fill_1 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_342 ();
 sg13g2_fill_2 FILLER_38_360 ();
 sg13g2_fill_1 FILLER_38_483 ();
 sg13g2_fill_1 FILLER_38_502 ();
 sg13g2_fill_2 FILLER_38_539 ();
 sg13g2_fill_2 FILLER_38_571 ();
 sg13g2_fill_1 FILLER_38_573 ();
 sg13g2_fill_2 FILLER_38_583 ();
 sg13g2_fill_2 FILLER_38_622 ();
 sg13g2_fill_1 FILLER_38_624 ();
 sg13g2_fill_2 FILLER_38_644 ();
 sg13g2_fill_1 FILLER_38_646 ();
 sg13g2_decap_4 FILLER_38_656 ();
 sg13g2_fill_2 FILLER_38_660 ();
 sg13g2_decap_4 FILLER_38_675 ();
 sg13g2_fill_2 FILLER_38_705 ();
 sg13g2_fill_2 FILLER_38_729 ();
 sg13g2_fill_1 FILLER_38_731 ();
 sg13g2_decap_8 FILLER_38_736 ();
 sg13g2_fill_1 FILLER_38_769 ();
 sg13g2_fill_2 FILLER_38_777 ();
 sg13g2_decap_8 FILLER_38_800 ();
 sg13g2_fill_1 FILLER_38_807 ();
 sg13g2_fill_2 FILLER_38_814 ();
 sg13g2_decap_8 FILLER_38_835 ();
 sg13g2_fill_2 FILLER_38_842 ();
 sg13g2_fill_1 FILLER_38_863 ();
 sg13g2_fill_1 FILLER_38_887 ();
 sg13g2_decap_8 FILLER_38_900 ();
 sg13g2_decap_8 FILLER_38_907 ();
 sg13g2_decap_8 FILLER_38_914 ();
 sg13g2_decap_8 FILLER_38_921 ();
 sg13g2_decap_8 FILLER_38_928 ();
 sg13g2_decap_8 FILLER_38_935 ();
 sg13g2_decap_8 FILLER_38_942 ();
 sg13g2_decap_8 FILLER_38_949 ();
 sg13g2_decap_8 FILLER_38_956 ();
 sg13g2_decap_8 FILLER_38_963 ();
 sg13g2_decap_8 FILLER_38_970 ();
 sg13g2_decap_8 FILLER_38_977 ();
 sg13g2_decap_8 FILLER_38_984 ();
 sg13g2_decap_8 FILLER_38_991 ();
 sg13g2_decap_8 FILLER_38_998 ();
 sg13g2_decap_8 FILLER_38_1005 ();
 sg13g2_decap_8 FILLER_38_1012 ();
 sg13g2_decap_8 FILLER_38_1019 ();
 sg13g2_decap_8 FILLER_38_1026 ();
 sg13g2_decap_8 FILLER_38_1033 ();
 sg13g2_decap_8 FILLER_38_1040 ();
 sg13g2_decap_8 FILLER_38_1047 ();
 sg13g2_decap_8 FILLER_38_1054 ();
 sg13g2_decap_8 FILLER_38_1061 ();
 sg13g2_decap_8 FILLER_38_1068 ();
 sg13g2_decap_8 FILLER_38_1075 ();
 sg13g2_decap_8 FILLER_38_1082 ();
 sg13g2_decap_8 FILLER_38_1089 ();
 sg13g2_decap_8 FILLER_38_1096 ();
 sg13g2_decap_8 FILLER_38_1103 ();
 sg13g2_decap_8 FILLER_38_1110 ();
 sg13g2_decap_8 FILLER_38_1117 ();
 sg13g2_decap_8 FILLER_38_1124 ();
 sg13g2_decap_8 FILLER_38_1131 ();
 sg13g2_decap_8 FILLER_38_1138 ();
 sg13g2_decap_8 FILLER_38_1145 ();
 sg13g2_decap_8 FILLER_38_1152 ();
 sg13g2_decap_8 FILLER_38_1159 ();
 sg13g2_decap_8 FILLER_38_1166 ();
 sg13g2_decap_8 FILLER_38_1173 ();
 sg13g2_decap_8 FILLER_38_1180 ();
 sg13g2_decap_8 FILLER_38_1187 ();
 sg13g2_decap_8 FILLER_38_1194 ();
 sg13g2_decap_8 FILLER_38_1201 ();
 sg13g2_decap_8 FILLER_38_1208 ();
 sg13g2_decap_8 FILLER_38_1215 ();
 sg13g2_decap_8 FILLER_38_1222 ();
 sg13g2_decap_8 FILLER_38_1229 ();
 sg13g2_decap_8 FILLER_38_1236 ();
 sg13g2_decap_8 FILLER_38_1243 ();
 sg13g2_decap_8 FILLER_38_1250 ();
 sg13g2_decap_8 FILLER_38_1257 ();
 sg13g2_decap_8 FILLER_38_1264 ();
 sg13g2_decap_8 FILLER_38_1271 ();
 sg13g2_decap_8 FILLER_38_1278 ();
 sg13g2_decap_8 FILLER_38_1285 ();
 sg13g2_decap_8 FILLER_38_1292 ();
 sg13g2_decap_8 FILLER_38_1299 ();
 sg13g2_decap_8 FILLER_38_1306 ();
 sg13g2_decap_8 FILLER_38_1313 ();
 sg13g2_decap_8 FILLER_38_1320 ();
 sg13g2_decap_8 FILLER_38_1327 ();
 sg13g2_decap_8 FILLER_38_1334 ();
 sg13g2_decap_8 FILLER_38_1341 ();
 sg13g2_decap_8 FILLER_38_1348 ();
 sg13g2_decap_8 FILLER_38_1355 ();
 sg13g2_decap_8 FILLER_38_1362 ();
 sg13g2_decap_8 FILLER_38_1369 ();
 sg13g2_decap_8 FILLER_38_1376 ();
 sg13g2_decap_8 FILLER_38_1383 ();
 sg13g2_decap_8 FILLER_38_1390 ();
 sg13g2_decap_8 FILLER_38_1397 ();
 sg13g2_decap_8 FILLER_38_1404 ();
 sg13g2_decap_8 FILLER_38_1411 ();
 sg13g2_decap_8 FILLER_38_1418 ();
 sg13g2_decap_8 FILLER_38_1425 ();
 sg13g2_decap_8 FILLER_38_1432 ();
 sg13g2_decap_8 FILLER_38_1439 ();
 sg13g2_decap_8 FILLER_38_1446 ();
 sg13g2_decap_8 FILLER_38_1453 ();
 sg13g2_decap_8 FILLER_38_1460 ();
 sg13g2_decap_8 FILLER_38_1467 ();
 sg13g2_decap_8 FILLER_38_1474 ();
 sg13g2_decap_8 FILLER_38_1481 ();
 sg13g2_decap_8 FILLER_38_1488 ();
 sg13g2_decap_8 FILLER_38_1495 ();
 sg13g2_decap_8 FILLER_38_1502 ();
 sg13g2_decap_8 FILLER_38_1509 ();
 sg13g2_decap_8 FILLER_38_1516 ();
 sg13g2_decap_8 FILLER_38_1523 ();
 sg13g2_decap_8 FILLER_38_1530 ();
 sg13g2_decap_8 FILLER_38_1537 ();
 sg13g2_decap_8 FILLER_38_1544 ();
 sg13g2_decap_8 FILLER_38_1551 ();
 sg13g2_decap_8 FILLER_38_1558 ();
 sg13g2_decap_8 FILLER_38_1565 ();
 sg13g2_decap_8 FILLER_38_1572 ();
 sg13g2_decap_8 FILLER_38_1579 ();
 sg13g2_decap_8 FILLER_38_1586 ();
 sg13g2_decap_8 FILLER_38_1593 ();
 sg13g2_decap_8 FILLER_38_1600 ();
 sg13g2_decap_8 FILLER_38_1607 ();
 sg13g2_decap_8 FILLER_38_1614 ();
 sg13g2_decap_8 FILLER_38_1621 ();
 sg13g2_decap_8 FILLER_38_1628 ();
 sg13g2_decap_8 FILLER_38_1635 ();
 sg13g2_decap_8 FILLER_38_1642 ();
 sg13g2_decap_8 FILLER_38_1649 ();
 sg13g2_decap_8 FILLER_38_1656 ();
 sg13g2_decap_8 FILLER_38_1663 ();
 sg13g2_decap_8 FILLER_38_1670 ();
 sg13g2_decap_8 FILLER_38_1677 ();
 sg13g2_decap_8 FILLER_38_1684 ();
 sg13g2_decap_8 FILLER_38_1691 ();
 sg13g2_decap_8 FILLER_38_1698 ();
 sg13g2_decap_8 FILLER_38_1705 ();
 sg13g2_decap_8 FILLER_38_1712 ();
 sg13g2_decap_8 FILLER_38_1719 ();
 sg13g2_decap_8 FILLER_38_1726 ();
 sg13g2_decap_8 FILLER_38_1733 ();
 sg13g2_decap_8 FILLER_38_1740 ();
 sg13g2_decap_8 FILLER_38_1747 ();
 sg13g2_decap_8 FILLER_38_1754 ();
 sg13g2_decap_8 FILLER_38_1761 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_4 FILLER_39_63 ();
 sg13g2_fill_1 FILLER_39_67 ();
 sg13g2_fill_2 FILLER_39_95 ();
 sg13g2_fill_1 FILLER_39_97 ();
 sg13g2_fill_2 FILLER_39_109 ();
 sg13g2_fill_1 FILLER_39_111 ();
 sg13g2_fill_1 FILLER_39_130 ();
 sg13g2_decap_8 FILLER_39_162 ();
 sg13g2_decap_4 FILLER_39_169 ();
 sg13g2_fill_2 FILLER_39_173 ();
 sg13g2_fill_1 FILLER_39_180 ();
 sg13g2_decap_8 FILLER_39_192 ();
 sg13g2_decap_4 FILLER_39_199 ();
 sg13g2_fill_1 FILLER_39_208 ();
 sg13g2_fill_1 FILLER_39_232 ();
 sg13g2_decap_8 FILLER_39_237 ();
 sg13g2_decap_4 FILLER_39_244 ();
 sg13g2_fill_1 FILLER_39_248 ();
 sg13g2_fill_2 FILLER_39_283 ();
 sg13g2_fill_1 FILLER_39_306 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_fill_2 FILLER_39_322 ();
 sg13g2_fill_2 FILLER_39_352 ();
 sg13g2_fill_1 FILLER_39_354 ();
 sg13g2_fill_1 FILLER_39_386 ();
 sg13g2_fill_1 FILLER_39_413 ();
 sg13g2_fill_1 FILLER_39_505 ();
 sg13g2_fill_2 FILLER_39_524 ();
 sg13g2_fill_2 FILLER_39_541 ();
 sg13g2_fill_1 FILLER_39_552 ();
 sg13g2_fill_2 FILLER_39_575 ();
 sg13g2_decap_4 FILLER_39_597 ();
 sg13g2_fill_1 FILLER_39_601 ();
 sg13g2_fill_2 FILLER_39_612 ();
 sg13g2_decap_8 FILLER_39_651 ();
 sg13g2_fill_2 FILLER_39_658 ();
 sg13g2_decap_8 FILLER_39_663 ();
 sg13g2_decap_8 FILLER_39_670 ();
 sg13g2_decap_8 FILLER_39_677 ();
 sg13g2_decap_4 FILLER_39_684 ();
 sg13g2_fill_1 FILLER_39_688 ();
 sg13g2_decap_4 FILLER_39_780 ();
 sg13g2_fill_1 FILLER_39_784 ();
 sg13g2_decap_4 FILLER_39_795 ();
 sg13g2_fill_1 FILLER_39_799 ();
 sg13g2_fill_2 FILLER_39_805 ();
 sg13g2_fill_2 FILLER_39_817 ();
 sg13g2_fill_1 FILLER_39_819 ();
 sg13g2_decap_8 FILLER_39_828 ();
 sg13g2_fill_2 FILLER_39_835 ();
 sg13g2_decap_4 FILLER_39_845 ();
 sg13g2_decap_8 FILLER_39_854 ();
 sg13g2_decap_8 FILLER_39_861 ();
 sg13g2_fill_2 FILLER_39_868 ();
 sg13g2_fill_1 FILLER_39_870 ();
 sg13g2_decap_8 FILLER_39_880 ();
 sg13g2_decap_8 FILLER_39_887 ();
 sg13g2_decap_8 FILLER_39_894 ();
 sg13g2_decap_8 FILLER_39_901 ();
 sg13g2_decap_8 FILLER_39_908 ();
 sg13g2_decap_8 FILLER_39_915 ();
 sg13g2_decap_8 FILLER_39_922 ();
 sg13g2_decap_8 FILLER_39_929 ();
 sg13g2_decap_8 FILLER_39_936 ();
 sg13g2_decap_8 FILLER_39_943 ();
 sg13g2_decap_8 FILLER_39_950 ();
 sg13g2_decap_8 FILLER_39_957 ();
 sg13g2_decap_8 FILLER_39_964 ();
 sg13g2_decap_8 FILLER_39_971 ();
 sg13g2_decap_8 FILLER_39_978 ();
 sg13g2_decap_8 FILLER_39_985 ();
 sg13g2_decap_8 FILLER_39_992 ();
 sg13g2_decap_8 FILLER_39_999 ();
 sg13g2_decap_8 FILLER_39_1006 ();
 sg13g2_decap_8 FILLER_39_1013 ();
 sg13g2_decap_8 FILLER_39_1020 ();
 sg13g2_decap_8 FILLER_39_1027 ();
 sg13g2_decap_8 FILLER_39_1034 ();
 sg13g2_decap_8 FILLER_39_1041 ();
 sg13g2_decap_8 FILLER_39_1048 ();
 sg13g2_decap_8 FILLER_39_1055 ();
 sg13g2_decap_8 FILLER_39_1062 ();
 sg13g2_decap_8 FILLER_39_1069 ();
 sg13g2_decap_8 FILLER_39_1076 ();
 sg13g2_decap_8 FILLER_39_1083 ();
 sg13g2_decap_8 FILLER_39_1090 ();
 sg13g2_decap_8 FILLER_39_1097 ();
 sg13g2_decap_8 FILLER_39_1104 ();
 sg13g2_decap_8 FILLER_39_1111 ();
 sg13g2_decap_8 FILLER_39_1118 ();
 sg13g2_decap_8 FILLER_39_1125 ();
 sg13g2_decap_8 FILLER_39_1132 ();
 sg13g2_decap_8 FILLER_39_1139 ();
 sg13g2_decap_8 FILLER_39_1146 ();
 sg13g2_decap_8 FILLER_39_1153 ();
 sg13g2_decap_8 FILLER_39_1160 ();
 sg13g2_decap_8 FILLER_39_1167 ();
 sg13g2_decap_8 FILLER_39_1174 ();
 sg13g2_decap_8 FILLER_39_1181 ();
 sg13g2_decap_8 FILLER_39_1188 ();
 sg13g2_decap_8 FILLER_39_1195 ();
 sg13g2_decap_8 FILLER_39_1202 ();
 sg13g2_decap_8 FILLER_39_1209 ();
 sg13g2_decap_8 FILLER_39_1216 ();
 sg13g2_decap_8 FILLER_39_1223 ();
 sg13g2_decap_8 FILLER_39_1230 ();
 sg13g2_decap_8 FILLER_39_1237 ();
 sg13g2_decap_8 FILLER_39_1244 ();
 sg13g2_decap_8 FILLER_39_1251 ();
 sg13g2_decap_8 FILLER_39_1258 ();
 sg13g2_decap_8 FILLER_39_1265 ();
 sg13g2_decap_8 FILLER_39_1272 ();
 sg13g2_decap_8 FILLER_39_1279 ();
 sg13g2_decap_8 FILLER_39_1286 ();
 sg13g2_decap_8 FILLER_39_1293 ();
 sg13g2_decap_8 FILLER_39_1300 ();
 sg13g2_decap_8 FILLER_39_1307 ();
 sg13g2_decap_8 FILLER_39_1314 ();
 sg13g2_decap_8 FILLER_39_1321 ();
 sg13g2_decap_8 FILLER_39_1328 ();
 sg13g2_decap_8 FILLER_39_1335 ();
 sg13g2_decap_8 FILLER_39_1342 ();
 sg13g2_decap_8 FILLER_39_1349 ();
 sg13g2_decap_8 FILLER_39_1356 ();
 sg13g2_decap_8 FILLER_39_1363 ();
 sg13g2_decap_8 FILLER_39_1370 ();
 sg13g2_decap_8 FILLER_39_1377 ();
 sg13g2_decap_8 FILLER_39_1384 ();
 sg13g2_decap_8 FILLER_39_1391 ();
 sg13g2_decap_8 FILLER_39_1398 ();
 sg13g2_decap_8 FILLER_39_1405 ();
 sg13g2_decap_8 FILLER_39_1412 ();
 sg13g2_decap_8 FILLER_39_1419 ();
 sg13g2_decap_8 FILLER_39_1426 ();
 sg13g2_decap_8 FILLER_39_1433 ();
 sg13g2_decap_8 FILLER_39_1440 ();
 sg13g2_decap_8 FILLER_39_1447 ();
 sg13g2_decap_8 FILLER_39_1454 ();
 sg13g2_decap_8 FILLER_39_1461 ();
 sg13g2_decap_8 FILLER_39_1468 ();
 sg13g2_decap_8 FILLER_39_1475 ();
 sg13g2_decap_8 FILLER_39_1482 ();
 sg13g2_decap_8 FILLER_39_1489 ();
 sg13g2_decap_8 FILLER_39_1496 ();
 sg13g2_decap_8 FILLER_39_1503 ();
 sg13g2_decap_8 FILLER_39_1510 ();
 sg13g2_decap_8 FILLER_39_1517 ();
 sg13g2_decap_8 FILLER_39_1524 ();
 sg13g2_decap_8 FILLER_39_1531 ();
 sg13g2_decap_8 FILLER_39_1538 ();
 sg13g2_decap_8 FILLER_39_1545 ();
 sg13g2_decap_8 FILLER_39_1552 ();
 sg13g2_decap_8 FILLER_39_1559 ();
 sg13g2_decap_8 FILLER_39_1566 ();
 sg13g2_decap_8 FILLER_39_1573 ();
 sg13g2_decap_8 FILLER_39_1580 ();
 sg13g2_decap_8 FILLER_39_1587 ();
 sg13g2_decap_8 FILLER_39_1594 ();
 sg13g2_decap_8 FILLER_39_1601 ();
 sg13g2_decap_8 FILLER_39_1608 ();
 sg13g2_decap_8 FILLER_39_1615 ();
 sg13g2_decap_8 FILLER_39_1622 ();
 sg13g2_decap_8 FILLER_39_1629 ();
 sg13g2_decap_8 FILLER_39_1636 ();
 sg13g2_decap_8 FILLER_39_1643 ();
 sg13g2_decap_8 FILLER_39_1650 ();
 sg13g2_decap_8 FILLER_39_1657 ();
 sg13g2_decap_8 FILLER_39_1664 ();
 sg13g2_decap_8 FILLER_39_1671 ();
 sg13g2_decap_8 FILLER_39_1678 ();
 sg13g2_decap_8 FILLER_39_1685 ();
 sg13g2_decap_8 FILLER_39_1692 ();
 sg13g2_decap_8 FILLER_39_1699 ();
 sg13g2_decap_8 FILLER_39_1706 ();
 sg13g2_decap_8 FILLER_39_1713 ();
 sg13g2_decap_8 FILLER_39_1720 ();
 sg13g2_decap_8 FILLER_39_1727 ();
 sg13g2_decap_8 FILLER_39_1734 ();
 sg13g2_decap_8 FILLER_39_1741 ();
 sg13g2_decap_8 FILLER_39_1748 ();
 sg13g2_decap_8 FILLER_39_1755 ();
 sg13g2_decap_4 FILLER_39_1762 ();
 sg13g2_fill_2 FILLER_39_1766 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_4 FILLER_40_70 ();
 sg13g2_fill_2 FILLER_40_74 ();
 sg13g2_fill_2 FILLER_40_102 ();
 sg13g2_fill_1 FILLER_40_104 ();
 sg13g2_fill_1 FILLER_40_142 ();
 sg13g2_fill_2 FILLER_40_169 ();
 sg13g2_decap_8 FILLER_40_202 ();
 sg13g2_decap_8 FILLER_40_223 ();
 sg13g2_fill_2 FILLER_40_230 ();
 sg13g2_fill_1 FILLER_40_232 ();
 sg13g2_fill_2 FILLER_40_253 ();
 sg13g2_decap_8 FILLER_40_279 ();
 sg13g2_fill_2 FILLER_40_286 ();
 sg13g2_fill_2 FILLER_40_312 ();
 sg13g2_fill_1 FILLER_40_340 ();
 sg13g2_fill_2 FILLER_40_376 ();
 sg13g2_fill_1 FILLER_40_378 ();
 sg13g2_fill_1 FILLER_40_398 ();
 sg13g2_decap_8 FILLER_40_407 ();
 sg13g2_decap_8 FILLER_40_414 ();
 sg13g2_decap_8 FILLER_40_421 ();
 sg13g2_decap_4 FILLER_40_428 ();
 sg13g2_fill_2 FILLER_40_436 ();
 sg13g2_fill_1 FILLER_40_438 ();
 sg13g2_decap_4 FILLER_40_457 ();
 sg13g2_fill_1 FILLER_40_478 ();
 sg13g2_fill_2 FILLER_40_541 ();
 sg13g2_fill_1 FILLER_40_543 ();
 sg13g2_fill_2 FILLER_40_564 ();
 sg13g2_fill_1 FILLER_40_566 ();
 sg13g2_fill_2 FILLER_40_583 ();
 sg13g2_fill_1 FILLER_40_585 ();
 sg13g2_fill_1 FILLER_40_609 ();
 sg13g2_fill_1 FILLER_40_638 ();
 sg13g2_decap_4 FILLER_40_666 ();
 sg13g2_fill_1 FILLER_40_670 ();
 sg13g2_decap_8 FILLER_40_696 ();
 sg13g2_decap_8 FILLER_40_703 ();
 sg13g2_fill_2 FILLER_40_710 ();
 sg13g2_fill_1 FILLER_40_712 ();
 sg13g2_decap_8 FILLER_40_717 ();
 sg13g2_decap_8 FILLER_40_724 ();
 sg13g2_decap_8 FILLER_40_731 ();
 sg13g2_decap_8 FILLER_40_738 ();
 sg13g2_fill_2 FILLER_40_745 ();
 sg13g2_fill_1 FILLER_40_747 ();
 sg13g2_fill_2 FILLER_40_761 ();
 sg13g2_fill_1 FILLER_40_763 ();
 sg13g2_decap_4 FILLER_40_788 ();
 sg13g2_decap_8 FILLER_40_817 ();
 sg13g2_fill_1 FILLER_40_824 ();
 sg13g2_decap_8 FILLER_40_829 ();
 sg13g2_decap_4 FILLER_40_836 ();
 sg13g2_decap_8 FILLER_40_844 ();
 sg13g2_decap_8 FILLER_40_851 ();
 sg13g2_decap_8 FILLER_40_858 ();
 sg13g2_decap_8 FILLER_40_865 ();
 sg13g2_decap_8 FILLER_40_872 ();
 sg13g2_decap_8 FILLER_40_879 ();
 sg13g2_decap_8 FILLER_40_886 ();
 sg13g2_decap_8 FILLER_40_893 ();
 sg13g2_decap_8 FILLER_40_900 ();
 sg13g2_decap_8 FILLER_40_907 ();
 sg13g2_decap_8 FILLER_40_914 ();
 sg13g2_decap_8 FILLER_40_921 ();
 sg13g2_decap_8 FILLER_40_928 ();
 sg13g2_decap_8 FILLER_40_935 ();
 sg13g2_decap_8 FILLER_40_942 ();
 sg13g2_decap_8 FILLER_40_949 ();
 sg13g2_decap_8 FILLER_40_956 ();
 sg13g2_decap_8 FILLER_40_963 ();
 sg13g2_decap_8 FILLER_40_970 ();
 sg13g2_decap_8 FILLER_40_977 ();
 sg13g2_decap_8 FILLER_40_984 ();
 sg13g2_decap_8 FILLER_40_991 ();
 sg13g2_decap_8 FILLER_40_998 ();
 sg13g2_decap_8 FILLER_40_1005 ();
 sg13g2_decap_8 FILLER_40_1012 ();
 sg13g2_decap_8 FILLER_40_1019 ();
 sg13g2_decap_8 FILLER_40_1026 ();
 sg13g2_decap_8 FILLER_40_1033 ();
 sg13g2_decap_8 FILLER_40_1040 ();
 sg13g2_decap_8 FILLER_40_1047 ();
 sg13g2_decap_8 FILLER_40_1054 ();
 sg13g2_decap_8 FILLER_40_1061 ();
 sg13g2_decap_8 FILLER_40_1068 ();
 sg13g2_decap_8 FILLER_40_1075 ();
 sg13g2_decap_8 FILLER_40_1082 ();
 sg13g2_decap_8 FILLER_40_1089 ();
 sg13g2_decap_8 FILLER_40_1096 ();
 sg13g2_decap_8 FILLER_40_1103 ();
 sg13g2_decap_8 FILLER_40_1110 ();
 sg13g2_decap_8 FILLER_40_1117 ();
 sg13g2_decap_8 FILLER_40_1124 ();
 sg13g2_decap_8 FILLER_40_1131 ();
 sg13g2_decap_8 FILLER_40_1138 ();
 sg13g2_decap_8 FILLER_40_1145 ();
 sg13g2_decap_8 FILLER_40_1152 ();
 sg13g2_decap_8 FILLER_40_1159 ();
 sg13g2_decap_8 FILLER_40_1166 ();
 sg13g2_decap_8 FILLER_40_1173 ();
 sg13g2_decap_8 FILLER_40_1180 ();
 sg13g2_decap_8 FILLER_40_1187 ();
 sg13g2_decap_8 FILLER_40_1194 ();
 sg13g2_decap_8 FILLER_40_1201 ();
 sg13g2_decap_8 FILLER_40_1208 ();
 sg13g2_decap_8 FILLER_40_1215 ();
 sg13g2_decap_8 FILLER_40_1222 ();
 sg13g2_decap_8 FILLER_40_1229 ();
 sg13g2_decap_8 FILLER_40_1236 ();
 sg13g2_decap_8 FILLER_40_1243 ();
 sg13g2_decap_8 FILLER_40_1250 ();
 sg13g2_decap_8 FILLER_40_1257 ();
 sg13g2_decap_8 FILLER_40_1264 ();
 sg13g2_decap_8 FILLER_40_1271 ();
 sg13g2_decap_8 FILLER_40_1278 ();
 sg13g2_decap_8 FILLER_40_1285 ();
 sg13g2_decap_8 FILLER_40_1292 ();
 sg13g2_decap_8 FILLER_40_1299 ();
 sg13g2_decap_8 FILLER_40_1306 ();
 sg13g2_decap_8 FILLER_40_1313 ();
 sg13g2_decap_8 FILLER_40_1320 ();
 sg13g2_decap_8 FILLER_40_1327 ();
 sg13g2_decap_8 FILLER_40_1334 ();
 sg13g2_decap_8 FILLER_40_1341 ();
 sg13g2_decap_8 FILLER_40_1348 ();
 sg13g2_decap_8 FILLER_40_1355 ();
 sg13g2_decap_8 FILLER_40_1362 ();
 sg13g2_decap_8 FILLER_40_1369 ();
 sg13g2_decap_8 FILLER_40_1376 ();
 sg13g2_decap_8 FILLER_40_1383 ();
 sg13g2_decap_8 FILLER_40_1390 ();
 sg13g2_decap_8 FILLER_40_1397 ();
 sg13g2_decap_8 FILLER_40_1404 ();
 sg13g2_decap_8 FILLER_40_1411 ();
 sg13g2_decap_8 FILLER_40_1418 ();
 sg13g2_decap_8 FILLER_40_1425 ();
 sg13g2_decap_8 FILLER_40_1432 ();
 sg13g2_decap_8 FILLER_40_1439 ();
 sg13g2_decap_8 FILLER_40_1446 ();
 sg13g2_decap_8 FILLER_40_1453 ();
 sg13g2_decap_8 FILLER_40_1460 ();
 sg13g2_decap_8 FILLER_40_1467 ();
 sg13g2_decap_8 FILLER_40_1474 ();
 sg13g2_decap_8 FILLER_40_1481 ();
 sg13g2_decap_8 FILLER_40_1488 ();
 sg13g2_decap_8 FILLER_40_1495 ();
 sg13g2_decap_8 FILLER_40_1502 ();
 sg13g2_decap_8 FILLER_40_1509 ();
 sg13g2_decap_8 FILLER_40_1516 ();
 sg13g2_decap_8 FILLER_40_1523 ();
 sg13g2_decap_8 FILLER_40_1530 ();
 sg13g2_decap_8 FILLER_40_1537 ();
 sg13g2_decap_8 FILLER_40_1544 ();
 sg13g2_decap_8 FILLER_40_1551 ();
 sg13g2_decap_8 FILLER_40_1558 ();
 sg13g2_decap_8 FILLER_40_1565 ();
 sg13g2_decap_8 FILLER_40_1572 ();
 sg13g2_decap_8 FILLER_40_1579 ();
 sg13g2_decap_8 FILLER_40_1586 ();
 sg13g2_decap_8 FILLER_40_1593 ();
 sg13g2_decap_8 FILLER_40_1600 ();
 sg13g2_decap_8 FILLER_40_1607 ();
 sg13g2_decap_8 FILLER_40_1614 ();
 sg13g2_decap_8 FILLER_40_1621 ();
 sg13g2_decap_8 FILLER_40_1628 ();
 sg13g2_decap_8 FILLER_40_1635 ();
 sg13g2_decap_8 FILLER_40_1642 ();
 sg13g2_decap_8 FILLER_40_1649 ();
 sg13g2_decap_8 FILLER_40_1656 ();
 sg13g2_decap_8 FILLER_40_1663 ();
 sg13g2_decap_8 FILLER_40_1670 ();
 sg13g2_decap_8 FILLER_40_1677 ();
 sg13g2_decap_8 FILLER_40_1684 ();
 sg13g2_decap_8 FILLER_40_1691 ();
 sg13g2_decap_8 FILLER_40_1698 ();
 sg13g2_decap_8 FILLER_40_1705 ();
 sg13g2_decap_8 FILLER_40_1712 ();
 sg13g2_decap_8 FILLER_40_1719 ();
 sg13g2_decap_8 FILLER_40_1726 ();
 sg13g2_decap_8 FILLER_40_1733 ();
 sg13g2_decap_8 FILLER_40_1740 ();
 sg13g2_decap_8 FILLER_40_1747 ();
 sg13g2_decap_8 FILLER_40_1754 ();
 sg13g2_decap_8 FILLER_40_1761 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_fill_1 FILLER_41_70 ();
 sg13g2_fill_2 FILLER_41_84 ();
 sg13g2_fill_2 FILLER_41_95 ();
 sg13g2_fill_1 FILLER_41_97 ();
 sg13g2_decap_4 FILLER_41_107 ();
 sg13g2_fill_2 FILLER_41_111 ();
 sg13g2_fill_2 FILLER_41_149 ();
 sg13g2_fill_2 FILLER_41_155 ();
 sg13g2_fill_1 FILLER_41_157 ();
 sg13g2_fill_1 FILLER_41_180 ();
 sg13g2_fill_2 FILLER_41_189 ();
 sg13g2_fill_1 FILLER_41_200 ();
 sg13g2_fill_2 FILLER_41_232 ();
 sg13g2_fill_2 FILLER_41_266 ();
 sg13g2_fill_1 FILLER_41_268 ();
 sg13g2_decap_4 FILLER_41_275 ();
 sg13g2_decap_8 FILLER_41_283 ();
 sg13g2_decap_8 FILLER_41_290 ();
 sg13g2_decap_4 FILLER_41_297 ();
 sg13g2_fill_1 FILLER_41_301 ();
 sg13g2_decap_4 FILLER_41_310 ();
 sg13g2_fill_1 FILLER_41_314 ();
 sg13g2_fill_1 FILLER_41_326 ();
 sg13g2_decap_8 FILLER_41_332 ();
 sg13g2_fill_2 FILLER_41_339 ();
 sg13g2_fill_1 FILLER_41_341 ();
 sg13g2_fill_2 FILLER_41_353 ();
 sg13g2_fill_2 FILLER_41_447 ();
 sg13g2_fill_2 FILLER_41_479 ();
 sg13g2_fill_2 FILLER_41_491 ();
 sg13g2_fill_1 FILLER_41_493 ();
 sg13g2_fill_1 FILLER_41_503 ();
 sg13g2_fill_1 FILLER_41_531 ();
 sg13g2_fill_2 FILLER_41_538 ();
 sg13g2_decap_4 FILLER_41_549 ();
 sg13g2_fill_2 FILLER_41_553 ();
 sg13g2_fill_1 FILLER_41_563 ();
 sg13g2_fill_1 FILLER_41_576 ();
 sg13g2_fill_2 FILLER_41_599 ();
 sg13g2_fill_1 FILLER_41_601 ();
 sg13g2_decap_8 FILLER_41_622 ();
 sg13g2_decap_8 FILLER_41_629 ();
 sg13g2_fill_1 FILLER_41_636 ();
 sg13g2_fill_2 FILLER_41_642 ();
 sg13g2_decap_4 FILLER_41_661 ();
 sg13g2_decap_8 FILLER_41_674 ();
 sg13g2_fill_2 FILLER_41_681 ();
 sg13g2_decap_8 FILLER_41_693 ();
 sg13g2_fill_2 FILLER_41_705 ();
 sg13g2_fill_1 FILLER_41_707 ();
 sg13g2_decap_8 FILLER_41_724 ();
 sg13g2_decap_8 FILLER_41_731 ();
 sg13g2_decap_4 FILLER_41_738 ();
 sg13g2_fill_1 FILLER_41_742 ();
 sg13g2_fill_2 FILLER_41_769 ();
 sg13g2_fill_1 FILLER_41_771 ();
 sg13g2_fill_2 FILLER_41_781 ();
 sg13g2_decap_8 FILLER_41_788 ();
 sg13g2_fill_2 FILLER_41_795 ();
 sg13g2_decap_4 FILLER_41_801 ();
 sg13g2_fill_1 FILLER_41_805 ();
 sg13g2_decap_8 FILLER_41_855 ();
 sg13g2_decap_8 FILLER_41_862 ();
 sg13g2_decap_8 FILLER_41_869 ();
 sg13g2_fill_2 FILLER_41_876 ();
 sg13g2_fill_1 FILLER_41_878 ();
 sg13g2_decap_8 FILLER_41_891 ();
 sg13g2_decap_8 FILLER_41_898 ();
 sg13g2_fill_2 FILLER_41_905 ();
 sg13g2_fill_1 FILLER_41_907 ();
 sg13g2_decap_8 FILLER_41_918 ();
 sg13g2_decap_8 FILLER_41_925 ();
 sg13g2_decap_8 FILLER_41_932 ();
 sg13g2_decap_8 FILLER_41_939 ();
 sg13g2_decap_8 FILLER_41_946 ();
 sg13g2_decap_8 FILLER_41_953 ();
 sg13g2_decap_8 FILLER_41_960 ();
 sg13g2_decap_8 FILLER_41_967 ();
 sg13g2_decap_8 FILLER_41_974 ();
 sg13g2_decap_8 FILLER_41_981 ();
 sg13g2_decap_8 FILLER_41_988 ();
 sg13g2_decap_8 FILLER_41_995 ();
 sg13g2_decap_8 FILLER_41_1002 ();
 sg13g2_decap_8 FILLER_41_1009 ();
 sg13g2_decap_8 FILLER_41_1016 ();
 sg13g2_decap_8 FILLER_41_1023 ();
 sg13g2_decap_8 FILLER_41_1030 ();
 sg13g2_decap_8 FILLER_41_1037 ();
 sg13g2_decap_8 FILLER_41_1044 ();
 sg13g2_decap_8 FILLER_41_1051 ();
 sg13g2_decap_8 FILLER_41_1058 ();
 sg13g2_decap_8 FILLER_41_1065 ();
 sg13g2_decap_8 FILLER_41_1072 ();
 sg13g2_decap_8 FILLER_41_1079 ();
 sg13g2_decap_8 FILLER_41_1086 ();
 sg13g2_decap_8 FILLER_41_1093 ();
 sg13g2_decap_8 FILLER_41_1100 ();
 sg13g2_decap_8 FILLER_41_1107 ();
 sg13g2_decap_8 FILLER_41_1114 ();
 sg13g2_decap_8 FILLER_41_1121 ();
 sg13g2_decap_8 FILLER_41_1128 ();
 sg13g2_decap_8 FILLER_41_1135 ();
 sg13g2_decap_8 FILLER_41_1142 ();
 sg13g2_decap_8 FILLER_41_1149 ();
 sg13g2_decap_8 FILLER_41_1156 ();
 sg13g2_decap_8 FILLER_41_1163 ();
 sg13g2_decap_8 FILLER_41_1170 ();
 sg13g2_decap_8 FILLER_41_1177 ();
 sg13g2_decap_8 FILLER_41_1184 ();
 sg13g2_decap_8 FILLER_41_1191 ();
 sg13g2_decap_8 FILLER_41_1198 ();
 sg13g2_decap_8 FILLER_41_1205 ();
 sg13g2_decap_8 FILLER_41_1212 ();
 sg13g2_decap_8 FILLER_41_1219 ();
 sg13g2_decap_8 FILLER_41_1226 ();
 sg13g2_decap_8 FILLER_41_1233 ();
 sg13g2_decap_8 FILLER_41_1240 ();
 sg13g2_decap_8 FILLER_41_1247 ();
 sg13g2_decap_8 FILLER_41_1254 ();
 sg13g2_decap_8 FILLER_41_1261 ();
 sg13g2_decap_8 FILLER_41_1268 ();
 sg13g2_decap_8 FILLER_41_1275 ();
 sg13g2_decap_8 FILLER_41_1282 ();
 sg13g2_decap_8 FILLER_41_1289 ();
 sg13g2_decap_8 FILLER_41_1296 ();
 sg13g2_decap_8 FILLER_41_1303 ();
 sg13g2_decap_8 FILLER_41_1310 ();
 sg13g2_decap_8 FILLER_41_1317 ();
 sg13g2_decap_8 FILLER_41_1324 ();
 sg13g2_decap_8 FILLER_41_1331 ();
 sg13g2_decap_8 FILLER_41_1338 ();
 sg13g2_decap_8 FILLER_41_1345 ();
 sg13g2_decap_8 FILLER_41_1352 ();
 sg13g2_decap_8 FILLER_41_1359 ();
 sg13g2_decap_8 FILLER_41_1366 ();
 sg13g2_decap_8 FILLER_41_1373 ();
 sg13g2_decap_8 FILLER_41_1380 ();
 sg13g2_decap_8 FILLER_41_1387 ();
 sg13g2_decap_8 FILLER_41_1394 ();
 sg13g2_decap_8 FILLER_41_1401 ();
 sg13g2_decap_8 FILLER_41_1408 ();
 sg13g2_decap_8 FILLER_41_1415 ();
 sg13g2_decap_8 FILLER_41_1422 ();
 sg13g2_decap_8 FILLER_41_1429 ();
 sg13g2_decap_8 FILLER_41_1436 ();
 sg13g2_decap_8 FILLER_41_1443 ();
 sg13g2_decap_8 FILLER_41_1450 ();
 sg13g2_decap_8 FILLER_41_1457 ();
 sg13g2_decap_8 FILLER_41_1464 ();
 sg13g2_decap_8 FILLER_41_1471 ();
 sg13g2_decap_8 FILLER_41_1478 ();
 sg13g2_decap_8 FILLER_41_1485 ();
 sg13g2_decap_8 FILLER_41_1492 ();
 sg13g2_decap_8 FILLER_41_1499 ();
 sg13g2_decap_8 FILLER_41_1506 ();
 sg13g2_decap_8 FILLER_41_1513 ();
 sg13g2_decap_8 FILLER_41_1520 ();
 sg13g2_decap_8 FILLER_41_1527 ();
 sg13g2_decap_8 FILLER_41_1534 ();
 sg13g2_decap_8 FILLER_41_1541 ();
 sg13g2_decap_8 FILLER_41_1548 ();
 sg13g2_decap_8 FILLER_41_1555 ();
 sg13g2_decap_8 FILLER_41_1562 ();
 sg13g2_decap_8 FILLER_41_1569 ();
 sg13g2_decap_8 FILLER_41_1576 ();
 sg13g2_decap_8 FILLER_41_1583 ();
 sg13g2_decap_8 FILLER_41_1590 ();
 sg13g2_decap_8 FILLER_41_1597 ();
 sg13g2_decap_8 FILLER_41_1604 ();
 sg13g2_decap_8 FILLER_41_1611 ();
 sg13g2_decap_8 FILLER_41_1618 ();
 sg13g2_decap_8 FILLER_41_1625 ();
 sg13g2_decap_8 FILLER_41_1632 ();
 sg13g2_decap_8 FILLER_41_1639 ();
 sg13g2_decap_8 FILLER_41_1646 ();
 sg13g2_decap_8 FILLER_41_1653 ();
 sg13g2_decap_8 FILLER_41_1660 ();
 sg13g2_decap_8 FILLER_41_1667 ();
 sg13g2_decap_8 FILLER_41_1674 ();
 sg13g2_decap_8 FILLER_41_1681 ();
 sg13g2_decap_8 FILLER_41_1688 ();
 sg13g2_decap_8 FILLER_41_1695 ();
 sg13g2_decap_8 FILLER_41_1702 ();
 sg13g2_decap_8 FILLER_41_1709 ();
 sg13g2_decap_8 FILLER_41_1716 ();
 sg13g2_decap_8 FILLER_41_1723 ();
 sg13g2_decap_8 FILLER_41_1730 ();
 sg13g2_decap_8 FILLER_41_1737 ();
 sg13g2_decap_8 FILLER_41_1744 ();
 sg13g2_decap_8 FILLER_41_1751 ();
 sg13g2_decap_8 FILLER_41_1758 ();
 sg13g2_fill_2 FILLER_41_1765 ();
 sg13g2_fill_1 FILLER_41_1767 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_4 FILLER_42_56 ();
 sg13g2_fill_1 FILLER_42_86 ();
 sg13g2_fill_2 FILLER_42_96 ();
 sg13g2_fill_1 FILLER_42_98 ();
 sg13g2_fill_2 FILLER_42_145 ();
 sg13g2_fill_2 FILLER_42_204 ();
 sg13g2_fill_2 FILLER_42_212 ();
 sg13g2_fill_1 FILLER_42_214 ();
 sg13g2_decap_8 FILLER_42_221 ();
 sg13g2_decap_4 FILLER_42_228 ();
 sg13g2_fill_2 FILLER_42_232 ();
 sg13g2_fill_2 FILLER_42_239 ();
 sg13g2_decap_8 FILLER_42_258 ();
 sg13g2_fill_2 FILLER_42_289 ();
 sg13g2_fill_1 FILLER_42_291 ();
 sg13g2_fill_1 FILLER_42_302 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_fill_1 FILLER_42_322 ();
 sg13g2_fill_2 FILLER_42_349 ();
 sg13g2_fill_1 FILLER_42_351 ();
 sg13g2_fill_2 FILLER_42_365 ();
 sg13g2_fill_1 FILLER_42_367 ();
 sg13g2_fill_2 FILLER_42_377 ();
 sg13g2_fill_1 FILLER_42_425 ();
 sg13g2_fill_1 FILLER_42_440 ();
 sg13g2_fill_2 FILLER_42_464 ();
 sg13g2_fill_1 FILLER_42_466 ();
 sg13g2_fill_2 FILLER_42_505 ();
 sg13g2_fill_1 FILLER_42_507 ();
 sg13g2_fill_2 FILLER_42_513 ();
 sg13g2_fill_1 FILLER_42_523 ();
 sg13g2_fill_1 FILLER_42_567 ();
 sg13g2_fill_2 FILLER_42_573 ();
 sg13g2_decap_8 FILLER_42_583 ();
 sg13g2_decap_4 FILLER_42_590 ();
 sg13g2_fill_2 FILLER_42_594 ();
 sg13g2_decap_4 FILLER_42_609 ();
 sg13g2_fill_1 FILLER_42_626 ();
 sg13g2_decap_8 FILLER_42_650 ();
 sg13g2_fill_1 FILLER_42_657 ();
 sg13g2_decap_4 FILLER_42_674 ();
 sg13g2_fill_1 FILLER_42_678 ();
 sg13g2_decap_8 FILLER_42_684 ();
 sg13g2_fill_2 FILLER_42_691 ();
 sg13g2_decap_4 FILLER_42_700 ();
 sg13g2_fill_1 FILLER_42_704 ();
 sg13g2_decap_8 FILLER_42_729 ();
 sg13g2_decap_8 FILLER_42_736 ();
 sg13g2_decap_8 FILLER_42_743 ();
 sg13g2_fill_2 FILLER_42_750 ();
 sg13g2_fill_1 FILLER_42_770 ();
 sg13g2_fill_2 FILLER_42_812 ();
 sg13g2_decap_4 FILLER_42_859 ();
 sg13g2_fill_2 FILLER_42_863 ();
 sg13g2_fill_1 FILLER_42_875 ();
 sg13g2_fill_2 FILLER_42_889 ();
 sg13g2_fill_2 FILLER_42_904 ();
 sg13g2_decap_8 FILLER_42_937 ();
 sg13g2_decap_8 FILLER_42_944 ();
 sg13g2_decap_8 FILLER_42_951 ();
 sg13g2_fill_2 FILLER_42_958 ();
 sg13g2_decap_8 FILLER_42_965 ();
 sg13g2_decap_8 FILLER_42_972 ();
 sg13g2_decap_8 FILLER_42_979 ();
 sg13g2_fill_2 FILLER_42_986 ();
 sg13g2_fill_1 FILLER_42_988 ();
 sg13g2_decap_8 FILLER_42_993 ();
 sg13g2_decap_8 FILLER_42_1000 ();
 sg13g2_decap_8 FILLER_42_1007 ();
 sg13g2_decap_8 FILLER_42_1014 ();
 sg13g2_decap_8 FILLER_42_1021 ();
 sg13g2_decap_8 FILLER_42_1028 ();
 sg13g2_decap_8 FILLER_42_1035 ();
 sg13g2_decap_8 FILLER_42_1042 ();
 sg13g2_decap_8 FILLER_42_1049 ();
 sg13g2_decap_8 FILLER_42_1056 ();
 sg13g2_decap_8 FILLER_42_1063 ();
 sg13g2_decap_8 FILLER_42_1070 ();
 sg13g2_decap_8 FILLER_42_1077 ();
 sg13g2_decap_8 FILLER_42_1084 ();
 sg13g2_decap_8 FILLER_42_1091 ();
 sg13g2_decap_8 FILLER_42_1098 ();
 sg13g2_decap_8 FILLER_42_1105 ();
 sg13g2_decap_8 FILLER_42_1112 ();
 sg13g2_decap_8 FILLER_42_1119 ();
 sg13g2_decap_8 FILLER_42_1126 ();
 sg13g2_decap_8 FILLER_42_1133 ();
 sg13g2_decap_8 FILLER_42_1140 ();
 sg13g2_decap_8 FILLER_42_1147 ();
 sg13g2_decap_8 FILLER_42_1154 ();
 sg13g2_decap_8 FILLER_42_1161 ();
 sg13g2_decap_8 FILLER_42_1168 ();
 sg13g2_decap_8 FILLER_42_1175 ();
 sg13g2_decap_8 FILLER_42_1182 ();
 sg13g2_decap_8 FILLER_42_1189 ();
 sg13g2_decap_8 FILLER_42_1196 ();
 sg13g2_decap_8 FILLER_42_1203 ();
 sg13g2_decap_8 FILLER_42_1210 ();
 sg13g2_decap_8 FILLER_42_1217 ();
 sg13g2_decap_8 FILLER_42_1224 ();
 sg13g2_decap_8 FILLER_42_1231 ();
 sg13g2_decap_8 FILLER_42_1238 ();
 sg13g2_decap_8 FILLER_42_1245 ();
 sg13g2_decap_8 FILLER_42_1252 ();
 sg13g2_decap_8 FILLER_42_1259 ();
 sg13g2_decap_8 FILLER_42_1266 ();
 sg13g2_decap_8 FILLER_42_1273 ();
 sg13g2_decap_8 FILLER_42_1280 ();
 sg13g2_decap_8 FILLER_42_1287 ();
 sg13g2_decap_8 FILLER_42_1294 ();
 sg13g2_decap_8 FILLER_42_1301 ();
 sg13g2_decap_8 FILLER_42_1308 ();
 sg13g2_decap_8 FILLER_42_1315 ();
 sg13g2_decap_8 FILLER_42_1322 ();
 sg13g2_decap_8 FILLER_42_1329 ();
 sg13g2_decap_8 FILLER_42_1336 ();
 sg13g2_decap_8 FILLER_42_1343 ();
 sg13g2_decap_8 FILLER_42_1350 ();
 sg13g2_decap_8 FILLER_42_1357 ();
 sg13g2_decap_8 FILLER_42_1364 ();
 sg13g2_decap_8 FILLER_42_1371 ();
 sg13g2_decap_8 FILLER_42_1378 ();
 sg13g2_decap_8 FILLER_42_1385 ();
 sg13g2_decap_8 FILLER_42_1392 ();
 sg13g2_decap_8 FILLER_42_1399 ();
 sg13g2_decap_8 FILLER_42_1406 ();
 sg13g2_decap_8 FILLER_42_1413 ();
 sg13g2_decap_8 FILLER_42_1420 ();
 sg13g2_decap_8 FILLER_42_1427 ();
 sg13g2_decap_8 FILLER_42_1434 ();
 sg13g2_decap_8 FILLER_42_1441 ();
 sg13g2_decap_8 FILLER_42_1448 ();
 sg13g2_decap_8 FILLER_42_1455 ();
 sg13g2_decap_8 FILLER_42_1462 ();
 sg13g2_decap_8 FILLER_42_1469 ();
 sg13g2_decap_8 FILLER_42_1476 ();
 sg13g2_decap_8 FILLER_42_1483 ();
 sg13g2_decap_8 FILLER_42_1490 ();
 sg13g2_decap_8 FILLER_42_1497 ();
 sg13g2_decap_8 FILLER_42_1504 ();
 sg13g2_decap_8 FILLER_42_1511 ();
 sg13g2_decap_8 FILLER_42_1518 ();
 sg13g2_decap_8 FILLER_42_1525 ();
 sg13g2_decap_8 FILLER_42_1532 ();
 sg13g2_decap_8 FILLER_42_1539 ();
 sg13g2_decap_8 FILLER_42_1546 ();
 sg13g2_decap_8 FILLER_42_1553 ();
 sg13g2_decap_8 FILLER_42_1560 ();
 sg13g2_decap_8 FILLER_42_1567 ();
 sg13g2_decap_8 FILLER_42_1574 ();
 sg13g2_decap_8 FILLER_42_1581 ();
 sg13g2_decap_8 FILLER_42_1588 ();
 sg13g2_decap_8 FILLER_42_1595 ();
 sg13g2_decap_8 FILLER_42_1602 ();
 sg13g2_decap_8 FILLER_42_1609 ();
 sg13g2_decap_8 FILLER_42_1616 ();
 sg13g2_decap_8 FILLER_42_1623 ();
 sg13g2_decap_8 FILLER_42_1630 ();
 sg13g2_decap_8 FILLER_42_1637 ();
 sg13g2_decap_8 FILLER_42_1644 ();
 sg13g2_decap_8 FILLER_42_1651 ();
 sg13g2_decap_8 FILLER_42_1658 ();
 sg13g2_decap_8 FILLER_42_1665 ();
 sg13g2_decap_8 FILLER_42_1672 ();
 sg13g2_decap_8 FILLER_42_1679 ();
 sg13g2_decap_8 FILLER_42_1686 ();
 sg13g2_decap_8 FILLER_42_1693 ();
 sg13g2_decap_8 FILLER_42_1700 ();
 sg13g2_decap_8 FILLER_42_1707 ();
 sg13g2_decap_8 FILLER_42_1714 ();
 sg13g2_decap_8 FILLER_42_1721 ();
 sg13g2_decap_8 FILLER_42_1728 ();
 sg13g2_decap_8 FILLER_42_1735 ();
 sg13g2_decap_8 FILLER_42_1742 ();
 sg13g2_decap_8 FILLER_42_1749 ();
 sg13g2_decap_8 FILLER_42_1756 ();
 sg13g2_decap_4 FILLER_42_1763 ();
 sg13g2_fill_1 FILLER_42_1767 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_fill_1 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_27 ();
 sg13g2_decap_8 FILLER_43_34 ();
 sg13g2_decap_8 FILLER_43_41 ();
 sg13g2_fill_2 FILLER_43_48 ();
 sg13g2_fill_1 FILLER_43_59 ();
 sg13g2_decap_8 FILLER_43_64 ();
 sg13g2_decap_8 FILLER_43_71 ();
 sg13g2_decap_4 FILLER_43_78 ();
 sg13g2_decap_4 FILLER_43_125 ();
 sg13g2_fill_2 FILLER_43_129 ();
 sg13g2_decap_8 FILLER_43_167 ();
 sg13g2_decap_8 FILLER_43_174 ();
 sg13g2_fill_1 FILLER_43_181 ();
 sg13g2_fill_2 FILLER_43_193 ();
 sg13g2_decap_4 FILLER_43_204 ();
 sg13g2_fill_1 FILLER_43_208 ();
 sg13g2_decap_4 FILLER_43_229 ();
 sg13g2_fill_2 FILLER_43_233 ();
 sg13g2_fill_2 FILLER_43_250 ();
 sg13g2_decap_8 FILLER_43_260 ();
 sg13g2_fill_1 FILLER_43_267 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_fill_1 FILLER_43_301 ();
 sg13g2_decap_8 FILLER_43_318 ();
 sg13g2_decap_4 FILLER_43_325 ();
 sg13g2_fill_1 FILLER_43_329 ();
 sg13g2_fill_2 FILLER_43_334 ();
 sg13g2_fill_1 FILLER_43_336 ();
 sg13g2_fill_2 FILLER_43_348 ();
 sg13g2_fill_1 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_382 ();
 sg13g2_decap_8 FILLER_43_389 ();
 sg13g2_fill_2 FILLER_43_396 ();
 sg13g2_fill_1 FILLER_43_398 ();
 sg13g2_fill_2 FILLER_43_478 ();
 sg13g2_fill_1 FILLER_43_480 ();
 sg13g2_decap_4 FILLER_43_526 ();
 sg13g2_fill_2 FILLER_43_530 ();
 sg13g2_fill_1 FILLER_43_543 ();
 sg13g2_fill_2 FILLER_43_549 ();
 sg13g2_decap_4 FILLER_43_572 ();
 sg13g2_decap_8 FILLER_43_589 ();
 sg13g2_decap_8 FILLER_43_596 ();
 sg13g2_fill_2 FILLER_43_603 ();
 sg13g2_fill_1 FILLER_43_605 ();
 sg13g2_fill_2 FILLER_43_614 ();
 sg13g2_fill_2 FILLER_43_621 ();
 sg13g2_fill_1 FILLER_43_628 ();
 sg13g2_decap_4 FILLER_43_642 ();
 sg13g2_decap_8 FILLER_43_654 ();
 sg13g2_fill_1 FILLER_43_661 ();
 sg13g2_fill_2 FILLER_43_671 ();
 sg13g2_fill_1 FILLER_43_673 ();
 sg13g2_fill_1 FILLER_43_684 ();
 sg13g2_fill_2 FILLER_43_694 ();
 sg13g2_fill_1 FILLER_43_711 ();
 sg13g2_decap_4 FILLER_43_736 ();
 sg13g2_decap_4 FILLER_43_771 ();
 sg13g2_fill_1 FILLER_43_775 ();
 sg13g2_fill_2 FILLER_43_792 ();
 sg13g2_fill_1 FILLER_43_794 ();
 sg13g2_fill_1 FILLER_43_804 ();
 sg13g2_fill_1 FILLER_43_838 ();
 sg13g2_fill_2 FILLER_43_859 ();
 sg13g2_fill_2 FILLER_43_876 ();
 sg13g2_fill_1 FILLER_43_878 ();
 sg13g2_decap_8 FILLER_43_892 ();
 sg13g2_fill_2 FILLER_43_904 ();
 sg13g2_fill_2 FILLER_43_927 ();
 sg13g2_fill_1 FILLER_43_934 ();
 sg13g2_fill_2 FILLER_43_945 ();
 sg13g2_fill_1 FILLER_43_947 ();
 sg13g2_fill_2 FILLER_43_968 ();
 sg13g2_fill_1 FILLER_43_970 ();
 sg13g2_decap_8 FILLER_43_1017 ();
 sg13g2_decap_8 FILLER_43_1024 ();
 sg13g2_decap_8 FILLER_43_1031 ();
 sg13g2_decap_8 FILLER_43_1038 ();
 sg13g2_decap_8 FILLER_43_1045 ();
 sg13g2_decap_8 FILLER_43_1052 ();
 sg13g2_decap_8 FILLER_43_1059 ();
 sg13g2_decap_8 FILLER_43_1066 ();
 sg13g2_decap_8 FILLER_43_1073 ();
 sg13g2_decap_8 FILLER_43_1080 ();
 sg13g2_decap_8 FILLER_43_1087 ();
 sg13g2_decap_8 FILLER_43_1094 ();
 sg13g2_decap_8 FILLER_43_1101 ();
 sg13g2_decap_8 FILLER_43_1108 ();
 sg13g2_decap_8 FILLER_43_1115 ();
 sg13g2_decap_8 FILLER_43_1122 ();
 sg13g2_decap_8 FILLER_43_1129 ();
 sg13g2_decap_8 FILLER_43_1136 ();
 sg13g2_decap_8 FILLER_43_1143 ();
 sg13g2_decap_8 FILLER_43_1150 ();
 sg13g2_decap_8 FILLER_43_1157 ();
 sg13g2_decap_8 FILLER_43_1164 ();
 sg13g2_decap_8 FILLER_43_1171 ();
 sg13g2_decap_8 FILLER_43_1178 ();
 sg13g2_decap_8 FILLER_43_1185 ();
 sg13g2_decap_8 FILLER_43_1192 ();
 sg13g2_decap_8 FILLER_43_1199 ();
 sg13g2_decap_8 FILLER_43_1206 ();
 sg13g2_decap_8 FILLER_43_1213 ();
 sg13g2_decap_8 FILLER_43_1220 ();
 sg13g2_decap_8 FILLER_43_1227 ();
 sg13g2_decap_8 FILLER_43_1234 ();
 sg13g2_decap_8 FILLER_43_1241 ();
 sg13g2_decap_8 FILLER_43_1248 ();
 sg13g2_decap_8 FILLER_43_1255 ();
 sg13g2_decap_8 FILLER_43_1262 ();
 sg13g2_decap_8 FILLER_43_1269 ();
 sg13g2_decap_8 FILLER_43_1276 ();
 sg13g2_decap_8 FILLER_43_1283 ();
 sg13g2_decap_8 FILLER_43_1290 ();
 sg13g2_decap_8 FILLER_43_1297 ();
 sg13g2_decap_8 FILLER_43_1304 ();
 sg13g2_decap_8 FILLER_43_1311 ();
 sg13g2_decap_8 FILLER_43_1318 ();
 sg13g2_decap_8 FILLER_43_1325 ();
 sg13g2_decap_8 FILLER_43_1332 ();
 sg13g2_decap_8 FILLER_43_1339 ();
 sg13g2_decap_8 FILLER_43_1346 ();
 sg13g2_decap_8 FILLER_43_1353 ();
 sg13g2_decap_8 FILLER_43_1360 ();
 sg13g2_decap_8 FILLER_43_1367 ();
 sg13g2_decap_8 FILLER_43_1374 ();
 sg13g2_decap_8 FILLER_43_1381 ();
 sg13g2_decap_8 FILLER_43_1388 ();
 sg13g2_decap_8 FILLER_43_1395 ();
 sg13g2_decap_8 FILLER_43_1402 ();
 sg13g2_decap_8 FILLER_43_1409 ();
 sg13g2_decap_8 FILLER_43_1416 ();
 sg13g2_decap_8 FILLER_43_1423 ();
 sg13g2_decap_8 FILLER_43_1430 ();
 sg13g2_decap_8 FILLER_43_1437 ();
 sg13g2_decap_8 FILLER_43_1444 ();
 sg13g2_decap_8 FILLER_43_1451 ();
 sg13g2_decap_8 FILLER_43_1458 ();
 sg13g2_decap_8 FILLER_43_1465 ();
 sg13g2_decap_8 FILLER_43_1472 ();
 sg13g2_decap_8 FILLER_43_1479 ();
 sg13g2_decap_8 FILLER_43_1486 ();
 sg13g2_decap_8 FILLER_43_1493 ();
 sg13g2_decap_8 FILLER_43_1500 ();
 sg13g2_decap_8 FILLER_43_1507 ();
 sg13g2_decap_8 FILLER_43_1514 ();
 sg13g2_decap_8 FILLER_43_1521 ();
 sg13g2_decap_8 FILLER_43_1528 ();
 sg13g2_decap_8 FILLER_43_1535 ();
 sg13g2_decap_8 FILLER_43_1542 ();
 sg13g2_decap_8 FILLER_43_1549 ();
 sg13g2_decap_8 FILLER_43_1556 ();
 sg13g2_decap_8 FILLER_43_1563 ();
 sg13g2_decap_8 FILLER_43_1570 ();
 sg13g2_decap_8 FILLER_43_1577 ();
 sg13g2_decap_8 FILLER_43_1584 ();
 sg13g2_decap_8 FILLER_43_1591 ();
 sg13g2_decap_8 FILLER_43_1598 ();
 sg13g2_decap_8 FILLER_43_1605 ();
 sg13g2_decap_8 FILLER_43_1612 ();
 sg13g2_decap_8 FILLER_43_1619 ();
 sg13g2_decap_8 FILLER_43_1626 ();
 sg13g2_decap_8 FILLER_43_1633 ();
 sg13g2_decap_8 FILLER_43_1640 ();
 sg13g2_decap_8 FILLER_43_1647 ();
 sg13g2_decap_8 FILLER_43_1654 ();
 sg13g2_decap_8 FILLER_43_1661 ();
 sg13g2_decap_8 FILLER_43_1668 ();
 sg13g2_decap_8 FILLER_43_1675 ();
 sg13g2_decap_8 FILLER_43_1682 ();
 sg13g2_decap_8 FILLER_43_1689 ();
 sg13g2_decap_8 FILLER_43_1696 ();
 sg13g2_decap_8 FILLER_43_1703 ();
 sg13g2_decap_8 FILLER_43_1710 ();
 sg13g2_decap_8 FILLER_43_1717 ();
 sg13g2_decap_8 FILLER_43_1724 ();
 sg13g2_decap_8 FILLER_43_1731 ();
 sg13g2_decap_8 FILLER_43_1738 ();
 sg13g2_decap_8 FILLER_43_1745 ();
 sg13g2_decap_8 FILLER_43_1752 ();
 sg13g2_decap_8 FILLER_43_1759 ();
 sg13g2_fill_2 FILLER_43_1766 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_fill_1 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_37 ();
 sg13g2_fill_1 FILLER_44_44 ();
 sg13g2_decap_4 FILLER_44_79 ();
 sg13g2_fill_1 FILLER_44_83 ();
 sg13g2_fill_1 FILLER_44_108 ();
 sg13g2_fill_2 FILLER_44_114 ();
 sg13g2_fill_1 FILLER_44_116 ();
 sg13g2_decap_4 FILLER_44_121 ();
 sg13g2_decap_4 FILLER_44_135 ();
 sg13g2_fill_2 FILLER_44_144 ();
 sg13g2_decap_8 FILLER_44_181 ();
 sg13g2_fill_2 FILLER_44_218 ();
 sg13g2_decap_4 FILLER_44_243 ();
 sg13g2_fill_2 FILLER_44_247 ();
 sg13g2_fill_1 FILLER_44_284 ();
 sg13g2_decap_8 FILLER_44_295 ();
 sg13g2_fill_2 FILLER_44_302 ();
 sg13g2_fill_1 FILLER_44_304 ();
 sg13g2_decap_8 FILLER_44_324 ();
 sg13g2_fill_1 FILLER_44_331 ();
 sg13g2_fill_2 FILLER_44_367 ();
 sg13g2_fill_1 FILLER_44_403 ();
 sg13g2_fill_2 FILLER_44_430 ();
 sg13g2_fill_1 FILLER_44_441 ();
 sg13g2_fill_1 FILLER_44_459 ();
 sg13g2_decap_4 FILLER_44_469 ();
 sg13g2_fill_1 FILLER_44_489 ();
 sg13g2_fill_1 FILLER_44_520 ();
 sg13g2_decap_8 FILLER_44_543 ();
 sg13g2_decap_4 FILLER_44_550 ();
 sg13g2_fill_2 FILLER_44_554 ();
 sg13g2_decap_4 FILLER_44_571 ();
 sg13g2_decap_8 FILLER_44_591 ();
 sg13g2_decap_4 FILLER_44_598 ();
 sg13g2_fill_2 FILLER_44_602 ();
 sg13g2_fill_2 FILLER_44_616 ();
 sg13g2_fill_1 FILLER_44_618 ();
 sg13g2_decap_4 FILLER_44_658 ();
 sg13g2_fill_1 FILLER_44_682 ();
 sg13g2_fill_2 FILLER_44_705 ();
 sg13g2_decap_8 FILLER_44_740 ();
 sg13g2_decap_4 FILLER_44_747 ();
 sg13g2_decap_4 FILLER_44_759 ();
 sg13g2_decap_4 FILLER_44_813 ();
 sg13g2_fill_1 FILLER_44_817 ();
 sg13g2_fill_2 FILLER_44_835 ();
 sg13g2_fill_1 FILLER_44_837 ();
 sg13g2_fill_2 FILLER_44_867 ();
 sg13g2_decap_4 FILLER_44_874 ();
 sg13g2_fill_1 FILLER_44_878 ();
 sg13g2_decap_8 FILLER_44_883 ();
 sg13g2_decap_8 FILLER_44_890 ();
 sg13g2_decap_8 FILLER_44_915 ();
 sg13g2_decap_4 FILLER_44_922 ();
 sg13g2_fill_2 FILLER_44_926 ();
 sg13g2_decap_4 FILLER_44_932 ();
 sg13g2_fill_1 FILLER_44_936 ();
 sg13g2_decap_4 FILLER_44_947 ();
 sg13g2_decap_8 FILLER_44_963 ();
 sg13g2_decap_4 FILLER_44_975 ();
 sg13g2_fill_1 FILLER_44_979 ();
 sg13g2_fill_1 FILLER_44_1001 ();
 sg13g2_decap_8 FILLER_44_1023 ();
 sg13g2_decap_8 FILLER_44_1030 ();
 sg13g2_decap_8 FILLER_44_1037 ();
 sg13g2_decap_8 FILLER_44_1044 ();
 sg13g2_decap_8 FILLER_44_1051 ();
 sg13g2_decap_8 FILLER_44_1058 ();
 sg13g2_decap_8 FILLER_44_1065 ();
 sg13g2_decap_8 FILLER_44_1072 ();
 sg13g2_decap_8 FILLER_44_1079 ();
 sg13g2_decap_8 FILLER_44_1086 ();
 sg13g2_decap_8 FILLER_44_1093 ();
 sg13g2_decap_8 FILLER_44_1100 ();
 sg13g2_decap_8 FILLER_44_1107 ();
 sg13g2_decap_8 FILLER_44_1114 ();
 sg13g2_decap_8 FILLER_44_1121 ();
 sg13g2_decap_8 FILLER_44_1128 ();
 sg13g2_decap_8 FILLER_44_1135 ();
 sg13g2_decap_8 FILLER_44_1142 ();
 sg13g2_decap_8 FILLER_44_1149 ();
 sg13g2_decap_8 FILLER_44_1156 ();
 sg13g2_decap_8 FILLER_44_1163 ();
 sg13g2_decap_8 FILLER_44_1170 ();
 sg13g2_decap_8 FILLER_44_1177 ();
 sg13g2_decap_8 FILLER_44_1184 ();
 sg13g2_decap_8 FILLER_44_1191 ();
 sg13g2_decap_8 FILLER_44_1198 ();
 sg13g2_decap_8 FILLER_44_1205 ();
 sg13g2_decap_8 FILLER_44_1212 ();
 sg13g2_decap_8 FILLER_44_1219 ();
 sg13g2_decap_8 FILLER_44_1226 ();
 sg13g2_decap_8 FILLER_44_1233 ();
 sg13g2_decap_8 FILLER_44_1240 ();
 sg13g2_decap_8 FILLER_44_1247 ();
 sg13g2_decap_8 FILLER_44_1254 ();
 sg13g2_decap_8 FILLER_44_1261 ();
 sg13g2_decap_8 FILLER_44_1268 ();
 sg13g2_decap_8 FILLER_44_1275 ();
 sg13g2_decap_8 FILLER_44_1282 ();
 sg13g2_decap_8 FILLER_44_1289 ();
 sg13g2_decap_8 FILLER_44_1296 ();
 sg13g2_decap_8 FILLER_44_1303 ();
 sg13g2_decap_8 FILLER_44_1310 ();
 sg13g2_decap_8 FILLER_44_1317 ();
 sg13g2_decap_8 FILLER_44_1324 ();
 sg13g2_decap_8 FILLER_44_1331 ();
 sg13g2_decap_8 FILLER_44_1338 ();
 sg13g2_decap_8 FILLER_44_1345 ();
 sg13g2_decap_8 FILLER_44_1352 ();
 sg13g2_decap_8 FILLER_44_1359 ();
 sg13g2_decap_8 FILLER_44_1366 ();
 sg13g2_decap_8 FILLER_44_1373 ();
 sg13g2_decap_8 FILLER_44_1380 ();
 sg13g2_decap_8 FILLER_44_1387 ();
 sg13g2_decap_8 FILLER_44_1394 ();
 sg13g2_decap_8 FILLER_44_1401 ();
 sg13g2_decap_8 FILLER_44_1408 ();
 sg13g2_decap_8 FILLER_44_1415 ();
 sg13g2_decap_8 FILLER_44_1422 ();
 sg13g2_decap_8 FILLER_44_1429 ();
 sg13g2_decap_8 FILLER_44_1436 ();
 sg13g2_decap_8 FILLER_44_1443 ();
 sg13g2_decap_8 FILLER_44_1450 ();
 sg13g2_decap_8 FILLER_44_1457 ();
 sg13g2_decap_8 FILLER_44_1464 ();
 sg13g2_decap_8 FILLER_44_1471 ();
 sg13g2_decap_8 FILLER_44_1478 ();
 sg13g2_decap_8 FILLER_44_1485 ();
 sg13g2_decap_8 FILLER_44_1492 ();
 sg13g2_decap_8 FILLER_44_1499 ();
 sg13g2_decap_8 FILLER_44_1506 ();
 sg13g2_decap_8 FILLER_44_1513 ();
 sg13g2_decap_8 FILLER_44_1520 ();
 sg13g2_decap_8 FILLER_44_1527 ();
 sg13g2_decap_8 FILLER_44_1534 ();
 sg13g2_decap_8 FILLER_44_1541 ();
 sg13g2_decap_8 FILLER_44_1548 ();
 sg13g2_decap_8 FILLER_44_1555 ();
 sg13g2_decap_8 FILLER_44_1562 ();
 sg13g2_decap_8 FILLER_44_1569 ();
 sg13g2_decap_8 FILLER_44_1576 ();
 sg13g2_decap_8 FILLER_44_1583 ();
 sg13g2_decap_8 FILLER_44_1590 ();
 sg13g2_decap_8 FILLER_44_1597 ();
 sg13g2_decap_8 FILLER_44_1604 ();
 sg13g2_decap_8 FILLER_44_1611 ();
 sg13g2_decap_8 FILLER_44_1618 ();
 sg13g2_decap_8 FILLER_44_1625 ();
 sg13g2_decap_8 FILLER_44_1632 ();
 sg13g2_decap_8 FILLER_44_1639 ();
 sg13g2_decap_8 FILLER_44_1646 ();
 sg13g2_decap_8 FILLER_44_1653 ();
 sg13g2_decap_8 FILLER_44_1660 ();
 sg13g2_decap_8 FILLER_44_1667 ();
 sg13g2_decap_8 FILLER_44_1674 ();
 sg13g2_decap_8 FILLER_44_1681 ();
 sg13g2_decap_8 FILLER_44_1688 ();
 sg13g2_decap_8 FILLER_44_1695 ();
 sg13g2_decap_8 FILLER_44_1702 ();
 sg13g2_decap_8 FILLER_44_1709 ();
 sg13g2_decap_8 FILLER_44_1716 ();
 sg13g2_decap_8 FILLER_44_1723 ();
 sg13g2_decap_8 FILLER_44_1730 ();
 sg13g2_decap_8 FILLER_44_1737 ();
 sg13g2_decap_8 FILLER_44_1744 ();
 sg13g2_decap_8 FILLER_44_1751 ();
 sg13g2_decap_8 FILLER_44_1758 ();
 sg13g2_fill_2 FILLER_44_1765 ();
 sg13g2_fill_1 FILLER_44_1767 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_27 ();
 sg13g2_decap_4 FILLER_45_38 ();
 sg13g2_fill_2 FILLER_45_57 ();
 sg13g2_fill_1 FILLER_45_74 ();
 sg13g2_decap_4 FILLER_45_85 ();
 sg13g2_decap_8 FILLER_45_93 ();
 sg13g2_fill_1 FILLER_45_107 ();
 sg13g2_fill_2 FILLER_45_121 ();
 sg13g2_fill_1 FILLER_45_123 ();
 sg13g2_fill_1 FILLER_45_131 ();
 sg13g2_fill_2 FILLER_45_153 ();
 sg13g2_fill_1 FILLER_45_155 ();
 sg13g2_fill_1 FILLER_45_202 ();
 sg13g2_fill_1 FILLER_45_233 ();
 sg13g2_decap_4 FILLER_45_253 ();
 sg13g2_fill_2 FILLER_45_262 ();
 sg13g2_fill_1 FILLER_45_264 ();
 sg13g2_fill_1 FILLER_45_270 ();
 sg13g2_decap_4 FILLER_45_280 ();
 sg13g2_fill_1 FILLER_45_284 ();
 sg13g2_fill_2 FILLER_45_300 ();
 sg13g2_fill_1 FILLER_45_302 ();
 sg13g2_fill_1 FILLER_45_313 ();
 sg13g2_fill_1 FILLER_45_324 ();
 sg13g2_fill_2 FILLER_45_361 ();
 sg13g2_fill_2 FILLER_45_387 ();
 sg13g2_fill_2 FILLER_45_394 ();
 sg13g2_fill_1 FILLER_45_417 ();
 sg13g2_fill_1 FILLER_45_431 ();
 sg13g2_decap_4 FILLER_45_458 ();
 sg13g2_fill_1 FILLER_45_462 ();
 sg13g2_decap_8 FILLER_45_504 ();
 sg13g2_fill_1 FILLER_45_511 ();
 sg13g2_fill_1 FILLER_45_521 ();
 sg13g2_fill_2 FILLER_45_535 ();
 sg13g2_fill_1 FILLER_45_537 ();
 sg13g2_decap_4 FILLER_45_552 ();
 sg13g2_fill_2 FILLER_45_575 ();
 sg13g2_fill_2 FILLER_45_588 ();
 sg13g2_fill_1 FILLER_45_590 ();
 sg13g2_fill_2 FILLER_45_596 ();
 sg13g2_fill_1 FILLER_45_603 ();
 sg13g2_decap_8 FILLER_45_609 ();
 sg13g2_decap_8 FILLER_45_616 ();
 sg13g2_fill_1 FILLER_45_623 ();
 sg13g2_fill_1 FILLER_45_635 ();
 sg13g2_decap_4 FILLER_45_654 ();
 sg13g2_fill_1 FILLER_45_658 ();
 sg13g2_decap_8 FILLER_45_664 ();
 sg13g2_fill_1 FILLER_45_671 ();
 sg13g2_decap_4 FILLER_45_696 ();
 sg13g2_fill_2 FILLER_45_700 ();
 sg13g2_decap_8 FILLER_45_730 ();
 sg13g2_fill_2 FILLER_45_737 ();
 sg13g2_fill_1 FILLER_45_739 ();
 sg13g2_decap_4 FILLER_45_766 ();
 sg13g2_fill_1 FILLER_45_770 ();
 sg13g2_decap_8 FILLER_45_775 ();
 sg13g2_decap_8 FILLER_45_782 ();
 sg13g2_fill_1 FILLER_45_789 ();
 sg13g2_fill_2 FILLER_45_807 ();
 sg13g2_fill_1 FILLER_45_809 ();
 sg13g2_fill_2 FILLER_45_836 ();
 sg13g2_fill_2 FILLER_45_848 ();
 sg13g2_fill_1 FILLER_45_850 ();
 sg13g2_fill_2 FILLER_45_859 ();
 sg13g2_fill_2 FILLER_45_875 ();
 sg13g2_fill_1 FILLER_45_877 ();
 sg13g2_fill_2 FILLER_45_890 ();
 sg13g2_fill_1 FILLER_45_892 ();
 sg13g2_decap_4 FILLER_45_926 ();
 sg13g2_fill_1 FILLER_45_930 ();
 sg13g2_decap_4 FILLER_45_943 ();
 sg13g2_fill_1 FILLER_45_947 ();
 sg13g2_decap_8 FILLER_45_961 ();
 sg13g2_fill_2 FILLER_45_976 ();
 sg13g2_decap_8 FILLER_45_983 ();
 sg13g2_fill_2 FILLER_45_990 ();
 sg13g2_fill_1 FILLER_45_992 ();
 sg13g2_fill_2 FILLER_45_998 ();
 sg13g2_fill_1 FILLER_45_1000 ();
 sg13g2_decap_8 FILLER_45_1030 ();
 sg13g2_decap_8 FILLER_45_1037 ();
 sg13g2_decap_8 FILLER_45_1044 ();
 sg13g2_decap_8 FILLER_45_1051 ();
 sg13g2_decap_8 FILLER_45_1058 ();
 sg13g2_decap_8 FILLER_45_1065 ();
 sg13g2_decap_8 FILLER_45_1072 ();
 sg13g2_decap_8 FILLER_45_1079 ();
 sg13g2_decap_8 FILLER_45_1086 ();
 sg13g2_decap_8 FILLER_45_1093 ();
 sg13g2_decap_8 FILLER_45_1100 ();
 sg13g2_decap_8 FILLER_45_1107 ();
 sg13g2_decap_8 FILLER_45_1114 ();
 sg13g2_decap_8 FILLER_45_1121 ();
 sg13g2_decap_8 FILLER_45_1128 ();
 sg13g2_decap_8 FILLER_45_1135 ();
 sg13g2_decap_8 FILLER_45_1142 ();
 sg13g2_decap_8 FILLER_45_1149 ();
 sg13g2_decap_8 FILLER_45_1156 ();
 sg13g2_decap_8 FILLER_45_1163 ();
 sg13g2_decap_8 FILLER_45_1170 ();
 sg13g2_decap_8 FILLER_45_1177 ();
 sg13g2_decap_8 FILLER_45_1184 ();
 sg13g2_decap_8 FILLER_45_1191 ();
 sg13g2_decap_8 FILLER_45_1198 ();
 sg13g2_decap_8 FILLER_45_1205 ();
 sg13g2_decap_8 FILLER_45_1212 ();
 sg13g2_decap_8 FILLER_45_1219 ();
 sg13g2_decap_8 FILLER_45_1226 ();
 sg13g2_decap_8 FILLER_45_1233 ();
 sg13g2_decap_8 FILLER_45_1240 ();
 sg13g2_decap_8 FILLER_45_1247 ();
 sg13g2_decap_8 FILLER_45_1254 ();
 sg13g2_decap_8 FILLER_45_1261 ();
 sg13g2_decap_8 FILLER_45_1268 ();
 sg13g2_decap_8 FILLER_45_1275 ();
 sg13g2_decap_8 FILLER_45_1282 ();
 sg13g2_decap_8 FILLER_45_1289 ();
 sg13g2_decap_8 FILLER_45_1296 ();
 sg13g2_decap_8 FILLER_45_1303 ();
 sg13g2_decap_8 FILLER_45_1310 ();
 sg13g2_decap_8 FILLER_45_1317 ();
 sg13g2_decap_8 FILLER_45_1324 ();
 sg13g2_decap_8 FILLER_45_1331 ();
 sg13g2_decap_8 FILLER_45_1338 ();
 sg13g2_decap_8 FILLER_45_1345 ();
 sg13g2_decap_8 FILLER_45_1352 ();
 sg13g2_decap_8 FILLER_45_1359 ();
 sg13g2_decap_8 FILLER_45_1366 ();
 sg13g2_decap_8 FILLER_45_1373 ();
 sg13g2_decap_8 FILLER_45_1380 ();
 sg13g2_decap_8 FILLER_45_1387 ();
 sg13g2_decap_8 FILLER_45_1394 ();
 sg13g2_decap_8 FILLER_45_1401 ();
 sg13g2_decap_8 FILLER_45_1408 ();
 sg13g2_decap_8 FILLER_45_1415 ();
 sg13g2_decap_8 FILLER_45_1422 ();
 sg13g2_decap_8 FILLER_45_1429 ();
 sg13g2_decap_8 FILLER_45_1436 ();
 sg13g2_decap_8 FILLER_45_1443 ();
 sg13g2_decap_8 FILLER_45_1450 ();
 sg13g2_decap_8 FILLER_45_1457 ();
 sg13g2_decap_8 FILLER_45_1464 ();
 sg13g2_decap_8 FILLER_45_1471 ();
 sg13g2_decap_8 FILLER_45_1478 ();
 sg13g2_decap_8 FILLER_45_1485 ();
 sg13g2_decap_8 FILLER_45_1492 ();
 sg13g2_decap_8 FILLER_45_1499 ();
 sg13g2_decap_8 FILLER_45_1506 ();
 sg13g2_decap_8 FILLER_45_1513 ();
 sg13g2_decap_8 FILLER_45_1520 ();
 sg13g2_decap_8 FILLER_45_1527 ();
 sg13g2_decap_8 FILLER_45_1534 ();
 sg13g2_decap_8 FILLER_45_1541 ();
 sg13g2_decap_8 FILLER_45_1548 ();
 sg13g2_decap_8 FILLER_45_1555 ();
 sg13g2_decap_8 FILLER_45_1562 ();
 sg13g2_decap_8 FILLER_45_1569 ();
 sg13g2_decap_8 FILLER_45_1576 ();
 sg13g2_decap_8 FILLER_45_1583 ();
 sg13g2_decap_8 FILLER_45_1590 ();
 sg13g2_decap_8 FILLER_45_1597 ();
 sg13g2_decap_8 FILLER_45_1604 ();
 sg13g2_decap_8 FILLER_45_1611 ();
 sg13g2_decap_8 FILLER_45_1618 ();
 sg13g2_decap_8 FILLER_45_1625 ();
 sg13g2_decap_8 FILLER_45_1632 ();
 sg13g2_decap_8 FILLER_45_1639 ();
 sg13g2_decap_8 FILLER_45_1646 ();
 sg13g2_decap_8 FILLER_45_1653 ();
 sg13g2_decap_8 FILLER_45_1660 ();
 sg13g2_decap_8 FILLER_45_1667 ();
 sg13g2_decap_8 FILLER_45_1674 ();
 sg13g2_decap_8 FILLER_45_1681 ();
 sg13g2_decap_8 FILLER_45_1688 ();
 sg13g2_decap_8 FILLER_45_1695 ();
 sg13g2_decap_8 FILLER_45_1702 ();
 sg13g2_decap_8 FILLER_45_1709 ();
 sg13g2_decap_8 FILLER_45_1716 ();
 sg13g2_decap_8 FILLER_45_1723 ();
 sg13g2_decap_8 FILLER_45_1730 ();
 sg13g2_decap_8 FILLER_45_1737 ();
 sg13g2_decap_8 FILLER_45_1744 ();
 sg13g2_decap_8 FILLER_45_1751 ();
 sg13g2_decap_8 FILLER_45_1758 ();
 sg13g2_fill_2 FILLER_45_1765 ();
 sg13g2_fill_1 FILLER_45_1767 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_4 ();
 sg13g2_decap_8 FILLER_46_36 ();
 sg13g2_decap_4 FILLER_46_43 ();
 sg13g2_fill_1 FILLER_46_47 ();
 sg13g2_fill_2 FILLER_46_54 ();
 sg13g2_fill_1 FILLER_46_56 ();
 sg13g2_fill_2 FILLER_46_61 ();
 sg13g2_fill_1 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_73 ();
 sg13g2_decap_8 FILLER_46_80 ();
 sg13g2_decap_8 FILLER_46_87 ();
 sg13g2_fill_2 FILLER_46_103 ();
 sg13g2_fill_1 FILLER_46_113 ();
 sg13g2_decap_8 FILLER_46_118 ();
 sg13g2_fill_2 FILLER_46_125 ();
 sg13g2_fill_2 FILLER_46_136 ();
 sg13g2_fill_1 FILLER_46_155 ();
 sg13g2_fill_1 FILLER_46_165 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_fill_1 FILLER_46_189 ();
 sg13g2_fill_2 FILLER_46_203 ();
 sg13g2_fill_1 FILLER_46_205 ();
 sg13g2_fill_2 FILLER_46_216 ();
 sg13g2_fill_2 FILLER_46_244 ();
 sg13g2_fill_1 FILLER_46_246 ();
 sg13g2_decap_4 FILLER_46_257 ();
 sg13g2_decap_8 FILLER_46_297 ();
 sg13g2_fill_2 FILLER_46_323 ();
 sg13g2_fill_1 FILLER_46_325 ();
 sg13g2_fill_2 FILLER_46_368 ();
 sg13g2_fill_2 FILLER_46_461 ();
 sg13g2_fill_1 FILLER_46_463 ();
 sg13g2_decap_8 FILLER_46_474 ();
 sg13g2_fill_2 FILLER_46_481 ();
 sg13g2_fill_1 FILLER_46_483 ();
 sg13g2_fill_2 FILLER_46_510 ();
 sg13g2_fill_1 FILLER_46_512 ();
 sg13g2_fill_2 FILLER_46_532 ();
 sg13g2_fill_1 FILLER_46_534 ();
 sg13g2_decap_8 FILLER_46_540 ();
 sg13g2_decap_8 FILLER_46_547 ();
 sg13g2_fill_2 FILLER_46_559 ();
 sg13g2_fill_1 FILLER_46_561 ();
 sg13g2_fill_1 FILLER_46_566 ();
 sg13g2_fill_2 FILLER_46_571 ();
 sg13g2_decap_4 FILLER_46_577 ();
 sg13g2_fill_2 FILLER_46_581 ();
 sg13g2_fill_2 FILLER_46_609 ();
 sg13g2_fill_1 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_627 ();
 sg13g2_fill_1 FILLER_46_634 ();
 sg13g2_fill_1 FILLER_46_638 ();
 sg13g2_decap_4 FILLER_46_643 ();
 sg13g2_fill_1 FILLER_46_647 ();
 sg13g2_fill_1 FILLER_46_653 ();
 sg13g2_fill_2 FILLER_46_663 ();
 sg13g2_decap_8 FILLER_46_670 ();
 sg13g2_fill_1 FILLER_46_677 ();
 sg13g2_fill_2 FILLER_46_698 ();
 sg13g2_decap_8 FILLER_46_724 ();
 sg13g2_fill_1 FILLER_46_731 ();
 sg13g2_fill_2 FILLER_46_819 ();
 sg13g2_decap_4 FILLER_46_851 ();
 sg13g2_fill_1 FILLER_46_855 ();
 sg13g2_decap_8 FILLER_46_866 ();
 sg13g2_fill_1 FILLER_46_893 ();
 sg13g2_fill_1 FILLER_46_898 ();
 sg13g2_fill_2 FILLER_46_909 ();
 sg13g2_fill_2 FILLER_46_915 ();
 sg13g2_fill_1 FILLER_46_917 ();
 sg13g2_fill_1 FILLER_46_928 ();
 sg13g2_fill_2 FILLER_46_940 ();
 sg13g2_fill_1 FILLER_46_942 ();
 sg13g2_fill_1 FILLER_46_960 ();
 sg13g2_fill_2 FILLER_46_986 ();
 sg13g2_fill_1 FILLER_46_988 ();
 sg13g2_decap_8 FILLER_46_997 ();
 sg13g2_decap_8 FILLER_46_1004 ();
 sg13g2_decap_8 FILLER_46_1011 ();
 sg13g2_decap_8 FILLER_46_1031 ();
 sg13g2_decap_8 FILLER_46_1038 ();
 sg13g2_decap_8 FILLER_46_1045 ();
 sg13g2_decap_8 FILLER_46_1052 ();
 sg13g2_decap_8 FILLER_46_1059 ();
 sg13g2_decap_8 FILLER_46_1066 ();
 sg13g2_decap_8 FILLER_46_1073 ();
 sg13g2_decap_8 FILLER_46_1080 ();
 sg13g2_decap_8 FILLER_46_1087 ();
 sg13g2_decap_8 FILLER_46_1094 ();
 sg13g2_decap_8 FILLER_46_1101 ();
 sg13g2_decap_8 FILLER_46_1108 ();
 sg13g2_decap_8 FILLER_46_1115 ();
 sg13g2_decap_8 FILLER_46_1122 ();
 sg13g2_decap_8 FILLER_46_1129 ();
 sg13g2_decap_8 FILLER_46_1136 ();
 sg13g2_decap_8 FILLER_46_1143 ();
 sg13g2_decap_8 FILLER_46_1150 ();
 sg13g2_decap_8 FILLER_46_1157 ();
 sg13g2_decap_8 FILLER_46_1164 ();
 sg13g2_decap_8 FILLER_46_1171 ();
 sg13g2_decap_8 FILLER_46_1178 ();
 sg13g2_decap_8 FILLER_46_1185 ();
 sg13g2_decap_8 FILLER_46_1192 ();
 sg13g2_decap_8 FILLER_46_1199 ();
 sg13g2_decap_8 FILLER_46_1206 ();
 sg13g2_decap_8 FILLER_46_1213 ();
 sg13g2_decap_8 FILLER_46_1220 ();
 sg13g2_decap_8 FILLER_46_1227 ();
 sg13g2_decap_8 FILLER_46_1234 ();
 sg13g2_decap_8 FILLER_46_1241 ();
 sg13g2_decap_8 FILLER_46_1248 ();
 sg13g2_decap_8 FILLER_46_1255 ();
 sg13g2_decap_8 FILLER_46_1262 ();
 sg13g2_decap_8 FILLER_46_1269 ();
 sg13g2_decap_8 FILLER_46_1276 ();
 sg13g2_decap_8 FILLER_46_1283 ();
 sg13g2_decap_8 FILLER_46_1290 ();
 sg13g2_decap_8 FILLER_46_1297 ();
 sg13g2_decap_8 FILLER_46_1304 ();
 sg13g2_decap_8 FILLER_46_1311 ();
 sg13g2_decap_8 FILLER_46_1318 ();
 sg13g2_decap_8 FILLER_46_1325 ();
 sg13g2_decap_8 FILLER_46_1332 ();
 sg13g2_decap_8 FILLER_46_1339 ();
 sg13g2_decap_8 FILLER_46_1346 ();
 sg13g2_decap_8 FILLER_46_1353 ();
 sg13g2_decap_8 FILLER_46_1360 ();
 sg13g2_decap_8 FILLER_46_1367 ();
 sg13g2_decap_8 FILLER_46_1374 ();
 sg13g2_decap_8 FILLER_46_1381 ();
 sg13g2_decap_8 FILLER_46_1388 ();
 sg13g2_decap_8 FILLER_46_1395 ();
 sg13g2_decap_8 FILLER_46_1402 ();
 sg13g2_decap_8 FILLER_46_1409 ();
 sg13g2_decap_8 FILLER_46_1416 ();
 sg13g2_decap_8 FILLER_46_1423 ();
 sg13g2_decap_8 FILLER_46_1430 ();
 sg13g2_decap_8 FILLER_46_1437 ();
 sg13g2_decap_8 FILLER_46_1444 ();
 sg13g2_decap_8 FILLER_46_1451 ();
 sg13g2_decap_8 FILLER_46_1458 ();
 sg13g2_decap_8 FILLER_46_1465 ();
 sg13g2_decap_8 FILLER_46_1472 ();
 sg13g2_decap_8 FILLER_46_1479 ();
 sg13g2_decap_8 FILLER_46_1486 ();
 sg13g2_decap_8 FILLER_46_1493 ();
 sg13g2_decap_8 FILLER_46_1500 ();
 sg13g2_decap_8 FILLER_46_1507 ();
 sg13g2_decap_8 FILLER_46_1514 ();
 sg13g2_decap_8 FILLER_46_1521 ();
 sg13g2_decap_8 FILLER_46_1528 ();
 sg13g2_decap_8 FILLER_46_1535 ();
 sg13g2_decap_8 FILLER_46_1542 ();
 sg13g2_decap_8 FILLER_46_1549 ();
 sg13g2_decap_8 FILLER_46_1556 ();
 sg13g2_decap_8 FILLER_46_1563 ();
 sg13g2_decap_8 FILLER_46_1570 ();
 sg13g2_decap_8 FILLER_46_1577 ();
 sg13g2_decap_8 FILLER_46_1584 ();
 sg13g2_decap_8 FILLER_46_1591 ();
 sg13g2_decap_8 FILLER_46_1598 ();
 sg13g2_decap_8 FILLER_46_1605 ();
 sg13g2_decap_8 FILLER_46_1612 ();
 sg13g2_decap_8 FILLER_46_1619 ();
 sg13g2_decap_8 FILLER_46_1626 ();
 sg13g2_decap_8 FILLER_46_1633 ();
 sg13g2_decap_8 FILLER_46_1640 ();
 sg13g2_decap_8 FILLER_46_1647 ();
 sg13g2_decap_8 FILLER_46_1654 ();
 sg13g2_decap_8 FILLER_46_1661 ();
 sg13g2_decap_8 FILLER_46_1668 ();
 sg13g2_decap_8 FILLER_46_1675 ();
 sg13g2_decap_8 FILLER_46_1682 ();
 sg13g2_decap_8 FILLER_46_1689 ();
 sg13g2_decap_8 FILLER_46_1696 ();
 sg13g2_decap_8 FILLER_46_1703 ();
 sg13g2_decap_8 FILLER_46_1710 ();
 sg13g2_decap_8 FILLER_46_1717 ();
 sg13g2_decap_8 FILLER_46_1724 ();
 sg13g2_decap_8 FILLER_46_1731 ();
 sg13g2_decap_8 FILLER_46_1738 ();
 sg13g2_decap_8 FILLER_46_1745 ();
 sg13g2_decap_8 FILLER_46_1752 ();
 sg13g2_decap_8 FILLER_46_1759 ();
 sg13g2_fill_2 FILLER_46_1766 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_7 ();
 sg13g2_fill_1 FILLER_47_12 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_fill_1 FILLER_47_65 ();
 sg13g2_fill_2 FILLER_47_82 ();
 sg13g2_fill_1 FILLER_47_84 ();
 sg13g2_decap_4 FILLER_47_127 ();
 sg13g2_fill_2 FILLER_47_131 ();
 sg13g2_fill_2 FILLER_47_149 ();
 sg13g2_fill_1 FILLER_47_151 ();
 sg13g2_fill_2 FILLER_47_188 ();
 sg13g2_decap_8 FILLER_47_237 ();
 sg13g2_fill_2 FILLER_47_244 ();
 sg13g2_fill_1 FILLER_47_246 ();
 sg13g2_fill_1 FILLER_47_286 ();
 sg13g2_decap_4 FILLER_47_320 ();
 sg13g2_decap_4 FILLER_47_331 ();
 sg13g2_fill_2 FILLER_47_335 ();
 sg13g2_decap_8 FILLER_47_460 ();
 sg13g2_decap_8 FILLER_47_467 ();
 sg13g2_fill_2 FILLER_47_474 ();
 sg13g2_fill_2 FILLER_47_484 ();
 sg13g2_fill_1 FILLER_47_486 ();
 sg13g2_decap_8 FILLER_47_501 ();
 sg13g2_decap_4 FILLER_47_508 ();
 sg13g2_fill_2 FILLER_47_512 ();
 sg13g2_decap_4 FILLER_47_528 ();
 sg13g2_fill_1 FILLER_47_532 ();
 sg13g2_fill_1 FILLER_47_536 ();
 sg13g2_fill_2 FILLER_47_559 ();
 sg13g2_fill_2 FILLER_47_571 ();
 sg13g2_fill_2 FILLER_47_585 ();
 sg13g2_fill_2 FILLER_47_597 ();
 sg13g2_decap_8 FILLER_47_604 ();
 sg13g2_decap_8 FILLER_47_611 ();
 sg13g2_decap_4 FILLER_47_623 ();
 sg13g2_fill_2 FILLER_47_627 ();
 sg13g2_fill_2 FILLER_47_654 ();
 sg13g2_fill_1 FILLER_47_656 ();
 sg13g2_decap_4 FILLER_47_662 ();
 sg13g2_decap_4 FILLER_47_670 ();
 sg13g2_fill_1 FILLER_47_682 ();
 sg13g2_decap_8 FILLER_47_703 ();
 sg13g2_decap_8 FILLER_47_720 ();
 sg13g2_fill_2 FILLER_47_737 ();
 sg13g2_fill_1 FILLER_47_739 ();
 sg13g2_fill_2 FILLER_47_784 ();
 sg13g2_fill_1 FILLER_47_786 ();
 sg13g2_decap_4 FILLER_47_795 ();
 sg13g2_fill_1 FILLER_47_803 ();
 sg13g2_decap_4 FILLER_47_844 ();
 sg13g2_decap_8 FILLER_47_869 ();
 sg13g2_fill_2 FILLER_47_884 ();
 sg13g2_fill_1 FILLER_47_894 ();
 sg13g2_decap_4 FILLER_47_942 ();
 sg13g2_fill_2 FILLER_47_970 ();
 sg13g2_decap_4 FILLER_47_980 ();
 sg13g2_fill_2 FILLER_47_984 ();
 sg13g2_fill_2 FILLER_47_997 ();
 sg13g2_fill_1 FILLER_47_999 ();
 sg13g2_decap_4 FILLER_47_1008 ();
 sg13g2_decap_8 FILLER_47_1030 ();
 sg13g2_decap_8 FILLER_47_1037 ();
 sg13g2_decap_8 FILLER_47_1044 ();
 sg13g2_decap_8 FILLER_47_1051 ();
 sg13g2_decap_8 FILLER_47_1058 ();
 sg13g2_decap_8 FILLER_47_1065 ();
 sg13g2_decap_8 FILLER_47_1072 ();
 sg13g2_decap_8 FILLER_47_1079 ();
 sg13g2_decap_8 FILLER_47_1086 ();
 sg13g2_decap_8 FILLER_47_1093 ();
 sg13g2_decap_8 FILLER_47_1100 ();
 sg13g2_decap_8 FILLER_47_1107 ();
 sg13g2_decap_8 FILLER_47_1114 ();
 sg13g2_decap_8 FILLER_47_1121 ();
 sg13g2_decap_8 FILLER_47_1128 ();
 sg13g2_decap_8 FILLER_47_1135 ();
 sg13g2_decap_8 FILLER_47_1142 ();
 sg13g2_decap_8 FILLER_47_1149 ();
 sg13g2_decap_8 FILLER_47_1156 ();
 sg13g2_decap_8 FILLER_47_1163 ();
 sg13g2_decap_8 FILLER_47_1170 ();
 sg13g2_decap_8 FILLER_47_1177 ();
 sg13g2_decap_8 FILLER_47_1184 ();
 sg13g2_decap_8 FILLER_47_1191 ();
 sg13g2_decap_8 FILLER_47_1198 ();
 sg13g2_decap_8 FILLER_47_1205 ();
 sg13g2_decap_8 FILLER_47_1212 ();
 sg13g2_decap_8 FILLER_47_1219 ();
 sg13g2_decap_8 FILLER_47_1226 ();
 sg13g2_decap_8 FILLER_47_1233 ();
 sg13g2_decap_8 FILLER_47_1240 ();
 sg13g2_decap_8 FILLER_47_1247 ();
 sg13g2_decap_8 FILLER_47_1254 ();
 sg13g2_decap_8 FILLER_47_1261 ();
 sg13g2_decap_8 FILLER_47_1268 ();
 sg13g2_decap_8 FILLER_47_1275 ();
 sg13g2_decap_8 FILLER_47_1282 ();
 sg13g2_decap_8 FILLER_47_1289 ();
 sg13g2_decap_8 FILLER_47_1296 ();
 sg13g2_decap_8 FILLER_47_1303 ();
 sg13g2_decap_8 FILLER_47_1310 ();
 sg13g2_decap_8 FILLER_47_1317 ();
 sg13g2_decap_8 FILLER_47_1324 ();
 sg13g2_decap_8 FILLER_47_1331 ();
 sg13g2_decap_8 FILLER_47_1338 ();
 sg13g2_decap_8 FILLER_47_1345 ();
 sg13g2_decap_8 FILLER_47_1352 ();
 sg13g2_decap_8 FILLER_47_1359 ();
 sg13g2_decap_8 FILLER_47_1366 ();
 sg13g2_decap_8 FILLER_47_1373 ();
 sg13g2_decap_8 FILLER_47_1380 ();
 sg13g2_decap_8 FILLER_47_1387 ();
 sg13g2_decap_8 FILLER_47_1394 ();
 sg13g2_decap_8 FILLER_47_1401 ();
 sg13g2_decap_8 FILLER_47_1408 ();
 sg13g2_decap_8 FILLER_47_1415 ();
 sg13g2_decap_8 FILLER_47_1422 ();
 sg13g2_decap_8 FILLER_47_1429 ();
 sg13g2_decap_8 FILLER_47_1436 ();
 sg13g2_decap_8 FILLER_47_1443 ();
 sg13g2_decap_8 FILLER_47_1450 ();
 sg13g2_decap_8 FILLER_47_1457 ();
 sg13g2_decap_8 FILLER_47_1464 ();
 sg13g2_decap_8 FILLER_47_1471 ();
 sg13g2_decap_8 FILLER_47_1478 ();
 sg13g2_decap_8 FILLER_47_1485 ();
 sg13g2_decap_8 FILLER_47_1492 ();
 sg13g2_decap_8 FILLER_47_1499 ();
 sg13g2_decap_8 FILLER_47_1506 ();
 sg13g2_decap_8 FILLER_47_1513 ();
 sg13g2_decap_8 FILLER_47_1520 ();
 sg13g2_decap_8 FILLER_47_1527 ();
 sg13g2_decap_8 FILLER_47_1534 ();
 sg13g2_decap_8 FILLER_47_1541 ();
 sg13g2_decap_8 FILLER_47_1548 ();
 sg13g2_decap_8 FILLER_47_1555 ();
 sg13g2_decap_8 FILLER_47_1562 ();
 sg13g2_decap_8 FILLER_47_1569 ();
 sg13g2_decap_8 FILLER_47_1576 ();
 sg13g2_decap_8 FILLER_47_1583 ();
 sg13g2_decap_8 FILLER_47_1590 ();
 sg13g2_decap_8 FILLER_47_1597 ();
 sg13g2_decap_8 FILLER_47_1604 ();
 sg13g2_decap_8 FILLER_47_1611 ();
 sg13g2_decap_8 FILLER_47_1618 ();
 sg13g2_decap_8 FILLER_47_1625 ();
 sg13g2_decap_8 FILLER_47_1632 ();
 sg13g2_decap_8 FILLER_47_1639 ();
 sg13g2_decap_8 FILLER_47_1646 ();
 sg13g2_decap_8 FILLER_47_1653 ();
 sg13g2_decap_8 FILLER_47_1660 ();
 sg13g2_decap_8 FILLER_47_1667 ();
 sg13g2_decap_8 FILLER_47_1674 ();
 sg13g2_decap_8 FILLER_47_1681 ();
 sg13g2_decap_8 FILLER_47_1688 ();
 sg13g2_decap_8 FILLER_47_1695 ();
 sg13g2_decap_8 FILLER_47_1702 ();
 sg13g2_decap_8 FILLER_47_1709 ();
 sg13g2_decap_8 FILLER_47_1716 ();
 sg13g2_decap_8 FILLER_47_1723 ();
 sg13g2_decap_8 FILLER_47_1730 ();
 sg13g2_decap_8 FILLER_47_1737 ();
 sg13g2_decap_8 FILLER_47_1744 ();
 sg13g2_decap_8 FILLER_47_1751 ();
 sg13g2_decap_8 FILLER_47_1758 ();
 sg13g2_fill_2 FILLER_47_1765 ();
 sg13g2_fill_1 FILLER_47_1767 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_37 ();
 sg13g2_fill_2 FILLER_48_44 ();
 sg13g2_fill_1 FILLER_48_57 ();
 sg13g2_decap_4 FILLER_48_63 ();
 sg13g2_fill_2 FILLER_48_67 ();
 sg13g2_fill_2 FILLER_48_92 ();
 sg13g2_fill_2 FILLER_48_102 ();
 sg13g2_fill_1 FILLER_48_108 ();
 sg13g2_decap_4 FILLER_48_114 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_fill_2 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_155 ();
 sg13g2_decap_8 FILLER_48_162 ();
 sg13g2_decap_4 FILLER_48_191 ();
 sg13g2_fill_1 FILLER_48_195 ();
 sg13g2_decap_4 FILLER_48_205 ();
 sg13g2_fill_2 FILLER_48_209 ();
 sg13g2_fill_2 FILLER_48_244 ();
 sg13g2_fill_2 FILLER_48_263 ();
 sg13g2_fill_1 FILLER_48_272 ();
 sg13g2_decap_4 FILLER_48_294 ();
 sg13g2_fill_1 FILLER_48_298 ();
 sg13g2_fill_2 FILLER_48_324 ();
 sg13g2_fill_1 FILLER_48_359 ();
 sg13g2_fill_2 FILLER_48_377 ();
 sg13g2_fill_2 FILLER_48_409 ();
 sg13g2_decap_8 FILLER_48_456 ();
 sg13g2_decap_4 FILLER_48_463 ();
 sg13g2_fill_1 FILLER_48_467 ();
 sg13g2_fill_2 FILLER_48_500 ();
 sg13g2_fill_1 FILLER_48_502 ();
 sg13g2_fill_2 FILLER_48_517 ();
 sg13g2_fill_1 FILLER_48_519 ();
 sg13g2_decap_8 FILLER_48_529 ();
 sg13g2_decap_8 FILLER_48_547 ();
 sg13g2_decap_4 FILLER_48_554 ();
 sg13g2_fill_1 FILLER_48_566 ();
 sg13g2_fill_2 FILLER_48_576 ();
 sg13g2_decap_8 FILLER_48_583 ();
 sg13g2_decap_4 FILLER_48_600 ();
 sg13g2_decap_8 FILLER_48_615 ();
 sg13g2_decap_4 FILLER_48_622 ();
 sg13g2_decap_4 FILLER_48_636 ();
 sg13g2_fill_2 FILLER_48_640 ();
 sg13g2_fill_2 FILLER_48_645 ();
 sg13g2_fill_1 FILLER_48_647 ();
 sg13g2_fill_2 FILLER_48_657 ();
 sg13g2_decap_4 FILLER_48_664 ();
 sg13g2_fill_1 FILLER_48_668 ();
 sg13g2_decap_4 FILLER_48_694 ();
 sg13g2_fill_1 FILLER_48_698 ();
 sg13g2_fill_2 FILLER_48_720 ();
 sg13g2_fill_1 FILLER_48_722 ();
 sg13g2_fill_1 FILLER_48_743 ();
 sg13g2_fill_2 FILLER_48_771 ();
 sg13g2_fill_1 FILLER_48_773 ();
 sg13g2_fill_1 FILLER_48_779 ();
 sg13g2_decap_4 FILLER_48_789 ();
 sg13g2_fill_2 FILLER_48_793 ();
 sg13g2_decap_4 FILLER_48_799 ();
 sg13g2_fill_1 FILLER_48_803 ();
 sg13g2_decap_4 FILLER_48_809 ();
 sg13g2_fill_2 FILLER_48_820 ();
 sg13g2_decap_4 FILLER_48_852 ();
 sg13g2_fill_2 FILLER_48_856 ();
 sg13g2_decap_8 FILLER_48_869 ();
 sg13g2_decap_8 FILLER_48_876 ();
 sg13g2_decap_8 FILLER_48_883 ();
 sg13g2_decap_8 FILLER_48_890 ();
 sg13g2_decap_4 FILLER_48_897 ();
 sg13g2_fill_1 FILLER_48_926 ();
 sg13g2_fill_2 FILLER_48_953 ();
 sg13g2_fill_2 FILLER_48_984 ();
 sg13g2_decap_4 FILLER_48_1010 ();
 sg13g2_decap_8 FILLER_48_1035 ();
 sg13g2_decap_8 FILLER_48_1042 ();
 sg13g2_decap_8 FILLER_48_1049 ();
 sg13g2_decap_8 FILLER_48_1056 ();
 sg13g2_decap_8 FILLER_48_1063 ();
 sg13g2_decap_8 FILLER_48_1070 ();
 sg13g2_decap_8 FILLER_48_1077 ();
 sg13g2_decap_8 FILLER_48_1084 ();
 sg13g2_decap_8 FILLER_48_1091 ();
 sg13g2_decap_8 FILLER_48_1098 ();
 sg13g2_decap_8 FILLER_48_1105 ();
 sg13g2_decap_8 FILLER_48_1112 ();
 sg13g2_decap_8 FILLER_48_1119 ();
 sg13g2_decap_8 FILLER_48_1126 ();
 sg13g2_decap_8 FILLER_48_1133 ();
 sg13g2_decap_8 FILLER_48_1140 ();
 sg13g2_decap_8 FILLER_48_1147 ();
 sg13g2_decap_8 FILLER_48_1154 ();
 sg13g2_decap_8 FILLER_48_1161 ();
 sg13g2_decap_8 FILLER_48_1168 ();
 sg13g2_decap_8 FILLER_48_1175 ();
 sg13g2_decap_8 FILLER_48_1182 ();
 sg13g2_decap_8 FILLER_48_1189 ();
 sg13g2_decap_8 FILLER_48_1196 ();
 sg13g2_decap_8 FILLER_48_1203 ();
 sg13g2_decap_8 FILLER_48_1210 ();
 sg13g2_decap_8 FILLER_48_1217 ();
 sg13g2_decap_8 FILLER_48_1224 ();
 sg13g2_decap_8 FILLER_48_1231 ();
 sg13g2_decap_8 FILLER_48_1238 ();
 sg13g2_decap_8 FILLER_48_1245 ();
 sg13g2_decap_8 FILLER_48_1252 ();
 sg13g2_decap_8 FILLER_48_1259 ();
 sg13g2_decap_8 FILLER_48_1266 ();
 sg13g2_decap_8 FILLER_48_1273 ();
 sg13g2_decap_8 FILLER_48_1280 ();
 sg13g2_decap_8 FILLER_48_1287 ();
 sg13g2_decap_8 FILLER_48_1294 ();
 sg13g2_decap_8 FILLER_48_1301 ();
 sg13g2_decap_8 FILLER_48_1308 ();
 sg13g2_decap_8 FILLER_48_1315 ();
 sg13g2_decap_8 FILLER_48_1322 ();
 sg13g2_decap_8 FILLER_48_1329 ();
 sg13g2_decap_8 FILLER_48_1336 ();
 sg13g2_decap_8 FILLER_48_1343 ();
 sg13g2_decap_8 FILLER_48_1350 ();
 sg13g2_decap_8 FILLER_48_1357 ();
 sg13g2_decap_8 FILLER_48_1364 ();
 sg13g2_decap_8 FILLER_48_1371 ();
 sg13g2_decap_8 FILLER_48_1378 ();
 sg13g2_decap_8 FILLER_48_1385 ();
 sg13g2_decap_8 FILLER_48_1392 ();
 sg13g2_decap_8 FILLER_48_1399 ();
 sg13g2_decap_8 FILLER_48_1406 ();
 sg13g2_decap_8 FILLER_48_1413 ();
 sg13g2_decap_8 FILLER_48_1420 ();
 sg13g2_decap_8 FILLER_48_1427 ();
 sg13g2_decap_8 FILLER_48_1434 ();
 sg13g2_decap_8 FILLER_48_1441 ();
 sg13g2_decap_8 FILLER_48_1448 ();
 sg13g2_decap_8 FILLER_48_1455 ();
 sg13g2_decap_8 FILLER_48_1462 ();
 sg13g2_decap_8 FILLER_48_1469 ();
 sg13g2_decap_8 FILLER_48_1476 ();
 sg13g2_decap_8 FILLER_48_1483 ();
 sg13g2_decap_8 FILLER_48_1490 ();
 sg13g2_decap_8 FILLER_48_1497 ();
 sg13g2_decap_8 FILLER_48_1504 ();
 sg13g2_decap_8 FILLER_48_1511 ();
 sg13g2_decap_8 FILLER_48_1518 ();
 sg13g2_decap_8 FILLER_48_1525 ();
 sg13g2_decap_8 FILLER_48_1532 ();
 sg13g2_decap_8 FILLER_48_1539 ();
 sg13g2_decap_8 FILLER_48_1546 ();
 sg13g2_decap_8 FILLER_48_1553 ();
 sg13g2_decap_8 FILLER_48_1560 ();
 sg13g2_decap_8 FILLER_48_1567 ();
 sg13g2_decap_8 FILLER_48_1574 ();
 sg13g2_decap_8 FILLER_48_1581 ();
 sg13g2_decap_8 FILLER_48_1588 ();
 sg13g2_decap_8 FILLER_48_1595 ();
 sg13g2_decap_8 FILLER_48_1602 ();
 sg13g2_decap_8 FILLER_48_1609 ();
 sg13g2_decap_8 FILLER_48_1616 ();
 sg13g2_decap_8 FILLER_48_1623 ();
 sg13g2_decap_8 FILLER_48_1630 ();
 sg13g2_decap_8 FILLER_48_1637 ();
 sg13g2_decap_8 FILLER_48_1644 ();
 sg13g2_decap_8 FILLER_48_1651 ();
 sg13g2_decap_8 FILLER_48_1658 ();
 sg13g2_decap_8 FILLER_48_1665 ();
 sg13g2_decap_8 FILLER_48_1672 ();
 sg13g2_decap_8 FILLER_48_1679 ();
 sg13g2_decap_8 FILLER_48_1686 ();
 sg13g2_decap_8 FILLER_48_1693 ();
 sg13g2_decap_8 FILLER_48_1700 ();
 sg13g2_decap_8 FILLER_48_1707 ();
 sg13g2_decap_8 FILLER_48_1714 ();
 sg13g2_decap_8 FILLER_48_1721 ();
 sg13g2_decap_8 FILLER_48_1728 ();
 sg13g2_decap_8 FILLER_48_1735 ();
 sg13g2_decap_8 FILLER_48_1742 ();
 sg13g2_decap_8 FILLER_48_1749 ();
 sg13g2_decap_8 FILLER_48_1756 ();
 sg13g2_decap_4 FILLER_48_1763 ();
 sg13g2_fill_1 FILLER_48_1767 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_7 ();
 sg13g2_fill_1 FILLER_49_9 ();
 sg13g2_decap_4 FILLER_49_31 ();
 sg13g2_fill_2 FILLER_49_35 ();
 sg13g2_fill_2 FILLER_49_78 ();
 sg13g2_fill_1 FILLER_49_80 ();
 sg13g2_fill_2 FILLER_49_91 ();
 sg13g2_fill_1 FILLER_49_93 ();
 sg13g2_fill_2 FILLER_49_99 ();
 sg13g2_decap_8 FILLER_49_114 ();
 sg13g2_fill_2 FILLER_49_121 ();
 sg13g2_fill_1 FILLER_49_123 ();
 sg13g2_fill_1 FILLER_49_146 ();
 sg13g2_decap_8 FILLER_49_152 ();
 sg13g2_fill_2 FILLER_49_159 ();
 sg13g2_fill_2 FILLER_49_169 ();
 sg13g2_fill_2 FILLER_49_179 ();
 sg13g2_fill_1 FILLER_49_181 ();
 sg13g2_fill_1 FILLER_49_192 ();
 sg13g2_fill_2 FILLER_49_211 ();
 sg13g2_fill_1 FILLER_49_213 ();
 sg13g2_fill_2 FILLER_49_338 ();
 sg13g2_fill_1 FILLER_49_349 ();
 sg13g2_fill_2 FILLER_49_387 ();
 sg13g2_fill_1 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_49_464 ();
 sg13g2_fill_2 FILLER_49_471 ();
 sg13g2_fill_1 FILLER_49_495 ();
 sg13g2_fill_1 FILLER_49_520 ();
 sg13g2_decap_8 FILLER_49_537 ();
 sg13g2_fill_2 FILLER_49_544 ();
 sg13g2_fill_1 FILLER_49_546 ();
 sg13g2_fill_1 FILLER_49_576 ();
 sg13g2_fill_1 FILLER_49_592 ();
 sg13g2_fill_2 FILLER_49_609 ();
 sg13g2_fill_1 FILLER_49_611 ();
 sg13g2_decap_4 FILLER_49_643 ();
 sg13g2_fill_2 FILLER_49_647 ();
 sg13g2_fill_2 FILLER_49_670 ();
 sg13g2_fill_2 FILLER_49_690 ();
 sg13g2_fill_1 FILLER_49_692 ();
 sg13g2_fill_2 FILLER_49_706 ();
 sg13g2_decap_8 FILLER_49_718 ();
 sg13g2_fill_2 FILLER_49_725 ();
 sg13g2_fill_1 FILLER_49_737 ();
 sg13g2_fill_1 FILLER_49_751 ();
 sg13g2_fill_1 FILLER_49_778 ();
 sg13g2_fill_1 FILLER_49_810 ();
 sg13g2_fill_1 FILLER_49_830 ();
 sg13g2_fill_2 FILLER_49_849 ();
 sg13g2_fill_1 FILLER_49_851 ();
 sg13g2_decap_8 FILLER_49_861 ();
 sg13g2_fill_2 FILLER_49_868 ();
 sg13g2_fill_1 FILLER_49_870 ();
 sg13g2_fill_2 FILLER_49_880 ();
 sg13g2_decap_8 FILLER_49_910 ();
 sg13g2_fill_2 FILLER_49_917 ();
 sg13g2_decap_8 FILLER_49_938 ();
 sg13g2_decap_8 FILLER_49_945 ();
 sg13g2_fill_1 FILLER_49_956 ();
 sg13g2_fill_2 FILLER_49_976 ();
 sg13g2_decap_4 FILLER_49_997 ();
 sg13g2_decap_4 FILLER_49_1006 ();
 sg13g2_decap_8 FILLER_49_1038 ();
 sg13g2_decap_8 FILLER_49_1045 ();
 sg13g2_decap_8 FILLER_49_1052 ();
 sg13g2_decap_8 FILLER_49_1059 ();
 sg13g2_decap_8 FILLER_49_1066 ();
 sg13g2_decap_8 FILLER_49_1073 ();
 sg13g2_decap_8 FILLER_49_1080 ();
 sg13g2_decap_8 FILLER_49_1087 ();
 sg13g2_decap_8 FILLER_49_1094 ();
 sg13g2_decap_8 FILLER_49_1101 ();
 sg13g2_decap_8 FILLER_49_1108 ();
 sg13g2_decap_8 FILLER_49_1115 ();
 sg13g2_decap_8 FILLER_49_1122 ();
 sg13g2_decap_8 FILLER_49_1129 ();
 sg13g2_decap_8 FILLER_49_1136 ();
 sg13g2_decap_8 FILLER_49_1143 ();
 sg13g2_decap_8 FILLER_49_1150 ();
 sg13g2_decap_8 FILLER_49_1157 ();
 sg13g2_decap_8 FILLER_49_1164 ();
 sg13g2_decap_8 FILLER_49_1171 ();
 sg13g2_decap_8 FILLER_49_1178 ();
 sg13g2_decap_8 FILLER_49_1185 ();
 sg13g2_decap_8 FILLER_49_1192 ();
 sg13g2_decap_8 FILLER_49_1199 ();
 sg13g2_decap_8 FILLER_49_1206 ();
 sg13g2_decap_8 FILLER_49_1213 ();
 sg13g2_decap_8 FILLER_49_1220 ();
 sg13g2_decap_8 FILLER_49_1227 ();
 sg13g2_decap_8 FILLER_49_1234 ();
 sg13g2_decap_8 FILLER_49_1241 ();
 sg13g2_decap_8 FILLER_49_1248 ();
 sg13g2_decap_8 FILLER_49_1255 ();
 sg13g2_decap_8 FILLER_49_1262 ();
 sg13g2_decap_8 FILLER_49_1269 ();
 sg13g2_decap_8 FILLER_49_1276 ();
 sg13g2_decap_8 FILLER_49_1283 ();
 sg13g2_decap_8 FILLER_49_1290 ();
 sg13g2_decap_8 FILLER_49_1297 ();
 sg13g2_decap_8 FILLER_49_1304 ();
 sg13g2_decap_8 FILLER_49_1311 ();
 sg13g2_decap_8 FILLER_49_1318 ();
 sg13g2_decap_8 FILLER_49_1325 ();
 sg13g2_decap_8 FILLER_49_1332 ();
 sg13g2_decap_8 FILLER_49_1339 ();
 sg13g2_decap_8 FILLER_49_1346 ();
 sg13g2_decap_8 FILLER_49_1353 ();
 sg13g2_decap_8 FILLER_49_1360 ();
 sg13g2_decap_8 FILLER_49_1367 ();
 sg13g2_decap_8 FILLER_49_1374 ();
 sg13g2_decap_8 FILLER_49_1381 ();
 sg13g2_decap_8 FILLER_49_1388 ();
 sg13g2_decap_8 FILLER_49_1395 ();
 sg13g2_decap_8 FILLER_49_1402 ();
 sg13g2_decap_8 FILLER_49_1409 ();
 sg13g2_decap_8 FILLER_49_1416 ();
 sg13g2_decap_8 FILLER_49_1423 ();
 sg13g2_decap_8 FILLER_49_1430 ();
 sg13g2_decap_8 FILLER_49_1437 ();
 sg13g2_decap_8 FILLER_49_1444 ();
 sg13g2_decap_8 FILLER_49_1451 ();
 sg13g2_decap_8 FILLER_49_1458 ();
 sg13g2_decap_8 FILLER_49_1465 ();
 sg13g2_decap_8 FILLER_49_1472 ();
 sg13g2_decap_8 FILLER_49_1479 ();
 sg13g2_decap_8 FILLER_49_1486 ();
 sg13g2_decap_8 FILLER_49_1493 ();
 sg13g2_decap_8 FILLER_49_1500 ();
 sg13g2_decap_8 FILLER_49_1507 ();
 sg13g2_decap_8 FILLER_49_1514 ();
 sg13g2_decap_8 FILLER_49_1521 ();
 sg13g2_decap_8 FILLER_49_1528 ();
 sg13g2_decap_8 FILLER_49_1535 ();
 sg13g2_decap_8 FILLER_49_1542 ();
 sg13g2_decap_8 FILLER_49_1549 ();
 sg13g2_decap_8 FILLER_49_1556 ();
 sg13g2_decap_8 FILLER_49_1563 ();
 sg13g2_decap_8 FILLER_49_1570 ();
 sg13g2_decap_8 FILLER_49_1577 ();
 sg13g2_decap_8 FILLER_49_1584 ();
 sg13g2_decap_8 FILLER_49_1591 ();
 sg13g2_decap_8 FILLER_49_1598 ();
 sg13g2_decap_8 FILLER_49_1605 ();
 sg13g2_decap_8 FILLER_49_1612 ();
 sg13g2_decap_8 FILLER_49_1619 ();
 sg13g2_decap_8 FILLER_49_1626 ();
 sg13g2_decap_8 FILLER_49_1633 ();
 sg13g2_decap_8 FILLER_49_1640 ();
 sg13g2_decap_8 FILLER_49_1647 ();
 sg13g2_decap_8 FILLER_49_1654 ();
 sg13g2_decap_8 FILLER_49_1661 ();
 sg13g2_decap_8 FILLER_49_1668 ();
 sg13g2_decap_8 FILLER_49_1675 ();
 sg13g2_decap_8 FILLER_49_1682 ();
 sg13g2_decap_8 FILLER_49_1689 ();
 sg13g2_decap_8 FILLER_49_1696 ();
 sg13g2_decap_8 FILLER_49_1703 ();
 sg13g2_decap_8 FILLER_49_1710 ();
 sg13g2_decap_8 FILLER_49_1717 ();
 sg13g2_decap_8 FILLER_49_1724 ();
 sg13g2_decap_8 FILLER_49_1731 ();
 sg13g2_decap_8 FILLER_49_1738 ();
 sg13g2_decap_8 FILLER_49_1745 ();
 sg13g2_decap_8 FILLER_49_1752 ();
 sg13g2_decap_8 FILLER_49_1759 ();
 sg13g2_fill_2 FILLER_49_1766 ();
 sg13g2_decap_4 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_28 ();
 sg13g2_fill_1 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_53 ();
 sg13g2_decap_8 FILLER_50_60 ();
 sg13g2_decap_4 FILLER_50_67 ();
 sg13g2_fill_1 FILLER_50_71 ();
 sg13g2_fill_1 FILLER_50_81 ();
 sg13g2_decap_4 FILLER_50_122 ();
 sg13g2_fill_1 FILLER_50_126 ();
 sg13g2_fill_2 FILLER_50_183 ();
 sg13g2_fill_2 FILLER_50_195 ();
 sg13g2_fill_1 FILLER_50_197 ();
 sg13g2_fill_1 FILLER_50_207 ();
 sg13g2_decap_8 FILLER_50_220 ();
 sg13g2_fill_1 FILLER_50_227 ();
 sg13g2_decap_8 FILLER_50_233 ();
 sg13g2_decap_4 FILLER_50_254 ();
 sg13g2_decap_4 FILLER_50_263 ();
 sg13g2_decap_8 FILLER_50_273 ();
 sg13g2_decap_8 FILLER_50_280 ();
 sg13g2_fill_2 FILLER_50_287 ();
 sg13g2_fill_1 FILLER_50_289 ();
 sg13g2_fill_2 FILLER_50_297 ();
 sg13g2_decap_4 FILLER_50_312 ();
 sg13g2_fill_1 FILLER_50_316 ();
 sg13g2_fill_2 FILLER_50_405 ();
 sg13g2_fill_1 FILLER_50_407 ();
 sg13g2_fill_1 FILLER_50_432 ();
 sg13g2_decap_8 FILLER_50_442 ();
 sg13g2_fill_1 FILLER_50_453 ();
 sg13g2_fill_2 FILLER_50_460 ();
 sg13g2_fill_1 FILLER_50_462 ();
 sg13g2_decap_8 FILLER_50_469 ();
 sg13g2_fill_1 FILLER_50_476 ();
 sg13g2_fill_1 FILLER_50_483 ();
 sg13g2_decap_8 FILLER_50_489 ();
 sg13g2_decap_4 FILLER_50_496 ();
 sg13g2_decap_8 FILLER_50_528 ();
 sg13g2_decap_8 FILLER_50_535 ();
 sg13g2_fill_1 FILLER_50_542 ();
 sg13g2_decap_8 FILLER_50_553 ();
 sg13g2_decap_8 FILLER_50_560 ();
 sg13g2_fill_1 FILLER_50_590 ();
 sg13g2_fill_1 FILLER_50_604 ();
 sg13g2_fill_2 FILLER_50_609 ();
 sg13g2_fill_1 FILLER_50_611 ();
 sg13g2_fill_2 FILLER_50_616 ();
 sg13g2_decap_8 FILLER_50_638 ();
 sg13g2_decap_4 FILLER_50_645 ();
 sg13g2_fill_1 FILLER_50_649 ();
 sg13g2_decap_4 FILLER_50_658 ();
 sg13g2_decap_8 FILLER_50_667 ();
 sg13g2_fill_1 FILLER_50_674 ();
 sg13g2_decap_4 FILLER_50_685 ();
 sg13g2_fill_2 FILLER_50_719 ();
 sg13g2_fill_1 FILLER_50_721 ();
 sg13g2_decap_8 FILLER_50_775 ();
 sg13g2_fill_2 FILLER_50_782 ();
 sg13g2_fill_2 FILLER_50_789 ();
 sg13g2_fill_1 FILLER_50_791 ();
 sg13g2_fill_2 FILLER_50_796 ();
 sg13g2_fill_2 FILLER_50_811 ();
 sg13g2_fill_1 FILLER_50_827 ();
 sg13g2_fill_1 FILLER_50_858 ();
 sg13g2_decap_8 FILLER_50_893 ();
 sg13g2_fill_2 FILLER_50_900 ();
 sg13g2_decap_8 FILLER_50_910 ();
 sg13g2_decap_8 FILLER_50_938 ();
 sg13g2_fill_1 FILLER_50_961 ();
 sg13g2_decap_8 FILLER_50_967 ();
 sg13g2_decap_8 FILLER_50_974 ();
 sg13g2_decap_8 FILLER_50_981 ();
 sg13g2_decap_8 FILLER_50_1003 ();
 sg13g2_decap_8 FILLER_50_1010 ();
 sg13g2_decap_8 FILLER_50_1043 ();
 sg13g2_decap_8 FILLER_50_1050 ();
 sg13g2_decap_8 FILLER_50_1057 ();
 sg13g2_decap_8 FILLER_50_1064 ();
 sg13g2_decap_8 FILLER_50_1071 ();
 sg13g2_decap_8 FILLER_50_1078 ();
 sg13g2_decap_8 FILLER_50_1085 ();
 sg13g2_decap_8 FILLER_50_1092 ();
 sg13g2_decap_8 FILLER_50_1099 ();
 sg13g2_decap_8 FILLER_50_1106 ();
 sg13g2_decap_8 FILLER_50_1113 ();
 sg13g2_decap_8 FILLER_50_1120 ();
 sg13g2_decap_8 FILLER_50_1127 ();
 sg13g2_decap_8 FILLER_50_1134 ();
 sg13g2_decap_8 FILLER_50_1141 ();
 sg13g2_decap_8 FILLER_50_1148 ();
 sg13g2_decap_8 FILLER_50_1155 ();
 sg13g2_decap_8 FILLER_50_1162 ();
 sg13g2_decap_8 FILLER_50_1169 ();
 sg13g2_decap_8 FILLER_50_1176 ();
 sg13g2_decap_8 FILLER_50_1183 ();
 sg13g2_decap_8 FILLER_50_1190 ();
 sg13g2_decap_8 FILLER_50_1197 ();
 sg13g2_decap_8 FILLER_50_1204 ();
 sg13g2_decap_8 FILLER_50_1211 ();
 sg13g2_decap_8 FILLER_50_1218 ();
 sg13g2_decap_8 FILLER_50_1225 ();
 sg13g2_decap_8 FILLER_50_1232 ();
 sg13g2_decap_8 FILLER_50_1239 ();
 sg13g2_decap_8 FILLER_50_1246 ();
 sg13g2_decap_8 FILLER_50_1253 ();
 sg13g2_decap_8 FILLER_50_1260 ();
 sg13g2_decap_8 FILLER_50_1267 ();
 sg13g2_decap_8 FILLER_50_1274 ();
 sg13g2_decap_8 FILLER_50_1281 ();
 sg13g2_decap_8 FILLER_50_1288 ();
 sg13g2_decap_8 FILLER_50_1295 ();
 sg13g2_decap_8 FILLER_50_1302 ();
 sg13g2_decap_8 FILLER_50_1309 ();
 sg13g2_decap_8 FILLER_50_1316 ();
 sg13g2_decap_8 FILLER_50_1323 ();
 sg13g2_decap_8 FILLER_50_1330 ();
 sg13g2_decap_8 FILLER_50_1337 ();
 sg13g2_decap_8 FILLER_50_1344 ();
 sg13g2_decap_8 FILLER_50_1351 ();
 sg13g2_decap_8 FILLER_50_1358 ();
 sg13g2_decap_8 FILLER_50_1365 ();
 sg13g2_decap_8 FILLER_50_1372 ();
 sg13g2_decap_8 FILLER_50_1379 ();
 sg13g2_decap_8 FILLER_50_1386 ();
 sg13g2_decap_8 FILLER_50_1393 ();
 sg13g2_decap_8 FILLER_50_1400 ();
 sg13g2_decap_8 FILLER_50_1407 ();
 sg13g2_decap_8 FILLER_50_1414 ();
 sg13g2_decap_8 FILLER_50_1421 ();
 sg13g2_decap_8 FILLER_50_1428 ();
 sg13g2_decap_8 FILLER_50_1435 ();
 sg13g2_decap_8 FILLER_50_1442 ();
 sg13g2_decap_8 FILLER_50_1449 ();
 sg13g2_decap_8 FILLER_50_1456 ();
 sg13g2_decap_8 FILLER_50_1463 ();
 sg13g2_decap_8 FILLER_50_1470 ();
 sg13g2_decap_8 FILLER_50_1477 ();
 sg13g2_decap_8 FILLER_50_1484 ();
 sg13g2_decap_8 FILLER_50_1491 ();
 sg13g2_decap_8 FILLER_50_1498 ();
 sg13g2_decap_8 FILLER_50_1505 ();
 sg13g2_decap_8 FILLER_50_1512 ();
 sg13g2_decap_8 FILLER_50_1519 ();
 sg13g2_decap_8 FILLER_50_1526 ();
 sg13g2_decap_8 FILLER_50_1533 ();
 sg13g2_decap_8 FILLER_50_1540 ();
 sg13g2_decap_8 FILLER_50_1547 ();
 sg13g2_decap_8 FILLER_50_1554 ();
 sg13g2_decap_8 FILLER_50_1561 ();
 sg13g2_decap_8 FILLER_50_1568 ();
 sg13g2_decap_8 FILLER_50_1575 ();
 sg13g2_decap_8 FILLER_50_1582 ();
 sg13g2_decap_8 FILLER_50_1589 ();
 sg13g2_decap_8 FILLER_50_1596 ();
 sg13g2_decap_8 FILLER_50_1603 ();
 sg13g2_decap_8 FILLER_50_1610 ();
 sg13g2_decap_8 FILLER_50_1617 ();
 sg13g2_decap_8 FILLER_50_1624 ();
 sg13g2_decap_8 FILLER_50_1631 ();
 sg13g2_decap_8 FILLER_50_1638 ();
 sg13g2_decap_8 FILLER_50_1645 ();
 sg13g2_decap_8 FILLER_50_1652 ();
 sg13g2_decap_8 FILLER_50_1659 ();
 sg13g2_decap_8 FILLER_50_1666 ();
 sg13g2_decap_8 FILLER_50_1673 ();
 sg13g2_decap_8 FILLER_50_1680 ();
 sg13g2_decap_8 FILLER_50_1687 ();
 sg13g2_decap_8 FILLER_50_1694 ();
 sg13g2_decap_8 FILLER_50_1701 ();
 sg13g2_decap_8 FILLER_50_1708 ();
 sg13g2_decap_8 FILLER_50_1715 ();
 sg13g2_decap_8 FILLER_50_1722 ();
 sg13g2_decap_8 FILLER_50_1729 ();
 sg13g2_decap_8 FILLER_50_1736 ();
 sg13g2_decap_8 FILLER_50_1743 ();
 sg13g2_decap_8 FILLER_50_1750 ();
 sg13g2_decap_8 FILLER_50_1757 ();
 sg13g2_decap_4 FILLER_50_1764 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_7 ();
 sg13g2_fill_1 FILLER_51_9 ();
 sg13g2_fill_1 FILLER_51_22 ();
 sg13g2_decap_4 FILLER_51_28 ();
 sg13g2_fill_1 FILLER_51_32 ();
 sg13g2_fill_1 FILLER_51_38 ();
 sg13g2_decap_4 FILLER_51_44 ();
 sg13g2_fill_2 FILLER_51_48 ();
 sg13g2_fill_2 FILLER_51_59 ();
 sg13g2_fill_2 FILLER_51_67 ();
 sg13g2_decap_8 FILLER_51_82 ();
 sg13g2_decap_8 FILLER_51_89 ();
 sg13g2_decap_8 FILLER_51_96 ();
 sg13g2_fill_1 FILLER_51_122 ();
 sg13g2_decap_4 FILLER_51_135 ();
 sg13g2_fill_1 FILLER_51_139 ();
 sg13g2_decap_8 FILLER_51_161 ();
 sg13g2_decap_8 FILLER_51_168 ();
 sg13g2_decap_4 FILLER_51_175 ();
 sg13g2_decap_4 FILLER_51_211 ();
 sg13g2_fill_2 FILLER_51_215 ();
 sg13g2_decap_4 FILLER_51_231 ();
 sg13g2_fill_1 FILLER_51_235 ();
 sg13g2_fill_2 FILLER_51_244 ();
 sg13g2_decap_4 FILLER_51_256 ();
 sg13g2_decap_4 FILLER_51_275 ();
 sg13g2_fill_2 FILLER_51_285 ();
 sg13g2_decap_8 FILLER_51_297 ();
 sg13g2_decap_8 FILLER_51_304 ();
 sg13g2_fill_1 FILLER_51_311 ();
 sg13g2_fill_2 FILLER_51_348 ();
 sg13g2_fill_1 FILLER_51_350 ();
 sg13g2_fill_1 FILLER_51_361 ();
 sg13g2_fill_2 FILLER_51_385 ();
 sg13g2_fill_1 FILLER_51_387 ();
 sg13g2_fill_2 FILLER_51_405 ();
 sg13g2_fill_1 FILLER_51_459 ();
 sg13g2_fill_1 FILLER_51_480 ();
 sg13g2_fill_1 FILLER_51_497 ();
 sg13g2_decap_8 FILLER_51_558 ();
 sg13g2_decap_4 FILLER_51_565 ();
 sg13g2_fill_2 FILLER_51_569 ();
 sg13g2_fill_2 FILLER_51_599 ();
 sg13g2_fill_2 FILLER_51_607 ();
 sg13g2_fill_2 FILLER_51_615 ();
 sg13g2_fill_1 FILLER_51_617 ();
 sg13g2_fill_2 FILLER_51_633 ();
 sg13g2_fill_1 FILLER_51_653 ();
 sg13g2_decap_8 FILLER_51_667 ();
 sg13g2_decap_8 FILLER_51_674 ();
 sg13g2_decap_4 FILLER_51_698 ();
 sg13g2_fill_2 FILLER_51_711 ();
 sg13g2_fill_1 FILLER_51_713 ();
 sg13g2_decap_4 FILLER_51_722 ();
 sg13g2_decap_8 FILLER_51_745 ();
 sg13g2_fill_2 FILLER_51_848 ();
 sg13g2_fill_1 FILLER_51_881 ();
 sg13g2_fill_2 FILLER_51_916 ();
 sg13g2_decap_8 FILLER_51_924 ();
 sg13g2_decap_8 FILLER_51_931 ();
 sg13g2_decap_8 FILLER_51_938 ();
 sg13g2_fill_1 FILLER_51_945 ();
 sg13g2_fill_2 FILLER_51_966 ();
 sg13g2_fill_1 FILLER_51_976 ();
 sg13g2_fill_1 FILLER_51_987 ();
 sg13g2_fill_1 FILLER_51_993 ();
 sg13g2_fill_2 FILLER_51_1005 ();
 sg13g2_fill_1 FILLER_51_1019 ();
 sg13g2_decap_8 FILLER_51_1043 ();
 sg13g2_decap_8 FILLER_51_1050 ();
 sg13g2_decap_8 FILLER_51_1057 ();
 sg13g2_decap_8 FILLER_51_1064 ();
 sg13g2_decap_8 FILLER_51_1071 ();
 sg13g2_decap_8 FILLER_51_1078 ();
 sg13g2_decap_8 FILLER_51_1085 ();
 sg13g2_decap_8 FILLER_51_1092 ();
 sg13g2_decap_8 FILLER_51_1099 ();
 sg13g2_decap_8 FILLER_51_1106 ();
 sg13g2_decap_8 FILLER_51_1113 ();
 sg13g2_decap_8 FILLER_51_1120 ();
 sg13g2_decap_8 FILLER_51_1127 ();
 sg13g2_decap_8 FILLER_51_1134 ();
 sg13g2_decap_8 FILLER_51_1141 ();
 sg13g2_decap_8 FILLER_51_1148 ();
 sg13g2_decap_8 FILLER_51_1155 ();
 sg13g2_decap_8 FILLER_51_1162 ();
 sg13g2_decap_8 FILLER_51_1169 ();
 sg13g2_decap_8 FILLER_51_1176 ();
 sg13g2_decap_8 FILLER_51_1183 ();
 sg13g2_decap_8 FILLER_51_1190 ();
 sg13g2_decap_8 FILLER_51_1197 ();
 sg13g2_decap_8 FILLER_51_1204 ();
 sg13g2_decap_8 FILLER_51_1211 ();
 sg13g2_decap_8 FILLER_51_1218 ();
 sg13g2_decap_8 FILLER_51_1225 ();
 sg13g2_decap_8 FILLER_51_1232 ();
 sg13g2_decap_8 FILLER_51_1239 ();
 sg13g2_decap_8 FILLER_51_1246 ();
 sg13g2_decap_8 FILLER_51_1253 ();
 sg13g2_decap_8 FILLER_51_1260 ();
 sg13g2_decap_8 FILLER_51_1267 ();
 sg13g2_decap_8 FILLER_51_1274 ();
 sg13g2_decap_8 FILLER_51_1281 ();
 sg13g2_decap_8 FILLER_51_1288 ();
 sg13g2_decap_8 FILLER_51_1295 ();
 sg13g2_decap_8 FILLER_51_1302 ();
 sg13g2_decap_8 FILLER_51_1309 ();
 sg13g2_decap_8 FILLER_51_1316 ();
 sg13g2_decap_8 FILLER_51_1323 ();
 sg13g2_decap_8 FILLER_51_1330 ();
 sg13g2_decap_8 FILLER_51_1337 ();
 sg13g2_decap_8 FILLER_51_1344 ();
 sg13g2_decap_8 FILLER_51_1351 ();
 sg13g2_decap_8 FILLER_51_1358 ();
 sg13g2_decap_8 FILLER_51_1365 ();
 sg13g2_decap_8 FILLER_51_1372 ();
 sg13g2_decap_8 FILLER_51_1379 ();
 sg13g2_decap_8 FILLER_51_1386 ();
 sg13g2_decap_8 FILLER_51_1393 ();
 sg13g2_decap_8 FILLER_51_1400 ();
 sg13g2_decap_8 FILLER_51_1407 ();
 sg13g2_decap_8 FILLER_51_1414 ();
 sg13g2_decap_8 FILLER_51_1421 ();
 sg13g2_decap_8 FILLER_51_1428 ();
 sg13g2_decap_8 FILLER_51_1435 ();
 sg13g2_decap_8 FILLER_51_1442 ();
 sg13g2_decap_8 FILLER_51_1449 ();
 sg13g2_decap_8 FILLER_51_1456 ();
 sg13g2_decap_8 FILLER_51_1463 ();
 sg13g2_decap_8 FILLER_51_1470 ();
 sg13g2_decap_8 FILLER_51_1477 ();
 sg13g2_decap_8 FILLER_51_1484 ();
 sg13g2_decap_8 FILLER_51_1491 ();
 sg13g2_decap_8 FILLER_51_1498 ();
 sg13g2_decap_8 FILLER_51_1505 ();
 sg13g2_decap_8 FILLER_51_1512 ();
 sg13g2_decap_8 FILLER_51_1519 ();
 sg13g2_decap_8 FILLER_51_1526 ();
 sg13g2_decap_8 FILLER_51_1533 ();
 sg13g2_decap_8 FILLER_51_1540 ();
 sg13g2_decap_8 FILLER_51_1547 ();
 sg13g2_decap_8 FILLER_51_1554 ();
 sg13g2_decap_8 FILLER_51_1561 ();
 sg13g2_decap_8 FILLER_51_1568 ();
 sg13g2_decap_8 FILLER_51_1575 ();
 sg13g2_decap_8 FILLER_51_1582 ();
 sg13g2_decap_8 FILLER_51_1589 ();
 sg13g2_decap_8 FILLER_51_1596 ();
 sg13g2_decap_8 FILLER_51_1603 ();
 sg13g2_decap_8 FILLER_51_1610 ();
 sg13g2_decap_8 FILLER_51_1617 ();
 sg13g2_decap_8 FILLER_51_1624 ();
 sg13g2_decap_8 FILLER_51_1631 ();
 sg13g2_decap_8 FILLER_51_1638 ();
 sg13g2_decap_8 FILLER_51_1645 ();
 sg13g2_decap_8 FILLER_51_1652 ();
 sg13g2_decap_8 FILLER_51_1659 ();
 sg13g2_decap_8 FILLER_51_1666 ();
 sg13g2_decap_8 FILLER_51_1673 ();
 sg13g2_decap_8 FILLER_51_1680 ();
 sg13g2_decap_8 FILLER_51_1687 ();
 sg13g2_decap_8 FILLER_51_1694 ();
 sg13g2_decap_8 FILLER_51_1701 ();
 sg13g2_decap_8 FILLER_51_1708 ();
 sg13g2_decap_8 FILLER_51_1715 ();
 sg13g2_decap_8 FILLER_51_1722 ();
 sg13g2_decap_8 FILLER_51_1729 ();
 sg13g2_decap_8 FILLER_51_1736 ();
 sg13g2_decap_8 FILLER_51_1743 ();
 sg13g2_decap_8 FILLER_51_1750 ();
 sg13g2_decap_8 FILLER_51_1757 ();
 sg13g2_decap_4 FILLER_51_1764 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_63 ();
 sg13g2_decap_4 FILLER_52_90 ();
 sg13g2_fill_2 FILLER_52_127 ();
 sg13g2_fill_1 FILLER_52_129 ();
 sg13g2_decap_8 FILLER_52_135 ();
 sg13g2_fill_2 FILLER_52_142 ();
 sg13g2_decap_4 FILLER_52_161 ();
 sg13g2_decap_8 FILLER_52_191 ();
 sg13g2_decap_4 FILLER_52_198 ();
 sg13g2_fill_2 FILLER_52_202 ();
 sg13g2_decap_4 FILLER_52_231 ();
 sg13g2_fill_1 FILLER_52_235 ();
 sg13g2_decap_4 FILLER_52_292 ();
 sg13g2_decap_8 FILLER_52_301 ();
 sg13g2_decap_4 FILLER_52_308 ();
 sg13g2_fill_2 FILLER_52_322 ();
 sg13g2_fill_1 FILLER_52_362 ();
 sg13g2_fill_2 FILLER_52_394 ();
 sg13g2_fill_1 FILLER_52_396 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_fill_2 FILLER_52_462 ();
 sg13g2_fill_2 FILLER_52_486 ();
 sg13g2_fill_1 FILLER_52_488 ();
 sg13g2_fill_1 FILLER_52_516 ();
 sg13g2_decap_8 FILLER_52_523 ();
 sg13g2_decap_8 FILLER_52_530 ();
 sg13g2_decap_8 FILLER_52_537 ();
 sg13g2_decap_8 FILLER_52_548 ();
 sg13g2_decap_4 FILLER_52_555 ();
 sg13g2_fill_2 FILLER_52_574 ();
 sg13g2_decap_4 FILLER_52_584 ();
 sg13g2_fill_1 FILLER_52_592 ();
 sg13g2_fill_1 FILLER_52_601 ();
 sg13g2_decap_4 FILLER_52_632 ();
 sg13g2_decap_4 FILLER_52_639 ();
 sg13g2_fill_1 FILLER_52_652 ();
 sg13g2_decap_4 FILLER_52_662 ();
 sg13g2_fill_2 FILLER_52_666 ();
 sg13g2_fill_1 FILLER_52_672 ();
 sg13g2_fill_1 FILLER_52_678 ();
 sg13g2_decap_4 FILLER_52_706 ();
 sg13g2_decap_8 FILLER_52_720 ();
 sg13g2_decap_8 FILLER_52_732 ();
 sg13g2_fill_1 FILLER_52_739 ();
 sg13g2_decap_8 FILLER_52_744 ();
 sg13g2_fill_2 FILLER_52_751 ();
 sg13g2_fill_1 FILLER_52_753 ();
 sg13g2_decap_8 FILLER_52_779 ();
 sg13g2_decap_4 FILLER_52_786 ();
 sg13g2_fill_1 FILLER_52_790 ();
 sg13g2_fill_1 FILLER_52_799 ();
 sg13g2_fill_1 FILLER_52_809 ();
 sg13g2_fill_2 FILLER_52_824 ();
 sg13g2_fill_1 FILLER_52_826 ();
 sg13g2_decap_8 FILLER_52_874 ();
 sg13g2_fill_2 FILLER_52_881 ();
 sg13g2_fill_1 FILLER_52_883 ();
 sg13g2_decap_8 FILLER_52_901 ();
 sg13g2_decap_8 FILLER_52_928 ();
 sg13g2_decap_4 FILLER_52_935 ();
 sg13g2_decap_8 FILLER_52_965 ();
 sg13g2_fill_2 FILLER_52_972 ();
 sg13g2_decap_8 FILLER_52_980 ();
 sg13g2_fill_1 FILLER_52_992 ();
 sg13g2_decap_8 FILLER_52_1027 ();
 sg13g2_decap_8 FILLER_52_1034 ();
 sg13g2_decap_8 FILLER_52_1041 ();
 sg13g2_decap_8 FILLER_52_1048 ();
 sg13g2_decap_8 FILLER_52_1055 ();
 sg13g2_decap_8 FILLER_52_1062 ();
 sg13g2_decap_8 FILLER_52_1069 ();
 sg13g2_decap_8 FILLER_52_1076 ();
 sg13g2_decap_8 FILLER_52_1083 ();
 sg13g2_decap_8 FILLER_52_1090 ();
 sg13g2_decap_8 FILLER_52_1097 ();
 sg13g2_decap_8 FILLER_52_1104 ();
 sg13g2_decap_8 FILLER_52_1111 ();
 sg13g2_decap_8 FILLER_52_1118 ();
 sg13g2_decap_8 FILLER_52_1125 ();
 sg13g2_decap_8 FILLER_52_1132 ();
 sg13g2_decap_8 FILLER_52_1139 ();
 sg13g2_decap_8 FILLER_52_1146 ();
 sg13g2_decap_8 FILLER_52_1153 ();
 sg13g2_decap_8 FILLER_52_1160 ();
 sg13g2_decap_8 FILLER_52_1167 ();
 sg13g2_decap_8 FILLER_52_1174 ();
 sg13g2_decap_8 FILLER_52_1181 ();
 sg13g2_decap_8 FILLER_52_1188 ();
 sg13g2_decap_8 FILLER_52_1195 ();
 sg13g2_decap_8 FILLER_52_1202 ();
 sg13g2_decap_8 FILLER_52_1209 ();
 sg13g2_decap_8 FILLER_52_1216 ();
 sg13g2_decap_8 FILLER_52_1223 ();
 sg13g2_decap_8 FILLER_52_1230 ();
 sg13g2_decap_8 FILLER_52_1237 ();
 sg13g2_decap_8 FILLER_52_1244 ();
 sg13g2_decap_8 FILLER_52_1251 ();
 sg13g2_decap_8 FILLER_52_1258 ();
 sg13g2_decap_8 FILLER_52_1265 ();
 sg13g2_decap_8 FILLER_52_1272 ();
 sg13g2_decap_8 FILLER_52_1279 ();
 sg13g2_decap_8 FILLER_52_1286 ();
 sg13g2_decap_8 FILLER_52_1293 ();
 sg13g2_decap_8 FILLER_52_1300 ();
 sg13g2_decap_8 FILLER_52_1307 ();
 sg13g2_decap_8 FILLER_52_1314 ();
 sg13g2_decap_8 FILLER_52_1321 ();
 sg13g2_decap_8 FILLER_52_1328 ();
 sg13g2_decap_8 FILLER_52_1335 ();
 sg13g2_decap_8 FILLER_52_1342 ();
 sg13g2_decap_8 FILLER_52_1349 ();
 sg13g2_decap_8 FILLER_52_1356 ();
 sg13g2_decap_8 FILLER_52_1363 ();
 sg13g2_decap_8 FILLER_52_1370 ();
 sg13g2_decap_8 FILLER_52_1377 ();
 sg13g2_decap_8 FILLER_52_1384 ();
 sg13g2_decap_8 FILLER_52_1391 ();
 sg13g2_decap_8 FILLER_52_1398 ();
 sg13g2_decap_8 FILLER_52_1405 ();
 sg13g2_decap_8 FILLER_52_1412 ();
 sg13g2_decap_8 FILLER_52_1419 ();
 sg13g2_decap_8 FILLER_52_1426 ();
 sg13g2_decap_8 FILLER_52_1433 ();
 sg13g2_decap_8 FILLER_52_1440 ();
 sg13g2_decap_8 FILLER_52_1447 ();
 sg13g2_decap_8 FILLER_52_1454 ();
 sg13g2_decap_8 FILLER_52_1461 ();
 sg13g2_decap_8 FILLER_52_1468 ();
 sg13g2_decap_8 FILLER_52_1475 ();
 sg13g2_decap_8 FILLER_52_1482 ();
 sg13g2_decap_8 FILLER_52_1489 ();
 sg13g2_decap_8 FILLER_52_1496 ();
 sg13g2_decap_8 FILLER_52_1503 ();
 sg13g2_decap_8 FILLER_52_1510 ();
 sg13g2_decap_8 FILLER_52_1517 ();
 sg13g2_decap_8 FILLER_52_1524 ();
 sg13g2_decap_8 FILLER_52_1531 ();
 sg13g2_decap_8 FILLER_52_1538 ();
 sg13g2_decap_8 FILLER_52_1545 ();
 sg13g2_decap_8 FILLER_52_1552 ();
 sg13g2_decap_8 FILLER_52_1559 ();
 sg13g2_decap_8 FILLER_52_1566 ();
 sg13g2_decap_8 FILLER_52_1573 ();
 sg13g2_decap_8 FILLER_52_1580 ();
 sg13g2_decap_8 FILLER_52_1587 ();
 sg13g2_decap_8 FILLER_52_1594 ();
 sg13g2_decap_8 FILLER_52_1601 ();
 sg13g2_decap_8 FILLER_52_1608 ();
 sg13g2_decap_8 FILLER_52_1615 ();
 sg13g2_decap_8 FILLER_52_1622 ();
 sg13g2_decap_8 FILLER_52_1629 ();
 sg13g2_decap_8 FILLER_52_1636 ();
 sg13g2_decap_8 FILLER_52_1643 ();
 sg13g2_decap_8 FILLER_52_1650 ();
 sg13g2_decap_8 FILLER_52_1657 ();
 sg13g2_decap_8 FILLER_52_1664 ();
 sg13g2_decap_8 FILLER_52_1671 ();
 sg13g2_decap_8 FILLER_52_1678 ();
 sg13g2_decap_8 FILLER_52_1685 ();
 sg13g2_decap_8 FILLER_52_1692 ();
 sg13g2_decap_8 FILLER_52_1699 ();
 sg13g2_decap_8 FILLER_52_1706 ();
 sg13g2_decap_8 FILLER_52_1713 ();
 sg13g2_decap_8 FILLER_52_1720 ();
 sg13g2_decap_8 FILLER_52_1727 ();
 sg13g2_decap_8 FILLER_52_1734 ();
 sg13g2_decap_8 FILLER_52_1741 ();
 sg13g2_decap_8 FILLER_52_1748 ();
 sg13g2_decap_8 FILLER_52_1755 ();
 sg13g2_decap_4 FILLER_52_1762 ();
 sg13g2_fill_2 FILLER_52_1766 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_9 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_fill_2 FILLER_53_35 ();
 sg13g2_fill_1 FILLER_53_46 ();
 sg13g2_decap_4 FILLER_53_57 ();
 sg13g2_fill_1 FILLER_53_61 ();
 sg13g2_decap_8 FILLER_53_88 ();
 sg13g2_fill_1 FILLER_53_95 ();
 sg13g2_fill_1 FILLER_53_100 ();
 sg13g2_fill_2 FILLER_53_104 ();
 sg13g2_fill_2 FILLER_53_111 ();
 sg13g2_decap_4 FILLER_53_123 ();
 sg13g2_fill_1 FILLER_53_127 ();
 sg13g2_fill_2 FILLER_53_151 ();
 sg13g2_decap_4 FILLER_53_202 ();
 sg13g2_fill_1 FILLER_53_206 ();
 sg13g2_decap_8 FILLER_53_216 ();
 sg13g2_decap_4 FILLER_53_223 ();
 sg13g2_fill_2 FILLER_53_227 ();
 sg13g2_fill_2 FILLER_53_233 ();
 sg13g2_decap_4 FILLER_53_243 ();
 sg13g2_fill_1 FILLER_53_247 ();
 sg13g2_decap_8 FILLER_53_253 ();
 sg13g2_fill_2 FILLER_53_260 ();
 sg13g2_decap_8 FILLER_53_267 ();
 sg13g2_decap_4 FILLER_53_274 ();
 sg13g2_fill_2 FILLER_53_311 ();
 sg13g2_fill_1 FILLER_53_313 ();
 sg13g2_decap_8 FILLER_53_320 ();
 sg13g2_decap_8 FILLER_53_327 ();
 sg13g2_decap_4 FILLER_53_334 ();
 sg13g2_fill_2 FILLER_53_338 ();
 sg13g2_decap_8 FILLER_53_350 ();
 sg13g2_decap_4 FILLER_53_357 ();
 sg13g2_fill_2 FILLER_53_373 ();
 sg13g2_fill_2 FILLER_53_383 ();
 sg13g2_fill_1 FILLER_53_385 ();
 sg13g2_fill_1 FILLER_53_390 ();
 sg13g2_fill_1 FILLER_53_405 ();
 sg13g2_fill_1 FILLER_53_416 ();
 sg13g2_fill_1 FILLER_53_475 ();
 sg13g2_fill_1 FILLER_53_523 ();
 sg13g2_fill_2 FILLER_53_530 ();
 sg13g2_fill_1 FILLER_53_532 ();
 sg13g2_fill_2 FILLER_53_559 ();
 sg13g2_fill_1 FILLER_53_561 ();
 sg13g2_decap_8 FILLER_53_568 ();
 sg13g2_decap_8 FILLER_53_575 ();
 sg13g2_decap_8 FILLER_53_582 ();
 sg13g2_decap_4 FILLER_53_595 ();
 sg13g2_fill_1 FILLER_53_599 ();
 sg13g2_decap_4 FILLER_53_611 ();
 sg13g2_fill_1 FILLER_53_615 ();
 sg13g2_decap_8 FILLER_53_625 ();
 sg13g2_decap_4 FILLER_53_632 ();
 sg13g2_fill_1 FILLER_53_636 ();
 sg13g2_decap_8 FILLER_53_666 ();
 sg13g2_decap_4 FILLER_53_673 ();
 sg13g2_fill_1 FILLER_53_677 ();
 sg13g2_decap_4 FILLER_53_682 ();
 sg13g2_fill_2 FILLER_53_686 ();
 sg13g2_decap_4 FILLER_53_695 ();
 sg13g2_fill_2 FILLER_53_699 ();
 sg13g2_decap_8 FILLER_53_716 ();
 sg13g2_fill_1 FILLER_53_723 ();
 sg13g2_fill_1 FILLER_53_755 ();
 sg13g2_fill_2 FILLER_53_775 ();
 sg13g2_decap_8 FILLER_53_787 ();
 sg13g2_fill_1 FILLER_53_794 ();
 sg13g2_fill_2 FILLER_53_803 ();
 sg13g2_decap_4 FILLER_53_810 ();
 sg13g2_fill_2 FILLER_53_814 ();
 sg13g2_fill_2 FILLER_53_859 ();
 sg13g2_decap_4 FILLER_53_876 ();
 sg13g2_fill_2 FILLER_53_901 ();
 sg13g2_fill_1 FILLER_53_903 ();
 sg13g2_decap_8 FILLER_53_928 ();
 sg13g2_fill_2 FILLER_53_935 ();
 sg13g2_fill_2 FILLER_53_952 ();
 sg13g2_fill_2 FILLER_53_958 ();
 sg13g2_fill_1 FILLER_53_969 ();
 sg13g2_decap_4 FILLER_53_975 ();
 sg13g2_fill_2 FILLER_53_979 ();
 sg13g2_fill_2 FILLER_53_1006 ();
 sg13g2_decap_8 FILLER_53_1037 ();
 sg13g2_decap_8 FILLER_53_1044 ();
 sg13g2_decap_8 FILLER_53_1051 ();
 sg13g2_decap_8 FILLER_53_1058 ();
 sg13g2_decap_8 FILLER_53_1065 ();
 sg13g2_decap_8 FILLER_53_1072 ();
 sg13g2_decap_8 FILLER_53_1079 ();
 sg13g2_decap_8 FILLER_53_1086 ();
 sg13g2_decap_8 FILLER_53_1093 ();
 sg13g2_decap_8 FILLER_53_1100 ();
 sg13g2_decap_8 FILLER_53_1107 ();
 sg13g2_decap_8 FILLER_53_1114 ();
 sg13g2_decap_8 FILLER_53_1121 ();
 sg13g2_decap_8 FILLER_53_1128 ();
 sg13g2_decap_8 FILLER_53_1135 ();
 sg13g2_decap_8 FILLER_53_1142 ();
 sg13g2_decap_8 FILLER_53_1149 ();
 sg13g2_decap_8 FILLER_53_1156 ();
 sg13g2_decap_8 FILLER_53_1163 ();
 sg13g2_decap_8 FILLER_53_1170 ();
 sg13g2_decap_8 FILLER_53_1177 ();
 sg13g2_decap_8 FILLER_53_1184 ();
 sg13g2_decap_8 FILLER_53_1191 ();
 sg13g2_decap_8 FILLER_53_1198 ();
 sg13g2_decap_8 FILLER_53_1205 ();
 sg13g2_decap_8 FILLER_53_1212 ();
 sg13g2_decap_8 FILLER_53_1219 ();
 sg13g2_decap_8 FILLER_53_1226 ();
 sg13g2_decap_8 FILLER_53_1233 ();
 sg13g2_decap_8 FILLER_53_1240 ();
 sg13g2_decap_8 FILLER_53_1247 ();
 sg13g2_decap_8 FILLER_53_1254 ();
 sg13g2_decap_8 FILLER_53_1261 ();
 sg13g2_decap_8 FILLER_53_1268 ();
 sg13g2_decap_8 FILLER_53_1275 ();
 sg13g2_decap_8 FILLER_53_1282 ();
 sg13g2_decap_8 FILLER_53_1289 ();
 sg13g2_decap_8 FILLER_53_1296 ();
 sg13g2_decap_8 FILLER_53_1303 ();
 sg13g2_decap_8 FILLER_53_1310 ();
 sg13g2_decap_8 FILLER_53_1317 ();
 sg13g2_decap_8 FILLER_53_1324 ();
 sg13g2_decap_8 FILLER_53_1331 ();
 sg13g2_decap_8 FILLER_53_1338 ();
 sg13g2_decap_8 FILLER_53_1345 ();
 sg13g2_decap_8 FILLER_53_1352 ();
 sg13g2_decap_8 FILLER_53_1359 ();
 sg13g2_decap_8 FILLER_53_1366 ();
 sg13g2_decap_8 FILLER_53_1373 ();
 sg13g2_decap_8 FILLER_53_1380 ();
 sg13g2_decap_8 FILLER_53_1387 ();
 sg13g2_decap_8 FILLER_53_1394 ();
 sg13g2_decap_8 FILLER_53_1401 ();
 sg13g2_decap_8 FILLER_53_1408 ();
 sg13g2_decap_8 FILLER_53_1415 ();
 sg13g2_decap_8 FILLER_53_1422 ();
 sg13g2_decap_8 FILLER_53_1429 ();
 sg13g2_decap_8 FILLER_53_1436 ();
 sg13g2_decap_8 FILLER_53_1443 ();
 sg13g2_decap_8 FILLER_53_1450 ();
 sg13g2_decap_8 FILLER_53_1457 ();
 sg13g2_decap_8 FILLER_53_1464 ();
 sg13g2_decap_8 FILLER_53_1471 ();
 sg13g2_decap_8 FILLER_53_1478 ();
 sg13g2_decap_8 FILLER_53_1485 ();
 sg13g2_decap_8 FILLER_53_1492 ();
 sg13g2_decap_8 FILLER_53_1499 ();
 sg13g2_decap_8 FILLER_53_1506 ();
 sg13g2_decap_8 FILLER_53_1513 ();
 sg13g2_decap_8 FILLER_53_1520 ();
 sg13g2_decap_8 FILLER_53_1527 ();
 sg13g2_decap_8 FILLER_53_1534 ();
 sg13g2_decap_8 FILLER_53_1541 ();
 sg13g2_decap_8 FILLER_53_1548 ();
 sg13g2_decap_8 FILLER_53_1555 ();
 sg13g2_decap_8 FILLER_53_1562 ();
 sg13g2_decap_8 FILLER_53_1569 ();
 sg13g2_decap_8 FILLER_53_1576 ();
 sg13g2_decap_8 FILLER_53_1583 ();
 sg13g2_decap_8 FILLER_53_1590 ();
 sg13g2_decap_8 FILLER_53_1597 ();
 sg13g2_decap_8 FILLER_53_1604 ();
 sg13g2_decap_8 FILLER_53_1611 ();
 sg13g2_decap_8 FILLER_53_1618 ();
 sg13g2_decap_8 FILLER_53_1625 ();
 sg13g2_decap_8 FILLER_53_1632 ();
 sg13g2_decap_8 FILLER_53_1639 ();
 sg13g2_decap_8 FILLER_53_1646 ();
 sg13g2_decap_8 FILLER_53_1653 ();
 sg13g2_decap_8 FILLER_53_1660 ();
 sg13g2_decap_8 FILLER_53_1667 ();
 sg13g2_decap_8 FILLER_53_1674 ();
 sg13g2_decap_8 FILLER_53_1681 ();
 sg13g2_decap_8 FILLER_53_1688 ();
 sg13g2_decap_8 FILLER_53_1695 ();
 sg13g2_decap_8 FILLER_53_1702 ();
 sg13g2_decap_8 FILLER_53_1709 ();
 sg13g2_decap_8 FILLER_53_1716 ();
 sg13g2_decap_8 FILLER_53_1723 ();
 sg13g2_decap_8 FILLER_53_1730 ();
 sg13g2_decap_8 FILLER_53_1737 ();
 sg13g2_decap_8 FILLER_53_1744 ();
 sg13g2_decap_8 FILLER_53_1751 ();
 sg13g2_decap_8 FILLER_53_1758 ();
 sg13g2_fill_2 FILLER_53_1765 ();
 sg13g2_fill_1 FILLER_53_1767 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_4 FILLER_54_7 ();
 sg13g2_fill_1 FILLER_54_11 ();
 sg13g2_fill_1 FILLER_54_33 ();
 sg13g2_decap_4 FILLER_54_63 ();
 sg13g2_fill_2 FILLER_54_86 ();
 sg13g2_fill_1 FILLER_54_88 ();
 sg13g2_fill_2 FILLER_54_101 ();
 sg13g2_decap_4 FILLER_54_121 ();
 sg13g2_fill_1 FILLER_54_125 ();
 sg13g2_fill_1 FILLER_54_147 ();
 sg13g2_fill_2 FILLER_54_161 ();
 sg13g2_fill_1 FILLER_54_163 ();
 sg13g2_decap_8 FILLER_54_168 ();
 sg13g2_decap_8 FILLER_54_175 ();
 sg13g2_decap_8 FILLER_54_182 ();
 sg13g2_fill_1 FILLER_54_189 ();
 sg13g2_fill_2 FILLER_54_199 ();
 sg13g2_fill_1 FILLER_54_201 ();
 sg13g2_fill_2 FILLER_54_210 ();
 sg13g2_fill_1 FILLER_54_212 ();
 sg13g2_fill_2 FILLER_54_266 ();
 sg13g2_fill_1 FILLER_54_268 ();
 sg13g2_fill_2 FILLER_54_312 ();
 sg13g2_decap_4 FILLER_54_329 ();
 sg13g2_fill_2 FILLER_54_333 ();
 sg13g2_decap_8 FILLER_54_351 ();
 sg13g2_fill_1 FILLER_54_358 ();
 sg13g2_decap_4 FILLER_54_364 ();
 sg13g2_fill_1 FILLER_54_368 ();
 sg13g2_fill_1 FILLER_54_391 ();
 sg13g2_fill_2 FILLER_54_412 ();
 sg13g2_fill_1 FILLER_54_444 ();
 sg13g2_fill_2 FILLER_54_489 ();
 sg13g2_fill_1 FILLER_54_491 ();
 sg13g2_fill_2 FILLER_54_532 ();
 sg13g2_fill_2 FILLER_54_556 ();
 sg13g2_fill_1 FILLER_54_558 ();
 sg13g2_fill_2 FILLER_54_571 ();
 sg13g2_fill_1 FILLER_54_600 ();
 sg13g2_fill_2 FILLER_54_622 ();
 sg13g2_fill_1 FILLER_54_624 ();
 sg13g2_fill_2 FILLER_54_635 ();
 sg13g2_fill_2 FILLER_54_649 ();
 sg13g2_fill_2 FILLER_54_664 ();
 sg13g2_fill_1 FILLER_54_666 ();
 sg13g2_fill_2 FILLER_54_682 ();
 sg13g2_decap_8 FILLER_54_723 ();
 sg13g2_decap_8 FILLER_54_730 ();
 sg13g2_fill_2 FILLER_54_741 ();
 sg13g2_fill_2 FILLER_54_767 ();
 sg13g2_fill_1 FILLER_54_769 ();
 sg13g2_fill_1 FILLER_54_775 ();
 sg13g2_fill_2 FILLER_54_789 ();
 sg13g2_fill_1 FILLER_54_791 ();
 sg13g2_fill_1 FILLER_54_816 ();
 sg13g2_decap_4 FILLER_54_823 ();
 sg13g2_decap_8 FILLER_54_857 ();
 sg13g2_decap_8 FILLER_54_864 ();
 sg13g2_fill_2 FILLER_54_871 ();
 sg13g2_fill_2 FILLER_54_881 ();
 sg13g2_fill_2 FILLER_54_888 ();
 sg13g2_fill_1 FILLER_54_890 ();
 sg13g2_decap_8 FILLER_54_901 ();
 sg13g2_decap_4 FILLER_54_908 ();
 sg13g2_fill_2 FILLER_54_912 ();
 sg13g2_decap_8 FILLER_54_936 ();
 sg13g2_fill_2 FILLER_54_943 ();
 sg13g2_fill_1 FILLER_54_945 ();
 sg13g2_fill_1 FILLER_54_965 ();
 sg13g2_decap_4 FILLER_54_977 ();
 sg13g2_fill_1 FILLER_54_981 ();
 sg13g2_fill_1 FILLER_54_990 ();
 sg13g2_fill_1 FILLER_54_1014 ();
 sg13g2_decap_8 FILLER_54_1044 ();
 sg13g2_decap_8 FILLER_54_1051 ();
 sg13g2_decap_8 FILLER_54_1058 ();
 sg13g2_decap_8 FILLER_54_1065 ();
 sg13g2_decap_8 FILLER_54_1072 ();
 sg13g2_decap_8 FILLER_54_1079 ();
 sg13g2_decap_8 FILLER_54_1086 ();
 sg13g2_decap_8 FILLER_54_1093 ();
 sg13g2_decap_8 FILLER_54_1100 ();
 sg13g2_decap_8 FILLER_54_1107 ();
 sg13g2_decap_8 FILLER_54_1114 ();
 sg13g2_decap_8 FILLER_54_1121 ();
 sg13g2_decap_8 FILLER_54_1128 ();
 sg13g2_decap_8 FILLER_54_1135 ();
 sg13g2_decap_8 FILLER_54_1142 ();
 sg13g2_decap_8 FILLER_54_1149 ();
 sg13g2_decap_8 FILLER_54_1156 ();
 sg13g2_decap_8 FILLER_54_1163 ();
 sg13g2_decap_8 FILLER_54_1170 ();
 sg13g2_decap_8 FILLER_54_1177 ();
 sg13g2_decap_8 FILLER_54_1184 ();
 sg13g2_decap_8 FILLER_54_1191 ();
 sg13g2_decap_8 FILLER_54_1198 ();
 sg13g2_decap_8 FILLER_54_1205 ();
 sg13g2_decap_8 FILLER_54_1212 ();
 sg13g2_decap_8 FILLER_54_1219 ();
 sg13g2_decap_8 FILLER_54_1226 ();
 sg13g2_decap_8 FILLER_54_1233 ();
 sg13g2_decap_8 FILLER_54_1240 ();
 sg13g2_decap_8 FILLER_54_1247 ();
 sg13g2_decap_8 FILLER_54_1254 ();
 sg13g2_decap_8 FILLER_54_1261 ();
 sg13g2_decap_8 FILLER_54_1268 ();
 sg13g2_decap_8 FILLER_54_1275 ();
 sg13g2_decap_8 FILLER_54_1282 ();
 sg13g2_decap_8 FILLER_54_1289 ();
 sg13g2_decap_8 FILLER_54_1296 ();
 sg13g2_decap_8 FILLER_54_1303 ();
 sg13g2_decap_8 FILLER_54_1310 ();
 sg13g2_decap_8 FILLER_54_1317 ();
 sg13g2_decap_8 FILLER_54_1324 ();
 sg13g2_decap_8 FILLER_54_1331 ();
 sg13g2_decap_8 FILLER_54_1338 ();
 sg13g2_decap_8 FILLER_54_1345 ();
 sg13g2_decap_8 FILLER_54_1352 ();
 sg13g2_decap_8 FILLER_54_1359 ();
 sg13g2_decap_8 FILLER_54_1366 ();
 sg13g2_decap_8 FILLER_54_1373 ();
 sg13g2_decap_8 FILLER_54_1380 ();
 sg13g2_decap_8 FILLER_54_1387 ();
 sg13g2_decap_8 FILLER_54_1394 ();
 sg13g2_decap_8 FILLER_54_1401 ();
 sg13g2_decap_8 FILLER_54_1408 ();
 sg13g2_decap_8 FILLER_54_1415 ();
 sg13g2_decap_8 FILLER_54_1422 ();
 sg13g2_decap_8 FILLER_54_1429 ();
 sg13g2_decap_8 FILLER_54_1436 ();
 sg13g2_decap_8 FILLER_54_1443 ();
 sg13g2_decap_8 FILLER_54_1450 ();
 sg13g2_decap_8 FILLER_54_1457 ();
 sg13g2_decap_8 FILLER_54_1464 ();
 sg13g2_decap_8 FILLER_54_1471 ();
 sg13g2_decap_8 FILLER_54_1478 ();
 sg13g2_decap_8 FILLER_54_1485 ();
 sg13g2_decap_8 FILLER_54_1492 ();
 sg13g2_decap_8 FILLER_54_1499 ();
 sg13g2_decap_8 FILLER_54_1506 ();
 sg13g2_decap_8 FILLER_54_1513 ();
 sg13g2_decap_8 FILLER_54_1520 ();
 sg13g2_decap_8 FILLER_54_1527 ();
 sg13g2_decap_8 FILLER_54_1534 ();
 sg13g2_decap_8 FILLER_54_1541 ();
 sg13g2_decap_8 FILLER_54_1548 ();
 sg13g2_decap_8 FILLER_54_1555 ();
 sg13g2_decap_8 FILLER_54_1562 ();
 sg13g2_decap_8 FILLER_54_1569 ();
 sg13g2_decap_8 FILLER_54_1576 ();
 sg13g2_decap_8 FILLER_54_1583 ();
 sg13g2_decap_8 FILLER_54_1590 ();
 sg13g2_decap_8 FILLER_54_1597 ();
 sg13g2_decap_8 FILLER_54_1604 ();
 sg13g2_decap_8 FILLER_54_1611 ();
 sg13g2_decap_8 FILLER_54_1618 ();
 sg13g2_decap_8 FILLER_54_1625 ();
 sg13g2_decap_8 FILLER_54_1632 ();
 sg13g2_decap_8 FILLER_54_1639 ();
 sg13g2_decap_8 FILLER_54_1646 ();
 sg13g2_decap_8 FILLER_54_1653 ();
 sg13g2_decap_8 FILLER_54_1660 ();
 sg13g2_decap_8 FILLER_54_1667 ();
 sg13g2_decap_8 FILLER_54_1674 ();
 sg13g2_decap_8 FILLER_54_1681 ();
 sg13g2_decap_8 FILLER_54_1688 ();
 sg13g2_decap_8 FILLER_54_1695 ();
 sg13g2_decap_8 FILLER_54_1702 ();
 sg13g2_decap_8 FILLER_54_1709 ();
 sg13g2_decap_8 FILLER_54_1716 ();
 sg13g2_decap_8 FILLER_54_1723 ();
 sg13g2_decap_8 FILLER_54_1730 ();
 sg13g2_decap_8 FILLER_54_1737 ();
 sg13g2_decap_8 FILLER_54_1744 ();
 sg13g2_decap_8 FILLER_54_1751 ();
 sg13g2_decap_8 FILLER_54_1758 ();
 sg13g2_fill_2 FILLER_54_1765 ();
 sg13g2_fill_1 FILLER_54_1767 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_36 ();
 sg13g2_fill_2 FILLER_55_58 ();
 sg13g2_fill_1 FILLER_55_60 ();
 sg13g2_decap_8 FILLER_55_90 ();
 sg13g2_fill_1 FILLER_55_97 ();
 sg13g2_decap_8 FILLER_55_123 ();
 sg13g2_fill_2 FILLER_55_130 ();
 sg13g2_decap_8 FILLER_55_136 ();
 sg13g2_fill_1 FILLER_55_143 ();
 sg13g2_fill_1 FILLER_55_156 ();
 sg13g2_fill_2 FILLER_55_193 ();
 sg13g2_fill_2 FILLER_55_226 ();
 sg13g2_fill_1 FILLER_55_228 ();
 sg13g2_decap_4 FILLER_55_235 ();
 sg13g2_fill_1 FILLER_55_239 ();
 sg13g2_decap_4 FILLER_55_253 ();
 sg13g2_decap_8 FILLER_55_268 ();
 sg13g2_decap_8 FILLER_55_275 ();
 sg13g2_fill_1 FILLER_55_290 ();
 sg13g2_fill_2 FILLER_55_296 ();
 sg13g2_fill_1 FILLER_55_298 ();
 sg13g2_fill_2 FILLER_55_304 ();
 sg13g2_decap_4 FILLER_55_319 ();
 sg13g2_fill_2 FILLER_55_369 ();
 sg13g2_fill_1 FILLER_55_371 ();
 sg13g2_decap_8 FILLER_55_387 ();
 sg13g2_fill_2 FILLER_55_394 ();
 sg13g2_fill_1 FILLER_55_396 ();
 sg13g2_fill_1 FILLER_55_411 ();
 sg13g2_fill_1 FILLER_55_429 ();
 sg13g2_decap_8 FILLER_55_439 ();
 sg13g2_decap_4 FILLER_55_446 ();
 sg13g2_decap_8 FILLER_55_455 ();
 sg13g2_decap_4 FILLER_55_462 ();
 sg13g2_fill_1 FILLER_55_466 ();
 sg13g2_decap_8 FILLER_55_474 ();
 sg13g2_fill_1 FILLER_55_495 ();
 sg13g2_decap_8 FILLER_55_501 ();
 sg13g2_fill_2 FILLER_55_508 ();
 sg13g2_fill_1 FILLER_55_510 ();
 sg13g2_decap_4 FILLER_55_515 ();
 sg13g2_decap_4 FILLER_55_531 ();
 sg13g2_fill_2 FILLER_55_539 ();
 sg13g2_fill_1 FILLER_55_558 ();
 sg13g2_decap_8 FILLER_55_563 ();
 sg13g2_decap_4 FILLER_55_570 ();
 sg13g2_fill_2 FILLER_55_574 ();
 sg13g2_decap_8 FILLER_55_596 ();
 sg13g2_decap_8 FILLER_55_603 ();
 sg13g2_decap_8 FILLER_55_610 ();
 sg13g2_decap_4 FILLER_55_626 ();
 sg13g2_fill_2 FILLER_55_635 ();
 sg13g2_fill_1 FILLER_55_647 ();
 sg13g2_fill_2 FILLER_55_665 ();
 sg13g2_decap_4 FILLER_55_681 ();
 sg13g2_fill_2 FILLER_55_685 ();
 sg13g2_decap_4 FILLER_55_711 ();
 sg13g2_fill_1 FILLER_55_715 ();
 sg13g2_fill_1 FILLER_55_752 ();
 sg13g2_fill_2 FILLER_55_762 ();
 sg13g2_fill_1 FILLER_55_764 ();
 sg13g2_fill_1 FILLER_55_785 ();
 sg13g2_fill_2 FILLER_55_803 ();
 sg13g2_decap_4 FILLER_55_811 ();
 sg13g2_fill_2 FILLER_55_815 ();
 sg13g2_decap_8 FILLER_55_828 ();
 sg13g2_fill_1 FILLER_55_853 ();
 sg13g2_decap_4 FILLER_55_862 ();
 sg13g2_fill_1 FILLER_55_866 ();
 sg13g2_decap_4 FILLER_55_879 ();
 sg13g2_fill_1 FILLER_55_883 ();
 sg13g2_fill_2 FILLER_55_893 ();
 sg13g2_fill_1 FILLER_55_895 ();
 sg13g2_decap_8 FILLER_55_904 ();
 sg13g2_decap_4 FILLER_55_933 ();
 sg13g2_decap_8 FILLER_55_948 ();
 sg13g2_fill_2 FILLER_55_955 ();
 sg13g2_decap_8 FILLER_55_966 ();
 sg13g2_fill_2 FILLER_55_973 ();
 sg13g2_fill_1 FILLER_55_975 ();
 sg13g2_fill_2 FILLER_55_984 ();
 sg13g2_decap_4 FILLER_55_991 ();
 sg13g2_decap_8 FILLER_55_1005 ();
 sg13g2_decap_4 FILLER_55_1012 ();
 sg13g2_decap_4 FILLER_55_1021 ();
 sg13g2_decap_8 FILLER_55_1035 ();
 sg13g2_decap_8 FILLER_55_1042 ();
 sg13g2_decap_8 FILLER_55_1049 ();
 sg13g2_decap_8 FILLER_55_1056 ();
 sg13g2_decap_8 FILLER_55_1063 ();
 sg13g2_decap_8 FILLER_55_1070 ();
 sg13g2_decap_8 FILLER_55_1077 ();
 sg13g2_decap_8 FILLER_55_1084 ();
 sg13g2_decap_8 FILLER_55_1091 ();
 sg13g2_decap_8 FILLER_55_1098 ();
 sg13g2_decap_8 FILLER_55_1105 ();
 sg13g2_decap_8 FILLER_55_1112 ();
 sg13g2_decap_8 FILLER_55_1119 ();
 sg13g2_decap_8 FILLER_55_1126 ();
 sg13g2_decap_8 FILLER_55_1133 ();
 sg13g2_decap_8 FILLER_55_1140 ();
 sg13g2_decap_8 FILLER_55_1147 ();
 sg13g2_decap_8 FILLER_55_1154 ();
 sg13g2_decap_8 FILLER_55_1161 ();
 sg13g2_decap_8 FILLER_55_1168 ();
 sg13g2_decap_8 FILLER_55_1175 ();
 sg13g2_decap_8 FILLER_55_1182 ();
 sg13g2_decap_8 FILLER_55_1189 ();
 sg13g2_decap_8 FILLER_55_1196 ();
 sg13g2_decap_8 FILLER_55_1203 ();
 sg13g2_decap_8 FILLER_55_1210 ();
 sg13g2_decap_8 FILLER_55_1217 ();
 sg13g2_decap_8 FILLER_55_1224 ();
 sg13g2_decap_8 FILLER_55_1231 ();
 sg13g2_decap_8 FILLER_55_1238 ();
 sg13g2_decap_8 FILLER_55_1245 ();
 sg13g2_decap_8 FILLER_55_1252 ();
 sg13g2_decap_8 FILLER_55_1259 ();
 sg13g2_decap_8 FILLER_55_1266 ();
 sg13g2_decap_8 FILLER_55_1273 ();
 sg13g2_decap_8 FILLER_55_1280 ();
 sg13g2_decap_8 FILLER_55_1287 ();
 sg13g2_decap_8 FILLER_55_1294 ();
 sg13g2_decap_8 FILLER_55_1301 ();
 sg13g2_decap_8 FILLER_55_1308 ();
 sg13g2_decap_8 FILLER_55_1315 ();
 sg13g2_decap_8 FILLER_55_1322 ();
 sg13g2_decap_8 FILLER_55_1329 ();
 sg13g2_decap_8 FILLER_55_1336 ();
 sg13g2_decap_8 FILLER_55_1343 ();
 sg13g2_decap_8 FILLER_55_1350 ();
 sg13g2_decap_8 FILLER_55_1357 ();
 sg13g2_decap_8 FILLER_55_1364 ();
 sg13g2_decap_8 FILLER_55_1371 ();
 sg13g2_decap_8 FILLER_55_1378 ();
 sg13g2_decap_8 FILLER_55_1385 ();
 sg13g2_decap_8 FILLER_55_1392 ();
 sg13g2_decap_8 FILLER_55_1399 ();
 sg13g2_decap_8 FILLER_55_1406 ();
 sg13g2_decap_8 FILLER_55_1413 ();
 sg13g2_decap_8 FILLER_55_1420 ();
 sg13g2_decap_8 FILLER_55_1427 ();
 sg13g2_decap_8 FILLER_55_1434 ();
 sg13g2_decap_8 FILLER_55_1441 ();
 sg13g2_decap_8 FILLER_55_1448 ();
 sg13g2_decap_8 FILLER_55_1455 ();
 sg13g2_decap_8 FILLER_55_1462 ();
 sg13g2_decap_8 FILLER_55_1469 ();
 sg13g2_decap_8 FILLER_55_1476 ();
 sg13g2_decap_8 FILLER_55_1483 ();
 sg13g2_decap_8 FILLER_55_1490 ();
 sg13g2_decap_8 FILLER_55_1497 ();
 sg13g2_decap_8 FILLER_55_1504 ();
 sg13g2_decap_8 FILLER_55_1511 ();
 sg13g2_decap_8 FILLER_55_1518 ();
 sg13g2_decap_8 FILLER_55_1525 ();
 sg13g2_decap_8 FILLER_55_1532 ();
 sg13g2_decap_8 FILLER_55_1539 ();
 sg13g2_decap_8 FILLER_55_1546 ();
 sg13g2_decap_8 FILLER_55_1553 ();
 sg13g2_decap_8 FILLER_55_1560 ();
 sg13g2_decap_8 FILLER_55_1567 ();
 sg13g2_decap_8 FILLER_55_1574 ();
 sg13g2_decap_8 FILLER_55_1581 ();
 sg13g2_decap_8 FILLER_55_1588 ();
 sg13g2_decap_8 FILLER_55_1595 ();
 sg13g2_decap_8 FILLER_55_1602 ();
 sg13g2_decap_8 FILLER_55_1609 ();
 sg13g2_decap_8 FILLER_55_1616 ();
 sg13g2_decap_8 FILLER_55_1623 ();
 sg13g2_decap_8 FILLER_55_1630 ();
 sg13g2_decap_8 FILLER_55_1637 ();
 sg13g2_decap_8 FILLER_55_1644 ();
 sg13g2_decap_8 FILLER_55_1651 ();
 sg13g2_decap_8 FILLER_55_1658 ();
 sg13g2_decap_8 FILLER_55_1665 ();
 sg13g2_decap_8 FILLER_55_1672 ();
 sg13g2_decap_8 FILLER_55_1679 ();
 sg13g2_decap_8 FILLER_55_1686 ();
 sg13g2_decap_8 FILLER_55_1693 ();
 sg13g2_decap_8 FILLER_55_1700 ();
 sg13g2_decap_8 FILLER_55_1707 ();
 sg13g2_decap_8 FILLER_55_1714 ();
 sg13g2_decap_8 FILLER_55_1721 ();
 sg13g2_decap_8 FILLER_55_1728 ();
 sg13g2_decap_8 FILLER_55_1735 ();
 sg13g2_decap_8 FILLER_55_1742 ();
 sg13g2_decap_8 FILLER_55_1749 ();
 sg13g2_decap_8 FILLER_55_1756 ();
 sg13g2_decap_4 FILLER_55_1763 ();
 sg13g2_fill_1 FILLER_55_1767 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_fill_2 FILLER_56_28 ();
 sg13g2_fill_1 FILLER_56_30 ();
 sg13g2_decap_8 FILLER_56_36 ();
 sg13g2_decap_8 FILLER_56_43 ();
 sg13g2_fill_2 FILLER_56_50 ();
 sg13g2_fill_1 FILLER_56_52 ();
 sg13g2_decap_4 FILLER_56_57 ();
 sg13g2_fill_1 FILLER_56_61 ();
 sg13g2_decap_4 FILLER_56_79 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_fill_2 FILLER_56_105 ();
 sg13g2_fill_1 FILLER_56_107 ();
 sg13g2_decap_4 FILLER_56_123 ();
 sg13g2_fill_2 FILLER_56_130 ();
 sg13g2_fill_1 FILLER_56_132 ();
 sg13g2_decap_8 FILLER_56_156 ();
 sg13g2_fill_1 FILLER_56_172 ();
 sg13g2_fill_1 FILLER_56_222 ();
 sg13g2_decap_8 FILLER_56_268 ();
 sg13g2_fill_2 FILLER_56_275 ();
 sg13g2_fill_1 FILLER_56_297 ();
 sg13g2_fill_2 FILLER_56_311 ();
 sg13g2_fill_2 FILLER_56_331 ();
 sg13g2_fill_1 FILLER_56_333 ();
 sg13g2_fill_2 FILLER_56_347 ();
 sg13g2_fill_2 FILLER_56_357 ();
 sg13g2_decap_4 FILLER_56_369 ();
 sg13g2_fill_2 FILLER_56_373 ();
 sg13g2_decap_8 FILLER_56_380 ();
 sg13g2_decap_4 FILLER_56_387 ();
 sg13g2_fill_1 FILLER_56_391 ();
 sg13g2_decap_8 FILLER_56_405 ();
 sg13g2_fill_2 FILLER_56_412 ();
 sg13g2_fill_1 FILLER_56_418 ();
 sg13g2_fill_1 FILLER_56_428 ();
 sg13g2_fill_1 FILLER_56_455 ();
 sg13g2_fill_2 FILLER_56_531 ();
 sg13g2_fill_1 FILLER_56_533 ();
 sg13g2_decap_4 FILLER_56_567 ();
 sg13g2_fill_2 FILLER_56_571 ();
 sg13g2_decap_8 FILLER_56_592 ();
 sg13g2_fill_1 FILLER_56_599 ();
 sg13g2_decap_8 FILLER_56_617 ();
 sg13g2_decap_8 FILLER_56_624 ();
 sg13g2_fill_2 FILLER_56_631 ();
 sg13g2_fill_1 FILLER_56_633 ();
 sg13g2_fill_1 FILLER_56_643 ();
 sg13g2_fill_2 FILLER_56_649 ();
 sg13g2_decap_8 FILLER_56_701 ();
 sg13g2_decap_8 FILLER_56_708 ();
 sg13g2_fill_2 FILLER_56_741 ();
 sg13g2_fill_1 FILLER_56_743 ();
 sg13g2_decap_8 FILLER_56_796 ();
 sg13g2_decap_8 FILLER_56_815 ();
 sg13g2_decap_4 FILLER_56_822 ();
 sg13g2_fill_2 FILLER_56_826 ();
 sg13g2_fill_1 FILLER_56_837 ();
 sg13g2_decap_4 FILLER_56_854 ();
 sg13g2_fill_1 FILLER_56_858 ();
 sg13g2_fill_1 FILLER_56_878 ();
 sg13g2_fill_2 FILLER_56_889 ();
 sg13g2_decap_8 FILLER_56_911 ();
 sg13g2_fill_1 FILLER_56_922 ();
 sg13g2_fill_1 FILLER_56_940 ();
 sg13g2_fill_1 FILLER_56_970 ();
 sg13g2_fill_2 FILLER_56_984 ();
 sg13g2_fill_1 FILLER_56_986 ();
 sg13g2_fill_1 FILLER_56_1002 ();
 sg13g2_decap_8 FILLER_56_1011 ();
 sg13g2_fill_2 FILLER_56_1018 ();
 sg13g2_fill_1 FILLER_56_1020 ();
 sg13g2_decap_8 FILLER_56_1026 ();
 sg13g2_decap_8 FILLER_56_1033 ();
 sg13g2_decap_8 FILLER_56_1040 ();
 sg13g2_decap_8 FILLER_56_1047 ();
 sg13g2_decap_8 FILLER_56_1054 ();
 sg13g2_decap_8 FILLER_56_1061 ();
 sg13g2_decap_8 FILLER_56_1068 ();
 sg13g2_decap_8 FILLER_56_1075 ();
 sg13g2_decap_8 FILLER_56_1082 ();
 sg13g2_decap_8 FILLER_56_1089 ();
 sg13g2_decap_8 FILLER_56_1096 ();
 sg13g2_decap_8 FILLER_56_1103 ();
 sg13g2_decap_8 FILLER_56_1110 ();
 sg13g2_decap_8 FILLER_56_1117 ();
 sg13g2_decap_8 FILLER_56_1124 ();
 sg13g2_decap_8 FILLER_56_1131 ();
 sg13g2_decap_8 FILLER_56_1138 ();
 sg13g2_decap_8 FILLER_56_1145 ();
 sg13g2_decap_8 FILLER_56_1152 ();
 sg13g2_decap_8 FILLER_56_1159 ();
 sg13g2_decap_8 FILLER_56_1166 ();
 sg13g2_decap_8 FILLER_56_1173 ();
 sg13g2_decap_8 FILLER_56_1180 ();
 sg13g2_decap_8 FILLER_56_1187 ();
 sg13g2_decap_8 FILLER_56_1194 ();
 sg13g2_decap_8 FILLER_56_1201 ();
 sg13g2_decap_8 FILLER_56_1208 ();
 sg13g2_decap_8 FILLER_56_1215 ();
 sg13g2_decap_8 FILLER_56_1222 ();
 sg13g2_decap_8 FILLER_56_1229 ();
 sg13g2_decap_8 FILLER_56_1236 ();
 sg13g2_decap_8 FILLER_56_1243 ();
 sg13g2_decap_8 FILLER_56_1250 ();
 sg13g2_decap_8 FILLER_56_1257 ();
 sg13g2_decap_8 FILLER_56_1264 ();
 sg13g2_decap_8 FILLER_56_1271 ();
 sg13g2_decap_8 FILLER_56_1278 ();
 sg13g2_decap_8 FILLER_56_1285 ();
 sg13g2_decap_8 FILLER_56_1292 ();
 sg13g2_decap_8 FILLER_56_1299 ();
 sg13g2_decap_8 FILLER_56_1306 ();
 sg13g2_decap_8 FILLER_56_1313 ();
 sg13g2_decap_8 FILLER_56_1320 ();
 sg13g2_decap_8 FILLER_56_1327 ();
 sg13g2_decap_8 FILLER_56_1334 ();
 sg13g2_decap_8 FILLER_56_1341 ();
 sg13g2_decap_8 FILLER_56_1348 ();
 sg13g2_decap_8 FILLER_56_1355 ();
 sg13g2_decap_8 FILLER_56_1362 ();
 sg13g2_decap_8 FILLER_56_1369 ();
 sg13g2_decap_8 FILLER_56_1376 ();
 sg13g2_decap_8 FILLER_56_1383 ();
 sg13g2_decap_8 FILLER_56_1390 ();
 sg13g2_decap_8 FILLER_56_1397 ();
 sg13g2_decap_8 FILLER_56_1404 ();
 sg13g2_decap_8 FILLER_56_1411 ();
 sg13g2_decap_8 FILLER_56_1418 ();
 sg13g2_decap_8 FILLER_56_1425 ();
 sg13g2_decap_8 FILLER_56_1432 ();
 sg13g2_decap_8 FILLER_56_1439 ();
 sg13g2_decap_8 FILLER_56_1446 ();
 sg13g2_decap_8 FILLER_56_1453 ();
 sg13g2_decap_8 FILLER_56_1460 ();
 sg13g2_decap_8 FILLER_56_1467 ();
 sg13g2_decap_8 FILLER_56_1474 ();
 sg13g2_decap_8 FILLER_56_1481 ();
 sg13g2_decap_8 FILLER_56_1488 ();
 sg13g2_decap_8 FILLER_56_1495 ();
 sg13g2_decap_8 FILLER_56_1502 ();
 sg13g2_decap_8 FILLER_56_1509 ();
 sg13g2_decap_8 FILLER_56_1516 ();
 sg13g2_decap_8 FILLER_56_1523 ();
 sg13g2_decap_8 FILLER_56_1530 ();
 sg13g2_decap_8 FILLER_56_1537 ();
 sg13g2_decap_8 FILLER_56_1544 ();
 sg13g2_decap_8 FILLER_56_1551 ();
 sg13g2_decap_8 FILLER_56_1558 ();
 sg13g2_decap_8 FILLER_56_1565 ();
 sg13g2_decap_8 FILLER_56_1572 ();
 sg13g2_decap_8 FILLER_56_1579 ();
 sg13g2_decap_8 FILLER_56_1586 ();
 sg13g2_decap_8 FILLER_56_1593 ();
 sg13g2_decap_8 FILLER_56_1600 ();
 sg13g2_decap_8 FILLER_56_1607 ();
 sg13g2_decap_8 FILLER_56_1614 ();
 sg13g2_decap_8 FILLER_56_1621 ();
 sg13g2_decap_8 FILLER_56_1628 ();
 sg13g2_decap_8 FILLER_56_1635 ();
 sg13g2_decap_8 FILLER_56_1642 ();
 sg13g2_decap_8 FILLER_56_1649 ();
 sg13g2_decap_8 FILLER_56_1656 ();
 sg13g2_decap_8 FILLER_56_1663 ();
 sg13g2_decap_8 FILLER_56_1670 ();
 sg13g2_decap_8 FILLER_56_1677 ();
 sg13g2_decap_8 FILLER_56_1684 ();
 sg13g2_decap_8 FILLER_56_1691 ();
 sg13g2_decap_8 FILLER_56_1698 ();
 sg13g2_decap_8 FILLER_56_1705 ();
 sg13g2_decap_8 FILLER_56_1712 ();
 sg13g2_decap_8 FILLER_56_1719 ();
 sg13g2_decap_8 FILLER_56_1726 ();
 sg13g2_decap_8 FILLER_56_1733 ();
 sg13g2_decap_8 FILLER_56_1740 ();
 sg13g2_decap_8 FILLER_56_1747 ();
 sg13g2_decap_8 FILLER_56_1754 ();
 sg13g2_decap_8 FILLER_56_1761 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_93 ();
 sg13g2_fill_2 FILLER_57_135 ();
 sg13g2_fill_1 FILLER_57_137 ();
 sg13g2_decap_8 FILLER_57_152 ();
 sg13g2_fill_1 FILLER_57_159 ();
 sg13g2_decap_4 FILLER_57_172 ();
 sg13g2_fill_2 FILLER_57_196 ();
 sg13g2_decap_8 FILLER_57_237 ();
 sg13g2_fill_1 FILLER_57_244 ();
 sg13g2_fill_2 FILLER_57_266 ();
 sg13g2_fill_2 FILLER_57_273 ();
 sg13g2_fill_1 FILLER_57_285 ();
 sg13g2_decap_4 FILLER_57_303 ();
 sg13g2_fill_1 FILLER_57_307 ();
 sg13g2_fill_2 FILLER_57_316 ();
 sg13g2_decap_4 FILLER_57_326 ();
 sg13g2_fill_1 FILLER_57_334 ();
 sg13g2_decap_4 FILLER_57_339 ();
 sg13g2_decap_8 FILLER_57_359 ();
 sg13g2_fill_2 FILLER_57_366 ();
 sg13g2_fill_1 FILLER_57_368 ();
 sg13g2_fill_1 FILLER_57_380 ();
 sg13g2_decap_8 FILLER_57_429 ();
 sg13g2_decap_4 FILLER_57_436 ();
 sg13g2_decap_4 FILLER_57_444 ();
 sg13g2_fill_2 FILLER_57_479 ();
 sg13g2_fill_1 FILLER_57_481 ();
 sg13g2_fill_2 FILLER_57_486 ();
 sg13g2_fill_1 FILLER_57_495 ();
 sg13g2_fill_2 FILLER_57_514 ();
 sg13g2_fill_2 FILLER_57_523 ();
 sg13g2_fill_1 FILLER_57_525 ();
 sg13g2_fill_2 FILLER_57_566 ();
 sg13g2_fill_1 FILLER_57_568 ();
 sg13g2_fill_2 FILLER_57_599 ();
 sg13g2_fill_1 FILLER_57_601 ();
 sg13g2_decap_4 FILLER_57_614 ();
 sg13g2_fill_1 FILLER_57_635 ();
 sg13g2_fill_1 FILLER_57_661 ();
 sg13g2_decap_4 FILLER_57_668 ();
 sg13g2_decap_4 FILLER_57_680 ();
 sg13g2_fill_1 FILLER_57_707 ();
 sg13g2_fill_1 FILLER_57_712 ();
 sg13g2_fill_1 FILLER_57_728 ();
 sg13g2_fill_2 FILLER_57_755 ();
 sg13g2_fill_2 FILLER_57_797 ();
 sg13g2_fill_1 FILLER_57_805 ();
 sg13g2_fill_2 FILLER_57_811 ();
 sg13g2_fill_1 FILLER_57_813 ();
 sg13g2_fill_2 FILLER_57_819 ();
 sg13g2_fill_1 FILLER_57_821 ();
 sg13g2_fill_2 FILLER_57_856 ();
 sg13g2_fill_1 FILLER_57_874 ();
 sg13g2_fill_1 FILLER_57_886 ();
 sg13g2_fill_2 FILLER_57_895 ();
 sg13g2_decap_4 FILLER_57_907 ();
 sg13g2_fill_1 FILLER_57_911 ();
 sg13g2_fill_1 FILLER_57_921 ();
 sg13g2_decap_8 FILLER_57_931 ();
 sg13g2_fill_1 FILLER_57_938 ();
 sg13g2_fill_2 FILLER_57_944 ();
 sg13g2_decap_8 FILLER_57_953 ();
 sg13g2_fill_2 FILLER_57_960 ();
 sg13g2_fill_1 FILLER_57_962 ();
 sg13g2_decap_4 FILLER_57_976 ();
 sg13g2_fill_2 FILLER_57_980 ();
 sg13g2_fill_1 FILLER_57_987 ();
 sg13g2_decap_8 FILLER_57_1012 ();
 sg13g2_decap_8 FILLER_57_1019 ();
 sg13g2_decap_8 FILLER_57_1026 ();
 sg13g2_decap_8 FILLER_57_1033 ();
 sg13g2_decap_8 FILLER_57_1040 ();
 sg13g2_decap_8 FILLER_57_1047 ();
 sg13g2_decap_8 FILLER_57_1054 ();
 sg13g2_decap_8 FILLER_57_1061 ();
 sg13g2_decap_8 FILLER_57_1068 ();
 sg13g2_decap_8 FILLER_57_1075 ();
 sg13g2_decap_8 FILLER_57_1082 ();
 sg13g2_decap_8 FILLER_57_1089 ();
 sg13g2_decap_8 FILLER_57_1096 ();
 sg13g2_decap_8 FILLER_57_1103 ();
 sg13g2_decap_8 FILLER_57_1110 ();
 sg13g2_decap_8 FILLER_57_1117 ();
 sg13g2_decap_8 FILLER_57_1124 ();
 sg13g2_decap_8 FILLER_57_1131 ();
 sg13g2_decap_8 FILLER_57_1138 ();
 sg13g2_decap_8 FILLER_57_1145 ();
 sg13g2_decap_8 FILLER_57_1152 ();
 sg13g2_decap_8 FILLER_57_1159 ();
 sg13g2_decap_8 FILLER_57_1166 ();
 sg13g2_decap_8 FILLER_57_1173 ();
 sg13g2_decap_8 FILLER_57_1180 ();
 sg13g2_decap_8 FILLER_57_1187 ();
 sg13g2_decap_8 FILLER_57_1194 ();
 sg13g2_decap_8 FILLER_57_1201 ();
 sg13g2_decap_8 FILLER_57_1208 ();
 sg13g2_decap_8 FILLER_57_1215 ();
 sg13g2_decap_8 FILLER_57_1222 ();
 sg13g2_decap_8 FILLER_57_1229 ();
 sg13g2_decap_8 FILLER_57_1236 ();
 sg13g2_decap_8 FILLER_57_1243 ();
 sg13g2_decap_8 FILLER_57_1250 ();
 sg13g2_decap_8 FILLER_57_1257 ();
 sg13g2_decap_8 FILLER_57_1264 ();
 sg13g2_decap_8 FILLER_57_1271 ();
 sg13g2_decap_8 FILLER_57_1278 ();
 sg13g2_decap_8 FILLER_57_1285 ();
 sg13g2_decap_8 FILLER_57_1292 ();
 sg13g2_decap_8 FILLER_57_1299 ();
 sg13g2_decap_8 FILLER_57_1306 ();
 sg13g2_decap_8 FILLER_57_1313 ();
 sg13g2_decap_8 FILLER_57_1320 ();
 sg13g2_decap_8 FILLER_57_1327 ();
 sg13g2_decap_8 FILLER_57_1334 ();
 sg13g2_decap_8 FILLER_57_1341 ();
 sg13g2_decap_8 FILLER_57_1348 ();
 sg13g2_decap_8 FILLER_57_1355 ();
 sg13g2_decap_8 FILLER_57_1362 ();
 sg13g2_decap_8 FILLER_57_1369 ();
 sg13g2_decap_8 FILLER_57_1376 ();
 sg13g2_decap_8 FILLER_57_1383 ();
 sg13g2_decap_8 FILLER_57_1390 ();
 sg13g2_decap_8 FILLER_57_1397 ();
 sg13g2_decap_8 FILLER_57_1404 ();
 sg13g2_decap_8 FILLER_57_1411 ();
 sg13g2_decap_8 FILLER_57_1418 ();
 sg13g2_decap_8 FILLER_57_1425 ();
 sg13g2_decap_8 FILLER_57_1432 ();
 sg13g2_decap_8 FILLER_57_1439 ();
 sg13g2_decap_8 FILLER_57_1446 ();
 sg13g2_decap_8 FILLER_57_1453 ();
 sg13g2_decap_8 FILLER_57_1460 ();
 sg13g2_decap_8 FILLER_57_1467 ();
 sg13g2_decap_8 FILLER_57_1474 ();
 sg13g2_decap_8 FILLER_57_1481 ();
 sg13g2_decap_8 FILLER_57_1488 ();
 sg13g2_decap_8 FILLER_57_1495 ();
 sg13g2_decap_8 FILLER_57_1502 ();
 sg13g2_decap_8 FILLER_57_1509 ();
 sg13g2_decap_8 FILLER_57_1516 ();
 sg13g2_decap_8 FILLER_57_1523 ();
 sg13g2_decap_8 FILLER_57_1530 ();
 sg13g2_decap_8 FILLER_57_1537 ();
 sg13g2_decap_8 FILLER_57_1544 ();
 sg13g2_decap_8 FILLER_57_1551 ();
 sg13g2_decap_8 FILLER_57_1558 ();
 sg13g2_decap_8 FILLER_57_1565 ();
 sg13g2_decap_8 FILLER_57_1572 ();
 sg13g2_decap_8 FILLER_57_1579 ();
 sg13g2_decap_8 FILLER_57_1586 ();
 sg13g2_decap_8 FILLER_57_1593 ();
 sg13g2_decap_8 FILLER_57_1600 ();
 sg13g2_decap_8 FILLER_57_1607 ();
 sg13g2_decap_8 FILLER_57_1614 ();
 sg13g2_decap_8 FILLER_57_1621 ();
 sg13g2_decap_8 FILLER_57_1628 ();
 sg13g2_decap_8 FILLER_57_1635 ();
 sg13g2_decap_8 FILLER_57_1642 ();
 sg13g2_decap_8 FILLER_57_1649 ();
 sg13g2_decap_8 FILLER_57_1656 ();
 sg13g2_decap_8 FILLER_57_1663 ();
 sg13g2_decap_8 FILLER_57_1670 ();
 sg13g2_decap_8 FILLER_57_1677 ();
 sg13g2_decap_8 FILLER_57_1684 ();
 sg13g2_decap_8 FILLER_57_1691 ();
 sg13g2_decap_8 FILLER_57_1698 ();
 sg13g2_decap_8 FILLER_57_1705 ();
 sg13g2_decap_8 FILLER_57_1712 ();
 sg13g2_decap_8 FILLER_57_1719 ();
 sg13g2_decap_8 FILLER_57_1726 ();
 sg13g2_decap_8 FILLER_57_1733 ();
 sg13g2_decap_8 FILLER_57_1740 ();
 sg13g2_decap_8 FILLER_57_1747 ();
 sg13g2_decap_8 FILLER_57_1754 ();
 sg13g2_decap_8 FILLER_57_1761 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_4 FILLER_58_7 ();
 sg13g2_fill_2 FILLER_58_11 ();
 sg13g2_fill_2 FILLER_58_30 ();
 sg13g2_fill_1 FILLER_58_36 ();
 sg13g2_fill_1 FILLER_58_73 ();
 sg13g2_fill_1 FILLER_58_87 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_fill_2 FILLER_58_105 ();
 sg13g2_fill_1 FILLER_58_120 ();
 sg13g2_fill_1 FILLER_58_193 ();
 sg13g2_fill_1 FILLER_58_207 ();
 sg13g2_decap_8 FILLER_58_237 ();
 sg13g2_decap_4 FILLER_58_244 ();
 sg13g2_decap_8 FILLER_58_253 ();
 sg13g2_fill_2 FILLER_58_288 ();
 sg13g2_fill_1 FILLER_58_295 ();
 sg13g2_fill_2 FILLER_58_325 ();
 sg13g2_decap_8 FILLER_58_335 ();
 sg13g2_fill_2 FILLER_58_342 ();
 sg13g2_fill_2 FILLER_58_363 ();
 sg13g2_decap_8 FILLER_58_391 ();
 sg13g2_fill_2 FILLER_58_398 ();
 sg13g2_fill_1 FILLER_58_400 ();
 sg13g2_decap_8 FILLER_58_409 ();
 sg13g2_fill_2 FILLER_58_441 ();
 sg13g2_decap_4 FILLER_58_448 ();
 sg13g2_fill_1 FILLER_58_476 ();
 sg13g2_decap_4 FILLER_58_481 ();
 sg13g2_fill_2 FILLER_58_553 ();
 sg13g2_fill_1 FILLER_58_555 ();
 sg13g2_fill_1 FILLER_58_562 ();
 sg13g2_fill_2 FILLER_58_571 ();
 sg13g2_fill_1 FILLER_58_573 ();
 sg13g2_decap_8 FILLER_58_599 ();
 sg13g2_decap_4 FILLER_58_606 ();
 sg13g2_fill_1 FILLER_58_610 ();
 sg13g2_fill_1 FILLER_58_616 ();
 sg13g2_decap_8 FILLER_58_622 ();
 sg13g2_fill_2 FILLER_58_629 ();
 sg13g2_fill_2 FILLER_58_650 ();
 sg13g2_fill_2 FILLER_58_673 ();
 sg13g2_fill_1 FILLER_58_675 ();
 sg13g2_decap_4 FILLER_58_681 ();
 sg13g2_fill_2 FILLER_58_685 ();
 sg13g2_decap_8 FILLER_58_701 ();
 sg13g2_fill_2 FILLER_58_708 ();
 sg13g2_fill_1 FILLER_58_719 ();
 sg13g2_fill_2 FILLER_58_747 ();
 sg13g2_fill_1 FILLER_58_749 ();
 sg13g2_decap_8 FILLER_58_771 ();
 sg13g2_decap_4 FILLER_58_778 ();
 sg13g2_fill_1 FILLER_58_788 ();
 sg13g2_fill_2 FILLER_58_794 ();
 sg13g2_fill_2 FILLER_58_801 ();
 sg13g2_fill_1 FILLER_58_803 ();
 sg13g2_decap_8 FILLER_58_829 ();
 sg13g2_fill_2 FILLER_58_836 ();
 sg13g2_fill_1 FILLER_58_838 ();
 sg13g2_decap_8 FILLER_58_844 ();
 sg13g2_decap_8 FILLER_58_851 ();
 sg13g2_fill_1 FILLER_58_858 ();
 sg13g2_fill_2 FILLER_58_882 ();
 sg13g2_fill_2 FILLER_58_902 ();
 sg13g2_fill_1 FILLER_58_904 ();
 sg13g2_fill_2 FILLER_58_913 ();
 sg13g2_fill_2 FILLER_58_933 ();
 sg13g2_fill_1 FILLER_58_935 ();
 sg13g2_fill_1 FILLER_58_941 ();
 sg13g2_decap_8 FILLER_58_952 ();
 sg13g2_fill_1 FILLER_58_959 ();
 sg13g2_fill_2 FILLER_58_984 ();
 sg13g2_fill_1 FILLER_58_986 ();
 sg13g2_decap_8 FILLER_58_1006 ();
 sg13g2_decap_8 FILLER_58_1013 ();
 sg13g2_decap_8 FILLER_58_1020 ();
 sg13g2_decap_8 FILLER_58_1027 ();
 sg13g2_decap_8 FILLER_58_1034 ();
 sg13g2_decap_8 FILLER_58_1041 ();
 sg13g2_decap_8 FILLER_58_1048 ();
 sg13g2_decap_8 FILLER_58_1055 ();
 sg13g2_decap_8 FILLER_58_1062 ();
 sg13g2_decap_8 FILLER_58_1069 ();
 sg13g2_decap_8 FILLER_58_1076 ();
 sg13g2_decap_8 FILLER_58_1083 ();
 sg13g2_decap_8 FILLER_58_1090 ();
 sg13g2_decap_8 FILLER_58_1097 ();
 sg13g2_decap_8 FILLER_58_1104 ();
 sg13g2_decap_8 FILLER_58_1111 ();
 sg13g2_decap_8 FILLER_58_1118 ();
 sg13g2_decap_8 FILLER_58_1125 ();
 sg13g2_decap_8 FILLER_58_1132 ();
 sg13g2_decap_8 FILLER_58_1139 ();
 sg13g2_decap_8 FILLER_58_1146 ();
 sg13g2_decap_8 FILLER_58_1153 ();
 sg13g2_decap_8 FILLER_58_1160 ();
 sg13g2_decap_8 FILLER_58_1167 ();
 sg13g2_decap_8 FILLER_58_1174 ();
 sg13g2_decap_8 FILLER_58_1181 ();
 sg13g2_decap_8 FILLER_58_1188 ();
 sg13g2_decap_8 FILLER_58_1195 ();
 sg13g2_decap_8 FILLER_58_1202 ();
 sg13g2_decap_8 FILLER_58_1209 ();
 sg13g2_decap_8 FILLER_58_1216 ();
 sg13g2_decap_8 FILLER_58_1223 ();
 sg13g2_decap_8 FILLER_58_1230 ();
 sg13g2_decap_8 FILLER_58_1237 ();
 sg13g2_decap_8 FILLER_58_1244 ();
 sg13g2_decap_8 FILLER_58_1251 ();
 sg13g2_decap_8 FILLER_58_1258 ();
 sg13g2_decap_8 FILLER_58_1265 ();
 sg13g2_decap_8 FILLER_58_1272 ();
 sg13g2_decap_8 FILLER_58_1279 ();
 sg13g2_decap_8 FILLER_58_1286 ();
 sg13g2_decap_8 FILLER_58_1293 ();
 sg13g2_decap_8 FILLER_58_1300 ();
 sg13g2_decap_8 FILLER_58_1307 ();
 sg13g2_decap_8 FILLER_58_1314 ();
 sg13g2_decap_8 FILLER_58_1321 ();
 sg13g2_decap_8 FILLER_58_1328 ();
 sg13g2_decap_8 FILLER_58_1335 ();
 sg13g2_decap_8 FILLER_58_1342 ();
 sg13g2_decap_8 FILLER_58_1349 ();
 sg13g2_decap_8 FILLER_58_1356 ();
 sg13g2_decap_8 FILLER_58_1363 ();
 sg13g2_decap_8 FILLER_58_1370 ();
 sg13g2_decap_8 FILLER_58_1377 ();
 sg13g2_decap_8 FILLER_58_1384 ();
 sg13g2_decap_8 FILLER_58_1391 ();
 sg13g2_decap_8 FILLER_58_1398 ();
 sg13g2_decap_8 FILLER_58_1405 ();
 sg13g2_decap_8 FILLER_58_1412 ();
 sg13g2_decap_8 FILLER_58_1419 ();
 sg13g2_decap_8 FILLER_58_1426 ();
 sg13g2_decap_8 FILLER_58_1433 ();
 sg13g2_decap_8 FILLER_58_1440 ();
 sg13g2_decap_8 FILLER_58_1447 ();
 sg13g2_decap_8 FILLER_58_1454 ();
 sg13g2_decap_8 FILLER_58_1461 ();
 sg13g2_decap_8 FILLER_58_1468 ();
 sg13g2_decap_8 FILLER_58_1475 ();
 sg13g2_decap_8 FILLER_58_1482 ();
 sg13g2_decap_8 FILLER_58_1489 ();
 sg13g2_decap_8 FILLER_58_1496 ();
 sg13g2_decap_8 FILLER_58_1503 ();
 sg13g2_decap_8 FILLER_58_1510 ();
 sg13g2_decap_8 FILLER_58_1517 ();
 sg13g2_decap_8 FILLER_58_1524 ();
 sg13g2_decap_8 FILLER_58_1531 ();
 sg13g2_decap_8 FILLER_58_1538 ();
 sg13g2_decap_8 FILLER_58_1545 ();
 sg13g2_decap_8 FILLER_58_1552 ();
 sg13g2_decap_8 FILLER_58_1559 ();
 sg13g2_decap_8 FILLER_58_1566 ();
 sg13g2_decap_8 FILLER_58_1573 ();
 sg13g2_decap_8 FILLER_58_1580 ();
 sg13g2_decap_8 FILLER_58_1587 ();
 sg13g2_decap_8 FILLER_58_1594 ();
 sg13g2_decap_8 FILLER_58_1601 ();
 sg13g2_decap_8 FILLER_58_1608 ();
 sg13g2_decap_8 FILLER_58_1615 ();
 sg13g2_decap_8 FILLER_58_1622 ();
 sg13g2_decap_8 FILLER_58_1629 ();
 sg13g2_decap_8 FILLER_58_1636 ();
 sg13g2_decap_8 FILLER_58_1643 ();
 sg13g2_decap_8 FILLER_58_1650 ();
 sg13g2_decap_8 FILLER_58_1657 ();
 sg13g2_decap_8 FILLER_58_1664 ();
 sg13g2_decap_8 FILLER_58_1671 ();
 sg13g2_decap_8 FILLER_58_1678 ();
 sg13g2_decap_8 FILLER_58_1685 ();
 sg13g2_decap_8 FILLER_58_1692 ();
 sg13g2_decap_8 FILLER_58_1699 ();
 sg13g2_decap_8 FILLER_58_1706 ();
 sg13g2_decap_8 FILLER_58_1713 ();
 sg13g2_decap_8 FILLER_58_1720 ();
 sg13g2_decap_8 FILLER_58_1727 ();
 sg13g2_decap_8 FILLER_58_1734 ();
 sg13g2_decap_8 FILLER_58_1741 ();
 sg13g2_decap_8 FILLER_58_1748 ();
 sg13g2_decap_8 FILLER_58_1755 ();
 sg13g2_decap_4 FILLER_58_1762 ();
 sg13g2_fill_2 FILLER_58_1766 ();
 sg13g2_decap_4 FILLER_59_0 ();
 sg13g2_decap_4 FILLER_59_44 ();
 sg13g2_fill_1 FILLER_59_52 ();
 sg13g2_fill_1 FILLER_59_57 ();
 sg13g2_decap_4 FILLER_59_68 ();
 sg13g2_fill_2 FILLER_59_72 ();
 sg13g2_decap_8 FILLER_59_110 ();
 sg13g2_fill_2 FILLER_59_134 ();
 sg13g2_fill_1 FILLER_59_153 ();
 sg13g2_decap_8 FILLER_59_267 ();
 sg13g2_fill_1 FILLER_59_274 ();
 sg13g2_fill_2 FILLER_59_327 ();
 sg13g2_fill_1 FILLER_59_329 ();
 sg13g2_decap_4 FILLER_59_335 ();
 sg13g2_fill_2 FILLER_59_339 ();
 sg13g2_decap_4 FILLER_59_345 ();
 sg13g2_fill_2 FILLER_59_349 ();
 sg13g2_fill_1 FILLER_59_375 ();
 sg13g2_fill_2 FILLER_59_380 ();
 sg13g2_fill_1 FILLER_59_382 ();
 sg13g2_fill_2 FILLER_59_388 ();
 sg13g2_decap_4 FILLER_59_399 ();
 sg13g2_fill_1 FILLER_59_403 ();
 sg13g2_fill_2 FILLER_59_430 ();
 sg13g2_decap_8 FILLER_59_478 ();
 sg13g2_decap_8 FILLER_59_485 ();
 sg13g2_fill_2 FILLER_59_492 ();
 sg13g2_fill_1 FILLER_59_507 ();
 sg13g2_fill_2 FILLER_59_520 ();
 sg13g2_fill_1 FILLER_59_527 ();
 sg13g2_decap_8 FILLER_59_538 ();
 sg13g2_decap_8 FILLER_59_545 ();
 sg13g2_decap_4 FILLER_59_552 ();
 sg13g2_fill_2 FILLER_59_560 ();
 sg13g2_fill_2 FILLER_59_572 ();
 sg13g2_fill_1 FILLER_59_574 ();
 sg13g2_decap_8 FILLER_59_593 ();
 sg13g2_decap_8 FILLER_59_600 ();
 sg13g2_fill_1 FILLER_59_607 ();
 sg13g2_decap_4 FILLER_59_634 ();
 sg13g2_fill_1 FILLER_59_638 ();
 sg13g2_fill_1 FILLER_59_696 ();
 sg13g2_fill_1 FILLER_59_723 ();
 sg13g2_fill_1 FILLER_59_778 ();
 sg13g2_fill_2 FILLER_59_787 ();
 sg13g2_fill_2 FILLER_59_828 ();
 sg13g2_decap_4 FILLER_59_848 ();
 sg13g2_fill_1 FILLER_59_852 ();
 sg13g2_fill_1 FILLER_59_865 ();
 sg13g2_decap_8 FILLER_59_884 ();
 sg13g2_fill_1 FILLER_59_891 ();
 sg13g2_decap_4 FILLER_59_905 ();
 sg13g2_fill_2 FILLER_59_909 ();
 sg13g2_fill_2 FILLER_59_929 ();
 sg13g2_decap_4 FILLER_59_952 ();
 sg13g2_fill_2 FILLER_59_956 ();
 sg13g2_decap_8 FILLER_59_981 ();
 sg13g2_decap_8 FILLER_59_988 ();
 sg13g2_decap_8 FILLER_59_995 ();
 sg13g2_decap_8 FILLER_59_1002 ();
 sg13g2_decap_8 FILLER_59_1009 ();
 sg13g2_decap_8 FILLER_59_1016 ();
 sg13g2_decap_8 FILLER_59_1023 ();
 sg13g2_decap_8 FILLER_59_1030 ();
 sg13g2_decap_8 FILLER_59_1037 ();
 sg13g2_decap_8 FILLER_59_1044 ();
 sg13g2_decap_8 FILLER_59_1051 ();
 sg13g2_decap_8 FILLER_59_1058 ();
 sg13g2_decap_8 FILLER_59_1065 ();
 sg13g2_decap_8 FILLER_59_1072 ();
 sg13g2_decap_8 FILLER_59_1079 ();
 sg13g2_decap_8 FILLER_59_1086 ();
 sg13g2_decap_8 FILLER_59_1093 ();
 sg13g2_decap_8 FILLER_59_1100 ();
 sg13g2_decap_8 FILLER_59_1107 ();
 sg13g2_decap_8 FILLER_59_1114 ();
 sg13g2_decap_8 FILLER_59_1121 ();
 sg13g2_decap_8 FILLER_59_1128 ();
 sg13g2_decap_8 FILLER_59_1135 ();
 sg13g2_decap_8 FILLER_59_1142 ();
 sg13g2_decap_8 FILLER_59_1149 ();
 sg13g2_decap_8 FILLER_59_1156 ();
 sg13g2_decap_8 FILLER_59_1163 ();
 sg13g2_decap_8 FILLER_59_1170 ();
 sg13g2_decap_8 FILLER_59_1177 ();
 sg13g2_decap_8 FILLER_59_1184 ();
 sg13g2_decap_8 FILLER_59_1191 ();
 sg13g2_decap_8 FILLER_59_1198 ();
 sg13g2_decap_8 FILLER_59_1205 ();
 sg13g2_decap_8 FILLER_59_1212 ();
 sg13g2_decap_8 FILLER_59_1219 ();
 sg13g2_decap_8 FILLER_59_1226 ();
 sg13g2_decap_8 FILLER_59_1233 ();
 sg13g2_decap_8 FILLER_59_1240 ();
 sg13g2_decap_8 FILLER_59_1247 ();
 sg13g2_decap_8 FILLER_59_1254 ();
 sg13g2_decap_8 FILLER_59_1261 ();
 sg13g2_decap_8 FILLER_59_1268 ();
 sg13g2_decap_8 FILLER_59_1275 ();
 sg13g2_decap_8 FILLER_59_1282 ();
 sg13g2_decap_8 FILLER_59_1289 ();
 sg13g2_decap_8 FILLER_59_1296 ();
 sg13g2_decap_8 FILLER_59_1303 ();
 sg13g2_decap_8 FILLER_59_1310 ();
 sg13g2_decap_8 FILLER_59_1317 ();
 sg13g2_decap_8 FILLER_59_1324 ();
 sg13g2_decap_8 FILLER_59_1331 ();
 sg13g2_decap_8 FILLER_59_1338 ();
 sg13g2_decap_8 FILLER_59_1345 ();
 sg13g2_decap_8 FILLER_59_1352 ();
 sg13g2_decap_8 FILLER_59_1359 ();
 sg13g2_decap_8 FILLER_59_1366 ();
 sg13g2_decap_8 FILLER_59_1373 ();
 sg13g2_decap_8 FILLER_59_1380 ();
 sg13g2_decap_8 FILLER_59_1387 ();
 sg13g2_decap_8 FILLER_59_1394 ();
 sg13g2_decap_8 FILLER_59_1401 ();
 sg13g2_decap_8 FILLER_59_1408 ();
 sg13g2_decap_8 FILLER_59_1415 ();
 sg13g2_decap_8 FILLER_59_1422 ();
 sg13g2_decap_8 FILLER_59_1429 ();
 sg13g2_decap_8 FILLER_59_1436 ();
 sg13g2_decap_8 FILLER_59_1443 ();
 sg13g2_decap_8 FILLER_59_1450 ();
 sg13g2_decap_8 FILLER_59_1457 ();
 sg13g2_decap_8 FILLER_59_1464 ();
 sg13g2_decap_8 FILLER_59_1471 ();
 sg13g2_decap_8 FILLER_59_1478 ();
 sg13g2_decap_8 FILLER_59_1485 ();
 sg13g2_decap_8 FILLER_59_1492 ();
 sg13g2_decap_8 FILLER_59_1499 ();
 sg13g2_decap_8 FILLER_59_1506 ();
 sg13g2_decap_8 FILLER_59_1513 ();
 sg13g2_decap_8 FILLER_59_1520 ();
 sg13g2_decap_8 FILLER_59_1527 ();
 sg13g2_decap_8 FILLER_59_1534 ();
 sg13g2_decap_8 FILLER_59_1541 ();
 sg13g2_decap_8 FILLER_59_1548 ();
 sg13g2_decap_8 FILLER_59_1555 ();
 sg13g2_decap_8 FILLER_59_1562 ();
 sg13g2_decap_8 FILLER_59_1569 ();
 sg13g2_decap_8 FILLER_59_1576 ();
 sg13g2_decap_8 FILLER_59_1583 ();
 sg13g2_decap_8 FILLER_59_1590 ();
 sg13g2_decap_8 FILLER_59_1597 ();
 sg13g2_decap_8 FILLER_59_1604 ();
 sg13g2_decap_8 FILLER_59_1611 ();
 sg13g2_decap_8 FILLER_59_1618 ();
 sg13g2_decap_8 FILLER_59_1625 ();
 sg13g2_decap_8 FILLER_59_1632 ();
 sg13g2_decap_8 FILLER_59_1639 ();
 sg13g2_decap_8 FILLER_59_1646 ();
 sg13g2_decap_8 FILLER_59_1653 ();
 sg13g2_decap_8 FILLER_59_1660 ();
 sg13g2_decap_8 FILLER_59_1667 ();
 sg13g2_decap_8 FILLER_59_1674 ();
 sg13g2_decap_8 FILLER_59_1681 ();
 sg13g2_decap_8 FILLER_59_1688 ();
 sg13g2_decap_8 FILLER_59_1695 ();
 sg13g2_decap_8 FILLER_59_1702 ();
 sg13g2_decap_8 FILLER_59_1709 ();
 sg13g2_decap_8 FILLER_59_1716 ();
 sg13g2_decap_8 FILLER_59_1723 ();
 sg13g2_decap_8 FILLER_59_1730 ();
 sg13g2_decap_8 FILLER_59_1737 ();
 sg13g2_decap_8 FILLER_59_1744 ();
 sg13g2_decap_8 FILLER_59_1751 ();
 sg13g2_decap_8 FILLER_59_1758 ();
 sg13g2_fill_2 FILLER_59_1765 ();
 sg13g2_fill_1 FILLER_59_1767 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_fill_2 FILLER_60_14 ();
 sg13g2_fill_1 FILLER_60_16 ();
 sg13g2_decap_4 FILLER_60_69 ();
 sg13g2_fill_2 FILLER_60_73 ();
 sg13g2_decap_4 FILLER_60_80 ();
 sg13g2_fill_1 FILLER_60_84 ();
 sg13g2_fill_2 FILLER_60_103 ();
 sg13g2_fill_1 FILLER_60_105 ();
 sg13g2_fill_2 FILLER_60_142 ();
 sg13g2_fill_1 FILLER_60_144 ();
 sg13g2_fill_2 FILLER_60_182 ();
 sg13g2_fill_1 FILLER_60_184 ();
 sg13g2_fill_2 FILLER_60_195 ();
 sg13g2_fill_1 FILLER_60_206 ();
 sg13g2_fill_1 FILLER_60_217 ();
 sg13g2_fill_2 FILLER_60_229 ();
 sg13g2_fill_2 FILLER_60_244 ();
 sg13g2_fill_1 FILLER_60_246 ();
 sg13g2_fill_1 FILLER_60_260 ();
 sg13g2_fill_1 FILLER_60_296 ();
 sg13g2_fill_2 FILLER_60_310 ();
 sg13g2_fill_1 FILLER_60_319 ();
 sg13g2_fill_2 FILLER_60_365 ();
 sg13g2_fill_1 FILLER_60_367 ();
 sg13g2_fill_2 FILLER_60_385 ();
 sg13g2_fill_1 FILLER_60_387 ();
 sg13g2_decap_8 FILLER_60_398 ();
 sg13g2_fill_2 FILLER_60_405 ();
 sg13g2_decap_4 FILLER_60_412 ();
 sg13g2_fill_2 FILLER_60_443 ();
 sg13g2_decap_4 FILLER_60_457 ();
 sg13g2_fill_2 FILLER_60_461 ();
 sg13g2_decap_8 FILLER_60_487 ();
 sg13g2_decap_8 FILLER_60_494 ();
 sg13g2_fill_1 FILLER_60_513 ();
 sg13g2_fill_2 FILLER_60_523 ();
 sg13g2_fill_2 FILLER_60_534 ();
 sg13g2_fill_1 FILLER_60_536 ();
 sg13g2_fill_1 FILLER_60_542 ();
 sg13g2_fill_1 FILLER_60_547 ();
 sg13g2_fill_2 FILLER_60_560 ();
 sg13g2_decap_8 FILLER_60_574 ();
 sg13g2_decap_4 FILLER_60_581 ();
 sg13g2_fill_2 FILLER_60_585 ();
 sg13g2_decap_4 FILLER_60_593 ();
 sg13g2_fill_1 FILLER_60_619 ();
 sg13g2_decap_4 FILLER_60_637 ();
 sg13g2_decap_4 FILLER_60_648 ();
 sg13g2_fill_2 FILLER_60_659 ();
 sg13g2_decap_8 FILLER_60_666 ();
 sg13g2_fill_2 FILLER_60_673 ();
 sg13g2_fill_1 FILLER_60_709 ();
 sg13g2_decap_8 FILLER_60_715 ();
 sg13g2_fill_2 FILLER_60_722 ();
 sg13g2_decap_4 FILLER_60_729 ();
 sg13g2_fill_1 FILLER_60_733 ();
 sg13g2_fill_2 FILLER_60_739 ();
 sg13g2_fill_1 FILLER_60_741 ();
 sg13g2_decap_4 FILLER_60_755 ();
 sg13g2_fill_1 FILLER_60_759 ();
 sg13g2_decap_8 FILLER_60_766 ();
 sg13g2_decap_8 FILLER_60_773 ();
 sg13g2_decap_8 FILLER_60_780 ();
 sg13g2_decap_8 FILLER_60_787 ();
 sg13g2_fill_1 FILLER_60_800 ();
 sg13g2_decap_8 FILLER_60_809 ();
 sg13g2_decap_8 FILLER_60_824 ();
 sg13g2_decap_4 FILLER_60_851 ();
 sg13g2_decap_8 FILLER_60_873 ();
 sg13g2_fill_2 FILLER_60_880 ();
 sg13g2_fill_1 FILLER_60_882 ();
 sg13g2_decap_4 FILLER_60_914 ();
 sg13g2_fill_1 FILLER_60_918 ();
 sg13g2_decap_8 FILLER_60_923 ();
 sg13g2_decap_8 FILLER_60_930 ();
 sg13g2_fill_2 FILLER_60_937 ();
 sg13g2_decap_4 FILLER_60_948 ();
 sg13g2_fill_1 FILLER_60_952 ();
 sg13g2_fill_2 FILLER_60_957 ();
 sg13g2_fill_1 FILLER_60_959 ();
 sg13g2_fill_1 FILLER_60_968 ();
 sg13g2_decap_8 FILLER_60_978 ();
 sg13g2_decap_8 FILLER_60_985 ();
 sg13g2_decap_8 FILLER_60_992 ();
 sg13g2_decap_8 FILLER_60_999 ();
 sg13g2_decap_8 FILLER_60_1006 ();
 sg13g2_decap_8 FILLER_60_1013 ();
 sg13g2_decap_8 FILLER_60_1020 ();
 sg13g2_decap_8 FILLER_60_1027 ();
 sg13g2_decap_8 FILLER_60_1034 ();
 sg13g2_decap_8 FILLER_60_1041 ();
 sg13g2_decap_8 FILLER_60_1048 ();
 sg13g2_decap_8 FILLER_60_1055 ();
 sg13g2_decap_8 FILLER_60_1062 ();
 sg13g2_decap_8 FILLER_60_1069 ();
 sg13g2_decap_8 FILLER_60_1076 ();
 sg13g2_decap_8 FILLER_60_1083 ();
 sg13g2_decap_8 FILLER_60_1090 ();
 sg13g2_decap_8 FILLER_60_1097 ();
 sg13g2_decap_8 FILLER_60_1104 ();
 sg13g2_decap_8 FILLER_60_1111 ();
 sg13g2_decap_8 FILLER_60_1118 ();
 sg13g2_decap_8 FILLER_60_1125 ();
 sg13g2_decap_8 FILLER_60_1132 ();
 sg13g2_decap_8 FILLER_60_1139 ();
 sg13g2_decap_8 FILLER_60_1146 ();
 sg13g2_decap_8 FILLER_60_1153 ();
 sg13g2_decap_8 FILLER_60_1160 ();
 sg13g2_decap_8 FILLER_60_1167 ();
 sg13g2_decap_8 FILLER_60_1174 ();
 sg13g2_decap_8 FILLER_60_1181 ();
 sg13g2_decap_8 FILLER_60_1188 ();
 sg13g2_decap_8 FILLER_60_1195 ();
 sg13g2_decap_8 FILLER_60_1202 ();
 sg13g2_decap_8 FILLER_60_1209 ();
 sg13g2_decap_8 FILLER_60_1216 ();
 sg13g2_decap_8 FILLER_60_1223 ();
 sg13g2_decap_8 FILLER_60_1230 ();
 sg13g2_decap_8 FILLER_60_1237 ();
 sg13g2_decap_8 FILLER_60_1244 ();
 sg13g2_decap_8 FILLER_60_1251 ();
 sg13g2_decap_8 FILLER_60_1258 ();
 sg13g2_decap_8 FILLER_60_1265 ();
 sg13g2_decap_8 FILLER_60_1272 ();
 sg13g2_decap_8 FILLER_60_1279 ();
 sg13g2_decap_8 FILLER_60_1286 ();
 sg13g2_decap_8 FILLER_60_1293 ();
 sg13g2_decap_8 FILLER_60_1300 ();
 sg13g2_decap_8 FILLER_60_1307 ();
 sg13g2_decap_8 FILLER_60_1314 ();
 sg13g2_decap_8 FILLER_60_1321 ();
 sg13g2_decap_8 FILLER_60_1328 ();
 sg13g2_decap_8 FILLER_60_1335 ();
 sg13g2_decap_8 FILLER_60_1342 ();
 sg13g2_decap_8 FILLER_60_1349 ();
 sg13g2_decap_8 FILLER_60_1356 ();
 sg13g2_decap_8 FILLER_60_1363 ();
 sg13g2_decap_8 FILLER_60_1370 ();
 sg13g2_decap_8 FILLER_60_1377 ();
 sg13g2_decap_8 FILLER_60_1384 ();
 sg13g2_decap_8 FILLER_60_1391 ();
 sg13g2_decap_8 FILLER_60_1398 ();
 sg13g2_decap_8 FILLER_60_1405 ();
 sg13g2_decap_8 FILLER_60_1412 ();
 sg13g2_decap_8 FILLER_60_1419 ();
 sg13g2_decap_8 FILLER_60_1426 ();
 sg13g2_decap_8 FILLER_60_1433 ();
 sg13g2_decap_8 FILLER_60_1440 ();
 sg13g2_decap_8 FILLER_60_1447 ();
 sg13g2_decap_8 FILLER_60_1454 ();
 sg13g2_decap_8 FILLER_60_1461 ();
 sg13g2_decap_8 FILLER_60_1468 ();
 sg13g2_decap_8 FILLER_60_1475 ();
 sg13g2_decap_8 FILLER_60_1482 ();
 sg13g2_decap_8 FILLER_60_1489 ();
 sg13g2_decap_8 FILLER_60_1496 ();
 sg13g2_decap_8 FILLER_60_1503 ();
 sg13g2_decap_8 FILLER_60_1510 ();
 sg13g2_decap_8 FILLER_60_1517 ();
 sg13g2_decap_8 FILLER_60_1524 ();
 sg13g2_decap_8 FILLER_60_1531 ();
 sg13g2_decap_8 FILLER_60_1538 ();
 sg13g2_decap_8 FILLER_60_1545 ();
 sg13g2_decap_8 FILLER_60_1552 ();
 sg13g2_decap_8 FILLER_60_1559 ();
 sg13g2_decap_8 FILLER_60_1566 ();
 sg13g2_decap_8 FILLER_60_1573 ();
 sg13g2_decap_8 FILLER_60_1580 ();
 sg13g2_decap_8 FILLER_60_1587 ();
 sg13g2_decap_8 FILLER_60_1594 ();
 sg13g2_decap_8 FILLER_60_1601 ();
 sg13g2_decap_8 FILLER_60_1608 ();
 sg13g2_decap_8 FILLER_60_1615 ();
 sg13g2_decap_8 FILLER_60_1622 ();
 sg13g2_decap_8 FILLER_60_1629 ();
 sg13g2_decap_8 FILLER_60_1636 ();
 sg13g2_decap_8 FILLER_60_1643 ();
 sg13g2_decap_8 FILLER_60_1650 ();
 sg13g2_decap_8 FILLER_60_1657 ();
 sg13g2_decap_8 FILLER_60_1664 ();
 sg13g2_decap_8 FILLER_60_1671 ();
 sg13g2_decap_8 FILLER_60_1678 ();
 sg13g2_decap_8 FILLER_60_1685 ();
 sg13g2_decap_8 FILLER_60_1692 ();
 sg13g2_decap_8 FILLER_60_1699 ();
 sg13g2_decap_8 FILLER_60_1706 ();
 sg13g2_decap_8 FILLER_60_1713 ();
 sg13g2_decap_8 FILLER_60_1720 ();
 sg13g2_decap_8 FILLER_60_1727 ();
 sg13g2_decap_8 FILLER_60_1734 ();
 sg13g2_decap_8 FILLER_60_1741 ();
 sg13g2_decap_8 FILLER_60_1748 ();
 sg13g2_decap_8 FILLER_60_1755 ();
 sg13g2_decap_4 FILLER_60_1762 ();
 sg13g2_fill_2 FILLER_60_1766 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_7 ();
 sg13g2_fill_1 FILLER_61_34 ();
 sg13g2_fill_2 FILLER_61_51 ();
 sg13g2_fill_2 FILLER_61_67 ();
 sg13g2_fill_2 FILLER_61_78 ();
 sg13g2_fill_1 FILLER_61_94 ();
 sg13g2_decap_8 FILLER_61_110 ();
 sg13g2_fill_2 FILLER_61_117 ();
 sg13g2_fill_2 FILLER_61_165 ();
 sg13g2_fill_2 FILLER_61_193 ();
 sg13g2_fill_1 FILLER_61_195 ();
 sg13g2_fill_2 FILLER_61_222 ();
 sg13g2_fill_1 FILLER_61_224 ();
 sg13g2_decap_4 FILLER_61_261 ();
 sg13g2_fill_1 FILLER_61_265 ();
 sg13g2_decap_4 FILLER_61_272 ();
 sg13g2_decap_4 FILLER_61_336 ();
 sg13g2_fill_1 FILLER_61_340 ();
 sg13g2_fill_1 FILLER_61_391 ();
 sg13g2_decap_4 FILLER_61_405 ();
 sg13g2_fill_1 FILLER_61_409 ();
 sg13g2_fill_1 FILLER_61_459 ();
 sg13g2_fill_1 FILLER_61_538 ();
 sg13g2_fill_1 FILLER_61_552 ();
 sg13g2_fill_2 FILLER_61_558 ();
 sg13g2_fill_1 FILLER_61_569 ();
 sg13g2_fill_1 FILLER_61_604 ();
 sg13g2_fill_2 FILLER_61_627 ();
 sg13g2_fill_1 FILLER_61_629 ();
 sg13g2_fill_2 FILLER_61_660 ();
 sg13g2_fill_1 FILLER_61_697 ();
 sg13g2_fill_1 FILLER_61_732 ();
 sg13g2_fill_2 FILLER_61_765 ();
 sg13g2_decap_4 FILLER_61_804 ();
 sg13g2_decap_8 FILLER_61_812 ();
 sg13g2_fill_1 FILLER_61_819 ();
 sg13g2_decap_4 FILLER_61_829 ();
 sg13g2_fill_1 FILLER_61_833 ();
 sg13g2_fill_2 FILLER_61_847 ();
 sg13g2_fill_1 FILLER_61_849 ();
 sg13g2_decap_8 FILLER_61_858 ();
 sg13g2_decap_4 FILLER_61_865 ();
 sg13g2_decap_8 FILLER_61_873 ();
 sg13g2_decap_8 FILLER_61_880 ();
 sg13g2_decap_4 FILLER_61_887 ();
 sg13g2_fill_1 FILLER_61_891 ();
 sg13g2_decap_8 FILLER_61_906 ();
 sg13g2_fill_1 FILLER_61_913 ();
 sg13g2_fill_2 FILLER_61_924 ();
 sg13g2_fill_1 FILLER_61_952 ();
 sg13g2_decap_8 FILLER_61_984 ();
 sg13g2_decap_8 FILLER_61_991 ();
 sg13g2_decap_8 FILLER_61_998 ();
 sg13g2_decap_8 FILLER_61_1005 ();
 sg13g2_decap_8 FILLER_61_1012 ();
 sg13g2_decap_8 FILLER_61_1019 ();
 sg13g2_decap_8 FILLER_61_1026 ();
 sg13g2_decap_8 FILLER_61_1033 ();
 sg13g2_decap_8 FILLER_61_1040 ();
 sg13g2_decap_8 FILLER_61_1047 ();
 sg13g2_decap_8 FILLER_61_1054 ();
 sg13g2_decap_8 FILLER_61_1061 ();
 sg13g2_decap_8 FILLER_61_1068 ();
 sg13g2_decap_8 FILLER_61_1075 ();
 sg13g2_decap_8 FILLER_61_1082 ();
 sg13g2_decap_8 FILLER_61_1089 ();
 sg13g2_decap_8 FILLER_61_1096 ();
 sg13g2_decap_8 FILLER_61_1103 ();
 sg13g2_decap_8 FILLER_61_1110 ();
 sg13g2_decap_8 FILLER_61_1117 ();
 sg13g2_decap_8 FILLER_61_1124 ();
 sg13g2_decap_8 FILLER_61_1131 ();
 sg13g2_decap_8 FILLER_61_1138 ();
 sg13g2_decap_8 FILLER_61_1145 ();
 sg13g2_decap_8 FILLER_61_1152 ();
 sg13g2_decap_8 FILLER_61_1159 ();
 sg13g2_decap_8 FILLER_61_1166 ();
 sg13g2_decap_8 FILLER_61_1173 ();
 sg13g2_decap_8 FILLER_61_1180 ();
 sg13g2_decap_8 FILLER_61_1187 ();
 sg13g2_decap_8 FILLER_61_1194 ();
 sg13g2_decap_8 FILLER_61_1201 ();
 sg13g2_decap_8 FILLER_61_1208 ();
 sg13g2_decap_8 FILLER_61_1215 ();
 sg13g2_decap_8 FILLER_61_1222 ();
 sg13g2_decap_8 FILLER_61_1229 ();
 sg13g2_decap_8 FILLER_61_1236 ();
 sg13g2_decap_8 FILLER_61_1243 ();
 sg13g2_decap_8 FILLER_61_1250 ();
 sg13g2_decap_8 FILLER_61_1257 ();
 sg13g2_decap_8 FILLER_61_1264 ();
 sg13g2_decap_8 FILLER_61_1271 ();
 sg13g2_decap_8 FILLER_61_1278 ();
 sg13g2_decap_8 FILLER_61_1285 ();
 sg13g2_decap_8 FILLER_61_1292 ();
 sg13g2_decap_8 FILLER_61_1299 ();
 sg13g2_decap_8 FILLER_61_1306 ();
 sg13g2_decap_8 FILLER_61_1313 ();
 sg13g2_decap_8 FILLER_61_1320 ();
 sg13g2_decap_8 FILLER_61_1327 ();
 sg13g2_decap_8 FILLER_61_1334 ();
 sg13g2_decap_8 FILLER_61_1341 ();
 sg13g2_decap_8 FILLER_61_1348 ();
 sg13g2_decap_8 FILLER_61_1355 ();
 sg13g2_decap_8 FILLER_61_1362 ();
 sg13g2_decap_8 FILLER_61_1369 ();
 sg13g2_decap_8 FILLER_61_1376 ();
 sg13g2_decap_8 FILLER_61_1383 ();
 sg13g2_decap_8 FILLER_61_1390 ();
 sg13g2_decap_8 FILLER_61_1397 ();
 sg13g2_decap_8 FILLER_61_1404 ();
 sg13g2_decap_8 FILLER_61_1411 ();
 sg13g2_decap_8 FILLER_61_1418 ();
 sg13g2_decap_8 FILLER_61_1425 ();
 sg13g2_decap_8 FILLER_61_1432 ();
 sg13g2_decap_8 FILLER_61_1439 ();
 sg13g2_decap_8 FILLER_61_1446 ();
 sg13g2_decap_8 FILLER_61_1453 ();
 sg13g2_decap_8 FILLER_61_1460 ();
 sg13g2_decap_8 FILLER_61_1467 ();
 sg13g2_decap_8 FILLER_61_1474 ();
 sg13g2_decap_8 FILLER_61_1481 ();
 sg13g2_decap_8 FILLER_61_1488 ();
 sg13g2_decap_8 FILLER_61_1495 ();
 sg13g2_decap_8 FILLER_61_1502 ();
 sg13g2_decap_8 FILLER_61_1509 ();
 sg13g2_decap_8 FILLER_61_1516 ();
 sg13g2_decap_8 FILLER_61_1523 ();
 sg13g2_decap_8 FILLER_61_1530 ();
 sg13g2_decap_8 FILLER_61_1537 ();
 sg13g2_decap_8 FILLER_61_1544 ();
 sg13g2_decap_8 FILLER_61_1551 ();
 sg13g2_decap_8 FILLER_61_1558 ();
 sg13g2_decap_8 FILLER_61_1565 ();
 sg13g2_decap_8 FILLER_61_1572 ();
 sg13g2_decap_8 FILLER_61_1579 ();
 sg13g2_decap_8 FILLER_61_1586 ();
 sg13g2_decap_8 FILLER_61_1593 ();
 sg13g2_decap_8 FILLER_61_1600 ();
 sg13g2_decap_8 FILLER_61_1607 ();
 sg13g2_decap_8 FILLER_61_1614 ();
 sg13g2_decap_8 FILLER_61_1621 ();
 sg13g2_decap_8 FILLER_61_1628 ();
 sg13g2_decap_8 FILLER_61_1635 ();
 sg13g2_decap_8 FILLER_61_1642 ();
 sg13g2_decap_8 FILLER_61_1649 ();
 sg13g2_decap_8 FILLER_61_1656 ();
 sg13g2_decap_8 FILLER_61_1663 ();
 sg13g2_decap_8 FILLER_61_1670 ();
 sg13g2_decap_8 FILLER_61_1677 ();
 sg13g2_decap_8 FILLER_61_1684 ();
 sg13g2_decap_8 FILLER_61_1691 ();
 sg13g2_decap_8 FILLER_61_1698 ();
 sg13g2_decap_8 FILLER_61_1705 ();
 sg13g2_decap_8 FILLER_61_1712 ();
 sg13g2_decap_8 FILLER_61_1719 ();
 sg13g2_decap_8 FILLER_61_1726 ();
 sg13g2_decap_8 FILLER_61_1733 ();
 sg13g2_decap_8 FILLER_61_1740 ();
 sg13g2_decap_8 FILLER_61_1747 ();
 sg13g2_decap_8 FILLER_61_1754 ();
 sg13g2_decap_8 FILLER_61_1761 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_7 ();
 sg13g2_fill_2 FILLER_62_53 ();
 sg13g2_decap_4 FILLER_62_121 ();
 sg13g2_fill_2 FILLER_62_200 ();
 sg13g2_fill_2 FILLER_62_215 ();
 sg13g2_fill_1 FILLER_62_239 ();
 sg13g2_decap_4 FILLER_62_256 ();
 sg13g2_fill_2 FILLER_62_260 ();
 sg13g2_fill_2 FILLER_62_279 ();
 sg13g2_fill_2 FILLER_62_295 ();
 sg13g2_fill_1 FILLER_62_315 ();
 sg13g2_fill_2 FILLER_62_342 ();
 sg13g2_fill_2 FILLER_62_352 ();
 sg13g2_fill_1 FILLER_62_354 ();
 sg13g2_fill_2 FILLER_62_425 ();
 sg13g2_decap_8 FILLER_62_488 ();
 sg13g2_decap_4 FILLER_62_495 ();
 sg13g2_fill_1 FILLER_62_544 ();
 sg13g2_fill_1 FILLER_62_555 ();
 sg13g2_fill_1 FILLER_62_567 ();
 sg13g2_fill_2 FILLER_62_633 ();
 sg13g2_fill_2 FILLER_62_676 ();
 sg13g2_fill_1 FILLER_62_678 ();
 sg13g2_fill_1 FILLER_62_692 ();
 sg13g2_fill_2 FILLER_62_727 ();
 sg13g2_fill_2 FILLER_62_734 ();
 sg13g2_fill_1 FILLER_62_736 ();
 sg13g2_fill_2 FILLER_62_746 ();
 sg13g2_fill_2 FILLER_62_761 ();
 sg13g2_fill_2 FILLER_62_849 ();
 sg13g2_fill_2 FILLER_62_890 ();
 sg13g2_fill_2 FILLER_62_928 ();
 sg13g2_fill_1 FILLER_62_930 ();
 sg13g2_fill_2 FILLER_62_944 ();
 sg13g2_fill_1 FILLER_62_946 ();
 sg13g2_decap_4 FILLER_62_963 ();
 sg13g2_fill_1 FILLER_62_967 ();
 sg13g2_fill_2 FILLER_62_972 ();
 sg13g2_fill_1 FILLER_62_974 ();
 sg13g2_decap_8 FILLER_62_979 ();
 sg13g2_decap_8 FILLER_62_986 ();
 sg13g2_decap_8 FILLER_62_993 ();
 sg13g2_decap_8 FILLER_62_1000 ();
 sg13g2_decap_8 FILLER_62_1007 ();
 sg13g2_decap_8 FILLER_62_1014 ();
 sg13g2_decap_8 FILLER_62_1021 ();
 sg13g2_decap_8 FILLER_62_1028 ();
 sg13g2_decap_8 FILLER_62_1035 ();
 sg13g2_decap_8 FILLER_62_1042 ();
 sg13g2_decap_8 FILLER_62_1049 ();
 sg13g2_decap_8 FILLER_62_1056 ();
 sg13g2_decap_8 FILLER_62_1063 ();
 sg13g2_decap_8 FILLER_62_1070 ();
 sg13g2_decap_8 FILLER_62_1077 ();
 sg13g2_decap_8 FILLER_62_1084 ();
 sg13g2_decap_8 FILLER_62_1091 ();
 sg13g2_decap_8 FILLER_62_1098 ();
 sg13g2_decap_8 FILLER_62_1105 ();
 sg13g2_decap_8 FILLER_62_1112 ();
 sg13g2_decap_8 FILLER_62_1119 ();
 sg13g2_decap_8 FILLER_62_1126 ();
 sg13g2_decap_8 FILLER_62_1133 ();
 sg13g2_decap_8 FILLER_62_1140 ();
 sg13g2_decap_8 FILLER_62_1147 ();
 sg13g2_decap_8 FILLER_62_1154 ();
 sg13g2_decap_8 FILLER_62_1161 ();
 sg13g2_decap_8 FILLER_62_1168 ();
 sg13g2_decap_8 FILLER_62_1175 ();
 sg13g2_decap_8 FILLER_62_1182 ();
 sg13g2_decap_8 FILLER_62_1189 ();
 sg13g2_decap_8 FILLER_62_1196 ();
 sg13g2_decap_8 FILLER_62_1203 ();
 sg13g2_decap_8 FILLER_62_1210 ();
 sg13g2_decap_8 FILLER_62_1217 ();
 sg13g2_decap_8 FILLER_62_1224 ();
 sg13g2_decap_8 FILLER_62_1231 ();
 sg13g2_decap_8 FILLER_62_1238 ();
 sg13g2_decap_8 FILLER_62_1245 ();
 sg13g2_decap_8 FILLER_62_1252 ();
 sg13g2_decap_8 FILLER_62_1259 ();
 sg13g2_decap_8 FILLER_62_1266 ();
 sg13g2_decap_8 FILLER_62_1273 ();
 sg13g2_decap_8 FILLER_62_1280 ();
 sg13g2_decap_8 FILLER_62_1287 ();
 sg13g2_decap_8 FILLER_62_1294 ();
 sg13g2_decap_8 FILLER_62_1301 ();
 sg13g2_decap_8 FILLER_62_1308 ();
 sg13g2_decap_8 FILLER_62_1315 ();
 sg13g2_decap_8 FILLER_62_1322 ();
 sg13g2_decap_8 FILLER_62_1329 ();
 sg13g2_decap_8 FILLER_62_1336 ();
 sg13g2_decap_8 FILLER_62_1343 ();
 sg13g2_decap_8 FILLER_62_1350 ();
 sg13g2_decap_8 FILLER_62_1357 ();
 sg13g2_decap_8 FILLER_62_1364 ();
 sg13g2_decap_8 FILLER_62_1371 ();
 sg13g2_decap_8 FILLER_62_1378 ();
 sg13g2_decap_8 FILLER_62_1385 ();
 sg13g2_decap_8 FILLER_62_1392 ();
 sg13g2_decap_8 FILLER_62_1399 ();
 sg13g2_decap_8 FILLER_62_1406 ();
 sg13g2_decap_8 FILLER_62_1413 ();
 sg13g2_decap_8 FILLER_62_1420 ();
 sg13g2_decap_8 FILLER_62_1427 ();
 sg13g2_decap_8 FILLER_62_1434 ();
 sg13g2_decap_8 FILLER_62_1441 ();
 sg13g2_decap_8 FILLER_62_1448 ();
 sg13g2_decap_8 FILLER_62_1455 ();
 sg13g2_decap_8 FILLER_62_1462 ();
 sg13g2_decap_8 FILLER_62_1469 ();
 sg13g2_decap_8 FILLER_62_1476 ();
 sg13g2_decap_8 FILLER_62_1483 ();
 sg13g2_decap_8 FILLER_62_1490 ();
 sg13g2_decap_8 FILLER_62_1497 ();
 sg13g2_decap_8 FILLER_62_1504 ();
 sg13g2_decap_8 FILLER_62_1511 ();
 sg13g2_decap_8 FILLER_62_1518 ();
 sg13g2_decap_8 FILLER_62_1525 ();
 sg13g2_decap_8 FILLER_62_1532 ();
 sg13g2_decap_8 FILLER_62_1539 ();
 sg13g2_decap_8 FILLER_62_1546 ();
 sg13g2_decap_8 FILLER_62_1553 ();
 sg13g2_decap_8 FILLER_62_1560 ();
 sg13g2_decap_8 FILLER_62_1567 ();
 sg13g2_decap_8 FILLER_62_1574 ();
 sg13g2_decap_8 FILLER_62_1581 ();
 sg13g2_decap_8 FILLER_62_1588 ();
 sg13g2_decap_8 FILLER_62_1595 ();
 sg13g2_decap_8 FILLER_62_1602 ();
 sg13g2_decap_8 FILLER_62_1609 ();
 sg13g2_decap_8 FILLER_62_1616 ();
 sg13g2_decap_8 FILLER_62_1623 ();
 sg13g2_decap_8 FILLER_62_1630 ();
 sg13g2_decap_8 FILLER_62_1637 ();
 sg13g2_decap_8 FILLER_62_1644 ();
 sg13g2_decap_8 FILLER_62_1651 ();
 sg13g2_decap_8 FILLER_62_1658 ();
 sg13g2_decap_8 FILLER_62_1665 ();
 sg13g2_decap_8 FILLER_62_1672 ();
 sg13g2_decap_8 FILLER_62_1679 ();
 sg13g2_decap_8 FILLER_62_1686 ();
 sg13g2_decap_8 FILLER_62_1693 ();
 sg13g2_decap_8 FILLER_62_1700 ();
 sg13g2_decap_8 FILLER_62_1707 ();
 sg13g2_decap_8 FILLER_62_1714 ();
 sg13g2_decap_8 FILLER_62_1721 ();
 sg13g2_decap_8 FILLER_62_1728 ();
 sg13g2_decap_8 FILLER_62_1735 ();
 sg13g2_decap_8 FILLER_62_1742 ();
 sg13g2_decap_8 FILLER_62_1749 ();
 sg13g2_decap_8 FILLER_62_1756 ();
 sg13g2_decap_4 FILLER_62_1763 ();
 sg13g2_fill_1 FILLER_62_1767 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_4 FILLER_63_14 ();
 sg13g2_fill_1 FILLER_63_18 ();
 sg13g2_decap_8 FILLER_63_23 ();
 sg13g2_fill_2 FILLER_63_101 ();
 sg13g2_fill_1 FILLER_63_103 ();
 sg13g2_decap_8 FILLER_63_117 ();
 sg13g2_fill_2 FILLER_63_154 ();
 sg13g2_fill_1 FILLER_63_156 ();
 sg13g2_decap_8 FILLER_63_170 ();
 sg13g2_fill_1 FILLER_63_177 ();
 sg13g2_decap_8 FILLER_63_182 ();
 sg13g2_fill_2 FILLER_63_189 ();
 sg13g2_fill_1 FILLER_63_191 ();
 sg13g2_decap_4 FILLER_63_254 ();
 sg13g2_fill_1 FILLER_63_258 ();
 sg13g2_fill_2 FILLER_63_263 ();
 sg13g2_decap_4 FILLER_63_271 ();
 sg13g2_fill_1 FILLER_63_286 ();
 sg13g2_fill_1 FILLER_63_305 ();
 sg13g2_fill_2 FILLER_63_360 ();
 sg13g2_fill_1 FILLER_63_376 ();
 sg13g2_fill_2 FILLER_63_390 ();
 sg13g2_fill_1 FILLER_63_392 ();
 sg13g2_fill_1 FILLER_63_402 ();
 sg13g2_fill_2 FILLER_63_412 ();
 sg13g2_fill_1 FILLER_63_460 ();
 sg13g2_fill_1 FILLER_63_475 ();
 sg13g2_fill_2 FILLER_63_549 ();
 sg13g2_fill_2 FILLER_63_576 ();
 sg13g2_fill_2 FILLER_63_598 ();
 sg13g2_fill_1 FILLER_63_600 ();
 sg13g2_fill_2 FILLER_63_606 ();
 sg13g2_fill_1 FILLER_63_608 ();
 sg13g2_fill_2 FILLER_63_629 ();
 sg13g2_fill_1 FILLER_63_631 ();
 sg13g2_fill_2 FILLER_63_677 ();
 sg13g2_fill_1 FILLER_63_679 ();
 sg13g2_fill_1 FILLER_63_728 ();
 sg13g2_fill_2 FILLER_63_749 ();
 sg13g2_fill_1 FILLER_63_751 ();
 sg13g2_fill_2 FILLER_63_761 ();
 sg13g2_decap_8 FILLER_63_767 ();
 sg13g2_fill_2 FILLER_63_788 ();
 sg13g2_decap_4 FILLER_63_803 ();
 sg13g2_fill_2 FILLER_63_807 ();
 sg13g2_decap_8 FILLER_63_814 ();
 sg13g2_fill_2 FILLER_63_821 ();
 sg13g2_fill_1 FILLER_63_842 ();
 sg13g2_fill_1 FILLER_63_851 ();
 sg13g2_fill_2 FILLER_63_858 ();
 sg13g2_decap_8 FILLER_63_895 ();
 sg13g2_decap_4 FILLER_63_902 ();
 sg13g2_fill_1 FILLER_63_906 ();
 sg13g2_fill_1 FILLER_63_956 ();
 sg13g2_fill_2 FILLER_63_961 ();
 sg13g2_fill_1 FILLER_63_963 ();
 sg13g2_decap_8 FILLER_63_990 ();
 sg13g2_decap_8 FILLER_63_997 ();
 sg13g2_decap_8 FILLER_63_1004 ();
 sg13g2_decap_8 FILLER_63_1011 ();
 sg13g2_decap_8 FILLER_63_1018 ();
 sg13g2_decap_8 FILLER_63_1025 ();
 sg13g2_decap_8 FILLER_63_1032 ();
 sg13g2_decap_8 FILLER_63_1039 ();
 sg13g2_decap_8 FILLER_63_1046 ();
 sg13g2_decap_8 FILLER_63_1053 ();
 sg13g2_decap_8 FILLER_63_1060 ();
 sg13g2_decap_8 FILLER_63_1067 ();
 sg13g2_decap_8 FILLER_63_1074 ();
 sg13g2_decap_8 FILLER_63_1081 ();
 sg13g2_decap_8 FILLER_63_1088 ();
 sg13g2_decap_8 FILLER_63_1095 ();
 sg13g2_decap_8 FILLER_63_1102 ();
 sg13g2_decap_8 FILLER_63_1109 ();
 sg13g2_decap_8 FILLER_63_1116 ();
 sg13g2_decap_8 FILLER_63_1123 ();
 sg13g2_decap_8 FILLER_63_1130 ();
 sg13g2_decap_8 FILLER_63_1137 ();
 sg13g2_decap_8 FILLER_63_1144 ();
 sg13g2_decap_8 FILLER_63_1151 ();
 sg13g2_decap_8 FILLER_63_1158 ();
 sg13g2_decap_8 FILLER_63_1165 ();
 sg13g2_decap_8 FILLER_63_1172 ();
 sg13g2_decap_8 FILLER_63_1179 ();
 sg13g2_decap_8 FILLER_63_1186 ();
 sg13g2_decap_8 FILLER_63_1193 ();
 sg13g2_decap_8 FILLER_63_1200 ();
 sg13g2_decap_8 FILLER_63_1207 ();
 sg13g2_decap_8 FILLER_63_1214 ();
 sg13g2_decap_8 FILLER_63_1221 ();
 sg13g2_decap_8 FILLER_63_1228 ();
 sg13g2_decap_8 FILLER_63_1235 ();
 sg13g2_decap_8 FILLER_63_1242 ();
 sg13g2_decap_8 FILLER_63_1249 ();
 sg13g2_decap_8 FILLER_63_1256 ();
 sg13g2_decap_8 FILLER_63_1263 ();
 sg13g2_decap_8 FILLER_63_1270 ();
 sg13g2_decap_8 FILLER_63_1277 ();
 sg13g2_decap_8 FILLER_63_1284 ();
 sg13g2_decap_8 FILLER_63_1291 ();
 sg13g2_decap_8 FILLER_63_1298 ();
 sg13g2_decap_8 FILLER_63_1305 ();
 sg13g2_decap_8 FILLER_63_1312 ();
 sg13g2_decap_8 FILLER_63_1319 ();
 sg13g2_decap_8 FILLER_63_1326 ();
 sg13g2_decap_8 FILLER_63_1333 ();
 sg13g2_decap_8 FILLER_63_1340 ();
 sg13g2_decap_8 FILLER_63_1347 ();
 sg13g2_decap_8 FILLER_63_1354 ();
 sg13g2_decap_8 FILLER_63_1361 ();
 sg13g2_decap_8 FILLER_63_1368 ();
 sg13g2_decap_8 FILLER_63_1375 ();
 sg13g2_decap_8 FILLER_63_1382 ();
 sg13g2_decap_8 FILLER_63_1389 ();
 sg13g2_decap_8 FILLER_63_1396 ();
 sg13g2_decap_8 FILLER_63_1403 ();
 sg13g2_decap_8 FILLER_63_1410 ();
 sg13g2_decap_8 FILLER_63_1417 ();
 sg13g2_decap_8 FILLER_63_1424 ();
 sg13g2_decap_8 FILLER_63_1431 ();
 sg13g2_decap_8 FILLER_63_1438 ();
 sg13g2_decap_8 FILLER_63_1445 ();
 sg13g2_decap_8 FILLER_63_1452 ();
 sg13g2_decap_8 FILLER_63_1459 ();
 sg13g2_decap_8 FILLER_63_1466 ();
 sg13g2_decap_8 FILLER_63_1473 ();
 sg13g2_decap_8 FILLER_63_1480 ();
 sg13g2_decap_8 FILLER_63_1487 ();
 sg13g2_decap_8 FILLER_63_1494 ();
 sg13g2_decap_8 FILLER_63_1501 ();
 sg13g2_decap_8 FILLER_63_1508 ();
 sg13g2_decap_8 FILLER_63_1515 ();
 sg13g2_decap_8 FILLER_63_1522 ();
 sg13g2_decap_8 FILLER_63_1529 ();
 sg13g2_decap_8 FILLER_63_1536 ();
 sg13g2_decap_8 FILLER_63_1543 ();
 sg13g2_decap_8 FILLER_63_1550 ();
 sg13g2_decap_8 FILLER_63_1557 ();
 sg13g2_decap_8 FILLER_63_1564 ();
 sg13g2_decap_8 FILLER_63_1571 ();
 sg13g2_decap_8 FILLER_63_1578 ();
 sg13g2_decap_8 FILLER_63_1585 ();
 sg13g2_decap_8 FILLER_63_1592 ();
 sg13g2_decap_8 FILLER_63_1599 ();
 sg13g2_decap_8 FILLER_63_1606 ();
 sg13g2_decap_8 FILLER_63_1613 ();
 sg13g2_decap_8 FILLER_63_1620 ();
 sg13g2_decap_8 FILLER_63_1627 ();
 sg13g2_decap_8 FILLER_63_1634 ();
 sg13g2_decap_8 FILLER_63_1641 ();
 sg13g2_decap_8 FILLER_63_1648 ();
 sg13g2_decap_8 FILLER_63_1655 ();
 sg13g2_decap_8 FILLER_63_1662 ();
 sg13g2_decap_8 FILLER_63_1669 ();
 sg13g2_decap_8 FILLER_63_1676 ();
 sg13g2_decap_8 FILLER_63_1683 ();
 sg13g2_decap_8 FILLER_63_1690 ();
 sg13g2_decap_8 FILLER_63_1697 ();
 sg13g2_decap_8 FILLER_63_1704 ();
 sg13g2_decap_8 FILLER_63_1711 ();
 sg13g2_decap_8 FILLER_63_1718 ();
 sg13g2_decap_8 FILLER_63_1725 ();
 sg13g2_decap_8 FILLER_63_1732 ();
 sg13g2_decap_8 FILLER_63_1739 ();
 sg13g2_decap_8 FILLER_63_1746 ();
 sg13g2_decap_8 FILLER_63_1753 ();
 sg13g2_decap_8 FILLER_63_1760 ();
 sg13g2_fill_1 FILLER_63_1767 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_fill_2 FILLER_64_42 ();
 sg13g2_fill_1 FILLER_64_44 ();
 sg13g2_fill_2 FILLER_64_53 ();
 sg13g2_decap_4 FILLER_64_81 ();
 sg13g2_fill_1 FILLER_64_85 ();
 sg13g2_fill_2 FILLER_64_96 ();
 sg13g2_fill_1 FILLER_64_98 ();
 sg13g2_fill_1 FILLER_64_179 ();
 sg13g2_fill_1 FILLER_64_192 ();
 sg13g2_fill_1 FILLER_64_246 ();
 sg13g2_fill_2 FILLER_64_318 ();
 sg13g2_fill_2 FILLER_64_338 ();
 sg13g2_fill_2 FILLER_64_346 ();
 sg13g2_fill_2 FILLER_64_396 ();
 sg13g2_fill_1 FILLER_64_438 ();
 sg13g2_fill_1 FILLER_64_470 ();
 sg13g2_fill_2 FILLER_64_516 ();
 sg13g2_fill_2 FILLER_64_528 ();
 sg13g2_fill_1 FILLER_64_530 ();
 sg13g2_fill_2 FILLER_64_560 ();
 sg13g2_fill_1 FILLER_64_562 ();
 sg13g2_decap_4 FILLER_64_581 ();
 sg13g2_fill_2 FILLER_64_596 ();
 sg13g2_fill_1 FILLER_64_613 ();
 sg13g2_fill_1 FILLER_64_627 ();
 sg13g2_fill_1 FILLER_64_657 ();
 sg13g2_fill_1 FILLER_64_708 ();
 sg13g2_fill_1 FILLER_64_713 ();
 sg13g2_fill_1 FILLER_64_805 ();
 sg13g2_fill_2 FILLER_64_842 ();
 sg13g2_decap_4 FILLER_64_871 ();
 sg13g2_fill_1 FILLER_64_875 ();
 sg13g2_fill_1 FILLER_64_889 ();
 sg13g2_decap_8 FILLER_64_906 ();
 sg13g2_decap_8 FILLER_64_921 ();
 sg13g2_fill_2 FILLER_64_928 ();
 sg13g2_fill_1 FILLER_64_930 ();
 sg13g2_decap_8 FILLER_64_993 ();
 sg13g2_decap_8 FILLER_64_1000 ();
 sg13g2_decap_8 FILLER_64_1007 ();
 sg13g2_decap_8 FILLER_64_1014 ();
 sg13g2_decap_8 FILLER_64_1021 ();
 sg13g2_decap_8 FILLER_64_1028 ();
 sg13g2_decap_8 FILLER_64_1035 ();
 sg13g2_decap_8 FILLER_64_1042 ();
 sg13g2_decap_8 FILLER_64_1049 ();
 sg13g2_decap_8 FILLER_64_1056 ();
 sg13g2_decap_8 FILLER_64_1063 ();
 sg13g2_decap_8 FILLER_64_1070 ();
 sg13g2_decap_8 FILLER_64_1077 ();
 sg13g2_decap_8 FILLER_64_1084 ();
 sg13g2_decap_8 FILLER_64_1091 ();
 sg13g2_decap_8 FILLER_64_1098 ();
 sg13g2_decap_8 FILLER_64_1105 ();
 sg13g2_decap_8 FILLER_64_1112 ();
 sg13g2_decap_8 FILLER_64_1119 ();
 sg13g2_decap_8 FILLER_64_1126 ();
 sg13g2_decap_8 FILLER_64_1133 ();
 sg13g2_decap_8 FILLER_64_1140 ();
 sg13g2_decap_8 FILLER_64_1147 ();
 sg13g2_decap_8 FILLER_64_1154 ();
 sg13g2_decap_8 FILLER_64_1161 ();
 sg13g2_decap_8 FILLER_64_1168 ();
 sg13g2_decap_8 FILLER_64_1175 ();
 sg13g2_decap_8 FILLER_64_1182 ();
 sg13g2_decap_8 FILLER_64_1189 ();
 sg13g2_decap_8 FILLER_64_1196 ();
 sg13g2_decap_8 FILLER_64_1203 ();
 sg13g2_decap_8 FILLER_64_1210 ();
 sg13g2_decap_8 FILLER_64_1217 ();
 sg13g2_decap_8 FILLER_64_1224 ();
 sg13g2_decap_8 FILLER_64_1231 ();
 sg13g2_decap_8 FILLER_64_1238 ();
 sg13g2_decap_8 FILLER_64_1245 ();
 sg13g2_decap_8 FILLER_64_1252 ();
 sg13g2_decap_8 FILLER_64_1259 ();
 sg13g2_decap_8 FILLER_64_1266 ();
 sg13g2_decap_8 FILLER_64_1273 ();
 sg13g2_decap_8 FILLER_64_1280 ();
 sg13g2_decap_8 FILLER_64_1287 ();
 sg13g2_decap_8 FILLER_64_1294 ();
 sg13g2_decap_8 FILLER_64_1301 ();
 sg13g2_decap_8 FILLER_64_1308 ();
 sg13g2_decap_8 FILLER_64_1315 ();
 sg13g2_decap_8 FILLER_64_1322 ();
 sg13g2_decap_8 FILLER_64_1329 ();
 sg13g2_decap_8 FILLER_64_1336 ();
 sg13g2_decap_8 FILLER_64_1343 ();
 sg13g2_decap_8 FILLER_64_1350 ();
 sg13g2_decap_8 FILLER_64_1357 ();
 sg13g2_decap_8 FILLER_64_1364 ();
 sg13g2_decap_8 FILLER_64_1371 ();
 sg13g2_decap_8 FILLER_64_1378 ();
 sg13g2_decap_8 FILLER_64_1385 ();
 sg13g2_decap_8 FILLER_64_1392 ();
 sg13g2_decap_8 FILLER_64_1399 ();
 sg13g2_decap_8 FILLER_64_1406 ();
 sg13g2_decap_8 FILLER_64_1413 ();
 sg13g2_decap_8 FILLER_64_1420 ();
 sg13g2_decap_8 FILLER_64_1427 ();
 sg13g2_decap_8 FILLER_64_1434 ();
 sg13g2_decap_8 FILLER_64_1441 ();
 sg13g2_decap_8 FILLER_64_1448 ();
 sg13g2_decap_8 FILLER_64_1455 ();
 sg13g2_decap_8 FILLER_64_1462 ();
 sg13g2_decap_8 FILLER_64_1469 ();
 sg13g2_decap_8 FILLER_64_1476 ();
 sg13g2_decap_8 FILLER_64_1483 ();
 sg13g2_decap_8 FILLER_64_1490 ();
 sg13g2_decap_8 FILLER_64_1497 ();
 sg13g2_decap_8 FILLER_64_1504 ();
 sg13g2_decap_8 FILLER_64_1511 ();
 sg13g2_decap_8 FILLER_64_1518 ();
 sg13g2_decap_8 FILLER_64_1525 ();
 sg13g2_decap_8 FILLER_64_1532 ();
 sg13g2_decap_8 FILLER_64_1539 ();
 sg13g2_decap_8 FILLER_64_1546 ();
 sg13g2_decap_8 FILLER_64_1553 ();
 sg13g2_decap_8 FILLER_64_1560 ();
 sg13g2_decap_8 FILLER_64_1567 ();
 sg13g2_decap_8 FILLER_64_1574 ();
 sg13g2_decap_8 FILLER_64_1581 ();
 sg13g2_decap_8 FILLER_64_1588 ();
 sg13g2_decap_8 FILLER_64_1595 ();
 sg13g2_decap_8 FILLER_64_1602 ();
 sg13g2_decap_8 FILLER_64_1609 ();
 sg13g2_decap_8 FILLER_64_1616 ();
 sg13g2_decap_8 FILLER_64_1623 ();
 sg13g2_decap_8 FILLER_64_1630 ();
 sg13g2_decap_8 FILLER_64_1637 ();
 sg13g2_decap_8 FILLER_64_1644 ();
 sg13g2_decap_8 FILLER_64_1651 ();
 sg13g2_decap_8 FILLER_64_1658 ();
 sg13g2_decap_8 FILLER_64_1665 ();
 sg13g2_decap_8 FILLER_64_1672 ();
 sg13g2_decap_8 FILLER_64_1679 ();
 sg13g2_decap_8 FILLER_64_1686 ();
 sg13g2_decap_8 FILLER_64_1693 ();
 sg13g2_decap_8 FILLER_64_1700 ();
 sg13g2_decap_8 FILLER_64_1707 ();
 sg13g2_decap_8 FILLER_64_1714 ();
 sg13g2_decap_8 FILLER_64_1721 ();
 sg13g2_decap_8 FILLER_64_1728 ();
 sg13g2_decap_8 FILLER_64_1735 ();
 sg13g2_decap_8 FILLER_64_1742 ();
 sg13g2_decap_8 FILLER_64_1749 ();
 sg13g2_decap_8 FILLER_64_1756 ();
 sg13g2_decap_4 FILLER_64_1763 ();
 sg13g2_fill_1 FILLER_64_1767 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_116 ();
 sg13g2_decap_8 FILLER_65_123 ();
 sg13g2_fill_1 FILLER_65_130 ();
 sg13g2_fill_1 FILLER_65_157 ();
 sg13g2_fill_1 FILLER_65_184 ();
 sg13g2_fill_1 FILLER_65_241 ();
 sg13g2_fill_1 FILLER_65_252 ();
 sg13g2_decap_4 FILLER_65_262 ();
 sg13g2_fill_2 FILLER_65_275 ();
 sg13g2_fill_2 FILLER_65_282 ();
 sg13g2_decap_8 FILLER_65_288 ();
 sg13g2_decap_4 FILLER_65_295 ();
 sg13g2_fill_1 FILLER_65_355 ();
 sg13g2_fill_1 FILLER_65_367 ();
 sg13g2_fill_2 FILLER_65_399 ();
 sg13g2_decap_8 FILLER_65_405 ();
 sg13g2_fill_1 FILLER_65_412 ();
 sg13g2_fill_1 FILLER_65_417 ();
 sg13g2_decap_4 FILLER_65_425 ();
 sg13g2_fill_2 FILLER_65_429 ();
 sg13g2_fill_2 FILLER_65_474 ();
 sg13g2_fill_2 FILLER_65_506 ();
 sg13g2_fill_2 FILLER_65_525 ();
 sg13g2_fill_1 FILLER_65_527 ();
 sg13g2_fill_1 FILLER_65_533 ();
 sg13g2_fill_2 FILLER_65_543 ();
 sg13g2_fill_2 FILLER_65_599 ();
 sg13g2_fill_1 FILLER_65_601 ();
 sg13g2_fill_2 FILLER_65_607 ();
 sg13g2_fill_1 FILLER_65_629 ();
 sg13g2_decap_8 FILLER_65_662 ();
 sg13g2_decap_4 FILLER_65_669 ();
 sg13g2_fill_1 FILLER_65_673 ();
 sg13g2_fill_1 FILLER_65_695 ();
 sg13g2_fill_1 FILLER_65_710 ();
 sg13g2_decap_4 FILLER_65_726 ();
 sg13g2_fill_2 FILLER_65_730 ();
 sg13g2_decap_8 FILLER_65_744 ();
 sg13g2_fill_2 FILLER_65_751 ();
 sg13g2_decap_4 FILLER_65_762 ();
 sg13g2_fill_1 FILLER_65_766 ();
 sg13g2_decap_8 FILLER_65_772 ();
 sg13g2_decap_8 FILLER_65_779 ();
 sg13g2_fill_2 FILLER_65_786 ();
 sg13g2_fill_1 FILLER_65_788 ();
 sg13g2_fill_1 FILLER_65_792 ();
 sg13g2_decap_4 FILLER_65_811 ();
 sg13g2_fill_2 FILLER_65_841 ();
 sg13g2_fill_1 FILLER_65_843 ();
 sg13g2_fill_1 FILLER_65_850 ();
 sg13g2_fill_2 FILLER_65_863 ();
 sg13g2_fill_1 FILLER_65_875 ();
 sg13g2_fill_2 FILLER_65_895 ();
 sg13g2_fill_1 FILLER_65_897 ();
 sg13g2_fill_1 FILLER_65_922 ();
 sg13g2_fill_2 FILLER_65_949 ();
 sg13g2_decap_4 FILLER_65_956 ();
 sg13g2_fill_2 FILLER_65_960 ();
 sg13g2_decap_8 FILLER_65_975 ();
 sg13g2_fill_1 FILLER_65_982 ();
 sg13g2_decap_8 FILLER_65_1003 ();
 sg13g2_decap_8 FILLER_65_1010 ();
 sg13g2_decap_8 FILLER_65_1017 ();
 sg13g2_decap_8 FILLER_65_1024 ();
 sg13g2_decap_8 FILLER_65_1031 ();
 sg13g2_decap_8 FILLER_65_1038 ();
 sg13g2_decap_8 FILLER_65_1045 ();
 sg13g2_decap_8 FILLER_65_1052 ();
 sg13g2_decap_8 FILLER_65_1059 ();
 sg13g2_decap_8 FILLER_65_1066 ();
 sg13g2_decap_8 FILLER_65_1073 ();
 sg13g2_decap_8 FILLER_65_1080 ();
 sg13g2_decap_8 FILLER_65_1087 ();
 sg13g2_decap_8 FILLER_65_1094 ();
 sg13g2_decap_8 FILLER_65_1101 ();
 sg13g2_decap_8 FILLER_65_1108 ();
 sg13g2_decap_8 FILLER_65_1115 ();
 sg13g2_decap_8 FILLER_65_1122 ();
 sg13g2_decap_8 FILLER_65_1129 ();
 sg13g2_decap_8 FILLER_65_1136 ();
 sg13g2_decap_8 FILLER_65_1143 ();
 sg13g2_decap_8 FILLER_65_1150 ();
 sg13g2_decap_8 FILLER_65_1157 ();
 sg13g2_decap_8 FILLER_65_1164 ();
 sg13g2_decap_8 FILLER_65_1171 ();
 sg13g2_decap_8 FILLER_65_1178 ();
 sg13g2_decap_8 FILLER_65_1185 ();
 sg13g2_decap_8 FILLER_65_1192 ();
 sg13g2_decap_8 FILLER_65_1199 ();
 sg13g2_decap_8 FILLER_65_1206 ();
 sg13g2_decap_8 FILLER_65_1213 ();
 sg13g2_decap_8 FILLER_65_1220 ();
 sg13g2_decap_8 FILLER_65_1227 ();
 sg13g2_decap_8 FILLER_65_1234 ();
 sg13g2_decap_8 FILLER_65_1241 ();
 sg13g2_decap_8 FILLER_65_1248 ();
 sg13g2_decap_8 FILLER_65_1255 ();
 sg13g2_decap_8 FILLER_65_1262 ();
 sg13g2_decap_8 FILLER_65_1269 ();
 sg13g2_decap_8 FILLER_65_1276 ();
 sg13g2_decap_8 FILLER_65_1283 ();
 sg13g2_decap_8 FILLER_65_1290 ();
 sg13g2_decap_8 FILLER_65_1297 ();
 sg13g2_decap_8 FILLER_65_1304 ();
 sg13g2_decap_8 FILLER_65_1311 ();
 sg13g2_decap_8 FILLER_65_1318 ();
 sg13g2_decap_8 FILLER_65_1325 ();
 sg13g2_decap_8 FILLER_65_1332 ();
 sg13g2_decap_8 FILLER_65_1339 ();
 sg13g2_decap_8 FILLER_65_1346 ();
 sg13g2_decap_8 FILLER_65_1353 ();
 sg13g2_decap_8 FILLER_65_1360 ();
 sg13g2_decap_8 FILLER_65_1367 ();
 sg13g2_decap_8 FILLER_65_1374 ();
 sg13g2_decap_8 FILLER_65_1381 ();
 sg13g2_decap_8 FILLER_65_1388 ();
 sg13g2_decap_8 FILLER_65_1395 ();
 sg13g2_decap_8 FILLER_65_1402 ();
 sg13g2_decap_8 FILLER_65_1409 ();
 sg13g2_decap_8 FILLER_65_1416 ();
 sg13g2_decap_8 FILLER_65_1423 ();
 sg13g2_decap_8 FILLER_65_1430 ();
 sg13g2_decap_8 FILLER_65_1437 ();
 sg13g2_decap_8 FILLER_65_1444 ();
 sg13g2_decap_8 FILLER_65_1451 ();
 sg13g2_decap_8 FILLER_65_1458 ();
 sg13g2_decap_8 FILLER_65_1465 ();
 sg13g2_decap_8 FILLER_65_1472 ();
 sg13g2_decap_8 FILLER_65_1479 ();
 sg13g2_decap_8 FILLER_65_1486 ();
 sg13g2_decap_8 FILLER_65_1493 ();
 sg13g2_decap_8 FILLER_65_1500 ();
 sg13g2_decap_8 FILLER_65_1507 ();
 sg13g2_decap_8 FILLER_65_1514 ();
 sg13g2_decap_8 FILLER_65_1521 ();
 sg13g2_decap_8 FILLER_65_1528 ();
 sg13g2_decap_8 FILLER_65_1535 ();
 sg13g2_decap_8 FILLER_65_1542 ();
 sg13g2_decap_8 FILLER_65_1549 ();
 sg13g2_decap_8 FILLER_65_1556 ();
 sg13g2_decap_8 FILLER_65_1563 ();
 sg13g2_decap_8 FILLER_65_1570 ();
 sg13g2_decap_8 FILLER_65_1577 ();
 sg13g2_decap_8 FILLER_65_1584 ();
 sg13g2_decap_8 FILLER_65_1591 ();
 sg13g2_decap_8 FILLER_65_1598 ();
 sg13g2_decap_8 FILLER_65_1605 ();
 sg13g2_decap_8 FILLER_65_1612 ();
 sg13g2_decap_8 FILLER_65_1619 ();
 sg13g2_decap_8 FILLER_65_1626 ();
 sg13g2_decap_8 FILLER_65_1633 ();
 sg13g2_decap_8 FILLER_65_1640 ();
 sg13g2_decap_8 FILLER_65_1647 ();
 sg13g2_decap_8 FILLER_65_1654 ();
 sg13g2_decap_8 FILLER_65_1661 ();
 sg13g2_decap_8 FILLER_65_1668 ();
 sg13g2_decap_8 FILLER_65_1675 ();
 sg13g2_decap_8 FILLER_65_1682 ();
 sg13g2_decap_8 FILLER_65_1689 ();
 sg13g2_decap_8 FILLER_65_1696 ();
 sg13g2_decap_8 FILLER_65_1703 ();
 sg13g2_decap_8 FILLER_65_1710 ();
 sg13g2_decap_8 FILLER_65_1717 ();
 sg13g2_decap_8 FILLER_65_1724 ();
 sg13g2_decap_8 FILLER_65_1731 ();
 sg13g2_decap_8 FILLER_65_1738 ();
 sg13g2_decap_8 FILLER_65_1745 ();
 sg13g2_decap_8 FILLER_65_1752 ();
 sg13g2_decap_8 FILLER_65_1759 ();
 sg13g2_fill_2 FILLER_65_1766 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_fill_2 FILLER_66_84 ();
 sg13g2_fill_1 FILLER_66_86 ();
 sg13g2_decap_4 FILLER_66_91 ();
 sg13g2_fill_2 FILLER_66_95 ();
 sg13g2_fill_2 FILLER_66_102 ();
 sg13g2_decap_8 FILLER_66_113 ();
 sg13g2_decap_8 FILLER_66_120 ();
 sg13g2_decap_8 FILLER_66_127 ();
 sg13g2_fill_2 FILLER_66_134 ();
 sg13g2_fill_1 FILLER_66_136 ();
 sg13g2_fill_1 FILLER_66_141 ();
 sg13g2_fill_2 FILLER_66_146 ();
 sg13g2_fill_1 FILLER_66_148 ();
 sg13g2_fill_2 FILLER_66_163 ();
 sg13g2_decap_4 FILLER_66_168 ();
 sg13g2_fill_2 FILLER_66_172 ();
 sg13g2_fill_2 FILLER_66_183 ();
 sg13g2_fill_1 FILLER_66_185 ();
 sg13g2_decap_4 FILLER_66_190 ();
 sg13g2_fill_2 FILLER_66_204 ();
 sg13g2_decap_4 FILLER_66_211 ();
 sg13g2_fill_2 FILLER_66_215 ();
 sg13g2_fill_2 FILLER_66_235 ();
 sg13g2_fill_1 FILLER_66_237 ();
 sg13g2_fill_2 FILLER_66_243 ();
 sg13g2_fill_1 FILLER_66_245 ();
 sg13g2_decap_8 FILLER_66_259 ();
 sg13g2_fill_2 FILLER_66_266 ();
 sg13g2_fill_1 FILLER_66_268 ();
 sg13g2_fill_2 FILLER_66_287 ();
 sg13g2_decap_8 FILLER_66_294 ();
 sg13g2_fill_2 FILLER_66_306 ();
 sg13g2_fill_1 FILLER_66_313 ();
 sg13g2_fill_1 FILLER_66_328 ();
 sg13g2_fill_1 FILLER_66_351 ();
 sg13g2_fill_1 FILLER_66_367 ();
 sg13g2_fill_2 FILLER_66_395 ();
 sg13g2_fill_2 FILLER_66_406 ();
 sg13g2_fill_1 FILLER_66_460 ();
 sg13g2_fill_2 FILLER_66_465 ();
 sg13g2_fill_2 FILLER_66_482 ();
 sg13g2_fill_2 FILLER_66_518 ();
 sg13g2_fill_2 FILLER_66_532 ();
 sg13g2_fill_1 FILLER_66_534 ();
 sg13g2_fill_2 FILLER_66_544 ();
 sg13g2_fill_1 FILLER_66_546 ();
 sg13g2_fill_1 FILLER_66_557 ();
 sg13g2_fill_1 FILLER_66_567 ();
 sg13g2_fill_1 FILLER_66_571 ();
 sg13g2_fill_2 FILLER_66_582 ();
 sg13g2_fill_1 FILLER_66_584 ();
 sg13g2_fill_2 FILLER_66_610 ();
 sg13g2_fill_1 FILLER_66_612 ();
 sg13g2_decap_8 FILLER_66_623 ();
 sg13g2_fill_1 FILLER_66_639 ();
 sg13g2_fill_1 FILLER_66_657 ();
 sg13g2_fill_1 FILLER_66_693 ();
 sg13g2_fill_1 FILLER_66_703 ();
 sg13g2_fill_2 FILLER_66_712 ();
 sg13g2_fill_2 FILLER_66_738 ();
 sg13g2_fill_1 FILLER_66_740 ();
 sg13g2_decap_8 FILLER_66_748 ();
 sg13g2_decap_4 FILLER_66_755 ();
 sg13g2_fill_1 FILLER_66_783 ();
 sg13g2_decap_4 FILLER_66_790 ();
 sg13g2_fill_2 FILLER_66_806 ();
 sg13g2_decap_4 FILLER_66_839 ();
 sg13g2_decap_8 FILLER_66_855 ();
 sg13g2_fill_1 FILLER_66_862 ();
 sg13g2_fill_2 FILLER_66_868 ();
 sg13g2_fill_2 FILLER_66_888 ();
 sg13g2_fill_1 FILLER_66_907 ();
 sg13g2_decap_4 FILLER_66_917 ();
 sg13g2_fill_1 FILLER_66_978 ();
 sg13g2_fill_1 FILLER_66_992 ();
 sg13g2_decap_4 FILLER_66_1006 ();
 sg13g2_fill_2 FILLER_66_1010 ();
 sg13g2_decap_8 FILLER_66_1023 ();
 sg13g2_decap_8 FILLER_66_1030 ();
 sg13g2_decap_8 FILLER_66_1037 ();
 sg13g2_decap_8 FILLER_66_1044 ();
 sg13g2_decap_8 FILLER_66_1051 ();
 sg13g2_decap_8 FILLER_66_1058 ();
 sg13g2_decap_8 FILLER_66_1065 ();
 sg13g2_decap_8 FILLER_66_1072 ();
 sg13g2_decap_8 FILLER_66_1079 ();
 sg13g2_decap_8 FILLER_66_1086 ();
 sg13g2_decap_8 FILLER_66_1093 ();
 sg13g2_decap_8 FILLER_66_1100 ();
 sg13g2_decap_8 FILLER_66_1107 ();
 sg13g2_decap_8 FILLER_66_1114 ();
 sg13g2_decap_8 FILLER_66_1121 ();
 sg13g2_decap_8 FILLER_66_1128 ();
 sg13g2_decap_8 FILLER_66_1135 ();
 sg13g2_decap_8 FILLER_66_1142 ();
 sg13g2_decap_8 FILLER_66_1149 ();
 sg13g2_decap_8 FILLER_66_1156 ();
 sg13g2_decap_8 FILLER_66_1163 ();
 sg13g2_decap_8 FILLER_66_1170 ();
 sg13g2_decap_8 FILLER_66_1177 ();
 sg13g2_decap_8 FILLER_66_1184 ();
 sg13g2_decap_8 FILLER_66_1191 ();
 sg13g2_decap_8 FILLER_66_1198 ();
 sg13g2_decap_8 FILLER_66_1205 ();
 sg13g2_decap_8 FILLER_66_1212 ();
 sg13g2_decap_8 FILLER_66_1219 ();
 sg13g2_decap_8 FILLER_66_1226 ();
 sg13g2_decap_8 FILLER_66_1233 ();
 sg13g2_decap_8 FILLER_66_1240 ();
 sg13g2_decap_8 FILLER_66_1247 ();
 sg13g2_decap_8 FILLER_66_1254 ();
 sg13g2_decap_8 FILLER_66_1261 ();
 sg13g2_decap_8 FILLER_66_1268 ();
 sg13g2_decap_8 FILLER_66_1275 ();
 sg13g2_decap_8 FILLER_66_1282 ();
 sg13g2_decap_8 FILLER_66_1289 ();
 sg13g2_decap_8 FILLER_66_1296 ();
 sg13g2_decap_8 FILLER_66_1303 ();
 sg13g2_decap_8 FILLER_66_1310 ();
 sg13g2_decap_8 FILLER_66_1317 ();
 sg13g2_decap_8 FILLER_66_1324 ();
 sg13g2_decap_8 FILLER_66_1331 ();
 sg13g2_decap_8 FILLER_66_1338 ();
 sg13g2_decap_8 FILLER_66_1345 ();
 sg13g2_decap_8 FILLER_66_1352 ();
 sg13g2_decap_8 FILLER_66_1359 ();
 sg13g2_decap_8 FILLER_66_1366 ();
 sg13g2_decap_8 FILLER_66_1373 ();
 sg13g2_decap_8 FILLER_66_1380 ();
 sg13g2_decap_8 FILLER_66_1387 ();
 sg13g2_decap_8 FILLER_66_1394 ();
 sg13g2_decap_8 FILLER_66_1401 ();
 sg13g2_decap_8 FILLER_66_1408 ();
 sg13g2_decap_8 FILLER_66_1415 ();
 sg13g2_decap_8 FILLER_66_1422 ();
 sg13g2_decap_8 FILLER_66_1429 ();
 sg13g2_decap_8 FILLER_66_1436 ();
 sg13g2_decap_8 FILLER_66_1443 ();
 sg13g2_decap_8 FILLER_66_1450 ();
 sg13g2_decap_8 FILLER_66_1457 ();
 sg13g2_decap_8 FILLER_66_1464 ();
 sg13g2_decap_8 FILLER_66_1471 ();
 sg13g2_decap_8 FILLER_66_1478 ();
 sg13g2_decap_8 FILLER_66_1485 ();
 sg13g2_decap_8 FILLER_66_1492 ();
 sg13g2_decap_8 FILLER_66_1499 ();
 sg13g2_decap_8 FILLER_66_1506 ();
 sg13g2_decap_8 FILLER_66_1513 ();
 sg13g2_decap_8 FILLER_66_1520 ();
 sg13g2_decap_8 FILLER_66_1527 ();
 sg13g2_decap_8 FILLER_66_1534 ();
 sg13g2_decap_8 FILLER_66_1541 ();
 sg13g2_decap_8 FILLER_66_1548 ();
 sg13g2_decap_8 FILLER_66_1555 ();
 sg13g2_decap_8 FILLER_66_1562 ();
 sg13g2_decap_8 FILLER_66_1569 ();
 sg13g2_decap_8 FILLER_66_1576 ();
 sg13g2_decap_8 FILLER_66_1583 ();
 sg13g2_decap_8 FILLER_66_1590 ();
 sg13g2_decap_8 FILLER_66_1597 ();
 sg13g2_decap_8 FILLER_66_1604 ();
 sg13g2_decap_8 FILLER_66_1611 ();
 sg13g2_decap_8 FILLER_66_1618 ();
 sg13g2_decap_8 FILLER_66_1625 ();
 sg13g2_decap_8 FILLER_66_1632 ();
 sg13g2_decap_8 FILLER_66_1639 ();
 sg13g2_decap_8 FILLER_66_1646 ();
 sg13g2_decap_8 FILLER_66_1653 ();
 sg13g2_decap_8 FILLER_66_1660 ();
 sg13g2_decap_8 FILLER_66_1667 ();
 sg13g2_decap_8 FILLER_66_1674 ();
 sg13g2_decap_8 FILLER_66_1681 ();
 sg13g2_decap_8 FILLER_66_1688 ();
 sg13g2_decap_8 FILLER_66_1695 ();
 sg13g2_decap_8 FILLER_66_1702 ();
 sg13g2_decap_8 FILLER_66_1709 ();
 sg13g2_decap_8 FILLER_66_1716 ();
 sg13g2_decap_8 FILLER_66_1723 ();
 sg13g2_decap_8 FILLER_66_1730 ();
 sg13g2_decap_8 FILLER_66_1737 ();
 sg13g2_decap_8 FILLER_66_1744 ();
 sg13g2_decap_8 FILLER_66_1751 ();
 sg13g2_decap_8 FILLER_66_1758 ();
 sg13g2_fill_2 FILLER_66_1765 ();
 sg13g2_fill_1 FILLER_66_1767 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_4 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_103 ();
 sg13g2_decap_8 FILLER_67_110 ();
 sg13g2_decap_8 FILLER_67_117 ();
 sg13g2_fill_2 FILLER_67_211 ();
 sg13g2_fill_2 FILLER_67_235 ();
 sg13g2_fill_2 FILLER_67_243 ();
 sg13g2_fill_1 FILLER_67_245 ();
 sg13g2_fill_1 FILLER_67_266 ();
 sg13g2_fill_2 FILLER_67_356 ();
 sg13g2_fill_2 FILLER_67_392 ();
 sg13g2_fill_1 FILLER_67_402 ();
 sg13g2_fill_1 FILLER_67_419 ();
 sg13g2_fill_2 FILLER_67_429 ();
 sg13g2_fill_2 FILLER_67_448 ();
 sg13g2_fill_1 FILLER_67_450 ();
 sg13g2_fill_2 FILLER_67_493 ();
 sg13g2_fill_1 FILLER_67_495 ();
 sg13g2_fill_2 FILLER_67_509 ();
 sg13g2_fill_1 FILLER_67_511 ();
 sg13g2_fill_2 FILLER_67_516 ();
 sg13g2_fill_1 FILLER_67_518 ();
 sg13g2_fill_2 FILLER_67_524 ();
 sg13g2_fill_1 FILLER_67_526 ();
 sg13g2_fill_1 FILLER_67_535 ();
 sg13g2_fill_2 FILLER_67_542 ();
 sg13g2_fill_1 FILLER_67_544 ();
 sg13g2_fill_2 FILLER_67_555 ();
 sg13g2_fill_1 FILLER_67_557 ();
 sg13g2_fill_2 FILLER_67_566 ();
 sg13g2_fill_2 FILLER_67_577 ();
 sg13g2_fill_1 FILLER_67_592 ();
 sg13g2_decap_4 FILLER_67_603 ();
 sg13g2_fill_2 FILLER_67_607 ();
 sg13g2_fill_1 FILLER_67_697 ();
 sg13g2_fill_1 FILLER_67_724 ();
 sg13g2_fill_2 FILLER_67_757 ();
 sg13g2_fill_1 FILLER_67_759 ();
 sg13g2_decap_4 FILLER_67_809 ();
 sg13g2_fill_1 FILLER_67_813 ();
 sg13g2_fill_2 FILLER_67_824 ();
 sg13g2_decap_8 FILLER_67_886 ();
 sg13g2_decap_8 FILLER_67_893 ();
 sg13g2_fill_2 FILLER_67_900 ();
 sg13g2_fill_1 FILLER_67_902 ();
 sg13g2_decap_4 FILLER_67_914 ();
 sg13g2_decap_8 FILLER_67_1002 ();
 sg13g2_decap_8 FILLER_67_1027 ();
 sg13g2_decap_8 FILLER_67_1034 ();
 sg13g2_decap_8 FILLER_67_1041 ();
 sg13g2_decap_8 FILLER_67_1048 ();
 sg13g2_decap_8 FILLER_67_1055 ();
 sg13g2_decap_8 FILLER_67_1062 ();
 sg13g2_decap_8 FILLER_67_1069 ();
 sg13g2_decap_8 FILLER_67_1076 ();
 sg13g2_decap_8 FILLER_67_1083 ();
 sg13g2_decap_8 FILLER_67_1090 ();
 sg13g2_decap_8 FILLER_67_1097 ();
 sg13g2_decap_8 FILLER_67_1104 ();
 sg13g2_decap_8 FILLER_67_1111 ();
 sg13g2_decap_8 FILLER_67_1118 ();
 sg13g2_decap_8 FILLER_67_1125 ();
 sg13g2_decap_8 FILLER_67_1132 ();
 sg13g2_decap_8 FILLER_67_1139 ();
 sg13g2_decap_8 FILLER_67_1146 ();
 sg13g2_decap_8 FILLER_67_1153 ();
 sg13g2_decap_8 FILLER_67_1160 ();
 sg13g2_decap_8 FILLER_67_1167 ();
 sg13g2_decap_8 FILLER_67_1174 ();
 sg13g2_decap_8 FILLER_67_1181 ();
 sg13g2_decap_8 FILLER_67_1188 ();
 sg13g2_decap_8 FILLER_67_1195 ();
 sg13g2_decap_8 FILLER_67_1202 ();
 sg13g2_decap_8 FILLER_67_1209 ();
 sg13g2_decap_8 FILLER_67_1216 ();
 sg13g2_decap_8 FILLER_67_1223 ();
 sg13g2_decap_8 FILLER_67_1230 ();
 sg13g2_decap_8 FILLER_67_1237 ();
 sg13g2_decap_8 FILLER_67_1244 ();
 sg13g2_decap_8 FILLER_67_1251 ();
 sg13g2_decap_8 FILLER_67_1258 ();
 sg13g2_decap_8 FILLER_67_1265 ();
 sg13g2_decap_8 FILLER_67_1272 ();
 sg13g2_decap_8 FILLER_67_1279 ();
 sg13g2_decap_8 FILLER_67_1286 ();
 sg13g2_decap_8 FILLER_67_1293 ();
 sg13g2_decap_8 FILLER_67_1300 ();
 sg13g2_decap_8 FILLER_67_1307 ();
 sg13g2_decap_8 FILLER_67_1314 ();
 sg13g2_decap_8 FILLER_67_1321 ();
 sg13g2_decap_8 FILLER_67_1328 ();
 sg13g2_decap_8 FILLER_67_1335 ();
 sg13g2_decap_8 FILLER_67_1342 ();
 sg13g2_decap_8 FILLER_67_1349 ();
 sg13g2_decap_8 FILLER_67_1356 ();
 sg13g2_decap_8 FILLER_67_1363 ();
 sg13g2_decap_8 FILLER_67_1370 ();
 sg13g2_decap_8 FILLER_67_1377 ();
 sg13g2_decap_8 FILLER_67_1384 ();
 sg13g2_decap_8 FILLER_67_1391 ();
 sg13g2_decap_8 FILLER_67_1398 ();
 sg13g2_decap_8 FILLER_67_1405 ();
 sg13g2_decap_8 FILLER_67_1412 ();
 sg13g2_decap_8 FILLER_67_1419 ();
 sg13g2_decap_8 FILLER_67_1426 ();
 sg13g2_decap_8 FILLER_67_1433 ();
 sg13g2_decap_8 FILLER_67_1440 ();
 sg13g2_decap_8 FILLER_67_1447 ();
 sg13g2_decap_8 FILLER_67_1454 ();
 sg13g2_decap_8 FILLER_67_1461 ();
 sg13g2_decap_8 FILLER_67_1468 ();
 sg13g2_decap_8 FILLER_67_1475 ();
 sg13g2_decap_8 FILLER_67_1482 ();
 sg13g2_decap_8 FILLER_67_1489 ();
 sg13g2_decap_8 FILLER_67_1496 ();
 sg13g2_decap_8 FILLER_67_1503 ();
 sg13g2_decap_8 FILLER_67_1510 ();
 sg13g2_decap_8 FILLER_67_1517 ();
 sg13g2_decap_8 FILLER_67_1524 ();
 sg13g2_decap_8 FILLER_67_1531 ();
 sg13g2_decap_8 FILLER_67_1538 ();
 sg13g2_decap_8 FILLER_67_1545 ();
 sg13g2_decap_8 FILLER_67_1552 ();
 sg13g2_decap_8 FILLER_67_1559 ();
 sg13g2_decap_8 FILLER_67_1566 ();
 sg13g2_decap_8 FILLER_67_1573 ();
 sg13g2_decap_8 FILLER_67_1580 ();
 sg13g2_decap_8 FILLER_67_1587 ();
 sg13g2_decap_8 FILLER_67_1594 ();
 sg13g2_decap_8 FILLER_67_1601 ();
 sg13g2_decap_8 FILLER_67_1608 ();
 sg13g2_decap_8 FILLER_67_1615 ();
 sg13g2_decap_8 FILLER_67_1622 ();
 sg13g2_decap_8 FILLER_67_1629 ();
 sg13g2_decap_8 FILLER_67_1636 ();
 sg13g2_decap_8 FILLER_67_1643 ();
 sg13g2_decap_8 FILLER_67_1650 ();
 sg13g2_decap_8 FILLER_67_1657 ();
 sg13g2_decap_8 FILLER_67_1664 ();
 sg13g2_decap_8 FILLER_67_1671 ();
 sg13g2_decap_8 FILLER_67_1678 ();
 sg13g2_decap_8 FILLER_67_1685 ();
 sg13g2_decap_8 FILLER_67_1692 ();
 sg13g2_decap_8 FILLER_67_1699 ();
 sg13g2_decap_8 FILLER_67_1706 ();
 sg13g2_decap_8 FILLER_67_1713 ();
 sg13g2_decap_8 FILLER_67_1720 ();
 sg13g2_decap_8 FILLER_67_1727 ();
 sg13g2_decap_8 FILLER_67_1734 ();
 sg13g2_decap_8 FILLER_67_1741 ();
 sg13g2_decap_8 FILLER_67_1748 ();
 sg13g2_decap_8 FILLER_67_1755 ();
 sg13g2_decap_4 FILLER_67_1762 ();
 sg13g2_fill_2 FILLER_67_1766 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_4 FILLER_68_126 ();
 sg13g2_fill_2 FILLER_68_130 ();
 sg13g2_decap_4 FILLER_68_135 ();
 sg13g2_decap_4 FILLER_68_143 ();
 sg13g2_fill_1 FILLER_68_178 ();
 sg13g2_decap_4 FILLER_68_192 ();
 sg13g2_fill_2 FILLER_68_196 ();
 sg13g2_decap_4 FILLER_68_210 ();
 sg13g2_fill_2 FILLER_68_224 ();
 sg13g2_fill_1 FILLER_68_226 ();
 sg13g2_decap_4 FILLER_68_233 ();
 sg13g2_decap_8 FILLER_68_245 ();
 sg13g2_fill_2 FILLER_68_252 ();
 sg13g2_decap_8 FILLER_68_258 ();
 sg13g2_fill_1 FILLER_68_265 ();
 sg13g2_fill_1 FILLER_68_275 ();
 sg13g2_fill_1 FILLER_68_337 ();
 sg13g2_fill_1 FILLER_68_382 ();
 sg13g2_fill_2 FILLER_68_388 ();
 sg13g2_fill_2 FILLER_68_396 ();
 sg13g2_fill_2 FILLER_68_424 ();
 sg13g2_fill_2 FILLER_68_443 ();
 sg13g2_fill_1 FILLER_68_450 ();
 sg13g2_fill_2 FILLER_68_460 ();
 sg13g2_fill_2 FILLER_68_477 ();
 sg13g2_decap_4 FILLER_68_511 ();
 sg13g2_fill_1 FILLER_68_533 ();
 sg13g2_fill_2 FILLER_68_541 ();
 sg13g2_fill_1 FILLER_68_543 ();
 sg13g2_fill_2 FILLER_68_569 ();
 sg13g2_fill_1 FILLER_68_571 ();
 sg13g2_fill_2 FILLER_68_581 ();
 sg13g2_fill_1 FILLER_68_583 ();
 sg13g2_decap_4 FILLER_68_617 ();
 sg13g2_decap_8 FILLER_68_631 ();
 sg13g2_decap_8 FILLER_68_638 ();
 sg13g2_decap_4 FILLER_68_658 ();
 sg13g2_fill_2 FILLER_68_662 ();
 sg13g2_fill_2 FILLER_68_694 ();
 sg13g2_decap_8 FILLER_68_706 ();
 sg13g2_fill_2 FILLER_68_713 ();
 sg13g2_fill_1 FILLER_68_715 ();
 sg13g2_fill_1 FILLER_68_720 ();
 sg13g2_fill_2 FILLER_68_740 ();
 sg13g2_fill_2 FILLER_68_746 ();
 sg13g2_fill_1 FILLER_68_748 ();
 sg13g2_decap_4 FILLER_68_754 ();
 sg13g2_fill_1 FILLER_68_769 ();
 sg13g2_decap_4 FILLER_68_785 ();
 sg13g2_fill_2 FILLER_68_789 ();
 sg13g2_decap_4 FILLER_68_801 ();
 sg13g2_decap_4 FILLER_68_814 ();
 sg13g2_fill_2 FILLER_68_821 ();
 sg13g2_fill_1 FILLER_68_823 ();
 sg13g2_decap_8 FILLER_68_829 ();
 sg13g2_decap_4 FILLER_68_836 ();
 sg13g2_decap_8 FILLER_68_846 ();
 sg13g2_fill_2 FILLER_68_853 ();
 sg13g2_fill_1 FILLER_68_855 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_fill_1 FILLER_68_875 ();
 sg13g2_fill_2 FILLER_68_889 ();
 sg13g2_fill_1 FILLER_68_891 ();
 sg13g2_fill_2 FILLER_68_921 ();
 sg13g2_fill_1 FILLER_68_923 ();
 sg13g2_fill_2 FILLER_68_958 ();
 sg13g2_fill_1 FILLER_68_960 ();
 sg13g2_decap_8 FILLER_68_978 ();
 sg13g2_fill_1 FILLER_68_985 ();
 sg13g2_fill_2 FILLER_68_1010 ();
 sg13g2_decap_8 FILLER_68_1017 ();
 sg13g2_decap_8 FILLER_68_1024 ();
 sg13g2_decap_8 FILLER_68_1031 ();
 sg13g2_decap_8 FILLER_68_1038 ();
 sg13g2_decap_8 FILLER_68_1045 ();
 sg13g2_decap_8 FILLER_68_1052 ();
 sg13g2_decap_8 FILLER_68_1059 ();
 sg13g2_decap_8 FILLER_68_1066 ();
 sg13g2_decap_8 FILLER_68_1073 ();
 sg13g2_decap_8 FILLER_68_1080 ();
 sg13g2_decap_8 FILLER_68_1087 ();
 sg13g2_decap_8 FILLER_68_1094 ();
 sg13g2_decap_8 FILLER_68_1101 ();
 sg13g2_decap_8 FILLER_68_1108 ();
 sg13g2_decap_8 FILLER_68_1115 ();
 sg13g2_decap_8 FILLER_68_1122 ();
 sg13g2_decap_8 FILLER_68_1129 ();
 sg13g2_decap_8 FILLER_68_1136 ();
 sg13g2_decap_8 FILLER_68_1143 ();
 sg13g2_decap_8 FILLER_68_1150 ();
 sg13g2_decap_8 FILLER_68_1157 ();
 sg13g2_decap_8 FILLER_68_1164 ();
 sg13g2_decap_8 FILLER_68_1171 ();
 sg13g2_decap_8 FILLER_68_1178 ();
 sg13g2_decap_8 FILLER_68_1185 ();
 sg13g2_decap_8 FILLER_68_1192 ();
 sg13g2_decap_8 FILLER_68_1199 ();
 sg13g2_decap_8 FILLER_68_1206 ();
 sg13g2_decap_8 FILLER_68_1213 ();
 sg13g2_decap_8 FILLER_68_1220 ();
 sg13g2_decap_8 FILLER_68_1227 ();
 sg13g2_decap_8 FILLER_68_1234 ();
 sg13g2_decap_8 FILLER_68_1241 ();
 sg13g2_decap_8 FILLER_68_1248 ();
 sg13g2_decap_8 FILLER_68_1255 ();
 sg13g2_decap_8 FILLER_68_1262 ();
 sg13g2_decap_8 FILLER_68_1269 ();
 sg13g2_decap_8 FILLER_68_1276 ();
 sg13g2_decap_8 FILLER_68_1283 ();
 sg13g2_decap_8 FILLER_68_1290 ();
 sg13g2_decap_8 FILLER_68_1297 ();
 sg13g2_decap_8 FILLER_68_1304 ();
 sg13g2_decap_8 FILLER_68_1311 ();
 sg13g2_decap_8 FILLER_68_1318 ();
 sg13g2_decap_8 FILLER_68_1325 ();
 sg13g2_decap_8 FILLER_68_1332 ();
 sg13g2_decap_8 FILLER_68_1339 ();
 sg13g2_decap_8 FILLER_68_1346 ();
 sg13g2_decap_8 FILLER_68_1353 ();
 sg13g2_decap_8 FILLER_68_1360 ();
 sg13g2_decap_8 FILLER_68_1367 ();
 sg13g2_decap_8 FILLER_68_1374 ();
 sg13g2_decap_8 FILLER_68_1381 ();
 sg13g2_decap_8 FILLER_68_1388 ();
 sg13g2_decap_8 FILLER_68_1395 ();
 sg13g2_decap_8 FILLER_68_1402 ();
 sg13g2_decap_8 FILLER_68_1409 ();
 sg13g2_decap_8 FILLER_68_1416 ();
 sg13g2_decap_8 FILLER_68_1423 ();
 sg13g2_decap_8 FILLER_68_1430 ();
 sg13g2_decap_8 FILLER_68_1437 ();
 sg13g2_decap_8 FILLER_68_1444 ();
 sg13g2_decap_8 FILLER_68_1451 ();
 sg13g2_decap_8 FILLER_68_1458 ();
 sg13g2_decap_8 FILLER_68_1465 ();
 sg13g2_decap_8 FILLER_68_1472 ();
 sg13g2_decap_8 FILLER_68_1479 ();
 sg13g2_decap_8 FILLER_68_1486 ();
 sg13g2_decap_8 FILLER_68_1493 ();
 sg13g2_decap_8 FILLER_68_1500 ();
 sg13g2_decap_8 FILLER_68_1507 ();
 sg13g2_decap_8 FILLER_68_1514 ();
 sg13g2_decap_8 FILLER_68_1521 ();
 sg13g2_decap_8 FILLER_68_1528 ();
 sg13g2_decap_8 FILLER_68_1535 ();
 sg13g2_decap_8 FILLER_68_1542 ();
 sg13g2_decap_8 FILLER_68_1549 ();
 sg13g2_decap_8 FILLER_68_1556 ();
 sg13g2_decap_8 FILLER_68_1563 ();
 sg13g2_decap_8 FILLER_68_1570 ();
 sg13g2_decap_8 FILLER_68_1577 ();
 sg13g2_decap_8 FILLER_68_1584 ();
 sg13g2_decap_8 FILLER_68_1591 ();
 sg13g2_decap_8 FILLER_68_1598 ();
 sg13g2_decap_8 FILLER_68_1605 ();
 sg13g2_decap_8 FILLER_68_1612 ();
 sg13g2_decap_8 FILLER_68_1619 ();
 sg13g2_decap_8 FILLER_68_1626 ();
 sg13g2_decap_8 FILLER_68_1633 ();
 sg13g2_decap_8 FILLER_68_1640 ();
 sg13g2_decap_8 FILLER_68_1647 ();
 sg13g2_decap_8 FILLER_68_1654 ();
 sg13g2_decap_8 FILLER_68_1661 ();
 sg13g2_decap_8 FILLER_68_1668 ();
 sg13g2_decap_8 FILLER_68_1675 ();
 sg13g2_decap_8 FILLER_68_1682 ();
 sg13g2_decap_8 FILLER_68_1689 ();
 sg13g2_decap_8 FILLER_68_1696 ();
 sg13g2_decap_8 FILLER_68_1703 ();
 sg13g2_decap_8 FILLER_68_1710 ();
 sg13g2_decap_8 FILLER_68_1717 ();
 sg13g2_decap_8 FILLER_68_1724 ();
 sg13g2_decap_8 FILLER_68_1731 ();
 sg13g2_decap_8 FILLER_68_1738 ();
 sg13g2_decap_8 FILLER_68_1745 ();
 sg13g2_decap_8 FILLER_68_1752 ();
 sg13g2_decap_8 FILLER_68_1759 ();
 sg13g2_fill_2 FILLER_68_1766 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_fill_2 FILLER_69_119 ();
 sg13g2_fill_1 FILLER_69_121 ();
 sg13g2_decap_4 FILLER_69_151 ();
 sg13g2_fill_2 FILLER_69_172 ();
 sg13g2_fill_2 FILLER_69_189 ();
 sg13g2_fill_1 FILLER_69_191 ();
 sg13g2_decap_4 FILLER_69_215 ();
 sg13g2_fill_1 FILLER_69_219 ();
 sg13g2_fill_1 FILLER_69_233 ();
 sg13g2_fill_2 FILLER_69_259 ();
 sg13g2_fill_1 FILLER_69_278 ();
 sg13g2_fill_1 FILLER_69_320 ();
 sg13g2_fill_2 FILLER_69_340 ();
 sg13g2_fill_1 FILLER_69_346 ();
 sg13g2_fill_1 FILLER_69_394 ();
 sg13g2_fill_2 FILLER_69_418 ();
 sg13g2_fill_1 FILLER_69_420 ();
 sg13g2_fill_1 FILLER_69_461 ();
 sg13g2_decap_8 FILLER_69_467 ();
 sg13g2_decap_4 FILLER_69_485 ();
 sg13g2_fill_1 FILLER_69_489 ();
 sg13g2_decap_4 FILLER_69_518 ();
 sg13g2_fill_1 FILLER_69_522 ();
 sg13g2_decap_8 FILLER_69_536 ();
 sg13g2_decap_4 FILLER_69_543 ();
 sg13g2_fill_2 FILLER_69_547 ();
 sg13g2_fill_1 FILLER_69_558 ();
 sg13g2_decap_4 FILLER_69_570 ();
 sg13g2_fill_2 FILLER_69_574 ();
 sg13g2_fill_1 FILLER_69_590 ();
 sg13g2_fill_2 FILLER_69_609 ();
 sg13g2_decap_8 FILLER_69_631 ();
 sg13g2_decap_4 FILLER_69_638 ();
 sg13g2_decap_4 FILLER_69_664 ();
 sg13g2_fill_1 FILLER_69_697 ();
 sg13g2_fill_2 FILLER_69_721 ();
 sg13g2_decap_8 FILLER_69_728 ();
 sg13g2_fill_2 FILLER_69_735 ();
 sg13g2_fill_2 FILLER_69_763 ();
 sg13g2_fill_1 FILLER_69_765 ();
 sg13g2_fill_1 FILLER_69_783 ();
 sg13g2_fill_1 FILLER_69_801 ();
 sg13g2_decap_4 FILLER_69_839 ();
 sg13g2_fill_2 FILLER_69_843 ();
 sg13g2_fill_1 FILLER_69_857 ();
 sg13g2_fill_2 FILLER_69_864 ();
 sg13g2_fill_2 FILLER_69_885 ();
 sg13g2_fill_1 FILLER_69_887 ();
 sg13g2_fill_1 FILLER_69_910 ();
 sg13g2_fill_2 FILLER_69_916 ();
 sg13g2_fill_1 FILLER_69_918 ();
 sg13g2_fill_1 FILLER_69_929 ();
 sg13g2_decap_4 FILLER_69_952 ();
 sg13g2_fill_2 FILLER_69_956 ();
 sg13g2_decap_4 FILLER_69_972 ();
 sg13g2_fill_1 FILLER_69_976 ();
 sg13g2_decap_8 FILLER_69_985 ();
 sg13g2_fill_2 FILLER_69_1004 ();
 sg13g2_fill_1 FILLER_69_1006 ();
 sg13g2_decap_8 FILLER_69_1025 ();
 sg13g2_decap_8 FILLER_69_1032 ();
 sg13g2_decap_8 FILLER_69_1039 ();
 sg13g2_decap_8 FILLER_69_1046 ();
 sg13g2_decap_8 FILLER_69_1053 ();
 sg13g2_decap_8 FILLER_69_1060 ();
 sg13g2_decap_8 FILLER_69_1067 ();
 sg13g2_decap_8 FILLER_69_1074 ();
 sg13g2_decap_8 FILLER_69_1081 ();
 sg13g2_decap_8 FILLER_69_1088 ();
 sg13g2_decap_8 FILLER_69_1095 ();
 sg13g2_decap_8 FILLER_69_1102 ();
 sg13g2_decap_8 FILLER_69_1109 ();
 sg13g2_decap_8 FILLER_69_1116 ();
 sg13g2_decap_8 FILLER_69_1123 ();
 sg13g2_decap_8 FILLER_69_1130 ();
 sg13g2_decap_8 FILLER_69_1137 ();
 sg13g2_decap_8 FILLER_69_1144 ();
 sg13g2_decap_8 FILLER_69_1151 ();
 sg13g2_decap_8 FILLER_69_1158 ();
 sg13g2_decap_8 FILLER_69_1165 ();
 sg13g2_decap_8 FILLER_69_1172 ();
 sg13g2_decap_8 FILLER_69_1179 ();
 sg13g2_decap_8 FILLER_69_1186 ();
 sg13g2_decap_8 FILLER_69_1193 ();
 sg13g2_decap_8 FILLER_69_1200 ();
 sg13g2_decap_8 FILLER_69_1207 ();
 sg13g2_decap_8 FILLER_69_1214 ();
 sg13g2_decap_8 FILLER_69_1221 ();
 sg13g2_decap_8 FILLER_69_1228 ();
 sg13g2_decap_8 FILLER_69_1235 ();
 sg13g2_decap_8 FILLER_69_1242 ();
 sg13g2_decap_8 FILLER_69_1249 ();
 sg13g2_decap_8 FILLER_69_1256 ();
 sg13g2_decap_8 FILLER_69_1263 ();
 sg13g2_decap_8 FILLER_69_1270 ();
 sg13g2_decap_8 FILLER_69_1277 ();
 sg13g2_decap_8 FILLER_69_1284 ();
 sg13g2_decap_8 FILLER_69_1291 ();
 sg13g2_decap_8 FILLER_69_1298 ();
 sg13g2_decap_8 FILLER_69_1305 ();
 sg13g2_decap_8 FILLER_69_1312 ();
 sg13g2_decap_8 FILLER_69_1319 ();
 sg13g2_decap_8 FILLER_69_1326 ();
 sg13g2_decap_8 FILLER_69_1333 ();
 sg13g2_decap_8 FILLER_69_1340 ();
 sg13g2_decap_8 FILLER_69_1347 ();
 sg13g2_decap_8 FILLER_69_1354 ();
 sg13g2_decap_8 FILLER_69_1361 ();
 sg13g2_decap_8 FILLER_69_1368 ();
 sg13g2_decap_8 FILLER_69_1375 ();
 sg13g2_decap_8 FILLER_69_1382 ();
 sg13g2_decap_8 FILLER_69_1389 ();
 sg13g2_decap_8 FILLER_69_1396 ();
 sg13g2_decap_8 FILLER_69_1403 ();
 sg13g2_decap_8 FILLER_69_1410 ();
 sg13g2_decap_8 FILLER_69_1417 ();
 sg13g2_decap_8 FILLER_69_1424 ();
 sg13g2_decap_8 FILLER_69_1431 ();
 sg13g2_decap_8 FILLER_69_1438 ();
 sg13g2_decap_8 FILLER_69_1445 ();
 sg13g2_decap_8 FILLER_69_1452 ();
 sg13g2_decap_8 FILLER_69_1459 ();
 sg13g2_decap_8 FILLER_69_1466 ();
 sg13g2_decap_8 FILLER_69_1473 ();
 sg13g2_decap_8 FILLER_69_1480 ();
 sg13g2_decap_8 FILLER_69_1487 ();
 sg13g2_decap_8 FILLER_69_1494 ();
 sg13g2_decap_8 FILLER_69_1501 ();
 sg13g2_decap_8 FILLER_69_1508 ();
 sg13g2_decap_8 FILLER_69_1515 ();
 sg13g2_decap_8 FILLER_69_1522 ();
 sg13g2_decap_8 FILLER_69_1529 ();
 sg13g2_decap_8 FILLER_69_1536 ();
 sg13g2_decap_8 FILLER_69_1543 ();
 sg13g2_decap_8 FILLER_69_1550 ();
 sg13g2_decap_8 FILLER_69_1557 ();
 sg13g2_decap_8 FILLER_69_1564 ();
 sg13g2_decap_8 FILLER_69_1571 ();
 sg13g2_decap_8 FILLER_69_1578 ();
 sg13g2_decap_8 FILLER_69_1585 ();
 sg13g2_decap_8 FILLER_69_1592 ();
 sg13g2_decap_8 FILLER_69_1599 ();
 sg13g2_decap_8 FILLER_69_1606 ();
 sg13g2_decap_8 FILLER_69_1613 ();
 sg13g2_decap_8 FILLER_69_1620 ();
 sg13g2_decap_8 FILLER_69_1627 ();
 sg13g2_decap_8 FILLER_69_1634 ();
 sg13g2_decap_8 FILLER_69_1641 ();
 sg13g2_decap_8 FILLER_69_1648 ();
 sg13g2_decap_8 FILLER_69_1655 ();
 sg13g2_decap_8 FILLER_69_1662 ();
 sg13g2_decap_8 FILLER_69_1669 ();
 sg13g2_decap_8 FILLER_69_1676 ();
 sg13g2_decap_8 FILLER_69_1683 ();
 sg13g2_decap_8 FILLER_69_1690 ();
 sg13g2_decap_8 FILLER_69_1697 ();
 sg13g2_decap_8 FILLER_69_1704 ();
 sg13g2_decap_8 FILLER_69_1711 ();
 sg13g2_decap_8 FILLER_69_1718 ();
 sg13g2_decap_8 FILLER_69_1725 ();
 sg13g2_decap_8 FILLER_69_1732 ();
 sg13g2_decap_8 FILLER_69_1739 ();
 sg13g2_decap_8 FILLER_69_1746 ();
 sg13g2_decap_8 FILLER_69_1753 ();
 sg13g2_decap_8 FILLER_69_1760 ();
 sg13g2_fill_1 FILLER_69_1767 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_4 FILLER_70_126 ();
 sg13g2_fill_2 FILLER_70_130 ();
 sg13g2_fill_1 FILLER_70_190 ();
 sg13g2_fill_1 FILLER_70_213 ();
 sg13g2_fill_2 FILLER_70_231 ();
 sg13g2_fill_2 FILLER_70_238 ();
 sg13g2_decap_8 FILLER_70_250 ();
 sg13g2_decap_8 FILLER_70_257 ();
 sg13g2_fill_2 FILLER_70_264 ();
 sg13g2_fill_1 FILLER_70_266 ();
 sg13g2_fill_2 FILLER_70_271 ();
 sg13g2_fill_1 FILLER_70_273 ();
 sg13g2_fill_2 FILLER_70_368 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_fill_2 FILLER_70_424 ();
 sg13g2_fill_2 FILLER_70_470 ();
 sg13g2_decap_4 FILLER_70_502 ();
 sg13g2_decap_4 FILLER_70_510 ();
 sg13g2_fill_2 FILLER_70_514 ();
 sg13g2_fill_1 FILLER_70_538 ();
 sg13g2_decap_4 FILLER_70_563 ();
 sg13g2_fill_1 FILLER_70_589 ();
 sg13g2_decap_4 FILLER_70_626 ();
 sg13g2_fill_1 FILLER_70_630 ();
 sg13g2_fill_2 FILLER_70_698 ();
 sg13g2_fill_1 FILLER_70_711 ();
 sg13g2_fill_2 FILLER_70_729 ();
 sg13g2_decap_4 FILLER_70_750 ();
 sg13g2_fill_2 FILLER_70_754 ();
 sg13g2_fill_2 FILLER_70_768 ();
 sg13g2_decap_4 FILLER_70_787 ();
 sg13g2_fill_1 FILLER_70_791 ();
 sg13g2_decap_8 FILLER_70_797 ();
 sg13g2_decap_8 FILLER_70_804 ();
 sg13g2_decap_8 FILLER_70_811 ();
 sg13g2_decap_4 FILLER_70_818 ();
 sg13g2_fill_2 FILLER_70_822 ();
 sg13g2_fill_1 FILLER_70_829 ();
 sg13g2_decap_8 FILLER_70_852 ();
 sg13g2_decap_8 FILLER_70_859 ();
 sg13g2_fill_1 FILLER_70_866 ();
 sg13g2_decap_4 FILLER_70_895 ();
 sg13g2_fill_2 FILLER_70_909 ();
 sg13g2_decap_8 FILLER_70_919 ();
 sg13g2_decap_8 FILLER_70_926 ();
 sg13g2_decap_8 FILLER_70_933 ();
 sg13g2_decap_8 FILLER_70_961 ();
 sg13g2_decap_8 FILLER_70_968 ();
 sg13g2_decap_8 FILLER_70_975 ();
 sg13g2_fill_2 FILLER_70_982 ();
 sg13g2_decap_4 FILLER_70_991 ();
 sg13g2_fill_1 FILLER_70_1003 ();
 sg13g2_decap_4 FILLER_70_1008 ();
 sg13g2_fill_1 FILLER_70_1012 ();
 sg13g2_decap_4 FILLER_70_1017 ();
 sg13g2_decap_8 FILLER_70_1036 ();
 sg13g2_decap_8 FILLER_70_1043 ();
 sg13g2_decap_8 FILLER_70_1050 ();
 sg13g2_decap_8 FILLER_70_1057 ();
 sg13g2_decap_8 FILLER_70_1064 ();
 sg13g2_decap_8 FILLER_70_1071 ();
 sg13g2_decap_8 FILLER_70_1078 ();
 sg13g2_decap_8 FILLER_70_1085 ();
 sg13g2_decap_8 FILLER_70_1092 ();
 sg13g2_decap_8 FILLER_70_1099 ();
 sg13g2_decap_8 FILLER_70_1106 ();
 sg13g2_decap_8 FILLER_70_1113 ();
 sg13g2_decap_8 FILLER_70_1120 ();
 sg13g2_decap_8 FILLER_70_1127 ();
 sg13g2_decap_8 FILLER_70_1134 ();
 sg13g2_decap_8 FILLER_70_1141 ();
 sg13g2_decap_8 FILLER_70_1148 ();
 sg13g2_decap_8 FILLER_70_1155 ();
 sg13g2_decap_8 FILLER_70_1162 ();
 sg13g2_decap_8 FILLER_70_1169 ();
 sg13g2_decap_8 FILLER_70_1176 ();
 sg13g2_decap_8 FILLER_70_1183 ();
 sg13g2_decap_8 FILLER_70_1190 ();
 sg13g2_decap_8 FILLER_70_1197 ();
 sg13g2_decap_8 FILLER_70_1204 ();
 sg13g2_decap_8 FILLER_70_1211 ();
 sg13g2_decap_8 FILLER_70_1218 ();
 sg13g2_decap_8 FILLER_70_1225 ();
 sg13g2_decap_8 FILLER_70_1232 ();
 sg13g2_decap_8 FILLER_70_1239 ();
 sg13g2_decap_8 FILLER_70_1246 ();
 sg13g2_decap_8 FILLER_70_1253 ();
 sg13g2_decap_8 FILLER_70_1260 ();
 sg13g2_decap_8 FILLER_70_1267 ();
 sg13g2_decap_8 FILLER_70_1274 ();
 sg13g2_decap_8 FILLER_70_1281 ();
 sg13g2_decap_8 FILLER_70_1288 ();
 sg13g2_decap_8 FILLER_70_1295 ();
 sg13g2_decap_8 FILLER_70_1302 ();
 sg13g2_decap_8 FILLER_70_1309 ();
 sg13g2_decap_8 FILLER_70_1316 ();
 sg13g2_decap_8 FILLER_70_1323 ();
 sg13g2_decap_8 FILLER_70_1330 ();
 sg13g2_decap_8 FILLER_70_1337 ();
 sg13g2_decap_8 FILLER_70_1344 ();
 sg13g2_decap_8 FILLER_70_1351 ();
 sg13g2_decap_8 FILLER_70_1358 ();
 sg13g2_decap_8 FILLER_70_1365 ();
 sg13g2_decap_8 FILLER_70_1372 ();
 sg13g2_decap_8 FILLER_70_1379 ();
 sg13g2_decap_8 FILLER_70_1386 ();
 sg13g2_decap_8 FILLER_70_1393 ();
 sg13g2_decap_8 FILLER_70_1400 ();
 sg13g2_decap_8 FILLER_70_1407 ();
 sg13g2_decap_8 FILLER_70_1414 ();
 sg13g2_decap_8 FILLER_70_1421 ();
 sg13g2_decap_8 FILLER_70_1428 ();
 sg13g2_decap_8 FILLER_70_1435 ();
 sg13g2_decap_8 FILLER_70_1442 ();
 sg13g2_decap_8 FILLER_70_1449 ();
 sg13g2_decap_8 FILLER_70_1456 ();
 sg13g2_decap_8 FILLER_70_1463 ();
 sg13g2_decap_8 FILLER_70_1470 ();
 sg13g2_decap_8 FILLER_70_1477 ();
 sg13g2_decap_8 FILLER_70_1484 ();
 sg13g2_decap_8 FILLER_70_1491 ();
 sg13g2_decap_8 FILLER_70_1498 ();
 sg13g2_decap_8 FILLER_70_1505 ();
 sg13g2_decap_8 FILLER_70_1512 ();
 sg13g2_decap_8 FILLER_70_1519 ();
 sg13g2_decap_8 FILLER_70_1526 ();
 sg13g2_decap_8 FILLER_70_1533 ();
 sg13g2_decap_8 FILLER_70_1540 ();
 sg13g2_decap_8 FILLER_70_1547 ();
 sg13g2_decap_8 FILLER_70_1554 ();
 sg13g2_decap_8 FILLER_70_1561 ();
 sg13g2_decap_8 FILLER_70_1568 ();
 sg13g2_decap_8 FILLER_70_1575 ();
 sg13g2_decap_8 FILLER_70_1582 ();
 sg13g2_decap_8 FILLER_70_1589 ();
 sg13g2_decap_8 FILLER_70_1596 ();
 sg13g2_decap_8 FILLER_70_1603 ();
 sg13g2_decap_8 FILLER_70_1610 ();
 sg13g2_decap_8 FILLER_70_1617 ();
 sg13g2_decap_8 FILLER_70_1624 ();
 sg13g2_decap_8 FILLER_70_1631 ();
 sg13g2_decap_8 FILLER_70_1638 ();
 sg13g2_decap_8 FILLER_70_1645 ();
 sg13g2_decap_8 FILLER_70_1652 ();
 sg13g2_decap_8 FILLER_70_1659 ();
 sg13g2_decap_8 FILLER_70_1666 ();
 sg13g2_decap_8 FILLER_70_1673 ();
 sg13g2_decap_8 FILLER_70_1680 ();
 sg13g2_decap_8 FILLER_70_1687 ();
 sg13g2_decap_8 FILLER_70_1694 ();
 sg13g2_decap_8 FILLER_70_1701 ();
 sg13g2_decap_8 FILLER_70_1708 ();
 sg13g2_decap_8 FILLER_70_1715 ();
 sg13g2_decap_8 FILLER_70_1722 ();
 sg13g2_decap_8 FILLER_70_1729 ();
 sg13g2_decap_8 FILLER_70_1736 ();
 sg13g2_decap_8 FILLER_70_1743 ();
 sg13g2_decap_8 FILLER_70_1750 ();
 sg13g2_decap_8 FILLER_70_1757 ();
 sg13g2_decap_4 FILLER_70_1764 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_4 FILLER_71_133 ();
 sg13g2_fill_2 FILLER_71_137 ();
 sg13g2_decap_4 FILLER_71_142 ();
 sg13g2_fill_1 FILLER_71_146 ();
 sg13g2_decap_8 FILLER_71_151 ();
 sg13g2_fill_2 FILLER_71_158 ();
 sg13g2_fill_1 FILLER_71_160 ();
 sg13g2_fill_1 FILLER_71_180 ();
 sg13g2_fill_2 FILLER_71_218 ();
 sg13g2_fill_1 FILLER_71_220 ();
 sg13g2_decap_4 FILLER_71_231 ();
 sg13g2_fill_2 FILLER_71_235 ();
 sg13g2_decap_4 FILLER_71_240 ();
 sg13g2_fill_1 FILLER_71_244 ();
 sg13g2_fill_2 FILLER_71_292 ();
 sg13g2_fill_1 FILLER_71_294 ();
 sg13g2_fill_1 FILLER_71_351 ();
 sg13g2_fill_1 FILLER_71_378 ();
 sg13g2_fill_2 FILLER_71_393 ();
 sg13g2_fill_1 FILLER_71_410 ();
 sg13g2_fill_1 FILLER_71_422 ();
 sg13g2_decap_4 FILLER_71_458 ();
 sg13g2_fill_2 FILLER_71_469 ();
 sg13g2_decap_4 FILLER_71_475 ();
 sg13g2_fill_2 FILLER_71_486 ();
 sg13g2_decap_4 FILLER_71_498 ();
 sg13g2_fill_1 FILLER_71_523 ();
 sg13g2_fill_1 FILLER_71_537 ();
 sg13g2_decap_4 FILLER_71_543 ();
 sg13g2_fill_2 FILLER_71_547 ();
 sg13g2_decap_8 FILLER_71_554 ();
 sg13g2_decap_4 FILLER_71_565 ();
 sg13g2_fill_2 FILLER_71_574 ();
 sg13g2_fill_1 FILLER_71_576 ();
 sg13g2_fill_2 FILLER_71_582 ();
 sg13g2_decap_4 FILLER_71_609 ();
 sg13g2_fill_1 FILLER_71_613 ();
 sg13g2_decap_8 FILLER_71_662 ();
 sg13g2_decap_4 FILLER_71_669 ();
 sg13g2_fill_2 FILLER_71_673 ();
 sg13g2_fill_2 FILLER_71_732 ();
 sg13g2_fill_2 FILLER_71_748 ();
 sg13g2_fill_1 FILLER_71_750 ();
 sg13g2_fill_2 FILLER_71_756 ();
 sg13g2_decap_4 FILLER_71_780 ();
 sg13g2_fill_1 FILLER_71_813 ();
 sg13g2_decap_8 FILLER_71_829 ();
 sg13g2_decap_4 FILLER_71_836 ();
 sg13g2_decap_4 FILLER_71_857 ();
 sg13g2_decap_4 FILLER_71_869 ();
 sg13g2_fill_1 FILLER_71_873 ();
 sg13g2_fill_2 FILLER_71_878 ();
 sg13g2_fill_1 FILLER_71_880 ();
 sg13g2_fill_1 FILLER_71_890 ();
 sg13g2_decap_8 FILLER_71_904 ();
 sg13g2_decap_4 FILLER_71_911 ();
 sg13g2_fill_2 FILLER_71_928 ();
 sg13g2_fill_2 FILLER_71_939 ();
 sg13g2_fill_2 FILLER_71_946 ();
 sg13g2_fill_1 FILLER_71_961 ();
 sg13g2_fill_2 FILLER_71_974 ();
 sg13g2_fill_1 FILLER_71_976 ();
 sg13g2_fill_2 FILLER_71_1006 ();
 sg13g2_fill_1 FILLER_71_1008 ();
 sg13g2_decap_8 FILLER_71_1043 ();
 sg13g2_decap_8 FILLER_71_1050 ();
 sg13g2_decap_8 FILLER_71_1057 ();
 sg13g2_decap_8 FILLER_71_1064 ();
 sg13g2_decap_8 FILLER_71_1071 ();
 sg13g2_decap_8 FILLER_71_1078 ();
 sg13g2_decap_8 FILLER_71_1085 ();
 sg13g2_decap_8 FILLER_71_1092 ();
 sg13g2_decap_8 FILLER_71_1099 ();
 sg13g2_decap_8 FILLER_71_1106 ();
 sg13g2_decap_8 FILLER_71_1113 ();
 sg13g2_decap_8 FILLER_71_1120 ();
 sg13g2_decap_8 FILLER_71_1127 ();
 sg13g2_decap_8 FILLER_71_1134 ();
 sg13g2_decap_8 FILLER_71_1141 ();
 sg13g2_decap_8 FILLER_71_1148 ();
 sg13g2_decap_8 FILLER_71_1155 ();
 sg13g2_decap_8 FILLER_71_1162 ();
 sg13g2_decap_8 FILLER_71_1169 ();
 sg13g2_decap_8 FILLER_71_1176 ();
 sg13g2_decap_8 FILLER_71_1183 ();
 sg13g2_decap_8 FILLER_71_1190 ();
 sg13g2_decap_8 FILLER_71_1197 ();
 sg13g2_decap_8 FILLER_71_1204 ();
 sg13g2_decap_8 FILLER_71_1211 ();
 sg13g2_decap_8 FILLER_71_1218 ();
 sg13g2_decap_8 FILLER_71_1225 ();
 sg13g2_decap_8 FILLER_71_1232 ();
 sg13g2_decap_8 FILLER_71_1239 ();
 sg13g2_decap_8 FILLER_71_1246 ();
 sg13g2_decap_8 FILLER_71_1253 ();
 sg13g2_decap_8 FILLER_71_1260 ();
 sg13g2_decap_8 FILLER_71_1267 ();
 sg13g2_decap_8 FILLER_71_1274 ();
 sg13g2_decap_8 FILLER_71_1281 ();
 sg13g2_decap_8 FILLER_71_1288 ();
 sg13g2_decap_8 FILLER_71_1295 ();
 sg13g2_decap_8 FILLER_71_1302 ();
 sg13g2_decap_8 FILLER_71_1309 ();
 sg13g2_decap_8 FILLER_71_1316 ();
 sg13g2_decap_8 FILLER_71_1323 ();
 sg13g2_decap_8 FILLER_71_1330 ();
 sg13g2_decap_8 FILLER_71_1337 ();
 sg13g2_decap_8 FILLER_71_1344 ();
 sg13g2_decap_8 FILLER_71_1351 ();
 sg13g2_decap_8 FILLER_71_1358 ();
 sg13g2_decap_8 FILLER_71_1365 ();
 sg13g2_decap_8 FILLER_71_1372 ();
 sg13g2_decap_8 FILLER_71_1379 ();
 sg13g2_decap_8 FILLER_71_1386 ();
 sg13g2_decap_8 FILLER_71_1393 ();
 sg13g2_decap_8 FILLER_71_1400 ();
 sg13g2_decap_8 FILLER_71_1407 ();
 sg13g2_decap_8 FILLER_71_1414 ();
 sg13g2_decap_8 FILLER_71_1421 ();
 sg13g2_decap_8 FILLER_71_1428 ();
 sg13g2_decap_8 FILLER_71_1435 ();
 sg13g2_decap_8 FILLER_71_1442 ();
 sg13g2_decap_8 FILLER_71_1449 ();
 sg13g2_decap_8 FILLER_71_1456 ();
 sg13g2_decap_8 FILLER_71_1463 ();
 sg13g2_decap_8 FILLER_71_1470 ();
 sg13g2_decap_8 FILLER_71_1477 ();
 sg13g2_decap_8 FILLER_71_1484 ();
 sg13g2_decap_8 FILLER_71_1491 ();
 sg13g2_decap_8 FILLER_71_1498 ();
 sg13g2_decap_8 FILLER_71_1505 ();
 sg13g2_decap_8 FILLER_71_1512 ();
 sg13g2_decap_8 FILLER_71_1519 ();
 sg13g2_decap_8 FILLER_71_1526 ();
 sg13g2_decap_8 FILLER_71_1533 ();
 sg13g2_decap_8 FILLER_71_1540 ();
 sg13g2_decap_8 FILLER_71_1547 ();
 sg13g2_decap_8 FILLER_71_1554 ();
 sg13g2_decap_8 FILLER_71_1561 ();
 sg13g2_decap_8 FILLER_71_1568 ();
 sg13g2_decap_8 FILLER_71_1575 ();
 sg13g2_decap_8 FILLER_71_1582 ();
 sg13g2_decap_8 FILLER_71_1589 ();
 sg13g2_decap_8 FILLER_71_1596 ();
 sg13g2_decap_8 FILLER_71_1603 ();
 sg13g2_decap_8 FILLER_71_1610 ();
 sg13g2_decap_8 FILLER_71_1617 ();
 sg13g2_decap_8 FILLER_71_1624 ();
 sg13g2_decap_8 FILLER_71_1631 ();
 sg13g2_decap_8 FILLER_71_1638 ();
 sg13g2_decap_8 FILLER_71_1645 ();
 sg13g2_decap_8 FILLER_71_1652 ();
 sg13g2_decap_8 FILLER_71_1659 ();
 sg13g2_decap_8 FILLER_71_1666 ();
 sg13g2_decap_8 FILLER_71_1673 ();
 sg13g2_decap_8 FILLER_71_1680 ();
 sg13g2_decap_8 FILLER_71_1687 ();
 sg13g2_decap_8 FILLER_71_1694 ();
 sg13g2_decap_8 FILLER_71_1701 ();
 sg13g2_decap_8 FILLER_71_1708 ();
 sg13g2_decap_8 FILLER_71_1715 ();
 sg13g2_decap_8 FILLER_71_1722 ();
 sg13g2_decap_8 FILLER_71_1729 ();
 sg13g2_decap_8 FILLER_71_1736 ();
 sg13g2_decap_8 FILLER_71_1743 ();
 sg13g2_decap_8 FILLER_71_1750 ();
 sg13g2_decap_8 FILLER_71_1757 ();
 sg13g2_decap_4 FILLER_71_1764 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_fill_2 FILLER_72_168 ();
 sg13g2_fill_2 FILLER_72_225 ();
 sg13g2_fill_1 FILLER_72_227 ();
 sg13g2_fill_2 FILLER_72_232 ();
 sg13g2_fill_1 FILLER_72_234 ();
 sg13g2_decap_8 FILLER_72_261 ();
 sg13g2_fill_2 FILLER_72_268 ();
 sg13g2_fill_1 FILLER_72_270 ();
 sg13g2_fill_2 FILLER_72_323 ();
 sg13g2_fill_1 FILLER_72_325 ();
 sg13g2_decap_8 FILLER_72_352 ();
 sg13g2_fill_2 FILLER_72_359 ();
 sg13g2_fill_1 FILLER_72_361 ();
 sg13g2_fill_2 FILLER_72_429 ();
 sg13g2_fill_2 FILLER_72_440 ();
 sg13g2_fill_2 FILLER_72_456 ();
 sg13g2_fill_1 FILLER_72_458 ();
 sg13g2_fill_1 FILLER_72_464 ();
 sg13g2_decap_4 FILLER_72_498 ();
 sg13g2_decap_4 FILLER_72_508 ();
 sg13g2_fill_1 FILLER_72_512 ();
 sg13g2_fill_2 FILLER_72_527 ();
 sg13g2_fill_1 FILLER_72_529 ();
 sg13g2_decap_4 FILLER_72_573 ();
 sg13g2_decap_8 FILLER_72_582 ();
 sg13g2_decap_4 FILLER_72_589 ();
 sg13g2_fill_2 FILLER_72_593 ();
 sg13g2_fill_2 FILLER_72_607 ();
 sg13g2_fill_2 FILLER_72_613 ();
 sg13g2_fill_2 FILLER_72_627 ();
 sg13g2_fill_2 FILLER_72_664 ();
 sg13g2_fill_1 FILLER_72_666 ();
 sg13g2_decap_4 FILLER_72_671 ();
 sg13g2_fill_2 FILLER_72_675 ();
 sg13g2_fill_2 FILLER_72_699 ();
 sg13g2_fill_2 FILLER_72_706 ();
 sg13g2_fill_2 FILLER_72_734 ();
 sg13g2_fill_1 FILLER_72_784 ();
 sg13g2_fill_2 FILLER_72_793 ();
 sg13g2_fill_2 FILLER_72_808 ();
 sg13g2_fill_1 FILLER_72_823 ();
 sg13g2_fill_2 FILLER_72_842 ();
 sg13g2_fill_1 FILLER_72_864 ();
 sg13g2_fill_2 FILLER_72_876 ();
 sg13g2_fill_1 FILLER_72_878 ();
 sg13g2_fill_2 FILLER_72_903 ();
 sg13g2_fill_1 FILLER_72_905 ();
 sg13g2_decap_4 FILLER_72_932 ();
 sg13g2_decap_4 FILLER_72_947 ();
 sg13g2_fill_2 FILLER_72_961 ();
 sg13g2_decap_4 FILLER_72_967 ();
 sg13g2_fill_2 FILLER_72_988 ();
 sg13g2_fill_2 FILLER_72_1036 ();
 sg13g2_decap_8 FILLER_72_1044 ();
 sg13g2_decap_8 FILLER_72_1051 ();
 sg13g2_decap_8 FILLER_72_1058 ();
 sg13g2_decap_8 FILLER_72_1065 ();
 sg13g2_decap_8 FILLER_72_1072 ();
 sg13g2_decap_8 FILLER_72_1079 ();
 sg13g2_decap_8 FILLER_72_1086 ();
 sg13g2_decap_8 FILLER_72_1093 ();
 sg13g2_decap_8 FILLER_72_1100 ();
 sg13g2_decap_8 FILLER_72_1107 ();
 sg13g2_decap_8 FILLER_72_1114 ();
 sg13g2_decap_8 FILLER_72_1121 ();
 sg13g2_decap_8 FILLER_72_1128 ();
 sg13g2_decap_8 FILLER_72_1135 ();
 sg13g2_decap_8 FILLER_72_1142 ();
 sg13g2_decap_8 FILLER_72_1149 ();
 sg13g2_decap_8 FILLER_72_1156 ();
 sg13g2_decap_8 FILLER_72_1163 ();
 sg13g2_decap_8 FILLER_72_1170 ();
 sg13g2_decap_8 FILLER_72_1177 ();
 sg13g2_decap_8 FILLER_72_1184 ();
 sg13g2_decap_8 FILLER_72_1191 ();
 sg13g2_decap_8 FILLER_72_1198 ();
 sg13g2_decap_8 FILLER_72_1205 ();
 sg13g2_decap_8 FILLER_72_1212 ();
 sg13g2_decap_8 FILLER_72_1219 ();
 sg13g2_decap_8 FILLER_72_1226 ();
 sg13g2_decap_8 FILLER_72_1233 ();
 sg13g2_decap_8 FILLER_72_1240 ();
 sg13g2_decap_8 FILLER_72_1247 ();
 sg13g2_decap_8 FILLER_72_1254 ();
 sg13g2_decap_8 FILLER_72_1261 ();
 sg13g2_decap_8 FILLER_72_1268 ();
 sg13g2_decap_8 FILLER_72_1275 ();
 sg13g2_decap_8 FILLER_72_1282 ();
 sg13g2_decap_8 FILLER_72_1289 ();
 sg13g2_decap_8 FILLER_72_1296 ();
 sg13g2_decap_8 FILLER_72_1303 ();
 sg13g2_decap_8 FILLER_72_1310 ();
 sg13g2_decap_8 FILLER_72_1317 ();
 sg13g2_decap_8 FILLER_72_1324 ();
 sg13g2_decap_8 FILLER_72_1331 ();
 sg13g2_decap_8 FILLER_72_1338 ();
 sg13g2_decap_8 FILLER_72_1345 ();
 sg13g2_decap_8 FILLER_72_1352 ();
 sg13g2_decap_8 FILLER_72_1359 ();
 sg13g2_decap_8 FILLER_72_1366 ();
 sg13g2_decap_8 FILLER_72_1373 ();
 sg13g2_decap_8 FILLER_72_1380 ();
 sg13g2_decap_8 FILLER_72_1387 ();
 sg13g2_decap_8 FILLER_72_1394 ();
 sg13g2_decap_8 FILLER_72_1401 ();
 sg13g2_decap_8 FILLER_72_1408 ();
 sg13g2_decap_8 FILLER_72_1415 ();
 sg13g2_decap_8 FILLER_72_1422 ();
 sg13g2_decap_8 FILLER_72_1429 ();
 sg13g2_decap_8 FILLER_72_1436 ();
 sg13g2_decap_8 FILLER_72_1443 ();
 sg13g2_decap_8 FILLER_72_1450 ();
 sg13g2_decap_8 FILLER_72_1457 ();
 sg13g2_decap_8 FILLER_72_1464 ();
 sg13g2_decap_8 FILLER_72_1471 ();
 sg13g2_decap_8 FILLER_72_1478 ();
 sg13g2_decap_8 FILLER_72_1485 ();
 sg13g2_decap_8 FILLER_72_1492 ();
 sg13g2_decap_8 FILLER_72_1499 ();
 sg13g2_decap_8 FILLER_72_1506 ();
 sg13g2_decap_8 FILLER_72_1513 ();
 sg13g2_decap_8 FILLER_72_1520 ();
 sg13g2_decap_8 FILLER_72_1527 ();
 sg13g2_decap_8 FILLER_72_1534 ();
 sg13g2_decap_8 FILLER_72_1541 ();
 sg13g2_decap_8 FILLER_72_1548 ();
 sg13g2_decap_8 FILLER_72_1555 ();
 sg13g2_decap_8 FILLER_72_1562 ();
 sg13g2_decap_8 FILLER_72_1569 ();
 sg13g2_decap_8 FILLER_72_1576 ();
 sg13g2_decap_8 FILLER_72_1583 ();
 sg13g2_decap_8 FILLER_72_1590 ();
 sg13g2_decap_8 FILLER_72_1597 ();
 sg13g2_decap_8 FILLER_72_1604 ();
 sg13g2_decap_8 FILLER_72_1611 ();
 sg13g2_decap_8 FILLER_72_1618 ();
 sg13g2_decap_8 FILLER_72_1625 ();
 sg13g2_decap_8 FILLER_72_1632 ();
 sg13g2_decap_8 FILLER_72_1639 ();
 sg13g2_decap_8 FILLER_72_1646 ();
 sg13g2_decap_8 FILLER_72_1653 ();
 sg13g2_decap_8 FILLER_72_1660 ();
 sg13g2_decap_8 FILLER_72_1667 ();
 sg13g2_decap_8 FILLER_72_1674 ();
 sg13g2_decap_8 FILLER_72_1681 ();
 sg13g2_decap_8 FILLER_72_1688 ();
 sg13g2_decap_8 FILLER_72_1695 ();
 sg13g2_decap_8 FILLER_72_1702 ();
 sg13g2_decap_8 FILLER_72_1709 ();
 sg13g2_decap_8 FILLER_72_1716 ();
 sg13g2_decap_8 FILLER_72_1723 ();
 sg13g2_decap_8 FILLER_72_1730 ();
 sg13g2_decap_8 FILLER_72_1737 ();
 sg13g2_decap_8 FILLER_72_1744 ();
 sg13g2_decap_8 FILLER_72_1751 ();
 sg13g2_decap_8 FILLER_72_1758 ();
 sg13g2_fill_2 FILLER_72_1765 ();
 sg13g2_fill_1 FILLER_72_1767 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_fill_2 FILLER_73_178 ();
 sg13g2_fill_1 FILLER_73_180 ();
 sg13g2_decap_8 FILLER_73_185 ();
 sg13g2_decap_4 FILLER_73_192 ();
 sg13g2_decap_4 FILLER_73_201 ();
 sg13g2_fill_2 FILLER_73_205 ();
 sg13g2_decap_4 FILLER_73_211 ();
 sg13g2_fill_2 FILLER_73_215 ();
 sg13g2_decap_4 FILLER_73_252 ();
 sg13g2_decap_8 FILLER_73_282 ();
 sg13g2_decap_8 FILLER_73_289 ();
 sg13g2_fill_1 FILLER_73_296 ();
 sg13g2_decap_4 FILLER_73_323 ();
 sg13g2_fill_2 FILLER_73_327 ();
 sg13g2_decap_8 FILLER_73_355 ();
 sg13g2_decap_8 FILLER_73_362 ();
 sg13g2_decap_8 FILLER_73_369 ();
 sg13g2_decap_8 FILLER_73_376 ();
 sg13g2_decap_8 FILLER_73_383 ();
 sg13g2_decap_8 FILLER_73_390 ();
 sg13g2_decap_4 FILLER_73_397 ();
 sg13g2_fill_1 FILLER_73_401 ();
 sg13g2_fill_1 FILLER_73_467 ();
 sg13g2_decap_8 FILLER_73_480 ();
 sg13g2_fill_1 FILLER_73_487 ();
 sg13g2_fill_2 FILLER_73_498 ();
 sg13g2_fill_2 FILLER_73_530 ();
 sg13g2_fill_1 FILLER_73_543 ();
 sg13g2_fill_2 FILLER_73_553 ();
 sg13g2_fill_2 FILLER_73_558 ();
 sg13g2_decap_8 FILLER_73_577 ();
 sg13g2_fill_1 FILLER_73_584 ();
 sg13g2_fill_2 FILLER_73_594 ();
 sg13g2_fill_1 FILLER_73_596 ();
 sg13g2_fill_1 FILLER_73_613 ();
 sg13g2_fill_2 FILLER_73_623 ();
 sg13g2_fill_1 FILLER_73_625 ();
 sg13g2_fill_2 FILLER_73_643 ();
 sg13g2_fill_1 FILLER_73_645 ();
 sg13g2_decap_8 FILLER_73_667 ();
 sg13g2_decap_4 FILLER_73_674 ();
 sg13g2_fill_1 FILLER_73_678 ();
 sg13g2_fill_2 FILLER_73_715 ();
 sg13g2_fill_1 FILLER_73_717 ();
 sg13g2_fill_2 FILLER_73_731 ();
 sg13g2_fill_1 FILLER_73_733 ();
 sg13g2_decap_4 FILLER_73_747 ();
 sg13g2_decap_8 FILLER_73_756 ();
 sg13g2_fill_1 FILLER_73_763 ();
 sg13g2_fill_2 FILLER_73_778 ();
 sg13g2_decap_8 FILLER_73_816 ();
 sg13g2_decap_8 FILLER_73_836 ();
 sg13g2_decap_8 FILLER_73_843 ();
 sg13g2_decap_4 FILLER_73_850 ();
 sg13g2_fill_1 FILLER_73_854 ();
 sg13g2_fill_1 FILLER_73_876 ();
 sg13g2_fill_2 FILLER_73_895 ();
 sg13g2_decap_8 FILLER_73_902 ();
 sg13g2_decap_8 FILLER_73_909 ();
 sg13g2_fill_1 FILLER_73_916 ();
 sg13g2_decap_4 FILLER_73_921 ();
 sg13g2_fill_2 FILLER_73_925 ();
 sg13g2_fill_1 FILLER_73_943 ();
 sg13g2_decap_4 FILLER_73_969 ();
 sg13g2_fill_1 FILLER_73_973 ();
 sg13g2_fill_1 FILLER_73_982 ();
 sg13g2_decap_8 FILLER_73_1002 ();
 sg13g2_fill_1 FILLER_73_1009 ();
 sg13g2_decap_8 FILLER_73_1031 ();
 sg13g2_decap_8 FILLER_73_1050 ();
 sg13g2_decap_8 FILLER_73_1057 ();
 sg13g2_decap_8 FILLER_73_1064 ();
 sg13g2_decap_8 FILLER_73_1071 ();
 sg13g2_decap_8 FILLER_73_1078 ();
 sg13g2_decap_8 FILLER_73_1085 ();
 sg13g2_decap_8 FILLER_73_1092 ();
 sg13g2_decap_8 FILLER_73_1099 ();
 sg13g2_decap_8 FILLER_73_1106 ();
 sg13g2_decap_8 FILLER_73_1113 ();
 sg13g2_decap_8 FILLER_73_1120 ();
 sg13g2_decap_8 FILLER_73_1127 ();
 sg13g2_decap_8 FILLER_73_1134 ();
 sg13g2_decap_8 FILLER_73_1141 ();
 sg13g2_decap_8 FILLER_73_1148 ();
 sg13g2_decap_8 FILLER_73_1155 ();
 sg13g2_decap_8 FILLER_73_1162 ();
 sg13g2_decap_8 FILLER_73_1169 ();
 sg13g2_decap_8 FILLER_73_1176 ();
 sg13g2_decap_8 FILLER_73_1183 ();
 sg13g2_decap_8 FILLER_73_1190 ();
 sg13g2_decap_8 FILLER_73_1197 ();
 sg13g2_decap_8 FILLER_73_1204 ();
 sg13g2_decap_8 FILLER_73_1211 ();
 sg13g2_decap_8 FILLER_73_1218 ();
 sg13g2_decap_8 FILLER_73_1225 ();
 sg13g2_decap_8 FILLER_73_1232 ();
 sg13g2_decap_8 FILLER_73_1239 ();
 sg13g2_decap_8 FILLER_73_1246 ();
 sg13g2_decap_8 FILLER_73_1253 ();
 sg13g2_decap_8 FILLER_73_1260 ();
 sg13g2_decap_8 FILLER_73_1267 ();
 sg13g2_decap_8 FILLER_73_1274 ();
 sg13g2_decap_8 FILLER_73_1281 ();
 sg13g2_decap_8 FILLER_73_1288 ();
 sg13g2_decap_8 FILLER_73_1295 ();
 sg13g2_decap_8 FILLER_73_1302 ();
 sg13g2_decap_8 FILLER_73_1309 ();
 sg13g2_decap_8 FILLER_73_1316 ();
 sg13g2_decap_8 FILLER_73_1323 ();
 sg13g2_decap_8 FILLER_73_1330 ();
 sg13g2_decap_8 FILLER_73_1337 ();
 sg13g2_decap_8 FILLER_73_1344 ();
 sg13g2_decap_8 FILLER_73_1351 ();
 sg13g2_decap_8 FILLER_73_1358 ();
 sg13g2_decap_8 FILLER_73_1365 ();
 sg13g2_decap_8 FILLER_73_1372 ();
 sg13g2_decap_8 FILLER_73_1379 ();
 sg13g2_decap_8 FILLER_73_1386 ();
 sg13g2_decap_8 FILLER_73_1393 ();
 sg13g2_decap_8 FILLER_73_1400 ();
 sg13g2_decap_8 FILLER_73_1407 ();
 sg13g2_decap_8 FILLER_73_1414 ();
 sg13g2_decap_8 FILLER_73_1421 ();
 sg13g2_decap_8 FILLER_73_1428 ();
 sg13g2_decap_8 FILLER_73_1435 ();
 sg13g2_decap_8 FILLER_73_1442 ();
 sg13g2_decap_8 FILLER_73_1449 ();
 sg13g2_decap_8 FILLER_73_1456 ();
 sg13g2_decap_8 FILLER_73_1463 ();
 sg13g2_decap_8 FILLER_73_1470 ();
 sg13g2_decap_8 FILLER_73_1477 ();
 sg13g2_decap_8 FILLER_73_1484 ();
 sg13g2_decap_8 FILLER_73_1491 ();
 sg13g2_decap_8 FILLER_73_1498 ();
 sg13g2_decap_8 FILLER_73_1505 ();
 sg13g2_decap_8 FILLER_73_1512 ();
 sg13g2_decap_8 FILLER_73_1519 ();
 sg13g2_decap_8 FILLER_73_1526 ();
 sg13g2_decap_8 FILLER_73_1533 ();
 sg13g2_decap_8 FILLER_73_1540 ();
 sg13g2_decap_8 FILLER_73_1547 ();
 sg13g2_decap_8 FILLER_73_1554 ();
 sg13g2_decap_8 FILLER_73_1561 ();
 sg13g2_decap_8 FILLER_73_1568 ();
 sg13g2_decap_8 FILLER_73_1575 ();
 sg13g2_decap_8 FILLER_73_1582 ();
 sg13g2_decap_8 FILLER_73_1589 ();
 sg13g2_decap_8 FILLER_73_1596 ();
 sg13g2_decap_8 FILLER_73_1603 ();
 sg13g2_decap_8 FILLER_73_1610 ();
 sg13g2_decap_8 FILLER_73_1617 ();
 sg13g2_decap_8 FILLER_73_1624 ();
 sg13g2_decap_8 FILLER_73_1631 ();
 sg13g2_decap_8 FILLER_73_1638 ();
 sg13g2_decap_8 FILLER_73_1645 ();
 sg13g2_decap_8 FILLER_73_1652 ();
 sg13g2_decap_8 FILLER_73_1659 ();
 sg13g2_decap_8 FILLER_73_1666 ();
 sg13g2_decap_8 FILLER_73_1673 ();
 sg13g2_decap_8 FILLER_73_1680 ();
 sg13g2_decap_8 FILLER_73_1687 ();
 sg13g2_decap_8 FILLER_73_1694 ();
 sg13g2_decap_8 FILLER_73_1701 ();
 sg13g2_decap_8 FILLER_73_1708 ();
 sg13g2_decap_8 FILLER_73_1715 ();
 sg13g2_decap_8 FILLER_73_1722 ();
 sg13g2_decap_8 FILLER_73_1729 ();
 sg13g2_decap_8 FILLER_73_1736 ();
 sg13g2_decap_8 FILLER_73_1743 ();
 sg13g2_decap_8 FILLER_73_1750 ();
 sg13g2_decap_8 FILLER_73_1757 ();
 sg13g2_decap_4 FILLER_73_1764 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_decap_8 FILLER_74_175 ();
 sg13g2_decap_8 FILLER_74_182 ();
 sg13g2_decap_8 FILLER_74_189 ();
 sg13g2_decap_8 FILLER_74_196 ();
 sg13g2_decap_8 FILLER_74_203 ();
 sg13g2_decap_8 FILLER_74_210 ();
 sg13g2_decap_8 FILLER_74_217 ();
 sg13g2_decap_8 FILLER_74_224 ();
 sg13g2_decap_8 FILLER_74_231 ();
 sg13g2_decap_8 FILLER_74_238 ();
 sg13g2_decap_8 FILLER_74_245 ();
 sg13g2_decap_4 FILLER_74_252 ();
 sg13g2_fill_1 FILLER_74_256 ();
 sg13g2_fill_2 FILLER_74_283 ();
 sg13g2_decap_4 FILLER_74_298 ();
 sg13g2_fill_1 FILLER_74_311 ();
 sg13g2_decap_8 FILLER_74_316 ();
 sg13g2_decap_8 FILLER_74_323 ();
 sg13g2_fill_2 FILLER_74_330 ();
 sg13g2_fill_2 FILLER_74_345 ();
 sg13g2_fill_2 FILLER_74_373 ();
 sg13g2_fill_1 FILLER_74_431 ();
 sg13g2_decap_8 FILLER_74_445 ();
 sg13g2_decap_8 FILLER_74_452 ();
 sg13g2_decap_4 FILLER_74_459 ();
 sg13g2_fill_2 FILLER_74_463 ();
 sg13g2_fill_1 FILLER_74_491 ();
 sg13g2_fill_2 FILLER_74_512 ();
 sg13g2_fill_2 FILLER_74_532 ();
 sg13g2_decap_8 FILLER_74_554 ();
 sg13g2_decap_4 FILLER_74_561 ();
 sg13g2_fill_1 FILLER_74_565 ();
 sg13g2_fill_1 FILLER_74_599 ();
 sg13g2_fill_1 FILLER_74_624 ();
 sg13g2_fill_1 FILLER_74_645 ();
 sg13g2_decap_8 FILLER_74_682 ();
 sg13g2_fill_1 FILLER_74_689 ();
 sg13g2_decap_4 FILLER_74_694 ();
 sg13g2_fill_1 FILLER_74_698 ();
 sg13g2_fill_2 FILLER_74_716 ();
 sg13g2_fill_1 FILLER_74_727 ();
 sg13g2_fill_1 FILLER_74_738 ();
 sg13g2_fill_2 FILLER_74_770 ();
 sg13g2_fill_1 FILLER_74_772 ();
 sg13g2_decap_8 FILLER_74_791 ();
 sg13g2_fill_2 FILLER_74_798 ();
 sg13g2_fill_2 FILLER_74_842 ();
 sg13g2_fill_1 FILLER_74_844 ();
 sg13g2_fill_1 FILLER_74_873 ();
 sg13g2_fill_2 FILLER_74_889 ();
 sg13g2_decap_8 FILLER_74_912 ();
 sg13g2_decap_4 FILLER_74_919 ();
 sg13g2_fill_1 FILLER_74_923 ();
 sg13g2_decap_8 FILLER_74_941 ();
 sg13g2_decap_8 FILLER_74_948 ();
 sg13g2_decap_4 FILLER_74_961 ();
 sg13g2_fill_1 FILLER_74_965 ();
 sg13g2_decap_4 FILLER_74_975 ();
 sg13g2_fill_2 FILLER_74_979 ();
 sg13g2_decap_8 FILLER_74_1028 ();
 sg13g2_fill_2 FILLER_74_1035 ();
 sg13g2_decap_8 FILLER_74_1049 ();
 sg13g2_decap_8 FILLER_74_1056 ();
 sg13g2_decap_8 FILLER_74_1063 ();
 sg13g2_decap_8 FILLER_74_1070 ();
 sg13g2_decap_8 FILLER_74_1077 ();
 sg13g2_decap_8 FILLER_74_1084 ();
 sg13g2_decap_8 FILLER_74_1091 ();
 sg13g2_decap_8 FILLER_74_1098 ();
 sg13g2_decap_8 FILLER_74_1105 ();
 sg13g2_decap_8 FILLER_74_1112 ();
 sg13g2_decap_8 FILLER_74_1119 ();
 sg13g2_decap_8 FILLER_74_1126 ();
 sg13g2_decap_8 FILLER_74_1133 ();
 sg13g2_decap_8 FILLER_74_1140 ();
 sg13g2_decap_8 FILLER_74_1147 ();
 sg13g2_decap_8 FILLER_74_1154 ();
 sg13g2_decap_8 FILLER_74_1161 ();
 sg13g2_decap_8 FILLER_74_1168 ();
 sg13g2_decap_8 FILLER_74_1175 ();
 sg13g2_decap_8 FILLER_74_1182 ();
 sg13g2_decap_8 FILLER_74_1189 ();
 sg13g2_decap_8 FILLER_74_1196 ();
 sg13g2_decap_8 FILLER_74_1203 ();
 sg13g2_decap_8 FILLER_74_1210 ();
 sg13g2_decap_8 FILLER_74_1217 ();
 sg13g2_decap_8 FILLER_74_1224 ();
 sg13g2_decap_8 FILLER_74_1231 ();
 sg13g2_decap_8 FILLER_74_1238 ();
 sg13g2_decap_8 FILLER_74_1245 ();
 sg13g2_decap_8 FILLER_74_1252 ();
 sg13g2_decap_8 FILLER_74_1259 ();
 sg13g2_decap_8 FILLER_74_1266 ();
 sg13g2_decap_8 FILLER_74_1273 ();
 sg13g2_decap_8 FILLER_74_1280 ();
 sg13g2_decap_8 FILLER_74_1287 ();
 sg13g2_decap_8 FILLER_74_1294 ();
 sg13g2_decap_8 FILLER_74_1301 ();
 sg13g2_decap_8 FILLER_74_1308 ();
 sg13g2_decap_8 FILLER_74_1315 ();
 sg13g2_decap_8 FILLER_74_1322 ();
 sg13g2_decap_8 FILLER_74_1329 ();
 sg13g2_decap_8 FILLER_74_1336 ();
 sg13g2_decap_8 FILLER_74_1343 ();
 sg13g2_decap_8 FILLER_74_1350 ();
 sg13g2_decap_8 FILLER_74_1357 ();
 sg13g2_decap_8 FILLER_74_1364 ();
 sg13g2_decap_8 FILLER_74_1371 ();
 sg13g2_decap_8 FILLER_74_1378 ();
 sg13g2_decap_8 FILLER_74_1385 ();
 sg13g2_decap_8 FILLER_74_1392 ();
 sg13g2_decap_8 FILLER_74_1399 ();
 sg13g2_decap_8 FILLER_74_1406 ();
 sg13g2_decap_8 FILLER_74_1413 ();
 sg13g2_decap_8 FILLER_74_1420 ();
 sg13g2_decap_8 FILLER_74_1427 ();
 sg13g2_decap_8 FILLER_74_1434 ();
 sg13g2_decap_8 FILLER_74_1441 ();
 sg13g2_decap_8 FILLER_74_1448 ();
 sg13g2_decap_8 FILLER_74_1455 ();
 sg13g2_decap_8 FILLER_74_1462 ();
 sg13g2_decap_8 FILLER_74_1469 ();
 sg13g2_decap_8 FILLER_74_1476 ();
 sg13g2_decap_8 FILLER_74_1483 ();
 sg13g2_decap_8 FILLER_74_1490 ();
 sg13g2_decap_8 FILLER_74_1497 ();
 sg13g2_decap_8 FILLER_74_1504 ();
 sg13g2_decap_8 FILLER_74_1511 ();
 sg13g2_decap_8 FILLER_74_1518 ();
 sg13g2_decap_8 FILLER_74_1525 ();
 sg13g2_decap_8 FILLER_74_1532 ();
 sg13g2_decap_8 FILLER_74_1539 ();
 sg13g2_decap_8 FILLER_74_1546 ();
 sg13g2_decap_8 FILLER_74_1553 ();
 sg13g2_decap_8 FILLER_74_1560 ();
 sg13g2_decap_8 FILLER_74_1567 ();
 sg13g2_decap_8 FILLER_74_1574 ();
 sg13g2_decap_8 FILLER_74_1581 ();
 sg13g2_decap_8 FILLER_74_1588 ();
 sg13g2_decap_8 FILLER_74_1595 ();
 sg13g2_decap_8 FILLER_74_1602 ();
 sg13g2_decap_8 FILLER_74_1609 ();
 sg13g2_decap_8 FILLER_74_1616 ();
 sg13g2_decap_8 FILLER_74_1623 ();
 sg13g2_decap_8 FILLER_74_1630 ();
 sg13g2_decap_8 FILLER_74_1637 ();
 sg13g2_decap_8 FILLER_74_1644 ();
 sg13g2_decap_8 FILLER_74_1651 ();
 sg13g2_decap_8 FILLER_74_1658 ();
 sg13g2_decap_8 FILLER_74_1665 ();
 sg13g2_decap_8 FILLER_74_1672 ();
 sg13g2_decap_8 FILLER_74_1679 ();
 sg13g2_decap_8 FILLER_74_1686 ();
 sg13g2_decap_8 FILLER_74_1693 ();
 sg13g2_decap_8 FILLER_74_1700 ();
 sg13g2_decap_8 FILLER_74_1707 ();
 sg13g2_decap_8 FILLER_74_1714 ();
 sg13g2_decap_8 FILLER_74_1721 ();
 sg13g2_decap_8 FILLER_74_1728 ();
 sg13g2_decap_8 FILLER_74_1735 ();
 sg13g2_decap_8 FILLER_74_1742 ();
 sg13g2_decap_8 FILLER_74_1749 ();
 sg13g2_decap_8 FILLER_74_1756 ();
 sg13g2_decap_4 FILLER_74_1763 ();
 sg13g2_fill_1 FILLER_74_1767 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_8 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_196 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_224 ();
 sg13g2_decap_8 FILLER_75_231 ();
 sg13g2_decap_8 FILLER_75_238 ();
 sg13g2_decap_8 FILLER_75_245 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_decap_8 FILLER_75_259 ();
 sg13g2_decap_8 FILLER_75_266 ();
 sg13g2_decap_8 FILLER_75_273 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_decap_8 FILLER_75_287 ();
 sg13g2_decap_8 FILLER_75_294 ();
 sg13g2_decap_8 FILLER_75_301 ();
 sg13g2_decap_8 FILLER_75_308 ();
 sg13g2_decap_8 FILLER_75_315 ();
 sg13g2_decap_8 FILLER_75_322 ();
 sg13g2_fill_2 FILLER_75_329 ();
 sg13g2_fill_1 FILLER_75_331 ();
 sg13g2_decap_8 FILLER_75_345 ();
 sg13g2_decap_8 FILLER_75_352 ();
 sg13g2_decap_4 FILLER_75_359 ();
 sg13g2_fill_1 FILLER_75_389 ();
 sg13g2_fill_2 FILLER_75_403 ();
 sg13g2_decap_8 FILLER_75_410 ();
 sg13g2_decap_8 FILLER_75_417 ();
 sg13g2_decap_8 FILLER_75_424 ();
 sg13g2_decap_8 FILLER_75_431 ();
 sg13g2_fill_1 FILLER_75_438 ();
 sg13g2_decap_8 FILLER_75_465 ();
 sg13g2_fill_2 FILLER_75_472 ();
 sg13g2_fill_1 FILLER_75_474 ();
 sg13g2_decap_8 FILLER_75_479 ();
 sg13g2_fill_1 FILLER_75_486 ();
 sg13g2_fill_1 FILLER_75_531 ();
 sg13g2_fill_1 FILLER_75_537 ();
 sg13g2_fill_2 FILLER_75_601 ();
 sg13g2_fill_2 FILLER_75_607 ();
 sg13g2_decap_4 FILLER_75_612 ();
 sg13g2_fill_1 FILLER_75_629 ();
 sg13g2_fill_1 FILLER_75_645 ();
 sg13g2_decap_4 FILLER_75_663 ();
 sg13g2_decap_8 FILLER_75_671 ();
 sg13g2_decap_8 FILLER_75_678 ();
 sg13g2_decap_8 FILLER_75_685 ();
 sg13g2_decap_4 FILLER_75_746 ();
 sg13g2_decap_8 FILLER_75_800 ();
 sg13g2_decap_4 FILLER_75_807 ();
 sg13g2_fill_2 FILLER_75_816 ();
 sg13g2_fill_1 FILLER_75_818 ();
 sg13g2_decap_8 FILLER_75_846 ();
 sg13g2_fill_1 FILLER_75_853 ();
 sg13g2_fill_1 FILLER_75_873 ();
 sg13g2_fill_2 FILLER_75_893 ();
 sg13g2_fill_1 FILLER_75_895 ();
 sg13g2_decap_8 FILLER_75_901 ();
 sg13g2_decap_8 FILLER_75_911 ();
 sg13g2_fill_1 FILLER_75_918 ();
 sg13g2_fill_1 FILLER_75_946 ();
 sg13g2_decap_8 FILLER_75_957 ();
 sg13g2_fill_1 FILLER_75_964 ();
 sg13g2_decap_8 FILLER_75_973 ();
 sg13g2_decap_4 FILLER_75_980 ();
 sg13g2_fill_2 FILLER_75_984 ();
 sg13g2_fill_2 FILLER_75_990 ();
 sg13g2_decap_8 FILLER_75_1002 ();
 sg13g2_decap_4 FILLER_75_1009 ();
 sg13g2_fill_2 FILLER_75_1013 ();
 sg13g2_decap_8 FILLER_75_1028 ();
 sg13g2_decap_8 FILLER_75_1052 ();
 sg13g2_decap_8 FILLER_75_1059 ();
 sg13g2_decap_8 FILLER_75_1066 ();
 sg13g2_decap_8 FILLER_75_1073 ();
 sg13g2_decap_8 FILLER_75_1080 ();
 sg13g2_decap_8 FILLER_75_1087 ();
 sg13g2_decap_8 FILLER_75_1094 ();
 sg13g2_decap_8 FILLER_75_1101 ();
 sg13g2_decap_8 FILLER_75_1108 ();
 sg13g2_decap_8 FILLER_75_1115 ();
 sg13g2_decap_8 FILLER_75_1122 ();
 sg13g2_decap_8 FILLER_75_1129 ();
 sg13g2_decap_8 FILLER_75_1136 ();
 sg13g2_decap_8 FILLER_75_1143 ();
 sg13g2_decap_8 FILLER_75_1150 ();
 sg13g2_decap_8 FILLER_75_1157 ();
 sg13g2_decap_8 FILLER_75_1164 ();
 sg13g2_decap_8 FILLER_75_1171 ();
 sg13g2_decap_8 FILLER_75_1178 ();
 sg13g2_decap_8 FILLER_75_1185 ();
 sg13g2_decap_8 FILLER_75_1192 ();
 sg13g2_decap_8 FILLER_75_1199 ();
 sg13g2_decap_8 FILLER_75_1206 ();
 sg13g2_decap_8 FILLER_75_1213 ();
 sg13g2_decap_8 FILLER_75_1220 ();
 sg13g2_decap_8 FILLER_75_1227 ();
 sg13g2_decap_8 FILLER_75_1234 ();
 sg13g2_decap_8 FILLER_75_1241 ();
 sg13g2_decap_8 FILLER_75_1248 ();
 sg13g2_decap_8 FILLER_75_1255 ();
 sg13g2_decap_8 FILLER_75_1262 ();
 sg13g2_decap_8 FILLER_75_1269 ();
 sg13g2_decap_8 FILLER_75_1276 ();
 sg13g2_decap_8 FILLER_75_1283 ();
 sg13g2_decap_8 FILLER_75_1290 ();
 sg13g2_decap_8 FILLER_75_1297 ();
 sg13g2_decap_8 FILLER_75_1304 ();
 sg13g2_decap_8 FILLER_75_1311 ();
 sg13g2_decap_8 FILLER_75_1318 ();
 sg13g2_decap_8 FILLER_75_1325 ();
 sg13g2_decap_8 FILLER_75_1332 ();
 sg13g2_decap_8 FILLER_75_1339 ();
 sg13g2_decap_8 FILLER_75_1346 ();
 sg13g2_decap_8 FILLER_75_1353 ();
 sg13g2_decap_8 FILLER_75_1360 ();
 sg13g2_decap_8 FILLER_75_1367 ();
 sg13g2_decap_8 FILLER_75_1374 ();
 sg13g2_decap_8 FILLER_75_1381 ();
 sg13g2_decap_8 FILLER_75_1388 ();
 sg13g2_decap_8 FILLER_75_1395 ();
 sg13g2_decap_8 FILLER_75_1402 ();
 sg13g2_decap_8 FILLER_75_1409 ();
 sg13g2_decap_8 FILLER_75_1416 ();
 sg13g2_decap_8 FILLER_75_1423 ();
 sg13g2_decap_8 FILLER_75_1430 ();
 sg13g2_decap_8 FILLER_75_1437 ();
 sg13g2_decap_8 FILLER_75_1444 ();
 sg13g2_decap_8 FILLER_75_1451 ();
 sg13g2_decap_8 FILLER_75_1458 ();
 sg13g2_decap_8 FILLER_75_1465 ();
 sg13g2_decap_8 FILLER_75_1472 ();
 sg13g2_decap_8 FILLER_75_1479 ();
 sg13g2_decap_8 FILLER_75_1486 ();
 sg13g2_decap_8 FILLER_75_1493 ();
 sg13g2_decap_8 FILLER_75_1500 ();
 sg13g2_decap_8 FILLER_75_1507 ();
 sg13g2_decap_8 FILLER_75_1514 ();
 sg13g2_decap_8 FILLER_75_1521 ();
 sg13g2_decap_8 FILLER_75_1528 ();
 sg13g2_decap_8 FILLER_75_1535 ();
 sg13g2_decap_8 FILLER_75_1542 ();
 sg13g2_decap_8 FILLER_75_1549 ();
 sg13g2_decap_8 FILLER_75_1556 ();
 sg13g2_decap_8 FILLER_75_1563 ();
 sg13g2_decap_8 FILLER_75_1570 ();
 sg13g2_decap_8 FILLER_75_1577 ();
 sg13g2_decap_8 FILLER_75_1584 ();
 sg13g2_decap_8 FILLER_75_1591 ();
 sg13g2_decap_8 FILLER_75_1598 ();
 sg13g2_decap_8 FILLER_75_1605 ();
 sg13g2_decap_8 FILLER_75_1612 ();
 sg13g2_decap_8 FILLER_75_1619 ();
 sg13g2_decap_8 FILLER_75_1626 ();
 sg13g2_decap_8 FILLER_75_1633 ();
 sg13g2_decap_8 FILLER_75_1640 ();
 sg13g2_decap_8 FILLER_75_1647 ();
 sg13g2_decap_8 FILLER_75_1654 ();
 sg13g2_decap_8 FILLER_75_1661 ();
 sg13g2_decap_8 FILLER_75_1668 ();
 sg13g2_decap_8 FILLER_75_1675 ();
 sg13g2_decap_8 FILLER_75_1682 ();
 sg13g2_decap_8 FILLER_75_1689 ();
 sg13g2_decap_8 FILLER_75_1696 ();
 sg13g2_decap_8 FILLER_75_1703 ();
 sg13g2_decap_8 FILLER_75_1710 ();
 sg13g2_decap_8 FILLER_75_1717 ();
 sg13g2_decap_8 FILLER_75_1724 ();
 sg13g2_decap_8 FILLER_75_1731 ();
 sg13g2_decap_8 FILLER_75_1738 ();
 sg13g2_decap_8 FILLER_75_1745 ();
 sg13g2_decap_8 FILLER_75_1752 ();
 sg13g2_decap_8 FILLER_75_1759 ();
 sg13g2_fill_2 FILLER_75_1766 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_8 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_decap_8 FILLER_76_273 ();
 sg13g2_decap_8 FILLER_76_280 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_392 ();
 sg13g2_fill_2 FILLER_76_399 ();
 sg13g2_decap_4 FILLER_76_427 ();
 sg13g2_fill_1 FILLER_76_431 ();
 sg13g2_decap_8 FILLER_76_458 ();
 sg13g2_decap_4 FILLER_76_465 ();
 sg13g2_fill_2 FILLER_76_469 ();
 sg13g2_fill_2 FILLER_76_484 ();
 sg13g2_fill_1 FILLER_76_486 ();
 sg13g2_fill_2 FILLER_76_519 ();
 sg13g2_fill_2 FILLER_76_530 ();
 sg13g2_fill_1 FILLER_76_575 ();
 sg13g2_fill_2 FILLER_76_611 ();
 sg13g2_fill_1 FILLER_76_613 ();
 sg13g2_decap_4 FILLER_76_644 ();
 sg13g2_fill_2 FILLER_76_684 ();
 sg13g2_fill_1 FILLER_76_748 ();
 sg13g2_decap_4 FILLER_76_797 ();
 sg13g2_fill_1 FILLER_76_801 ();
 sg13g2_fill_1 FILLER_76_831 ();
 sg13g2_fill_1 FILLER_76_841 ();
 sg13g2_fill_1 FILLER_76_851 ();
 sg13g2_fill_2 FILLER_76_856 ();
 sg13g2_decap_4 FILLER_76_863 ();
 sg13g2_fill_1 FILLER_76_867 ();
 sg13g2_fill_2 FILLER_76_876 ();
 sg13g2_fill_1 FILLER_76_878 ();
 sg13g2_decap_8 FILLER_76_888 ();
 sg13g2_decap_8 FILLER_76_895 ();
 sg13g2_fill_1 FILLER_76_902 ();
 sg13g2_decap_8 FILLER_76_923 ();
 sg13g2_fill_1 FILLER_76_930 ();
 sg13g2_decap_8 FILLER_76_939 ();
 sg13g2_decap_4 FILLER_76_957 ();
 sg13g2_fill_2 FILLER_76_964 ();
 sg13g2_decap_8 FILLER_76_983 ();
 sg13g2_fill_2 FILLER_76_990 ();
 sg13g2_fill_1 FILLER_76_996 ();
 sg13g2_fill_1 FILLER_76_1010 ();
 sg13g2_fill_1 FILLER_76_1017 ();
 sg13g2_fill_2 FILLER_76_1028 ();
 sg13g2_fill_1 FILLER_76_1030 ();
 sg13g2_decap_8 FILLER_76_1052 ();
 sg13g2_decap_8 FILLER_76_1059 ();
 sg13g2_decap_8 FILLER_76_1066 ();
 sg13g2_decap_8 FILLER_76_1073 ();
 sg13g2_decap_8 FILLER_76_1080 ();
 sg13g2_decap_8 FILLER_76_1087 ();
 sg13g2_decap_8 FILLER_76_1094 ();
 sg13g2_decap_8 FILLER_76_1101 ();
 sg13g2_decap_8 FILLER_76_1108 ();
 sg13g2_decap_8 FILLER_76_1115 ();
 sg13g2_decap_8 FILLER_76_1122 ();
 sg13g2_decap_8 FILLER_76_1129 ();
 sg13g2_decap_8 FILLER_76_1136 ();
 sg13g2_decap_8 FILLER_76_1143 ();
 sg13g2_decap_8 FILLER_76_1150 ();
 sg13g2_decap_8 FILLER_76_1157 ();
 sg13g2_decap_8 FILLER_76_1164 ();
 sg13g2_decap_8 FILLER_76_1171 ();
 sg13g2_decap_8 FILLER_76_1178 ();
 sg13g2_decap_8 FILLER_76_1185 ();
 sg13g2_decap_8 FILLER_76_1192 ();
 sg13g2_decap_8 FILLER_76_1199 ();
 sg13g2_decap_8 FILLER_76_1206 ();
 sg13g2_decap_8 FILLER_76_1213 ();
 sg13g2_decap_8 FILLER_76_1220 ();
 sg13g2_decap_8 FILLER_76_1227 ();
 sg13g2_decap_8 FILLER_76_1234 ();
 sg13g2_decap_8 FILLER_76_1241 ();
 sg13g2_decap_8 FILLER_76_1248 ();
 sg13g2_decap_8 FILLER_76_1255 ();
 sg13g2_decap_8 FILLER_76_1262 ();
 sg13g2_decap_8 FILLER_76_1269 ();
 sg13g2_decap_8 FILLER_76_1276 ();
 sg13g2_decap_8 FILLER_76_1283 ();
 sg13g2_decap_8 FILLER_76_1290 ();
 sg13g2_decap_8 FILLER_76_1297 ();
 sg13g2_decap_8 FILLER_76_1304 ();
 sg13g2_decap_8 FILLER_76_1311 ();
 sg13g2_decap_8 FILLER_76_1318 ();
 sg13g2_decap_8 FILLER_76_1325 ();
 sg13g2_decap_8 FILLER_76_1332 ();
 sg13g2_decap_8 FILLER_76_1339 ();
 sg13g2_decap_8 FILLER_76_1346 ();
 sg13g2_decap_8 FILLER_76_1353 ();
 sg13g2_decap_8 FILLER_76_1360 ();
 sg13g2_decap_8 FILLER_76_1367 ();
 sg13g2_decap_8 FILLER_76_1374 ();
 sg13g2_decap_8 FILLER_76_1381 ();
 sg13g2_decap_8 FILLER_76_1388 ();
 sg13g2_decap_8 FILLER_76_1395 ();
 sg13g2_decap_8 FILLER_76_1402 ();
 sg13g2_decap_8 FILLER_76_1409 ();
 sg13g2_decap_8 FILLER_76_1416 ();
 sg13g2_decap_8 FILLER_76_1423 ();
 sg13g2_decap_8 FILLER_76_1430 ();
 sg13g2_decap_8 FILLER_76_1437 ();
 sg13g2_decap_8 FILLER_76_1444 ();
 sg13g2_decap_8 FILLER_76_1451 ();
 sg13g2_decap_8 FILLER_76_1458 ();
 sg13g2_decap_8 FILLER_76_1465 ();
 sg13g2_decap_8 FILLER_76_1472 ();
 sg13g2_decap_8 FILLER_76_1479 ();
 sg13g2_decap_8 FILLER_76_1486 ();
 sg13g2_decap_8 FILLER_76_1493 ();
 sg13g2_decap_8 FILLER_76_1500 ();
 sg13g2_decap_8 FILLER_76_1507 ();
 sg13g2_decap_8 FILLER_76_1514 ();
 sg13g2_decap_8 FILLER_76_1521 ();
 sg13g2_decap_8 FILLER_76_1528 ();
 sg13g2_decap_8 FILLER_76_1535 ();
 sg13g2_decap_8 FILLER_76_1542 ();
 sg13g2_decap_8 FILLER_76_1549 ();
 sg13g2_decap_8 FILLER_76_1556 ();
 sg13g2_decap_8 FILLER_76_1563 ();
 sg13g2_decap_8 FILLER_76_1570 ();
 sg13g2_decap_8 FILLER_76_1577 ();
 sg13g2_decap_8 FILLER_76_1584 ();
 sg13g2_decap_8 FILLER_76_1591 ();
 sg13g2_decap_8 FILLER_76_1598 ();
 sg13g2_decap_8 FILLER_76_1605 ();
 sg13g2_decap_8 FILLER_76_1612 ();
 sg13g2_decap_8 FILLER_76_1619 ();
 sg13g2_decap_8 FILLER_76_1626 ();
 sg13g2_decap_8 FILLER_76_1633 ();
 sg13g2_decap_8 FILLER_76_1640 ();
 sg13g2_decap_8 FILLER_76_1647 ();
 sg13g2_decap_8 FILLER_76_1654 ();
 sg13g2_decap_8 FILLER_76_1661 ();
 sg13g2_decap_8 FILLER_76_1668 ();
 sg13g2_decap_8 FILLER_76_1675 ();
 sg13g2_decap_8 FILLER_76_1682 ();
 sg13g2_decap_8 FILLER_76_1689 ();
 sg13g2_decap_8 FILLER_76_1696 ();
 sg13g2_decap_8 FILLER_76_1703 ();
 sg13g2_decap_8 FILLER_76_1710 ();
 sg13g2_decap_8 FILLER_76_1717 ();
 sg13g2_decap_8 FILLER_76_1724 ();
 sg13g2_decap_8 FILLER_76_1731 ();
 sg13g2_decap_8 FILLER_76_1738 ();
 sg13g2_decap_8 FILLER_76_1745 ();
 sg13g2_decap_8 FILLER_76_1752 ();
 sg13g2_decap_8 FILLER_76_1759 ();
 sg13g2_fill_2 FILLER_76_1766 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_8 FILLER_77_245 ();
 sg13g2_decap_8 FILLER_77_252 ();
 sg13g2_decap_8 FILLER_77_259 ();
 sg13g2_decap_8 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_273 ();
 sg13g2_decap_8 FILLER_77_280 ();
 sg13g2_decap_8 FILLER_77_287 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_decap_8 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_364 ();
 sg13g2_decap_8 FILLER_77_371 ();
 sg13g2_fill_2 FILLER_77_378 ();
 sg13g2_fill_1 FILLER_77_380 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_decap_4 FILLER_77_492 ();
 sg13g2_fill_2 FILLER_77_526 ();
 sg13g2_fill_2 FILLER_77_558 ();
 sg13g2_fill_1 FILLER_77_568 ();
 sg13g2_fill_2 FILLER_77_595 ();
 sg13g2_fill_1 FILLER_77_597 ();
 sg13g2_fill_1 FILLER_77_607 ();
 sg13g2_fill_2 FILLER_77_673 ();
 sg13g2_fill_1 FILLER_77_675 ();
 sg13g2_fill_1 FILLER_77_702 ();
 sg13g2_decap_4 FILLER_77_770 ();
 sg13g2_decap_4 FILLER_77_800 ();
 sg13g2_fill_2 FILLER_77_828 ();
 sg13g2_fill_1 FILLER_77_849 ();
 sg13g2_fill_1 FILLER_77_882 ();
 sg13g2_decap_4 FILLER_77_904 ();
 sg13g2_fill_1 FILLER_77_934 ();
 sg13g2_decap_8 FILLER_77_960 ();
 sg13g2_decap_8 FILLER_77_980 ();
 sg13g2_decap_4 FILLER_77_987 ();
 sg13g2_fill_1 FILLER_77_991 ();
 sg13g2_fill_1 FILLER_77_1007 ();
 sg13g2_fill_1 FILLER_77_1033 ();
 sg13g2_decap_8 FILLER_77_1054 ();
 sg13g2_decap_8 FILLER_77_1061 ();
 sg13g2_decap_8 FILLER_77_1068 ();
 sg13g2_decap_8 FILLER_77_1075 ();
 sg13g2_decap_8 FILLER_77_1082 ();
 sg13g2_decap_8 FILLER_77_1089 ();
 sg13g2_decap_8 FILLER_77_1096 ();
 sg13g2_decap_8 FILLER_77_1103 ();
 sg13g2_decap_8 FILLER_77_1110 ();
 sg13g2_decap_8 FILLER_77_1117 ();
 sg13g2_decap_8 FILLER_77_1124 ();
 sg13g2_decap_8 FILLER_77_1131 ();
 sg13g2_decap_8 FILLER_77_1138 ();
 sg13g2_decap_8 FILLER_77_1145 ();
 sg13g2_decap_8 FILLER_77_1152 ();
 sg13g2_decap_8 FILLER_77_1159 ();
 sg13g2_decap_8 FILLER_77_1166 ();
 sg13g2_decap_8 FILLER_77_1173 ();
 sg13g2_decap_8 FILLER_77_1180 ();
 sg13g2_decap_8 FILLER_77_1187 ();
 sg13g2_decap_8 FILLER_77_1194 ();
 sg13g2_decap_8 FILLER_77_1201 ();
 sg13g2_decap_8 FILLER_77_1208 ();
 sg13g2_decap_8 FILLER_77_1215 ();
 sg13g2_decap_8 FILLER_77_1222 ();
 sg13g2_decap_8 FILLER_77_1229 ();
 sg13g2_decap_8 FILLER_77_1236 ();
 sg13g2_decap_8 FILLER_77_1243 ();
 sg13g2_decap_8 FILLER_77_1250 ();
 sg13g2_decap_8 FILLER_77_1257 ();
 sg13g2_decap_8 FILLER_77_1264 ();
 sg13g2_decap_8 FILLER_77_1271 ();
 sg13g2_decap_8 FILLER_77_1278 ();
 sg13g2_decap_8 FILLER_77_1285 ();
 sg13g2_decap_8 FILLER_77_1292 ();
 sg13g2_decap_8 FILLER_77_1299 ();
 sg13g2_decap_8 FILLER_77_1306 ();
 sg13g2_decap_8 FILLER_77_1313 ();
 sg13g2_decap_8 FILLER_77_1320 ();
 sg13g2_decap_8 FILLER_77_1327 ();
 sg13g2_decap_8 FILLER_77_1334 ();
 sg13g2_decap_8 FILLER_77_1341 ();
 sg13g2_decap_8 FILLER_77_1348 ();
 sg13g2_decap_8 FILLER_77_1355 ();
 sg13g2_decap_8 FILLER_77_1362 ();
 sg13g2_decap_8 FILLER_77_1369 ();
 sg13g2_decap_8 FILLER_77_1376 ();
 sg13g2_decap_8 FILLER_77_1383 ();
 sg13g2_decap_8 FILLER_77_1390 ();
 sg13g2_decap_8 FILLER_77_1397 ();
 sg13g2_decap_8 FILLER_77_1404 ();
 sg13g2_decap_8 FILLER_77_1411 ();
 sg13g2_decap_8 FILLER_77_1418 ();
 sg13g2_decap_8 FILLER_77_1425 ();
 sg13g2_decap_8 FILLER_77_1432 ();
 sg13g2_decap_8 FILLER_77_1439 ();
 sg13g2_decap_8 FILLER_77_1446 ();
 sg13g2_decap_8 FILLER_77_1453 ();
 sg13g2_decap_8 FILLER_77_1460 ();
 sg13g2_decap_8 FILLER_77_1467 ();
 sg13g2_decap_8 FILLER_77_1474 ();
 sg13g2_decap_8 FILLER_77_1481 ();
 sg13g2_decap_8 FILLER_77_1488 ();
 sg13g2_decap_8 FILLER_77_1495 ();
 sg13g2_decap_8 FILLER_77_1502 ();
 sg13g2_decap_8 FILLER_77_1509 ();
 sg13g2_decap_8 FILLER_77_1516 ();
 sg13g2_decap_8 FILLER_77_1523 ();
 sg13g2_decap_8 FILLER_77_1530 ();
 sg13g2_decap_8 FILLER_77_1537 ();
 sg13g2_decap_8 FILLER_77_1544 ();
 sg13g2_decap_8 FILLER_77_1551 ();
 sg13g2_decap_8 FILLER_77_1558 ();
 sg13g2_decap_8 FILLER_77_1565 ();
 sg13g2_decap_8 FILLER_77_1572 ();
 sg13g2_decap_8 FILLER_77_1579 ();
 sg13g2_decap_8 FILLER_77_1586 ();
 sg13g2_decap_8 FILLER_77_1593 ();
 sg13g2_decap_8 FILLER_77_1600 ();
 sg13g2_decap_8 FILLER_77_1607 ();
 sg13g2_decap_8 FILLER_77_1614 ();
 sg13g2_decap_8 FILLER_77_1621 ();
 sg13g2_decap_8 FILLER_77_1628 ();
 sg13g2_decap_8 FILLER_77_1635 ();
 sg13g2_decap_8 FILLER_77_1642 ();
 sg13g2_decap_8 FILLER_77_1649 ();
 sg13g2_decap_8 FILLER_77_1656 ();
 sg13g2_decap_8 FILLER_77_1663 ();
 sg13g2_decap_8 FILLER_77_1670 ();
 sg13g2_decap_8 FILLER_77_1677 ();
 sg13g2_decap_8 FILLER_77_1684 ();
 sg13g2_decap_8 FILLER_77_1691 ();
 sg13g2_decap_8 FILLER_77_1698 ();
 sg13g2_decap_8 FILLER_77_1705 ();
 sg13g2_decap_8 FILLER_77_1712 ();
 sg13g2_decap_8 FILLER_77_1719 ();
 sg13g2_decap_8 FILLER_77_1726 ();
 sg13g2_decap_8 FILLER_77_1733 ();
 sg13g2_decap_8 FILLER_77_1740 ();
 sg13g2_decap_8 FILLER_77_1747 ();
 sg13g2_decap_8 FILLER_77_1754 ();
 sg13g2_decap_8 FILLER_77_1761 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_decap_8 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_259 ();
 sg13g2_decap_8 FILLER_78_266 ();
 sg13g2_decap_8 FILLER_78_273 ();
 sg13g2_decap_8 FILLER_78_280 ();
 sg13g2_decap_8 FILLER_78_287 ();
 sg13g2_decap_8 FILLER_78_294 ();
 sg13g2_decap_8 FILLER_78_301 ();
 sg13g2_decap_8 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_decap_8 FILLER_78_322 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_357 ();
 sg13g2_decap_8 FILLER_78_364 ();
 sg13g2_decap_8 FILLER_78_371 ();
 sg13g2_decap_8 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_decap_8 FILLER_78_406 ();
 sg13g2_decap_8 FILLER_78_413 ();
 sg13g2_decap_8 FILLER_78_420 ();
 sg13g2_decap_8 FILLER_78_427 ();
 sg13g2_decap_8 FILLER_78_434 ();
 sg13g2_decap_8 FILLER_78_441 ();
 sg13g2_decap_8 FILLER_78_448 ();
 sg13g2_decap_8 FILLER_78_455 ();
 sg13g2_decap_8 FILLER_78_462 ();
 sg13g2_decap_8 FILLER_78_469 ();
 sg13g2_fill_2 FILLER_78_476 ();
 sg13g2_decap_8 FILLER_78_495 ();
 sg13g2_decap_8 FILLER_78_572 ();
 sg13g2_fill_1 FILLER_78_579 ();
 sg13g2_fill_2 FILLER_78_584 ();
 sg13g2_fill_1 FILLER_78_621 ();
 sg13g2_fill_1 FILLER_78_626 ();
 sg13g2_decap_8 FILLER_78_636 ();
 sg13g2_fill_1 FILLER_78_643 ();
 sg13g2_decap_8 FILLER_78_657 ();
 sg13g2_decap_4 FILLER_78_664 ();
 sg13g2_fill_2 FILLER_78_668 ();
 sg13g2_decap_8 FILLER_78_675 ();
 sg13g2_decap_8 FILLER_78_682 ();
 sg13g2_decap_8 FILLER_78_689 ();
 sg13g2_fill_2 FILLER_78_696 ();
 sg13g2_decap_4 FILLER_78_724 ();
 sg13g2_fill_1 FILLER_78_728 ();
 sg13g2_decap_8 FILLER_78_738 ();
 sg13g2_fill_2 FILLER_78_758 ();
 sg13g2_fill_1 FILLER_78_760 ();
 sg13g2_decap_8 FILLER_78_796 ();
 sg13g2_fill_2 FILLER_78_803 ();
 sg13g2_fill_1 FILLER_78_815 ();
 sg13g2_decap_8 FILLER_78_826 ();
 sg13g2_fill_2 FILLER_78_833 ();
 sg13g2_fill_2 FILLER_78_839 ();
 sg13g2_fill_1 FILLER_78_841 ();
 sg13g2_decap_8 FILLER_78_851 ();
 sg13g2_fill_1 FILLER_78_863 ();
 sg13g2_decap_4 FILLER_78_869 ();
 sg13g2_fill_1 FILLER_78_873 ();
 sg13g2_fill_1 FILLER_78_882 ();
 sg13g2_decap_8 FILLER_78_895 ();
 sg13g2_decap_4 FILLER_78_902 ();
 sg13g2_fill_1 FILLER_78_906 ();
 sg13g2_decap_4 FILLER_78_932 ();
 sg13g2_fill_2 FILLER_78_936 ();
 sg13g2_fill_2 FILLER_78_958 ();
 sg13g2_fill_1 FILLER_78_960 ();
 sg13g2_decap_8 FILLER_78_1003 ();
 sg13g2_decap_4 FILLER_78_1010 ();
 sg13g2_fill_1 FILLER_78_1014 ();
 sg13g2_decap_8 FILLER_78_1033 ();
 sg13g2_decap_8 FILLER_78_1040 ();
 sg13g2_decap_8 FILLER_78_1047 ();
 sg13g2_decap_8 FILLER_78_1054 ();
 sg13g2_decap_8 FILLER_78_1061 ();
 sg13g2_decap_8 FILLER_78_1068 ();
 sg13g2_decap_8 FILLER_78_1075 ();
 sg13g2_decap_8 FILLER_78_1082 ();
 sg13g2_decap_8 FILLER_78_1089 ();
 sg13g2_decap_8 FILLER_78_1096 ();
 sg13g2_decap_8 FILLER_78_1103 ();
 sg13g2_decap_8 FILLER_78_1110 ();
 sg13g2_decap_8 FILLER_78_1117 ();
 sg13g2_decap_8 FILLER_78_1124 ();
 sg13g2_decap_8 FILLER_78_1131 ();
 sg13g2_decap_8 FILLER_78_1138 ();
 sg13g2_decap_8 FILLER_78_1145 ();
 sg13g2_decap_8 FILLER_78_1152 ();
 sg13g2_decap_8 FILLER_78_1159 ();
 sg13g2_decap_8 FILLER_78_1166 ();
 sg13g2_decap_8 FILLER_78_1173 ();
 sg13g2_decap_8 FILLER_78_1180 ();
 sg13g2_decap_8 FILLER_78_1187 ();
 sg13g2_decap_8 FILLER_78_1194 ();
 sg13g2_decap_8 FILLER_78_1201 ();
 sg13g2_decap_8 FILLER_78_1208 ();
 sg13g2_decap_8 FILLER_78_1215 ();
 sg13g2_decap_8 FILLER_78_1222 ();
 sg13g2_decap_8 FILLER_78_1229 ();
 sg13g2_decap_8 FILLER_78_1236 ();
 sg13g2_decap_8 FILLER_78_1243 ();
 sg13g2_decap_8 FILLER_78_1250 ();
 sg13g2_decap_8 FILLER_78_1257 ();
 sg13g2_decap_8 FILLER_78_1264 ();
 sg13g2_decap_8 FILLER_78_1271 ();
 sg13g2_decap_8 FILLER_78_1278 ();
 sg13g2_decap_8 FILLER_78_1285 ();
 sg13g2_decap_8 FILLER_78_1292 ();
 sg13g2_decap_8 FILLER_78_1299 ();
 sg13g2_decap_8 FILLER_78_1306 ();
 sg13g2_decap_8 FILLER_78_1313 ();
 sg13g2_decap_8 FILLER_78_1320 ();
 sg13g2_decap_8 FILLER_78_1327 ();
 sg13g2_decap_8 FILLER_78_1334 ();
 sg13g2_decap_8 FILLER_78_1341 ();
 sg13g2_decap_8 FILLER_78_1348 ();
 sg13g2_decap_8 FILLER_78_1355 ();
 sg13g2_decap_8 FILLER_78_1362 ();
 sg13g2_decap_8 FILLER_78_1369 ();
 sg13g2_decap_8 FILLER_78_1376 ();
 sg13g2_decap_8 FILLER_78_1383 ();
 sg13g2_decap_8 FILLER_78_1390 ();
 sg13g2_decap_8 FILLER_78_1397 ();
 sg13g2_decap_8 FILLER_78_1404 ();
 sg13g2_decap_8 FILLER_78_1411 ();
 sg13g2_decap_8 FILLER_78_1418 ();
 sg13g2_decap_8 FILLER_78_1425 ();
 sg13g2_decap_8 FILLER_78_1432 ();
 sg13g2_decap_8 FILLER_78_1439 ();
 sg13g2_decap_8 FILLER_78_1446 ();
 sg13g2_decap_8 FILLER_78_1453 ();
 sg13g2_decap_8 FILLER_78_1460 ();
 sg13g2_decap_8 FILLER_78_1467 ();
 sg13g2_decap_8 FILLER_78_1474 ();
 sg13g2_decap_8 FILLER_78_1481 ();
 sg13g2_decap_8 FILLER_78_1488 ();
 sg13g2_decap_8 FILLER_78_1495 ();
 sg13g2_decap_8 FILLER_78_1502 ();
 sg13g2_decap_8 FILLER_78_1509 ();
 sg13g2_decap_8 FILLER_78_1516 ();
 sg13g2_decap_8 FILLER_78_1523 ();
 sg13g2_decap_8 FILLER_78_1530 ();
 sg13g2_decap_8 FILLER_78_1537 ();
 sg13g2_decap_8 FILLER_78_1544 ();
 sg13g2_decap_8 FILLER_78_1551 ();
 sg13g2_decap_8 FILLER_78_1558 ();
 sg13g2_decap_8 FILLER_78_1565 ();
 sg13g2_decap_8 FILLER_78_1572 ();
 sg13g2_decap_8 FILLER_78_1579 ();
 sg13g2_decap_8 FILLER_78_1586 ();
 sg13g2_decap_8 FILLER_78_1593 ();
 sg13g2_decap_8 FILLER_78_1600 ();
 sg13g2_decap_8 FILLER_78_1607 ();
 sg13g2_decap_8 FILLER_78_1614 ();
 sg13g2_decap_8 FILLER_78_1621 ();
 sg13g2_decap_8 FILLER_78_1628 ();
 sg13g2_decap_8 FILLER_78_1635 ();
 sg13g2_decap_8 FILLER_78_1642 ();
 sg13g2_decap_8 FILLER_78_1649 ();
 sg13g2_decap_8 FILLER_78_1656 ();
 sg13g2_decap_8 FILLER_78_1663 ();
 sg13g2_decap_8 FILLER_78_1670 ();
 sg13g2_decap_8 FILLER_78_1677 ();
 sg13g2_decap_8 FILLER_78_1684 ();
 sg13g2_decap_8 FILLER_78_1691 ();
 sg13g2_decap_8 FILLER_78_1698 ();
 sg13g2_decap_8 FILLER_78_1705 ();
 sg13g2_decap_8 FILLER_78_1712 ();
 sg13g2_decap_8 FILLER_78_1719 ();
 sg13g2_decap_8 FILLER_78_1726 ();
 sg13g2_decap_8 FILLER_78_1733 ();
 sg13g2_decap_8 FILLER_78_1740 ();
 sg13g2_decap_8 FILLER_78_1747 ();
 sg13g2_decap_8 FILLER_78_1754 ();
 sg13g2_decap_8 FILLER_78_1761 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_decap_8 FILLER_79_245 ();
 sg13g2_decap_8 FILLER_79_252 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_decap_8 FILLER_79_266 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_decap_8 FILLER_79_280 ();
 sg13g2_decap_8 FILLER_79_287 ();
 sg13g2_decap_8 FILLER_79_294 ();
 sg13g2_decap_8 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_decap_8 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_79_329 ();
 sg13g2_decap_8 FILLER_79_336 ();
 sg13g2_decap_8 FILLER_79_343 ();
 sg13g2_decap_8 FILLER_79_350 ();
 sg13g2_decap_8 FILLER_79_357 ();
 sg13g2_decap_8 FILLER_79_364 ();
 sg13g2_decap_8 FILLER_79_371 ();
 sg13g2_decap_8 FILLER_79_378 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_decap_8 FILLER_79_406 ();
 sg13g2_decap_8 FILLER_79_413 ();
 sg13g2_decap_8 FILLER_79_420 ();
 sg13g2_decap_8 FILLER_79_427 ();
 sg13g2_decap_8 FILLER_79_434 ();
 sg13g2_decap_8 FILLER_79_441 ();
 sg13g2_decap_8 FILLER_79_448 ();
 sg13g2_decap_8 FILLER_79_455 ();
 sg13g2_decap_8 FILLER_79_462 ();
 sg13g2_decap_8 FILLER_79_469 ();
 sg13g2_decap_8 FILLER_79_476 ();
 sg13g2_decap_8 FILLER_79_483 ();
 sg13g2_decap_8 FILLER_79_490 ();
 sg13g2_decap_8 FILLER_79_497 ();
 sg13g2_decap_8 FILLER_79_504 ();
 sg13g2_fill_1 FILLER_79_511 ();
 sg13g2_fill_1 FILLER_79_521 ();
 sg13g2_fill_2 FILLER_79_535 ();
 sg13g2_fill_1 FILLER_79_537 ();
 sg13g2_decap_4 FILLER_79_543 ();
 sg13g2_fill_2 FILLER_79_547 ();
 sg13g2_decap_4 FILLER_79_553 ();
 sg13g2_fill_2 FILLER_79_557 ();
 sg13g2_fill_2 FILLER_79_608 ();
 sg13g2_fill_1 FILLER_79_610 ();
 sg13g2_decap_8 FILLER_79_637 ();
 sg13g2_decap_8 FILLER_79_644 ();
 sg13g2_decap_8 FILLER_79_651 ();
 sg13g2_decap_8 FILLER_79_658 ();
 sg13g2_decap_8 FILLER_79_665 ();
 sg13g2_decap_8 FILLER_79_672 ();
 sg13g2_decap_8 FILLER_79_679 ();
 sg13g2_decap_8 FILLER_79_686 ();
 sg13g2_decap_8 FILLER_79_693 ();
 sg13g2_decap_8 FILLER_79_700 ();
 sg13g2_fill_2 FILLER_79_707 ();
 sg13g2_decap_8 FILLER_79_713 ();
 sg13g2_decap_8 FILLER_79_720 ();
 sg13g2_fill_2 FILLER_79_727 ();
 sg13g2_decap_8 FILLER_79_755 ();
 sg13g2_fill_2 FILLER_79_762 ();
 sg13g2_fill_1 FILLER_79_764 ();
 sg13g2_fill_1 FILLER_79_819 ();
 sg13g2_fill_1 FILLER_79_846 ();
 sg13g2_fill_2 FILLER_79_871 ();
 sg13g2_fill_1 FILLER_79_873 ();
 sg13g2_fill_2 FILLER_79_882 ();
 sg13g2_fill_2 FILLER_79_985 ();
 sg13g2_fill_1 FILLER_79_987 ();
 sg13g2_fill_1 FILLER_79_1012 ();
 sg13g2_decap_8 FILLER_79_1037 ();
 sg13g2_decap_8 FILLER_79_1044 ();
 sg13g2_decap_8 FILLER_79_1051 ();
 sg13g2_decap_8 FILLER_79_1058 ();
 sg13g2_decap_8 FILLER_79_1065 ();
 sg13g2_decap_8 FILLER_79_1072 ();
 sg13g2_decap_8 FILLER_79_1079 ();
 sg13g2_decap_8 FILLER_79_1086 ();
 sg13g2_decap_8 FILLER_79_1093 ();
 sg13g2_decap_8 FILLER_79_1100 ();
 sg13g2_decap_8 FILLER_79_1107 ();
 sg13g2_decap_8 FILLER_79_1114 ();
 sg13g2_decap_8 FILLER_79_1121 ();
 sg13g2_decap_8 FILLER_79_1128 ();
 sg13g2_decap_8 FILLER_79_1135 ();
 sg13g2_decap_8 FILLER_79_1142 ();
 sg13g2_decap_8 FILLER_79_1149 ();
 sg13g2_decap_8 FILLER_79_1156 ();
 sg13g2_decap_8 FILLER_79_1163 ();
 sg13g2_decap_8 FILLER_79_1170 ();
 sg13g2_decap_8 FILLER_79_1177 ();
 sg13g2_decap_8 FILLER_79_1184 ();
 sg13g2_decap_8 FILLER_79_1191 ();
 sg13g2_decap_8 FILLER_79_1198 ();
 sg13g2_decap_8 FILLER_79_1205 ();
 sg13g2_decap_8 FILLER_79_1212 ();
 sg13g2_decap_8 FILLER_79_1219 ();
 sg13g2_decap_8 FILLER_79_1226 ();
 sg13g2_decap_8 FILLER_79_1233 ();
 sg13g2_decap_8 FILLER_79_1240 ();
 sg13g2_decap_8 FILLER_79_1247 ();
 sg13g2_decap_8 FILLER_79_1254 ();
 sg13g2_decap_8 FILLER_79_1261 ();
 sg13g2_decap_8 FILLER_79_1268 ();
 sg13g2_decap_8 FILLER_79_1275 ();
 sg13g2_decap_8 FILLER_79_1282 ();
 sg13g2_decap_8 FILLER_79_1289 ();
 sg13g2_decap_8 FILLER_79_1296 ();
 sg13g2_decap_8 FILLER_79_1303 ();
 sg13g2_decap_8 FILLER_79_1310 ();
 sg13g2_decap_8 FILLER_79_1317 ();
 sg13g2_decap_8 FILLER_79_1324 ();
 sg13g2_decap_8 FILLER_79_1331 ();
 sg13g2_decap_8 FILLER_79_1338 ();
 sg13g2_decap_8 FILLER_79_1345 ();
 sg13g2_decap_8 FILLER_79_1352 ();
 sg13g2_decap_8 FILLER_79_1359 ();
 sg13g2_decap_8 FILLER_79_1366 ();
 sg13g2_decap_8 FILLER_79_1373 ();
 sg13g2_decap_8 FILLER_79_1380 ();
 sg13g2_decap_8 FILLER_79_1387 ();
 sg13g2_decap_8 FILLER_79_1394 ();
 sg13g2_decap_8 FILLER_79_1401 ();
 sg13g2_decap_8 FILLER_79_1408 ();
 sg13g2_decap_8 FILLER_79_1415 ();
 sg13g2_decap_8 FILLER_79_1422 ();
 sg13g2_decap_8 FILLER_79_1429 ();
 sg13g2_decap_8 FILLER_79_1436 ();
 sg13g2_decap_8 FILLER_79_1443 ();
 sg13g2_decap_8 FILLER_79_1450 ();
 sg13g2_decap_8 FILLER_79_1457 ();
 sg13g2_decap_8 FILLER_79_1464 ();
 sg13g2_decap_8 FILLER_79_1471 ();
 sg13g2_decap_8 FILLER_79_1478 ();
 sg13g2_decap_8 FILLER_79_1485 ();
 sg13g2_decap_8 FILLER_79_1492 ();
 sg13g2_decap_8 FILLER_79_1499 ();
 sg13g2_decap_8 FILLER_79_1506 ();
 sg13g2_decap_8 FILLER_79_1513 ();
 sg13g2_decap_8 FILLER_79_1520 ();
 sg13g2_decap_8 FILLER_79_1527 ();
 sg13g2_decap_8 FILLER_79_1534 ();
 sg13g2_decap_8 FILLER_79_1541 ();
 sg13g2_decap_8 FILLER_79_1548 ();
 sg13g2_decap_8 FILLER_79_1555 ();
 sg13g2_decap_8 FILLER_79_1562 ();
 sg13g2_decap_8 FILLER_79_1569 ();
 sg13g2_decap_8 FILLER_79_1576 ();
 sg13g2_decap_8 FILLER_79_1583 ();
 sg13g2_decap_8 FILLER_79_1590 ();
 sg13g2_decap_8 FILLER_79_1597 ();
 sg13g2_decap_8 FILLER_79_1604 ();
 sg13g2_decap_8 FILLER_79_1611 ();
 sg13g2_decap_8 FILLER_79_1618 ();
 sg13g2_decap_8 FILLER_79_1625 ();
 sg13g2_decap_8 FILLER_79_1632 ();
 sg13g2_decap_8 FILLER_79_1639 ();
 sg13g2_decap_8 FILLER_79_1646 ();
 sg13g2_decap_8 FILLER_79_1653 ();
 sg13g2_decap_8 FILLER_79_1660 ();
 sg13g2_decap_8 FILLER_79_1667 ();
 sg13g2_decap_8 FILLER_79_1674 ();
 sg13g2_decap_8 FILLER_79_1681 ();
 sg13g2_decap_8 FILLER_79_1688 ();
 sg13g2_decap_8 FILLER_79_1695 ();
 sg13g2_decap_8 FILLER_79_1702 ();
 sg13g2_decap_8 FILLER_79_1709 ();
 sg13g2_decap_8 FILLER_79_1716 ();
 sg13g2_decap_8 FILLER_79_1723 ();
 sg13g2_decap_8 FILLER_79_1730 ();
 sg13g2_decap_8 FILLER_79_1737 ();
 sg13g2_decap_8 FILLER_79_1744 ();
 sg13g2_decap_8 FILLER_79_1751 ();
 sg13g2_decap_8 FILLER_79_1758 ();
 sg13g2_fill_2 FILLER_79_1765 ();
 sg13g2_fill_1 FILLER_79_1767 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_8 FILLER_80_229 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_decap_4 FILLER_80_243 ();
 sg13g2_fill_1 FILLER_80_247 ();
 sg13g2_decap_4 FILLER_80_252 ();
 sg13g2_decap_4 FILLER_80_260 ();
 sg13g2_decap_4 FILLER_80_268 ();
 sg13g2_decap_4 FILLER_80_276 ();
 sg13g2_decap_4 FILLER_80_284 ();
 sg13g2_decap_4 FILLER_80_292 ();
 sg13g2_decap_4 FILLER_80_300 ();
 sg13g2_decap_4 FILLER_80_308 ();
 sg13g2_decap_4 FILLER_80_316 ();
 sg13g2_decap_4 FILLER_80_324 ();
 sg13g2_decap_4 FILLER_80_332 ();
 sg13g2_decap_4 FILLER_80_340 ();
 sg13g2_decap_4 FILLER_80_348 ();
 sg13g2_decap_4 FILLER_80_356 ();
 sg13g2_decap_4 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_372 ();
 sg13g2_decap_8 FILLER_80_379 ();
 sg13g2_decap_8 FILLER_80_386 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_8 FILLER_80_400 ();
 sg13g2_decap_8 FILLER_80_407 ();
 sg13g2_decap_8 FILLER_80_414 ();
 sg13g2_decap_8 FILLER_80_421 ();
 sg13g2_decap_8 FILLER_80_428 ();
 sg13g2_decap_8 FILLER_80_435 ();
 sg13g2_decap_8 FILLER_80_442 ();
 sg13g2_decap_8 FILLER_80_449 ();
 sg13g2_decap_8 FILLER_80_456 ();
 sg13g2_decap_8 FILLER_80_463 ();
 sg13g2_decap_8 FILLER_80_470 ();
 sg13g2_decap_8 FILLER_80_477 ();
 sg13g2_decap_8 FILLER_80_484 ();
 sg13g2_decap_8 FILLER_80_491 ();
 sg13g2_decap_8 FILLER_80_498 ();
 sg13g2_decap_8 FILLER_80_505 ();
 sg13g2_decap_8 FILLER_80_512 ();
 sg13g2_decap_8 FILLER_80_519 ();
 sg13g2_decap_8 FILLER_80_526 ();
 sg13g2_decap_8 FILLER_80_533 ();
 sg13g2_decap_8 FILLER_80_540 ();
 sg13g2_decap_8 FILLER_80_547 ();
 sg13g2_decap_8 FILLER_80_554 ();
 sg13g2_decap_8 FILLER_80_561 ();
 sg13g2_decap_8 FILLER_80_568 ();
 sg13g2_decap_4 FILLER_80_575 ();
 sg13g2_fill_1 FILLER_80_579 ();
 sg13g2_decap_8 FILLER_80_593 ();
 sg13g2_decap_8 FILLER_80_600 ();
 sg13g2_decap_8 FILLER_80_607 ();
 sg13g2_decap_8 FILLER_80_614 ();
 sg13g2_decap_8 FILLER_80_634 ();
 sg13g2_decap_8 FILLER_80_641 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_669 ();
 sg13g2_decap_8 FILLER_80_676 ();
 sg13g2_decap_8 FILLER_80_683 ();
 sg13g2_decap_8 FILLER_80_690 ();
 sg13g2_decap_8 FILLER_80_697 ();
 sg13g2_decap_8 FILLER_80_704 ();
 sg13g2_decap_8 FILLER_80_711 ();
 sg13g2_decap_8 FILLER_80_718 ();
 sg13g2_decap_8 FILLER_80_725 ();
 sg13g2_decap_8 FILLER_80_732 ();
 sg13g2_fill_1 FILLER_80_739 ();
 sg13g2_decap_8 FILLER_80_744 ();
 sg13g2_decap_8 FILLER_80_751 ();
 sg13g2_decap_8 FILLER_80_758 ();
 sg13g2_decap_8 FILLER_80_765 ();
 sg13g2_decap_4 FILLER_80_772 ();
 sg13g2_fill_2 FILLER_80_776 ();
 sg13g2_decap_8 FILLER_80_786 ();
 sg13g2_fill_1 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_807 ();
 sg13g2_decap_8 FILLER_80_814 ();
 sg13g2_decap_4 FILLER_80_821 ();
 sg13g2_decap_8 FILLER_80_842 ();
 sg13g2_decap_8 FILLER_80_849 ();
 sg13g2_fill_1 FILLER_80_856 ();
 sg13g2_decap_8 FILLER_80_861 ();
 sg13g2_fill_2 FILLER_80_868 ();
 sg13g2_fill_1 FILLER_80_870 ();
 sg13g2_decap_4 FILLER_80_875 ();
 sg13g2_fill_1 FILLER_80_879 ();
 sg13g2_decap_8 FILLER_80_884 ();
 sg13g2_fill_1 FILLER_80_891 ();
 sg13g2_decap_8 FILLER_80_895 ();
 sg13g2_decap_4 FILLER_80_902 ();
 sg13g2_decap_8 FILLER_80_926 ();
 sg13g2_decap_8 FILLER_80_933 ();
 sg13g2_decap_8 FILLER_80_940 ();
 sg13g2_fill_1 FILLER_80_947 ();
 sg13g2_decap_8 FILLER_80_956 ();
 sg13g2_fill_2 FILLER_80_963 ();
 sg13g2_fill_1 FILLER_80_965 ();
 sg13g2_fill_1 FILLER_80_970 ();
 sg13g2_decap_8 FILLER_80_979 ();
 sg13g2_fill_1 FILLER_80_986 ();
 sg13g2_decap_8 FILLER_80_1008 ();
 sg13g2_fill_2 FILLER_80_1015 ();
 sg13g2_fill_2 FILLER_80_1021 ();
 sg13g2_decap_8 FILLER_80_1033 ();
 sg13g2_decap_8 FILLER_80_1040 ();
 sg13g2_decap_8 FILLER_80_1047 ();
 sg13g2_decap_8 FILLER_80_1054 ();
 sg13g2_decap_8 FILLER_80_1061 ();
 sg13g2_decap_8 FILLER_80_1068 ();
 sg13g2_decap_8 FILLER_80_1075 ();
 sg13g2_decap_8 FILLER_80_1082 ();
 sg13g2_decap_8 FILLER_80_1089 ();
 sg13g2_decap_8 FILLER_80_1096 ();
 sg13g2_decap_8 FILLER_80_1103 ();
 sg13g2_decap_8 FILLER_80_1110 ();
 sg13g2_decap_8 FILLER_80_1117 ();
 sg13g2_decap_8 FILLER_80_1124 ();
 sg13g2_decap_8 FILLER_80_1131 ();
 sg13g2_decap_8 FILLER_80_1138 ();
 sg13g2_decap_8 FILLER_80_1145 ();
 sg13g2_decap_8 FILLER_80_1152 ();
 sg13g2_decap_8 FILLER_80_1159 ();
 sg13g2_decap_8 FILLER_80_1166 ();
 sg13g2_decap_8 FILLER_80_1173 ();
 sg13g2_decap_8 FILLER_80_1180 ();
 sg13g2_decap_8 FILLER_80_1187 ();
 sg13g2_decap_8 FILLER_80_1194 ();
 sg13g2_decap_8 FILLER_80_1201 ();
 sg13g2_decap_8 FILLER_80_1208 ();
 sg13g2_decap_8 FILLER_80_1215 ();
 sg13g2_decap_8 FILLER_80_1222 ();
 sg13g2_decap_8 FILLER_80_1229 ();
 sg13g2_decap_8 FILLER_80_1236 ();
 sg13g2_decap_8 FILLER_80_1243 ();
 sg13g2_decap_8 FILLER_80_1250 ();
 sg13g2_decap_8 FILLER_80_1257 ();
 sg13g2_decap_8 FILLER_80_1264 ();
 sg13g2_decap_8 FILLER_80_1271 ();
 sg13g2_decap_8 FILLER_80_1278 ();
 sg13g2_decap_8 FILLER_80_1285 ();
 sg13g2_decap_8 FILLER_80_1292 ();
 sg13g2_decap_8 FILLER_80_1299 ();
 sg13g2_decap_8 FILLER_80_1306 ();
 sg13g2_decap_8 FILLER_80_1313 ();
 sg13g2_decap_8 FILLER_80_1320 ();
 sg13g2_decap_8 FILLER_80_1327 ();
 sg13g2_decap_8 FILLER_80_1334 ();
 sg13g2_decap_8 FILLER_80_1341 ();
 sg13g2_decap_8 FILLER_80_1348 ();
 sg13g2_decap_8 FILLER_80_1355 ();
 sg13g2_decap_8 FILLER_80_1362 ();
 sg13g2_decap_8 FILLER_80_1369 ();
 sg13g2_decap_8 FILLER_80_1376 ();
 sg13g2_decap_8 FILLER_80_1383 ();
 sg13g2_decap_8 FILLER_80_1390 ();
 sg13g2_decap_8 FILLER_80_1397 ();
 sg13g2_decap_8 FILLER_80_1404 ();
 sg13g2_decap_8 FILLER_80_1411 ();
 sg13g2_decap_8 FILLER_80_1418 ();
 sg13g2_decap_8 FILLER_80_1425 ();
 sg13g2_decap_8 FILLER_80_1432 ();
 sg13g2_decap_8 FILLER_80_1439 ();
 sg13g2_decap_8 FILLER_80_1446 ();
 sg13g2_decap_8 FILLER_80_1453 ();
 sg13g2_decap_8 FILLER_80_1460 ();
 sg13g2_decap_8 FILLER_80_1467 ();
 sg13g2_decap_8 FILLER_80_1474 ();
 sg13g2_decap_8 FILLER_80_1481 ();
 sg13g2_decap_8 FILLER_80_1488 ();
 sg13g2_decap_8 FILLER_80_1495 ();
 sg13g2_decap_8 FILLER_80_1502 ();
 sg13g2_decap_8 FILLER_80_1509 ();
 sg13g2_decap_8 FILLER_80_1516 ();
 sg13g2_decap_8 FILLER_80_1523 ();
 sg13g2_decap_8 FILLER_80_1530 ();
 sg13g2_decap_8 FILLER_80_1537 ();
 sg13g2_decap_8 FILLER_80_1544 ();
 sg13g2_decap_8 FILLER_80_1551 ();
 sg13g2_decap_8 FILLER_80_1558 ();
 sg13g2_decap_8 FILLER_80_1565 ();
 sg13g2_decap_8 FILLER_80_1572 ();
 sg13g2_decap_8 FILLER_80_1579 ();
 sg13g2_decap_8 FILLER_80_1586 ();
 sg13g2_decap_8 FILLER_80_1593 ();
 sg13g2_decap_8 FILLER_80_1600 ();
 sg13g2_decap_8 FILLER_80_1607 ();
 sg13g2_decap_8 FILLER_80_1614 ();
 sg13g2_decap_8 FILLER_80_1621 ();
 sg13g2_decap_8 FILLER_80_1628 ();
 sg13g2_decap_8 FILLER_80_1635 ();
 sg13g2_decap_8 FILLER_80_1642 ();
 sg13g2_decap_8 FILLER_80_1649 ();
 sg13g2_decap_8 FILLER_80_1656 ();
 sg13g2_decap_8 FILLER_80_1663 ();
 sg13g2_decap_8 FILLER_80_1670 ();
 sg13g2_decap_8 FILLER_80_1677 ();
 sg13g2_decap_8 FILLER_80_1684 ();
 sg13g2_decap_8 FILLER_80_1691 ();
 sg13g2_decap_8 FILLER_80_1698 ();
 sg13g2_decap_8 FILLER_80_1705 ();
 sg13g2_decap_8 FILLER_80_1712 ();
 sg13g2_decap_8 FILLER_80_1719 ();
 sg13g2_decap_8 FILLER_80_1726 ();
 sg13g2_decap_8 FILLER_80_1733 ();
 sg13g2_decap_8 FILLER_80_1740 ();
 sg13g2_decap_8 FILLER_80_1747 ();
 sg13g2_decap_8 FILLER_80_1754 ();
 sg13g2_decap_8 FILLER_80_1761 ();
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net25;
 assign uio_out[1] = net26;
 assign uio_out[2] = net27;
 assign uio_out[3] = net28;
 assign uio_out[4] = net29;
 assign uio_out[5] = net30;
 assign uio_out[6] = net31;
 assign uio_out[7] = net32;
endmodule

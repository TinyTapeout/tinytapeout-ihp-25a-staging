module tt_um_quarren42_demoscene_top (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire clknet_0_clk;
 wire b;
 wire \bitmap_xofs[0] ;
 wire \bitmap_xofs[1] ;
 wire \bitmap_xofs[2] ;
 wire \bitmap_xofs[3] ;
 wire \bitmap_xofs[4] ;
 wire \bitmap_yofs[0] ;
 wire \bitmap_yofs[1] ;
 wire \bitmap_yofs[2] ;
 wire \bitmap_yofs[3] ;
 wire \bitmap_yofs[4] ;
 wire \bitsTemp[10] ;
 wire \bitsTemp[11] ;
 wire \bitsTemp[12] ;
 wire \bitsTemp[13] ;
 wire \bitsTemp[14] ;
 wire \bitsTemp[15] ;
 wire \bitsTemp[16] ;
 wire \bitsTemp[17] ;
 wire \bitsTemp[18] ;
 wire \bitsTemp[19] ;
 wire \bitsTemp[1] ;
 wire \bitsTemp[20] ;
 wire \bitsTemp[21] ;
 wire \bitsTemp[22] ;
 wire \bitsTemp[23] ;
 wire \bitsTemp[24] ;
 wire \bitsTemp[25] ;
 wire \bitsTemp[26] ;
 wire \bitsTemp[27] ;
 wire \bitsTemp[28] ;
 wire \bitsTemp[29] ;
 wire \bitsTemp[2] ;
 wire \bitsTemp[30] ;
 wire \bitsTemp[31] ;
 wire \bitsTemp[3] ;
 wire \bitsTemp[4] ;
 wire \bitsTemp[8] ;
 wire \bitsTemp[9] ;
 wire bmpOnH;
 wire bmpOnV;
 wire g;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire r;
 wire test_b_h;
 wire test_b_v;
 wire test_g_h;
 wire test_g_v;
 wire test_h;
 wire test_v;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire \v_offset[0] ;
 wire \v_offset[1] ;
 wire \v_offset[2] ;
 wire \v_offset[3] ;
 wire \v_offset[4] ;
 wire \v_offset[5] ;
 wire \v_offset[6] ;
 wire \v_offset[7] ;
 wire \v_offset[8] ;
 wire \v_offset[9] ;
 wire v_offset_rev_flag;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net1;
 wire net2;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;

 sg13g2_inv_1 _0990_ (.Y(_0116_),
    .A(net284));
 sg13g2_inv_2 _0991_ (.Y(_0117_),
    .A(\bitmap_xofs[1] ));
 sg13g2_inv_1 _0992_ (.Y(_0118_),
    .A(net281));
 sg13g2_inv_1 _0993_ (.Y(_0119_),
    .A(net277));
 sg13g2_inv_1 _0994_ (.Y(_0120_),
    .A(net264));
 sg13g2_inv_2 _0995_ (.Y(_0121_),
    .A(net101));
 sg13g2_inv_2 _0996_ (.Y(_0122_),
    .A(\hvsync_gen.vpos[2] ));
 sg13g2_inv_1 _0997_ (.Y(_0123_),
    .A(net272));
 sg13g2_inv_2 _0998_ (.Y(_0124_),
    .A(\hvsync_gen.vpos[9] ));
 sg13g2_inv_2 _0999_ (.Y(_0125_),
    .A(net253));
 sg13g2_inv_2 _1000_ (.Y(_0126_),
    .A(net248));
 sg13g2_inv_1 _1001_ (.Y(_0127_),
    .A(net251));
 sg13g2_inv_1 _1002_ (.Y(_0128_),
    .A(net245));
 sg13g2_inv_2 _1003_ (.Y(_0129_),
    .A(\v_offset[9] ));
 sg13g2_inv_1 _1004_ (.Y(_0130_),
    .A(net81));
 sg13g2_inv_2 _1005_ (.Y(_0131_),
    .A(_0035_));
 sg13g2_inv_2 _1006_ (.Y(_0132_),
    .A(_0039_));
 sg13g2_inv_1 _1007_ (.Y(_0133_),
    .A(net86));
 sg13g2_inv_1 _1008_ (.Y(_0134_),
    .A(_0043_));
 sg13g2_inv_2 _1009_ (.Y(_0135_),
    .A(net87));
 sg13g2_inv_1 _1010_ (.Y(_0136_),
    .A(net269));
 sg13g2_inv_1 _1011_ (.Y(_0137_),
    .A(_0053_));
 sg13g2_inv_1 _1012_ (.Y(_0138_),
    .A(\bitsTemp[1] ));
 sg13g2_inv_1 _1013_ (.Y(_0139_),
    .A(net229));
 sg13g2_nand3_1 _1014_ (.B(net266),
    .C(net267),
    .A(net263),
    .Y(_0140_));
 sg13g2_nand2_1 _1015_ (.Y(_0141_),
    .A(net103),
    .B(_0124_));
 sg13g2_nand3b_1 _1016_ (.B(net271),
    .C(_0122_),
    .Y(_0142_),
    .A_N(\bitmap_yofs[0] ));
 sg13g2_nor4_1 _1017_ (.A(_0123_),
    .B(net84),
    .C(_0141_),
    .D(_0142_),
    .Y(_0031_));
 sg13g2_nand2_2 _1018_ (.Y(_0143_),
    .A(net276),
    .B(net274));
 sg13g2_nor2_1 _1019_ (.A(\bitmap_xofs[1] ),
    .B(net283),
    .Y(_0144_));
 sg13g2_nand2_1 _1020_ (.Y(_0145_),
    .A(net260),
    .B(net259));
 sg13g2_nand3_1 _1021_ (.B(net274),
    .C(_0145_),
    .A(net279),
    .Y(_0146_));
 sg13g2_and2_1 _1022_ (.A(\bitmap_xofs[1] ),
    .B(net283),
    .X(_0147_));
 sg13g2_inv_1 _1023_ (.Y(_0148_),
    .A(net258));
 sg13g2_nand3_1 _1024_ (.B(net281),
    .C(net258),
    .A(net278),
    .Y(_0149_));
 sg13g2_nand3_1 _1025_ (.B(net274),
    .C(_0149_),
    .A(_0119_),
    .Y(_0150_));
 sg13g2_a22oi_1 _1026_ (.Y(_0030_),
    .B1(_0150_),
    .B2(_0130_),
    .A2(_0146_),
    .A1(_0143_));
 sg13g2_or2_1 _1027_ (.X(_0151_),
    .B(net238),
    .A(net236));
 sg13g2_nor2_2 _1028_ (.A(net254),
    .B(net257),
    .Y(_0152_));
 sg13g2_o21ai_1 _1029_ (.B1(net250),
    .Y(_0153_),
    .A1(net253),
    .A2(net256));
 sg13g2_and2_1 _1030_ (.A(net247),
    .B(net251),
    .X(_0154_));
 sg13g2_nand2_2 _1031_ (.Y(_0155_),
    .A(net248),
    .B(net251));
 sg13g2_nor2_1 _1032_ (.A(_0152_),
    .B(_0155_),
    .Y(_0156_));
 sg13g2_nor2b_1 _1033_ (.A(net245),
    .B_N(net242),
    .Y(_0157_));
 sg13g2_o21ai_1 _1034_ (.B1(_0157_),
    .Y(_0158_),
    .A1(net228),
    .A2(_0155_));
 sg13g2_a21o_2 _1035_ (.A2(_0158_),
    .A1(_0131_),
    .B1(_0151_),
    .X(_0159_));
 sg13g2_nor2b_1 _1036_ (.A(_0036_),
    .B_N(_0159_),
    .Y(_0160_));
 sg13g2_xnor2_1 _1037_ (.Y(_0161_),
    .A(_0036_),
    .B(_0159_));
 sg13g2_xor2_1 _1038_ (.B(_0159_),
    .A(_0036_),
    .X(_0162_));
 sg13g2_nand2_1 _1039_ (.Y(_0163_),
    .A(net241),
    .B(_0158_));
 sg13g2_a21oi_1 _1040_ (.A1(net244),
    .A2(_0158_),
    .Y(_0164_),
    .B1(_0132_));
 sg13g2_xnor2_1 _1041_ (.Y(_0165_),
    .A(_0038_),
    .B(_0164_));
 sg13g2_a22oi_1 _1042_ (.Y(_0166_),
    .B1(_0165_),
    .B2(_0133_),
    .A2(_0161_),
    .A1(net277));
 sg13g2_nor2_1 _1043_ (.A(_0133_),
    .B(_0165_),
    .Y(_0167_));
 sg13g2_xnor2_1 _1044_ (.Y(_0168_),
    .A(_0132_),
    .B(_0163_));
 sg13g2_xnor2_1 _1045_ (.Y(_0169_),
    .A(_0039_),
    .B(_0163_));
 sg13g2_nand2_1 _1046_ (.Y(_0170_),
    .A(net282),
    .B(_0169_));
 sg13g2_o21ai_1 _1047_ (.B1(_0041_),
    .Y(_0171_),
    .A1(net228),
    .A2(_0155_));
 sg13g2_xnor2_1 _1048_ (.Y(_0172_),
    .A(_0131_),
    .B(_0171_));
 sg13g2_nor2_1 _1049_ (.A(_0117_),
    .B(_0172_),
    .Y(_0173_));
 sg13g2_o21ai_1 _1050_ (.B1(_0171_),
    .Y(_0174_),
    .A1(_0041_),
    .A2(_0155_));
 sg13g2_inv_1 _1051_ (.Y(_0175_),
    .A(_0174_));
 sg13g2_xnor2_1 _1052_ (.Y(_0176_),
    .A(_0041_),
    .B(_0156_));
 sg13g2_xnor2_1 _1053_ (.Y(_0177_),
    .A(_0042_),
    .B(_0172_));
 sg13g2_a21oi_1 _1054_ (.A1(_0043_),
    .A2(_0176_),
    .Y(_0178_),
    .B1(_0177_));
 sg13g2_xnor2_1 _1055_ (.Y(_0179_),
    .A(net247),
    .B(_0153_));
 sg13g2_nor2_1 _1056_ (.A(net284),
    .B(_0179_),
    .Y(_0180_));
 sg13g2_nor2_1 _1057_ (.A(net254),
    .B(net251),
    .Y(_0181_));
 sg13g2_xnor2_1 _1058_ (.Y(_0182_),
    .A(net251),
    .B(net228));
 sg13g2_xnor2_1 _1059_ (.Y(_0183_),
    .A(net285),
    .B(_0182_));
 sg13g2_and2_1 _1060_ (.A(net284),
    .B(_0179_),
    .X(_0184_));
 sg13g2_or3_1 _1061_ (.A(_0180_),
    .B(_0183_),
    .C(_0184_),
    .X(_0185_));
 sg13g2_nand2_2 _1062_ (.Y(_0186_),
    .A(net254),
    .B(net256));
 sg13g2_xnor2_1 _1063_ (.Y(_0187_),
    .A(net253),
    .B(net256));
 sg13g2_nand2b_1 _1064_ (.Y(_0188_),
    .B(net256),
    .A_N(\hvsync_gen.hpos[0] ));
 sg13g2_xnor2_1 _1065_ (.Y(_0189_),
    .A(_0045_),
    .B(net227));
 sg13g2_a22oi_1 _1066_ (.Y(_0190_),
    .B1(_0188_),
    .B2(_0189_),
    .A2(net227),
    .A1(\hvsync_gen.hpos[1] ));
 sg13g2_or2_1 _1067_ (.X(_0191_),
    .B(_0190_),
    .A(_0185_));
 sg13g2_nor2_1 _1068_ (.A(_0043_),
    .B(_0176_),
    .Y(_0192_));
 sg13g2_nand2b_1 _1069_ (.Y(_0193_),
    .B(_0182_),
    .A_N(_0044_));
 sg13g2_nor2_1 _1070_ (.A(_0180_),
    .B(_0193_),
    .Y(_0194_));
 sg13g2_nor3_1 _1071_ (.A(_0184_),
    .B(_0192_),
    .C(_0194_),
    .Y(_0195_));
 sg13g2_a221oi_1 _1072_ (.B2(_0195_),
    .C1(_0177_),
    .B1(_0191_),
    .A1(_0043_),
    .Y(_0196_),
    .A2(_0176_));
 sg13g2_xnor2_1 _1073_ (.Y(_0197_),
    .A(_0040_),
    .B(_0169_));
 sg13g2_o21ai_1 _1074_ (.B1(_0197_),
    .Y(_0198_),
    .A1(_0173_),
    .A2(_0196_));
 sg13g2_a21oi_1 _1075_ (.A1(_0170_),
    .A2(_0198_),
    .Y(_0199_),
    .B1(_0167_));
 sg13g2_nand2b_1 _1076_ (.Y(_0200_),
    .B(_0166_),
    .A_N(_0199_));
 sg13g2_xnor2_1 _1077_ (.Y(_0201_),
    .A(\v_offset[9] ),
    .B(_0160_));
 sg13g2_xnor2_1 _1078_ (.Y(_0202_),
    .A(net275),
    .B(_0201_));
 sg13g2_a21oi_1 _1079_ (.A1(_0119_),
    .A2(_0162_),
    .Y(_0203_),
    .B1(_0202_));
 sg13g2_a22oi_1 _1080_ (.Y(_0204_),
    .B1(_0203_),
    .B2(_0200_),
    .A2(_0201_),
    .A1(_0130_));
 sg13g2_a21o_2 _1081_ (.A2(net250),
    .A1(net247),
    .B1(net246),
    .X(_0205_));
 sg13g2_xor2_1 _1082_ (.B(_0205_),
    .A(net241),
    .X(_0206_));
 sg13g2_xnor2_1 _1083_ (.Y(_0207_),
    .A(net241),
    .B(_0205_));
 sg13g2_nor2b_1 _1084_ (.A(\hvsync_gen.hpos[1] ),
    .B_N(net256),
    .Y(_0208_));
 sg13g2_xor2_1 _1085_ (.B(net256),
    .A(net287),
    .X(_0209_));
 sg13g2_xor2_1 _1086_ (.B(net253),
    .A(net287),
    .X(_0210_));
 sg13g2_nor2b_1 _1087_ (.A(_0210_),
    .B_N(_0188_),
    .Y(_0211_));
 sg13g2_a221oi_1 _1088_ (.B2(net286),
    .C1(_0211_),
    .B1(net250),
    .A1(net287),
    .Y(_0212_),
    .A2(_0125_));
 sg13g2_nor2_1 _1089_ (.A(net286),
    .B(net250),
    .Y(_0213_));
 sg13g2_nor2_2 _1090_ (.A(net248),
    .B(net252),
    .Y(_0214_));
 sg13g2_nor2_1 _1091_ (.A(_0154_),
    .B(_0214_),
    .Y(_0215_));
 sg13g2_nor3_1 _1092_ (.A(net284),
    .B(_0154_),
    .C(_0214_),
    .Y(_0216_));
 sg13g2_nor3_1 _1093_ (.A(_0212_),
    .B(_0213_),
    .C(_0216_),
    .Y(_0217_));
 sg13g2_xnor2_1 _1094_ (.Y(_0218_),
    .A(_0041_),
    .B(_0154_));
 sg13g2_inv_1 _1095_ (.Y(_0219_),
    .A(_0218_));
 sg13g2_o21ai_1 _1096_ (.B1(\hvsync_gen.hpos[3] ),
    .Y(_0220_),
    .A1(_0154_),
    .A2(_0214_));
 sg13g2_o21ai_1 _1097_ (.B1(_0220_),
    .Y(_0221_),
    .A1(_0043_),
    .A2(_0219_));
 sg13g2_xnor2_1 _1098_ (.Y(_0222_),
    .A(_0042_),
    .B(_0206_));
 sg13g2_a21oi_1 _1099_ (.A1(_0043_),
    .A2(_0219_),
    .Y(_0223_),
    .B1(_0222_));
 sg13g2_o21ai_1 _1100_ (.B1(_0223_),
    .Y(_0224_),
    .A1(_0217_),
    .A2(_0221_));
 sg13g2_o21ai_1 _1101_ (.B1(_0224_),
    .Y(_0225_),
    .A1(_0117_),
    .A2(_0206_));
 sg13g2_a21oi_2 _1102_ (.B1(net240),
    .Y(_0226_),
    .A2(_0205_),
    .A1(net241));
 sg13g2_nand3_1 _1103_ (.B(net240),
    .C(_0205_),
    .A(net241),
    .Y(_0227_));
 sg13g2_nand2b_2 _1104_ (.Y(_0228_),
    .B(_0227_),
    .A_N(_0226_));
 sg13g2_xnor2_1 _1105_ (.Y(_0229_),
    .A(net282),
    .B(_0228_));
 sg13g2_nor2b_1 _1106_ (.A(_0226_),
    .B_N(net237),
    .Y(_0230_));
 sg13g2_xnor2_1 _1107_ (.Y(_0231_),
    .A(net237),
    .B(_0226_));
 sg13g2_nand2b_1 _1108_ (.Y(_0232_),
    .B(net279),
    .A_N(_0231_));
 sg13g2_o21ai_1 _1109_ (.B1(_0232_),
    .Y(_0233_),
    .A1(_0040_),
    .A2(_0228_));
 sg13g2_a21oi_1 _1110_ (.A1(_0225_),
    .A2(_0229_),
    .Y(_0234_),
    .B1(_0233_));
 sg13g2_xnor2_1 _1111_ (.Y(_0235_),
    .A(_0036_),
    .B(_0230_));
 sg13g2_nor2b_1 _1112_ (.A(net279),
    .B_N(_0231_),
    .Y(_0236_));
 sg13g2_xor2_1 _1113_ (.B(_0235_),
    .A(_0046_),
    .X(_0237_));
 sg13g2_nor3_1 _1114_ (.A(_0234_),
    .B(_0236_),
    .C(_0237_),
    .Y(_0238_));
 sg13g2_nor2_1 _1115_ (.A(net233),
    .B(_0230_),
    .Y(_0239_));
 sg13g2_nor2_1 _1116_ (.A(_0129_),
    .B(_0239_),
    .Y(_0240_));
 sg13g2_nor2_2 _1117_ (.A(\v_offset[9] ),
    .B(net231),
    .Y(_0241_));
 sg13g2_xnor2_1 _1118_ (.Y(_0242_),
    .A(_0129_),
    .B(_0239_));
 sg13g2_a221oi_1 _1119_ (.B2(net274),
    .C1(_0238_),
    .B1(_0242_),
    .A1(net276),
    .Y(_0243_),
    .A2(_0235_));
 sg13g2_a21oi_1 _1120_ (.A1(_0129_),
    .A2(_0239_),
    .Y(_0244_),
    .B1(net274));
 sg13g2_nor3_1 _1121_ (.A(_0240_),
    .B(_0243_),
    .C(_0244_),
    .Y(_0245_));
 sg13g2_a21oi_2 _1122_ (.B1(\v_offset[9] ),
    .Y(_0246_),
    .A2(_0159_),
    .A1(net233));
 sg13g2_inv_1 _1123_ (.Y(_0247_),
    .A(_0246_));
 sg13g2_or2_1 _1124_ (.X(_0248_),
    .B(net256),
    .A(\hvsync_gen.hpos[0] ));
 sg13g2_xnor2_1 _1125_ (.Y(_0249_),
    .A(\hvsync_gen.hpos[0] ),
    .B(net256));
 sg13g2_nand2_1 _1126_ (.Y(_0250_),
    .A(_0189_),
    .B(_0249_));
 sg13g2_nor4_1 _1127_ (.A(_0167_),
    .B(_0185_),
    .C(_0192_),
    .D(_0250_),
    .Y(_0251_));
 sg13g2_nand3_1 _1128_ (.B(_0197_),
    .C(_0251_),
    .A(_0178_),
    .Y(_0252_));
 sg13g2_nand2_1 _1129_ (.Y(_0253_),
    .A(_0166_),
    .B(_0203_));
 sg13g2_o21ai_1 _1130_ (.B1(_0246_),
    .Y(_0254_),
    .A1(_0252_),
    .A2(_0253_));
 sg13g2_nor3_1 _1131_ (.A(_0204_),
    .B(_0245_),
    .C(_0254_),
    .Y(_0006_));
 sg13g2_nor2_1 _1132_ (.A(_0125_),
    .B(_0127_),
    .Y(_0255_));
 sg13g2_nand2_2 _1133_ (.Y(_0256_),
    .A(net255),
    .B(net252));
 sg13g2_nor2_2 _1134_ (.A(net249),
    .B(net245),
    .Y(_0257_));
 sg13g2_nand2_2 _1135_ (.Y(_0258_),
    .A(_0256_),
    .B(_0257_));
 sg13g2_xnor2_1 _1136_ (.Y(_0259_),
    .A(_0131_),
    .B(_0258_));
 sg13g2_inv_1 _1137_ (.Y(_0260_),
    .A(_0259_));
 sg13g2_xnor2_1 _1138_ (.Y(_0261_),
    .A(net255),
    .B(net252));
 sg13g2_nand2b_1 _1139_ (.Y(_0262_),
    .B(net257),
    .A_N(\hvsync_gen.vpos[0] ));
 sg13g2_nor2b_1 _1140_ (.A(\hvsync_gen.vpos[1] ),
    .B_N(net257),
    .Y(_0263_));
 sg13g2_xnor2_1 _1141_ (.Y(_0264_),
    .A(\hvsync_gen.vpos[1] ),
    .B(net257));
 sg13g2_xor2_1 _1142_ (.B(net255),
    .A(\hvsync_gen.vpos[1] ),
    .X(_0265_));
 sg13g2_nand2_1 _1143_ (.Y(_0266_),
    .A(_0262_),
    .B(_0265_));
 sg13g2_o21ai_1 _1144_ (.B1(_0266_),
    .Y(_0267_),
    .A1(_0123_),
    .A2(_0125_));
 sg13g2_xnor2_1 _1145_ (.Y(_0268_),
    .A(_0053_),
    .B(_0261_));
 sg13g2_a22oi_1 _1146_ (.Y(_0269_),
    .B1(_0267_),
    .B2(_0268_),
    .A2(_0261_),
    .A1(\hvsync_gen.vpos[2] ));
 sg13g2_xnor2_1 _1147_ (.Y(_0270_),
    .A(_0126_),
    .B(_0256_));
 sg13g2_a21oi_1 _1148_ (.A1(_0121_),
    .A2(_0270_),
    .Y(_0271_),
    .B1(_0269_));
 sg13g2_nand2b_1 _1149_ (.Y(_0272_),
    .B(\hvsync_gen.vpos[3] ),
    .A_N(_0270_));
 sg13g2_nand2_1 _1150_ (.Y(_0273_),
    .A(_0055_),
    .B(_0256_));
 sg13g2_xor2_1 _1151_ (.B(_0273_),
    .A(_0041_),
    .X(_0274_));
 sg13g2_o21ai_1 _1152_ (.B1(_0272_),
    .Y(_0275_),
    .A1(net269),
    .A2(_0274_));
 sg13g2_or2_1 _1153_ (.X(_0276_),
    .B(_0275_),
    .A(_0271_));
 sg13g2_xnor2_1 _1154_ (.Y(_0277_),
    .A(_0050_),
    .B(_0259_));
 sg13g2_a21oi_1 _1155_ (.A1(net269),
    .A2(_0274_),
    .Y(_0278_),
    .B1(_0277_));
 sg13g2_a22oi_1 _1156_ (.Y(_0279_),
    .B1(_0276_),
    .B2(_0278_),
    .A2(_0260_),
    .A1(net268));
 sg13g2_nor2_1 _1157_ (.A(net242),
    .B(_0258_),
    .Y(_0280_));
 sg13g2_xnor2_1 _1158_ (.Y(_0281_),
    .A(_0132_),
    .B(_0280_));
 sg13g2_xor2_1 _1159_ (.B(_0281_),
    .A(_0033_),
    .X(_0282_));
 sg13g2_nor2_2 _1160_ (.A(net243),
    .B(net238),
    .Y(_0283_));
 sg13g2_nand3_1 _1161_ (.B(_0257_),
    .C(_0283_),
    .A(_0256_),
    .Y(_0284_));
 sg13g2_xnor2_1 _1162_ (.Y(_0285_),
    .A(_0038_),
    .B(_0284_));
 sg13g2_a22oi_1 _1163_ (.Y(_0286_),
    .B1(_0285_),
    .B2(net263),
    .A2(_0281_),
    .A1(net266));
 sg13g2_o21ai_1 _1164_ (.B1(_0286_),
    .Y(_0287_),
    .A1(_0279_),
    .A2(_0282_));
 sg13g2_nor2_1 _1165_ (.A(net236),
    .B(_0284_),
    .Y(_0288_));
 sg13g2_o21ai_1 _1166_ (.B1(net231),
    .Y(_0289_),
    .A1(net234),
    .A2(_0284_));
 sg13g2_inv_1 _1167_ (.Y(_0290_),
    .A(_0289_));
 sg13g2_nor2_1 _1168_ (.A(net231),
    .B(_0151_),
    .Y(_0291_));
 sg13g2_a21oi_1 _1169_ (.A1(_0280_),
    .A2(_0291_),
    .Y(_0292_),
    .B1(_0290_));
 sg13g2_nand2b_1 _1170_ (.Y(_0293_),
    .B(_0120_),
    .A_N(_0285_));
 sg13g2_xor2_1 _1171_ (.B(_0292_),
    .A(_0049_),
    .X(_0294_));
 sg13g2_nand3_1 _1172_ (.B(_0293_),
    .C(_0294_),
    .A(_0287_),
    .Y(_0295_));
 sg13g2_nor2b_1 _1173_ (.A(_0292_),
    .B_N(\bitmap_yofs[4] ),
    .Y(_0296_));
 sg13g2_nor2_1 _1174_ (.A(_0124_),
    .B(\v_offset[9] ),
    .Y(_0297_));
 sg13g2_a21oi_1 _1175_ (.A1(_0289_),
    .A2(_0297_),
    .Y(_0298_),
    .B1(_0296_));
 sg13g2_nand2_1 _1176_ (.Y(_0299_),
    .A(_0124_),
    .B(\v_offset[9] ));
 sg13g2_a21oi_1 _1177_ (.A1(_0289_),
    .A2(_0299_),
    .Y(_0300_),
    .B1(_0297_));
 sg13g2_a21oi_1 _1178_ (.A1(_0295_),
    .A2(_0298_),
    .Y(_0301_),
    .B1(_0300_));
 sg13g2_nand2_2 _1179_ (.Y(_0302_),
    .A(_0186_),
    .B(_0214_));
 sg13g2_a21oi_2 _1180_ (.B1(net242),
    .Y(_0303_),
    .A2(_0302_),
    .A1(net246));
 sg13g2_nand2_2 _1181_ (.Y(_0304_),
    .A(net235),
    .B(net239));
 sg13g2_o21ai_1 _1182_ (.B1(_0036_),
    .Y(_0305_),
    .A1(_0303_),
    .A2(_0304_));
 sg13g2_xor2_1 _1183_ (.B(_0305_),
    .A(_0048_),
    .X(_0306_));
 sg13g2_or3_1 _1184_ (.A(_0036_),
    .B(_0303_),
    .C(_0304_),
    .X(_0307_));
 sg13g2_and2_1 _1185_ (.A(_0305_),
    .B(_0307_),
    .X(_0308_));
 sg13g2_xnor2_1 _1186_ (.Y(_0309_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_0306_));
 sg13g2_a21o_1 _1187_ (.A2(_0308_),
    .A1(_0049_),
    .B1(_0309_),
    .X(_0310_));
 sg13g2_nor2_1 _1188_ (.A(_0049_),
    .B(_0308_),
    .Y(_0311_));
 sg13g2_nor2_1 _1189_ (.A(_0039_),
    .B(_0303_),
    .Y(_0312_));
 sg13g2_xor2_1 _1190_ (.B(_0312_),
    .A(net234),
    .X(_0313_));
 sg13g2_a21oi_1 _1191_ (.A1(net263),
    .A2(_0313_),
    .Y(_0314_),
    .B1(_0311_));
 sg13g2_nand2_1 _1192_ (.Y(_0315_),
    .A(_0052_),
    .B(_0186_));
 sg13g2_xnor2_1 _1193_ (.Y(_0316_),
    .A(_0126_),
    .B(_0315_));
 sg13g2_nand2b_1 _1194_ (.Y(_0317_),
    .B(\hvsync_gen.vpos[3] ),
    .A_N(_0316_));
 sg13g2_xnor2_1 _1195_ (.Y(_0318_),
    .A(net246),
    .B(_0302_));
 sg13g2_inv_1 _1196_ (.Y(_0319_),
    .A(_0318_));
 sg13g2_o21ai_1 _1197_ (.B1(_0317_),
    .Y(_0320_),
    .A1(net269),
    .A2(_0318_));
 sg13g2_nand2_1 _1198_ (.Y(_0321_),
    .A(_0121_),
    .B(_0316_));
 sg13g2_xor2_1 _1199_ (.B(_0186_),
    .A(_0052_),
    .X(_0322_));
 sg13g2_nor2_1 _1200_ (.A(_0122_),
    .B(_0322_),
    .Y(_0323_));
 sg13g2_and2_1 _1201_ (.A(_0054_),
    .B(_0187_),
    .X(_0324_));
 sg13g2_nand2_1 _1202_ (.Y(_0325_),
    .A(_0054_),
    .B(net227));
 sg13g2_nor2_1 _1203_ (.A(_0054_),
    .B(net227),
    .Y(_0326_));
 sg13g2_a21o_1 _1204_ (.A2(_0325_),
    .A1(_0262_),
    .B1(_0326_),
    .X(_0327_));
 sg13g2_xnor2_1 _1205_ (.Y(_0328_),
    .A(_0053_),
    .B(_0322_));
 sg13g2_a21oi_1 _1206_ (.A1(_0121_),
    .A2(_0316_),
    .Y(_0329_),
    .B1(_0328_));
 sg13g2_a221oi_1 _1207_ (.B2(_0329_),
    .C1(_0320_),
    .B1(_0327_),
    .A1(_0321_),
    .Y(_0330_),
    .A2(_0323_));
 sg13g2_xnor2_1 _1208_ (.Y(_0331_),
    .A(net239),
    .B(_0303_));
 sg13g2_xnor2_1 _1209_ (.Y(_0332_),
    .A(_0033_),
    .B(_0331_));
 sg13g2_a21oi_1 _1210_ (.A1(_0186_),
    .A2(_0214_),
    .Y(_0333_),
    .B1(_0041_));
 sg13g2_xnor2_1 _1211_ (.Y(_0334_),
    .A(_0035_),
    .B(_0333_));
 sg13g2_a22oi_1 _1212_ (.Y(_0335_),
    .B1(_0334_),
    .B2(_0050_),
    .A2(_0318_),
    .A1(net269));
 sg13g2_o21ai_1 _1213_ (.B1(_0335_),
    .Y(_0336_),
    .A1(_0050_),
    .A2(_0334_));
 sg13g2_nand2b_1 _1214_ (.Y(_0337_),
    .B(_0332_),
    .A_N(_0336_));
 sg13g2_nor2b_1 _1215_ (.A(_0334_),
    .B_N(net268),
    .Y(_0338_));
 sg13g2_a22oi_1 _1216_ (.Y(_0339_),
    .B1(_0332_),
    .B2(_0338_),
    .A2(_0331_),
    .A1(net266));
 sg13g2_o21ai_1 _1217_ (.B1(_0339_),
    .Y(_0340_),
    .A1(_0330_),
    .A2(_0337_));
 sg13g2_o21ai_1 _1218_ (.B1(_0340_),
    .Y(_0341_),
    .A1(net263),
    .A2(_0313_));
 sg13g2_a21oi_1 _1219_ (.A1(_0314_),
    .A2(_0341_),
    .Y(_0342_),
    .B1(_0310_));
 sg13g2_a21oi_1 _1220_ (.A1(_0135_),
    .A2(_0306_),
    .Y(_0343_),
    .B1(_0342_));
 sg13g2_o21ai_1 _1221_ (.B1(_0241_),
    .Y(_0344_),
    .A1(_0303_),
    .A2(_0304_));
 sg13g2_xnor2_1 _1222_ (.Y(_0345_),
    .A(\hvsync_gen.vpos[0] ),
    .B(net257));
 sg13g2_nor3_1 _1223_ (.A(_0320_),
    .B(_0324_),
    .C(_0326_),
    .Y(_0346_));
 sg13g2_o21ai_1 _1224_ (.B1(_0346_),
    .Y(_0347_),
    .A1(net263),
    .A2(_0313_));
 sg13g2_nand3_1 _1225_ (.B(_0329_),
    .C(_0345_),
    .A(_0314_),
    .Y(_0348_));
 sg13g2_nor4_1 _1226_ (.A(_0310_),
    .B(_0337_),
    .C(_0347_),
    .D(_0348_),
    .Y(_0349_));
 sg13g2_nor4_1 _1227_ (.A(_0301_),
    .B(_0343_),
    .C(_0344_),
    .D(_0349_),
    .Y(_0007_));
 sg13g2_nor2b_2 _1228_ (.A(net251),
    .B_N(net248),
    .Y(_0350_));
 sg13g2_nand2b_2 _1229_ (.Y(_0351_),
    .B(_0350_),
    .A_N(_0186_));
 sg13g2_nand2_1 _1230_ (.Y(_0352_),
    .A(_0218_),
    .B(_0351_));
 sg13g2_nand3_1 _1231_ (.B(_0218_),
    .C(_0351_),
    .A(_0207_),
    .Y(_0353_));
 sg13g2_nor3_2 _1232_ (.A(_0228_),
    .B(_0231_),
    .C(_0353_),
    .Y(_0354_));
 sg13g2_nand2_1 _1233_ (.Y(_0355_),
    .A(_0235_),
    .B(_0354_));
 sg13g2_xnor2_1 _1234_ (.Y(_0356_),
    .A(_0242_),
    .B(_0355_));
 sg13g2_nand2_1 _1235_ (.Y(_0357_),
    .A(net274),
    .B(_0356_));
 sg13g2_xor2_1 _1236_ (.B(_0353_),
    .A(_0228_),
    .X(_0358_));
 sg13g2_nand3_1 _1237_ (.B(_0302_),
    .C(_0351_),
    .A(_0155_),
    .Y(_0359_));
 sg13g2_nand2b_1 _1238_ (.Y(_0360_),
    .B(_0116_),
    .A_N(_0359_));
 sg13g2_xnor2_1 _1239_ (.Y(_0361_),
    .A(_0127_),
    .B(_0186_));
 sg13g2_nand2b_1 _1240_ (.Y(_0362_),
    .B(net286),
    .A_N(_0361_));
 sg13g2_a22oi_1 _1241_ (.Y(_0363_),
    .B1(_0189_),
    .B2(_0248_),
    .A2(net227),
    .A1(net287));
 sg13g2_xnor2_1 _1242_ (.Y(_0364_),
    .A(net250),
    .B(_0044_));
 sg13g2_xor2_1 _1243_ (.B(_0364_),
    .A(_0186_),
    .X(_0365_));
 sg13g2_o21ai_1 _1244_ (.B1(_0362_),
    .Y(_0366_),
    .A1(_0363_),
    .A2(_0365_));
 sg13g2_mux2_1 _1245_ (.A0(_0041_),
    .A1(_0218_),
    .S(_0351_),
    .X(_0367_));
 sg13g2_inv_1 _1246_ (.Y(_0368_),
    .A(_0367_));
 sg13g2_and2_1 _1247_ (.A(\hvsync_gen.hpos[3] ),
    .B(_0359_),
    .X(_0369_));
 sg13g2_a221oi_1 _1248_ (.B2(_0134_),
    .C1(_0369_),
    .B1(_0368_),
    .A1(_0360_),
    .Y(_0370_),
    .A2(_0366_));
 sg13g2_a22oi_1 _1249_ (.Y(_0371_),
    .B1(_0367_),
    .B2(_0043_),
    .A2(_0352_),
    .A1(_0222_));
 sg13g2_o21ai_1 _1250_ (.B1(_0371_),
    .Y(_0372_),
    .A1(_0222_),
    .A2(_0352_));
 sg13g2_a21oi_1 _1251_ (.A1(_0206_),
    .A2(_0352_),
    .Y(_0373_),
    .B1(_0117_));
 sg13g2_nand2_1 _1252_ (.Y(_0374_),
    .A(_0353_),
    .B(_0373_));
 sg13g2_o21ai_1 _1253_ (.B1(_0374_),
    .Y(_0375_),
    .A1(_0370_),
    .A2(_0372_));
 sg13g2_xnor2_1 _1254_ (.Y(_0376_),
    .A(_0040_),
    .B(_0358_));
 sg13g2_a22oi_1 _1255_ (.Y(_0377_),
    .B1(_0375_),
    .B2(_0376_),
    .A2(_0358_),
    .A1(net282));
 sg13g2_o21ai_1 _1256_ (.B1(_0231_),
    .Y(_0378_),
    .A1(_0228_),
    .A2(_0353_));
 sg13g2_nor2b_1 _1257_ (.A(_0354_),
    .B_N(_0378_),
    .Y(_0379_));
 sg13g2_nor2_1 _1258_ (.A(net279),
    .B(_0379_),
    .Y(_0380_));
 sg13g2_xnor2_1 _1259_ (.Y(_0381_),
    .A(_0235_),
    .B(_0354_));
 sg13g2_nor2_1 _1260_ (.A(_0046_),
    .B(_0381_),
    .Y(_0382_));
 sg13g2_a21oi_1 _1261_ (.A1(net279),
    .A2(_0379_),
    .Y(_0383_),
    .B1(_0382_));
 sg13g2_o21ai_1 _1262_ (.B1(_0383_),
    .Y(_0384_),
    .A1(_0377_),
    .A2(_0380_));
 sg13g2_nand2_1 _1263_ (.Y(_0385_),
    .A(net94),
    .B(_0381_));
 sg13g2_xnor2_1 _1264_ (.Y(_0386_),
    .A(_0034_),
    .B(_0356_));
 sg13g2_nand3_1 _1265_ (.B(_0385_),
    .C(_0386_),
    .A(_0384_),
    .Y(_0387_));
 sg13g2_a22oi_1 _1266_ (.Y(_0388_),
    .B1(_0357_),
    .B2(_0387_),
    .A2(_0355_),
    .A1(_0240_));
 sg13g2_nor2_2 _1267_ (.A(_0035_),
    .B(_0174_),
    .Y(_0389_));
 sg13g2_nand2_1 _1268_ (.Y(_0390_),
    .A(_0168_),
    .B(_0389_));
 sg13g2_nand3b_1 _1269_ (.B(_0168_),
    .C(_0389_),
    .Y(_0391_),
    .A_N(_0165_));
 sg13g2_nor2_1 _1270_ (.A(_0161_),
    .B(_0391_),
    .Y(_0392_));
 sg13g2_nor3_1 _1271_ (.A(_0161_),
    .B(_0201_),
    .C(_0391_),
    .Y(_0393_));
 sg13g2_xnor2_1 _1272_ (.Y(_0394_),
    .A(_0201_),
    .B(_0392_));
 sg13g2_xnor2_1 _1273_ (.Y(_0395_),
    .A(_0034_),
    .B(_0394_));
 sg13g2_inv_1 _1274_ (.Y(_0396_),
    .A(_0395_));
 sg13g2_xnor2_1 _1275_ (.Y(_0397_),
    .A(_0162_),
    .B(_0391_));
 sg13g2_nor2_1 _1276_ (.A(net94),
    .B(_0397_),
    .Y(_0398_));
 sg13g2_xnor2_1 _1277_ (.Y(_0399_),
    .A(_0165_),
    .B(_0390_));
 sg13g2_or2_1 _1278_ (.X(_0400_),
    .B(_0399_),
    .A(net280));
 sg13g2_nand2_1 _1279_ (.Y(_0401_),
    .A(_0046_),
    .B(_0397_));
 sg13g2_nand3b_1 _1280_ (.B(_0400_),
    .C(_0401_),
    .Y(_0402_),
    .A_N(_0398_));
 sg13g2_nor2_1 _1281_ (.A(_0395_),
    .B(_0402_),
    .Y(_0403_));
 sg13g2_nor2b_1 _1282_ (.A(_0216_),
    .B_N(_0220_),
    .Y(_0404_));
 sg13g2_nor2_1 _1283_ (.A(_0364_),
    .B(_0404_),
    .Y(_0405_));
 sg13g2_xor2_1 _1284_ (.B(net227),
    .A(_0067_),
    .X(_0406_));
 sg13g2_xor2_1 _1285_ (.B(_0189_),
    .A(_0067_),
    .X(_0407_));
 sg13g2_a22oi_1 _1286_ (.Y(_0408_),
    .B1(_0407_),
    .B2(_0248_),
    .A2(_0406_),
    .A1(net287));
 sg13g2_nand2b_1 _1287_ (.Y(_0409_),
    .B(_0405_),
    .A_N(_0408_));
 sg13g2_or2_1 _1288_ (.X(_0410_),
    .B(net285),
    .A(net284));
 sg13g2_nor3_1 _1289_ (.A(_0116_),
    .B(net247),
    .C(_0213_),
    .Y(_0411_));
 sg13g2_o21ai_1 _1290_ (.B1(_0410_),
    .Y(_0412_),
    .A1(_0350_),
    .A2(_0411_));
 sg13g2_nand2_1 _1291_ (.Y(_0413_),
    .A(\bitmap_xofs[0] ),
    .B(_0218_));
 sg13g2_nand3_1 _1292_ (.B(_0412_),
    .C(_0413_),
    .A(_0409_),
    .Y(_0414_));
 sg13g2_xor2_1 _1293_ (.B(_0389_),
    .A(_0197_),
    .X(_0415_));
 sg13g2_or2_1 _1294_ (.X(_0416_),
    .B(_0218_),
    .A(net283));
 sg13g2_xnor2_1 _1295_ (.Y(_0417_),
    .A(_0175_),
    .B(_0177_));
 sg13g2_nand3_1 _1296_ (.B(_0416_),
    .C(_0417_),
    .A(_0415_),
    .Y(_0418_));
 sg13g2_nand2b_1 _1297_ (.Y(_0419_),
    .B(_0414_),
    .A_N(_0418_));
 sg13g2_o21ai_1 _1298_ (.B1(_0197_),
    .Y(_0420_),
    .A1(_0172_),
    .A2(_0175_));
 sg13g2_nand3_1 _1299_ (.B(_0415_),
    .C(_0420_),
    .A(\bitmap_xofs[1] ),
    .Y(_0421_));
 sg13g2_nand2_1 _1300_ (.Y(_0422_),
    .A(net280),
    .B(_0399_));
 sg13g2_or2_1 _1301_ (.X(_0423_),
    .B(_0389_),
    .A(_0168_));
 sg13g2_a21o_1 _1302_ (.A2(_0423_),
    .A1(_0390_),
    .B1(net260),
    .X(_0424_));
 sg13g2_nand4_1 _1303_ (.B(_0421_),
    .C(_0422_),
    .A(_0419_),
    .Y(_0425_),
    .D(_0424_));
 sg13g2_nor2b_1 _1304_ (.A(_0394_),
    .B_N(net275),
    .Y(_0426_));
 sg13g2_a221oi_1 _1305_ (.B2(_0425_),
    .C1(_0426_),
    .B1(_0403_),
    .A1(_0396_),
    .Y(_0427_),
    .A2(_0398_));
 sg13g2_a21oi_1 _1306_ (.A1(\bitmap_xofs[0] ),
    .A2(_0218_),
    .Y(_0428_),
    .B1(_0249_));
 sg13g2_nand4_1 _1307_ (.B(_0407_),
    .C(_0422_),
    .A(_0405_),
    .Y(_0429_),
    .D(_0428_));
 sg13g2_nor4_1 _1308_ (.A(_0395_),
    .B(_0402_),
    .C(_0418_),
    .D(_0429_),
    .Y(_0430_));
 sg13g2_xnor2_1 _1309_ (.Y(_0431_),
    .A(_0246_),
    .B(_0393_));
 sg13g2_nor4_1 _1310_ (.A(_0388_),
    .B(_0427_),
    .C(_0430_),
    .D(_0431_),
    .Y(_0004_));
 sg13g2_nand2_1 _1311_ (.Y(_0432_),
    .A(net243),
    .B(_0258_));
 sg13g2_a21oi_2 _1312_ (.B1(net239),
    .Y(_0433_),
    .A2(_0258_),
    .A1(net243));
 sg13g2_nor2_1 _1313_ (.A(_0038_),
    .B(_0433_),
    .Y(_0434_));
 sg13g2_xnor2_1 _1314_ (.Y(_0435_),
    .A(net231),
    .B(_0434_));
 sg13g2_o21ai_1 _1315_ (.B1(_0049_),
    .Y(_0436_),
    .A1(_0120_),
    .A2(_0435_));
 sg13g2_nand2_1 _1316_ (.Y(_0437_),
    .A(_0120_),
    .B(_0435_));
 sg13g2_xnor2_1 _1317_ (.Y(_0438_),
    .A(net234),
    .B(_0433_));
 sg13g2_xor2_1 _1318_ (.B(_0433_),
    .A(net234),
    .X(_0439_));
 sg13g2_nand2_1 _1319_ (.Y(_0440_),
    .A(net266),
    .B(_0438_));
 sg13g2_xnor2_1 _1320_ (.Y(_0441_),
    .A(_0132_),
    .B(_0432_));
 sg13g2_nor2b_1 _1321_ (.A(_0441_),
    .B_N(net268),
    .Y(_0442_));
 sg13g2_and3_1 _1322_ (.X(_0443_),
    .A(_0128_),
    .B(_0055_),
    .C(_0256_));
 sg13g2_a21oi_1 _1323_ (.A1(_0055_),
    .A2(_0256_),
    .Y(_0444_),
    .B1(_0128_));
 sg13g2_o21ai_1 _1324_ (.B1(net271),
    .Y(_0445_),
    .A1(_0443_),
    .A2(_0444_));
 sg13g2_xor2_1 _1325_ (.B(_0256_),
    .A(_0055_),
    .X(_0446_));
 sg13g2_xnor2_1 _1326_ (.Y(_0447_),
    .A(_0137_),
    .B(_0446_));
 sg13g2_or3_1 _1327_ (.A(net271),
    .B(_0443_),
    .C(_0444_),
    .X(_0448_));
 sg13g2_nand3_1 _1328_ (.B(_0447_),
    .C(_0448_),
    .A(_0445_),
    .Y(_0449_));
 sg13g2_nor2_1 _1329_ (.A(\hvsync_gen.vpos[0] ),
    .B(_0125_),
    .Y(_0450_));
 sg13g2_xnor2_1 _1330_ (.Y(_0451_),
    .A(_0054_),
    .B(_0261_));
 sg13g2_or2_1 _1331_ (.X(_0452_),
    .B(_0451_),
    .A(_0450_));
 sg13g2_o21ai_1 _1332_ (.B1(_0452_),
    .Y(_0453_),
    .A1(_0123_),
    .A2(_0261_));
 sg13g2_nand4_1 _1333_ (.B(_0447_),
    .C(_0448_),
    .A(_0445_),
    .Y(_0454_),
    .D(_0453_));
 sg13g2_o21ai_1 _1334_ (.B1(_0445_),
    .Y(_0455_),
    .A1(_0122_),
    .A2(_0446_));
 sg13g2_a22oi_1 _1335_ (.Y(_0456_),
    .B1(_0448_),
    .B2(_0455_),
    .A2(_0260_),
    .A1(_0136_));
 sg13g2_xnor2_1 _1336_ (.Y(_0457_),
    .A(_0050_),
    .B(_0441_));
 sg13g2_xnor2_1 _1337_ (.Y(_0458_),
    .A(net270),
    .B(_0259_));
 sg13g2_a221oi_1 _1338_ (.B2(_0456_),
    .C1(_0457_),
    .B1(_0454_),
    .A1(net269),
    .Y(_0459_),
    .A2(_0259_));
 sg13g2_xnor2_1 _1339_ (.Y(_0460_),
    .A(_0033_),
    .B(_0438_));
 sg13g2_o21ai_1 _1340_ (.B1(_0460_),
    .Y(_0461_),
    .A1(_0442_),
    .A2(_0459_));
 sg13g2_a22oi_1 _1341_ (.Y(_0462_),
    .B1(_0440_),
    .B2(_0461_),
    .A2(_0435_),
    .A1(_0120_));
 sg13g2_nand2_1 _1342_ (.Y(_0463_),
    .A(net235),
    .B(net231));
 sg13g2_o21ai_1 _1343_ (.B1(_0048_),
    .Y(_0464_),
    .A1(_0433_),
    .A2(_0463_));
 sg13g2_xnor2_1 _1344_ (.Y(_0465_),
    .A(_0135_),
    .B(_0464_));
 sg13g2_o21ai_1 _1345_ (.B1(_0465_),
    .Y(_0466_),
    .A1(_0436_),
    .A2(_0462_));
 sg13g2_nor2b_1 _1346_ (.A(net255),
    .B_N(net273),
    .Y(_0467_));
 sg13g2_nor4_1 _1347_ (.A(_0449_),
    .B(_0450_),
    .C(_0451_),
    .D(_0467_),
    .Y(_0468_));
 sg13g2_nand4_1 _1348_ (.B(_0437_),
    .C(_0460_),
    .A(_0047_),
    .Y(_0469_),
    .D(_0468_));
 sg13g2_or4_1 _1349_ (.A(_0436_),
    .B(_0457_),
    .C(_0458_),
    .D(_0469_),
    .X(_0470_));
 sg13g2_nand2b_1 _1350_ (.Y(_0471_),
    .B(_0470_),
    .A_N(_0464_));
 sg13g2_a21oi_1 _1351_ (.A1(net239),
    .A2(net231),
    .Y(_0472_),
    .B1(net235));
 sg13g2_nand2b_1 _1352_ (.Y(_0473_),
    .B(_0463_),
    .A_N(_0472_));
 sg13g2_nor2b_1 _1353_ (.A(_0291_),
    .B_N(_0473_),
    .Y(_0474_));
 sg13g2_nand2_1 _1354_ (.Y(_0475_),
    .A(net234),
    .B(_0283_));
 sg13g2_nand2b_1 _1355_ (.Y(_0476_),
    .B(net238),
    .A_N(net242));
 sg13g2_nor2b_1 _1356_ (.A(net242),
    .B_N(net245),
    .Y(_0477_));
 sg13g2_nor2_1 _1357_ (.A(net242),
    .B(net245),
    .Y(_0478_));
 sg13g2_o21ai_1 _1358_ (.B1(_0476_),
    .Y(_0479_),
    .A1(net238),
    .A2(_0477_));
 sg13g2_inv_1 _1359_ (.Y(_0480_),
    .A(_0479_));
 sg13g2_nand2_1 _1360_ (.Y(_0481_),
    .A(net238),
    .B(_0478_));
 sg13g2_nand2_1 _1361_ (.Y(_0482_),
    .A(_0479_),
    .B(_0481_));
 sg13g2_nor3_1 _1362_ (.A(_0157_),
    .B(_0257_),
    .C(_0477_),
    .Y(_0483_));
 sg13g2_nand2_1 _1363_ (.Y(_0484_),
    .A(net242),
    .B(_0257_));
 sg13g2_nand2b_1 _1364_ (.Y(_0485_),
    .B(_0484_),
    .A_N(_0483_));
 sg13g2_xor2_1 _1365_ (.B(net245),
    .A(net247),
    .X(_0486_));
 sg13g2_nor2_1 _1366_ (.A(_0214_),
    .B(_0486_),
    .Y(_0487_));
 sg13g2_a21oi_1 _1367_ (.A1(_0484_),
    .A2(_0487_),
    .Y(_0488_),
    .B1(_0483_));
 sg13g2_o21ai_1 _1368_ (.B1(_0479_),
    .Y(_0489_),
    .A1(_0482_),
    .A2(_0488_));
 sg13g2_a21oi_1 _1369_ (.A1(_0151_),
    .A2(_0304_),
    .Y(_0490_),
    .B1(_0283_));
 sg13g2_mux2_1 _1370_ (.A0(net249),
    .A1(_0215_),
    .S(_0256_),
    .X(_0491_));
 sg13g2_nor2_1 _1371_ (.A(net228),
    .B(_0261_),
    .Y(_0492_));
 sg13g2_nor4_2 _1372_ (.A(net228),
    .B(_0181_),
    .C(_0215_),
    .Y(_0493_),
    .D(_0255_));
 sg13g2_or2_2 _1373_ (.X(_0494_),
    .B(_0493_),
    .A(_0156_));
 sg13g2_a221oi_1 _1374_ (.B2(_0439_),
    .C1(_0490_),
    .B1(_0494_),
    .A1(_0475_),
    .Y(_0495_),
    .A2(_0489_));
 sg13g2_o21ai_1 _1375_ (.B1(_0473_),
    .Y(_0496_),
    .A1(_0291_),
    .A2(_0495_));
 sg13g2_nor2b_1 _1376_ (.A(net235),
    .B_N(net232),
    .Y(_0497_));
 sg13g2_xnor2_1 _1377_ (.Y(_0498_),
    .A(_0129_),
    .B(_0497_));
 sg13g2_nand2_1 _1378_ (.Y(_0499_),
    .A(_0496_),
    .B(_0498_));
 sg13g2_nand3_1 _1379_ (.B(_0463_),
    .C(_0499_),
    .A(_0129_),
    .Y(_0500_));
 sg13g2_xnor2_1 _1380_ (.Y(_0501_),
    .A(_0474_),
    .B(_0495_));
 sg13g2_or2_1 _1381_ (.X(_0502_),
    .B(_0501_),
    .A(_0049_));
 sg13g2_a21oi_1 _1382_ (.A1(net245),
    .A2(_0214_),
    .Y(_0503_),
    .B1(_0487_));
 sg13g2_a21oi_1 _1383_ (.A1(_0494_),
    .A2(_0503_),
    .Y(_0504_),
    .B1(_0487_));
 sg13g2_xnor2_1 _1384_ (.Y(_0505_),
    .A(_0485_),
    .B(_0504_));
 sg13g2_xor2_1 _1385_ (.B(_0503_),
    .A(_0494_),
    .X(_0506_));
 sg13g2_or2_1 _1386_ (.X(_0507_),
    .B(_0506_),
    .A(net269));
 sg13g2_and2_1 _1387_ (.A(net269),
    .B(_0506_),
    .X(_0508_));
 sg13g2_xnor2_1 _1388_ (.Y(_0509_),
    .A(_0491_),
    .B(_0492_));
 sg13g2_a21o_1 _1389_ (.A2(net228),
    .A1(_0127_),
    .B1(_0492_),
    .X(_0510_));
 sg13g2_or2_1 _1390_ (.X(_0511_),
    .B(_0510_),
    .A(_0137_));
 sg13g2_a21oi_1 _1391_ (.A1(_0137_),
    .A2(_0510_),
    .Y(_0512_),
    .B1(_0327_));
 sg13g2_a21oi_1 _1392_ (.A1(_0121_),
    .A2(_0509_),
    .Y(_0513_),
    .B1(_0512_));
 sg13g2_nor2_1 _1393_ (.A(_0121_),
    .B(_0509_),
    .Y(_0514_));
 sg13g2_a21oi_1 _1394_ (.A1(_0511_),
    .A2(_0513_),
    .Y(_0515_),
    .B1(_0514_));
 sg13g2_a21oi_1 _1395_ (.A1(_0507_),
    .A2(_0515_),
    .Y(_0516_),
    .B1(_0508_));
 sg13g2_xnor2_1 _1396_ (.Y(_0517_),
    .A(_0050_),
    .B(_0505_));
 sg13g2_a22oi_1 _1397_ (.Y(_0518_),
    .B1(_0516_),
    .B2(_0517_),
    .A2(_0505_),
    .A1(net268));
 sg13g2_o21ai_1 _1398_ (.B1(_0207_),
    .Y(_0519_),
    .A1(_0156_),
    .A2(_0493_));
 sg13g2_nand2_1 _1399_ (.Y(_0520_),
    .A(_0488_),
    .B(_0519_));
 sg13g2_xor2_1 _1400_ (.B(_0520_),
    .A(_0482_),
    .X(_0521_));
 sg13g2_xor2_1 _1401_ (.B(_0521_),
    .A(_0033_),
    .X(_0522_));
 sg13g2_a21oi_1 _1402_ (.A1(net234),
    .A2(_0283_),
    .Y(_0523_),
    .B1(_0490_));
 sg13g2_a21oi_1 _1403_ (.A1(_0481_),
    .A2(_0520_),
    .Y(_0524_),
    .B1(_0480_));
 sg13g2_xor2_1 _1404_ (.B(_0524_),
    .A(_0523_),
    .X(_0525_));
 sg13g2_a22oi_1 _1405_ (.Y(_0526_),
    .B1(_0525_),
    .B2(net264),
    .A2(_0521_),
    .A1(net265));
 sg13g2_o21ai_1 _1406_ (.B1(_0526_),
    .Y(_0527_),
    .A1(_0518_),
    .A2(_0522_));
 sg13g2_xnor2_1 _1407_ (.Y(_0528_),
    .A(_0496_),
    .B(_0498_));
 sg13g2_nand2_1 _1408_ (.Y(_0529_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_0528_));
 sg13g2_xnor2_1 _1409_ (.Y(_0530_),
    .A(_0135_),
    .B(_0528_));
 sg13g2_o21ai_1 _1410_ (.B1(_0529_),
    .Y(_0531_),
    .A1(_0502_),
    .A2(_0530_));
 sg13g2_nand2b_1 _1411_ (.Y(_0532_),
    .B(_0531_),
    .A_N(_0500_));
 sg13g2_xor2_1 _1412_ (.B(_0501_),
    .A(_0049_),
    .X(_0533_));
 sg13g2_o21ai_1 _1413_ (.B1(_0533_),
    .Y(_0534_),
    .A1(net263),
    .A2(_0525_));
 sg13g2_nor3_1 _1414_ (.A(_0500_),
    .B(_0530_),
    .C(_0534_),
    .Y(_0535_));
 sg13g2_a221oi_1 _1415_ (.B2(_0535_),
    .C1(_0471_),
    .B1(_0527_),
    .A1(_0124_),
    .Y(_0536_),
    .A2(_0466_));
 sg13g2_and2_1 _1416_ (.A(_0532_),
    .B(_0536_),
    .X(_0005_));
 sg13g2_nand2b_1 _1417_ (.Y(_0537_),
    .B(net275),
    .A_N(net233));
 sg13g2_xor2_1 _1418_ (.B(net233),
    .A(net275),
    .X(_0538_));
 sg13g2_nand2b_1 _1419_ (.Y(_0539_),
    .B(net277),
    .A_N(net237));
 sg13g2_nand2_1 _1420_ (.Y(_0540_),
    .A(_0119_),
    .B(net237));
 sg13g2_nand2b_1 _1421_ (.Y(_0541_),
    .B(net280),
    .A_N(net240));
 sg13g2_nand2b_1 _1422_ (.Y(_0542_),
    .B(_0540_),
    .A_N(_0541_));
 sg13g2_nand2_1 _1423_ (.Y(_0543_),
    .A(net260),
    .B(net241));
 sg13g2_nor2_1 _1424_ (.A(net283),
    .B(_0126_),
    .Y(_0544_));
 sg13g2_nor2_1 _1425_ (.A(_0116_),
    .B(net250),
    .Y(_0545_));
 sg13g2_nand2b_1 _1426_ (.Y(_0546_),
    .B(net286),
    .A_N(net253));
 sg13g2_nor2b_1 _1427_ (.A(net285),
    .B_N(net253),
    .Y(_0547_));
 sg13g2_xnor2_1 _1428_ (.Y(_0548_),
    .A(net285),
    .B(net253));
 sg13g2_o21ai_1 _1429_ (.B1(_0546_),
    .Y(_0549_),
    .A1(_0208_),
    .A2(_0547_));
 sg13g2_xnor2_1 _1430_ (.Y(_0550_),
    .A(\hvsync_gen.hpos[3] ),
    .B(net250));
 sg13g2_a21oi_1 _1431_ (.A1(_0549_),
    .A2(_0550_),
    .Y(_0551_),
    .B1(_0545_));
 sg13g2_a221oi_1 _1432_ (.B2(_0550_),
    .C1(_0545_),
    .B1(_0549_),
    .A1(net283),
    .Y(_0552_),
    .A2(_0126_));
 sg13g2_nor2_1 _1433_ (.A(_0117_),
    .B(net246),
    .Y(_0553_));
 sg13g2_xnor2_1 _1434_ (.Y(_0554_),
    .A(\bitmap_xofs[1] ),
    .B(net246));
 sg13g2_inv_1 _1435_ (.Y(_0555_),
    .A(_0554_));
 sg13g2_nor3_1 _1436_ (.A(_0544_),
    .B(_0552_),
    .C(_0555_),
    .Y(_0556_));
 sg13g2_nor2_1 _1437_ (.A(net260),
    .B(net241),
    .Y(_0557_));
 sg13g2_xnor2_1 _1438_ (.Y(_0558_),
    .A(net282),
    .B(net241));
 sg13g2_nand2_1 _1439_ (.Y(_0559_),
    .A(_0554_),
    .B(_0558_));
 sg13g2_nor3_1 _1440_ (.A(_0544_),
    .B(_0552_),
    .C(_0559_),
    .Y(_0560_));
 sg13g2_a21oi_1 _1441_ (.A1(_0543_),
    .A2(_0553_),
    .Y(_0561_),
    .B1(_0557_));
 sg13g2_nor2b_1 _1442_ (.A(_0560_),
    .B_N(_0561_),
    .Y(_0562_));
 sg13g2_nand3_1 _1443_ (.B(_0542_),
    .C(_0561_),
    .A(_0539_),
    .Y(_0563_));
 sg13g2_nor2b_1 _1444_ (.A(net280),
    .B_N(net240),
    .Y(_0564_));
 sg13g2_nand2_1 _1445_ (.Y(_0565_),
    .A(_0539_),
    .B(_0564_));
 sg13g2_and2_1 _1446_ (.A(_0540_),
    .B(_0565_),
    .X(_0566_));
 sg13g2_o21ai_1 _1447_ (.B1(_0566_),
    .Y(_0567_),
    .A1(_0560_),
    .A2(_0563_));
 sg13g2_o21ai_1 _1448_ (.B1(_0537_),
    .Y(_0568_),
    .A1(_0538_),
    .A2(_0567_));
 sg13g2_nand2_1 _1449_ (.Y(_0569_),
    .A(_0048_),
    .B(_0568_));
 sg13g2_and3_1 _1450_ (.X(_0570_),
    .A(_0048_),
    .B(_0247_),
    .C(_0568_));
 sg13g2_nor2_1 _1451_ (.A(_0048_),
    .B(_0568_),
    .Y(_0571_));
 sg13g2_xor2_1 _1452_ (.B(_0567_),
    .A(_0538_),
    .X(_0572_));
 sg13g2_nor2_1 _1453_ (.A(_0201_),
    .B(_0572_),
    .Y(_0573_));
 sg13g2_nor3_1 _1454_ (.A(_0570_),
    .B(_0571_),
    .C(_0573_),
    .Y(_0574_));
 sg13g2_and2_1 _1455_ (.A(_0539_),
    .B(_0540_),
    .X(_0575_));
 sg13g2_xnor2_1 _1456_ (.Y(_0576_),
    .A(net280),
    .B(net240));
 sg13g2_o21ai_1 _1457_ (.B1(_0541_),
    .Y(_0577_),
    .A1(_0562_),
    .A2(_0564_));
 sg13g2_xnor2_1 _1458_ (.Y(_0578_),
    .A(_0575_),
    .B(_0577_));
 sg13g2_or2_1 _1459_ (.X(_0579_),
    .B(_0578_),
    .A(_0162_));
 sg13g2_nand2_1 _1460_ (.Y(_0580_),
    .A(_0201_),
    .B(_0572_));
 sg13g2_nand2_1 _1461_ (.Y(_0581_),
    .A(_0579_),
    .B(_0580_));
 sg13g2_a22oi_1 _1462_ (.Y(_0582_),
    .B1(_0578_),
    .B2(_0162_),
    .A2(_0569_),
    .A1(_0246_));
 sg13g2_and4_1 _1463_ (.A(_0574_),
    .B(_0579_),
    .C(_0580_),
    .D(_0582_),
    .X(_0583_));
 sg13g2_xnor2_1 _1464_ (.Y(_0584_),
    .A(_0562_),
    .B(_0576_));
 sg13g2_or2_1 _1465_ (.X(_0585_),
    .B(_0584_),
    .A(_0165_));
 sg13g2_inv_1 _1466_ (.Y(_0586_),
    .A(_0585_));
 sg13g2_nor2_1 _1467_ (.A(_0553_),
    .B(_0556_),
    .Y(_0587_));
 sg13g2_xnor2_1 _1468_ (.Y(_0588_),
    .A(_0558_),
    .B(_0587_));
 sg13g2_a22oi_1 _1469_ (.Y(_0589_),
    .B1(_0588_),
    .B2(_0169_),
    .A2(_0584_),
    .A1(_0165_));
 sg13g2_o21ai_1 _1470_ (.B1(_0555_),
    .Y(_0590_),
    .A1(_0544_),
    .A2(_0552_));
 sg13g2_nand2b_1 _1471_ (.Y(_0591_),
    .B(_0590_),
    .A_N(_0556_));
 sg13g2_and2_1 _1472_ (.A(_0172_),
    .B(_0591_),
    .X(_0592_));
 sg13g2_xor2_1 _1473_ (.B(net247),
    .A(\bitmap_xofs[0] ),
    .X(_0593_));
 sg13g2_xnor2_1 _1474_ (.Y(_0594_),
    .A(_0551_),
    .B(_0593_));
 sg13g2_or2_1 _1475_ (.X(_0595_),
    .B(_0594_),
    .A(_0176_));
 sg13g2_o21ai_1 _1476_ (.B1(_0595_),
    .Y(_0596_),
    .A1(_0172_),
    .A2(_0591_));
 sg13g2_or2_1 _1477_ (.X(_0597_),
    .B(_0588_),
    .A(_0169_));
 sg13g2_nand3b_1 _1478_ (.B(_0596_),
    .C(_0597_),
    .Y(_0598_),
    .A_N(_0592_));
 sg13g2_a21oi_1 _1479_ (.A1(_0589_),
    .A2(_0598_),
    .Y(_0599_),
    .B1(_0586_));
 sg13g2_and2_1 _1480_ (.A(_0176_),
    .B(_0594_),
    .X(_0600_));
 sg13g2_nor3_1 _1481_ (.A(_0592_),
    .B(_0596_),
    .C(_0600_),
    .Y(_0601_));
 sg13g2_nand4_1 _1482_ (.B(_0589_),
    .C(_0597_),
    .A(_0585_),
    .Y(_0602_),
    .D(_0601_));
 sg13g2_xor2_1 _1483_ (.B(_0550_),
    .A(_0549_),
    .X(_0603_));
 sg13g2_or2_1 _1484_ (.X(_0604_),
    .B(_0603_),
    .A(_0179_));
 sg13g2_xnor2_1 _1485_ (.Y(_0605_),
    .A(_0208_),
    .B(_0548_));
 sg13g2_a22oi_1 _1486_ (.Y(_0606_),
    .B1(_0605_),
    .B2(_0182_),
    .A2(_0603_),
    .A1(_0179_));
 sg13g2_a21oi_1 _1487_ (.A1(net227),
    .A2(_0209_),
    .Y(_0607_),
    .B1(_0211_));
 sg13g2_nor2_1 _1488_ (.A(_0182_),
    .B(_0605_),
    .Y(_0608_));
 sg13g2_o21ai_1 _1489_ (.B1(_0606_),
    .Y(_0609_),
    .A1(_0607_),
    .A2(_0608_));
 sg13g2_nand2_1 _1490_ (.Y(_0610_),
    .A(_0604_),
    .B(_0606_));
 sg13g2_nand2_1 _1491_ (.Y(_0611_),
    .A(_0604_),
    .B(_0609_));
 sg13g2_nor2_1 _1492_ (.A(_0602_),
    .B(_0611_),
    .Y(_0612_));
 sg13g2_o21ai_1 _1493_ (.B1(_0583_),
    .Y(_0613_),
    .A1(_0599_),
    .A2(_0612_));
 sg13g2_a22oi_1 _1494_ (.Y(_0614_),
    .B1(_0574_),
    .B2(_0581_),
    .A2(_0569_),
    .A1(_0246_));
 sg13g2_nand2b_1 _1495_ (.Y(_0615_),
    .B(_0249_),
    .A_N(_0210_));
 sg13g2_nor4_2 _1496_ (.A(_0602_),
    .B(_0608_),
    .C(_0610_),
    .Y(_0616_),
    .D(_0615_));
 sg13g2_a221oi_1 _1497_ (.B2(_0583_),
    .C1(_0245_),
    .B1(_0616_),
    .A1(_0613_),
    .Y(_0002_),
    .A2(_0614_));
 sg13g2_nor2_1 _1498_ (.A(_0124_),
    .B(net231),
    .Y(_0617_));
 sg13g2_xnor2_1 _1499_ (.Y(_0618_),
    .A(\hvsync_gen.vpos[9] ),
    .B(net231));
 sg13g2_nor2b_1 _1500_ (.A(net234),
    .B_N(\bitmap_yofs[4] ),
    .Y(_0619_));
 sg13g2_inv_1 _1501_ (.Y(_0620_),
    .A(_0619_));
 sg13g2_nor2b_1 _1502_ (.A(net263),
    .B_N(net239),
    .Y(_0621_));
 sg13g2_nor2b_1 _1503_ (.A(\bitmap_yofs[4] ),
    .B_N(net234),
    .Y(_0622_));
 sg13g2_nand2b_1 _1504_ (.Y(_0623_),
    .B(net263),
    .A_N(net239));
 sg13g2_nor2b_1 _1505_ (.A(net243),
    .B_N(net265),
    .Y(_0624_));
 sg13g2_nand2b_1 _1506_ (.Y(_0625_),
    .B(net243),
    .A_N(net265));
 sg13g2_nor2b_1 _1507_ (.A(net245),
    .B_N(net267),
    .Y(_0626_));
 sg13g2_nor2_1 _1508_ (.A(\bitmap_yofs[0] ),
    .B(_0126_),
    .Y(_0627_));
 sg13g2_nor2_1 _1509_ (.A(_0121_),
    .B(net252),
    .Y(_0628_));
 sg13g2_nand2b_1 _1510_ (.Y(_0629_),
    .B(\hvsync_gen.vpos[2] ),
    .A_N(net255));
 sg13g2_nor2b_1 _1511_ (.A(\hvsync_gen.vpos[2] ),
    .B_N(net255),
    .Y(_0630_));
 sg13g2_xnor2_1 _1512_ (.Y(_0631_),
    .A(\hvsync_gen.vpos[2] ),
    .B(net255));
 sg13g2_o21ai_1 _1513_ (.B1(_0629_),
    .Y(_0632_),
    .A1(_0263_),
    .A2(_0630_));
 sg13g2_xnor2_1 _1514_ (.Y(_0633_),
    .A(net271),
    .B(net252));
 sg13g2_a21oi_1 _1515_ (.A1(_0632_),
    .A2(_0633_),
    .Y(_0634_),
    .B1(_0628_));
 sg13g2_a221oi_1 _1516_ (.B2(_0633_),
    .C1(_0628_),
    .B1(_0632_),
    .A1(\bitmap_yofs[0] ),
    .Y(_0635_),
    .A2(_0126_));
 sg13g2_nor2_1 _1517_ (.A(_0627_),
    .B(_0635_),
    .Y(_0636_));
 sg13g2_xnor2_1 _1518_ (.Y(_0637_),
    .A(net267),
    .B(\v_offset[4] ));
 sg13g2_a21oi_1 _1519_ (.A1(_0636_),
    .A2(_0637_),
    .Y(_0638_),
    .B1(_0626_));
 sg13g2_nor2b_1 _1520_ (.A(_0624_),
    .B_N(_0625_),
    .Y(_0639_));
 sg13g2_nand2_1 _1521_ (.Y(_0640_),
    .A(_0637_),
    .B(_0639_));
 sg13g2_or3_1 _1522_ (.A(_0627_),
    .B(_0635_),
    .C(_0640_),
    .X(_0641_));
 sg13g2_a21o_1 _1523_ (.A2(_0626_),
    .A1(_0625_),
    .B1(_0624_),
    .X(_0642_));
 sg13g2_nor2b_1 _1524_ (.A(_0642_),
    .B_N(_0641_),
    .Y(_0643_));
 sg13g2_nor2_1 _1525_ (.A(_0622_),
    .B(_0623_),
    .Y(_0644_));
 sg13g2_nor3_1 _1526_ (.A(_0619_),
    .B(_0642_),
    .C(_0644_),
    .Y(_0645_));
 sg13g2_a221oi_1 _1527_ (.B2(_0645_),
    .C1(_0622_),
    .B1(_0641_),
    .A1(_0620_),
    .Y(_0646_),
    .A2(_0621_));
 sg13g2_a21oi_1 _1528_ (.A1(_0618_),
    .A2(_0646_),
    .Y(_0647_),
    .B1(_0617_));
 sg13g2_nand2b_1 _1529_ (.Y(_0648_),
    .B(_0048_),
    .A_N(_0647_));
 sg13g2_nand2b_1 _1530_ (.Y(_0649_),
    .B(_0648_),
    .A_N(_0344_));
 sg13g2_nand2b_1 _1531_ (.Y(_0650_),
    .B(_0344_),
    .A_N(_0648_));
 sg13g2_xor2_1 _1532_ (.B(_0646_),
    .A(_0618_),
    .X(_0651_));
 sg13g2_nand2b_1 _1533_ (.Y(_0652_),
    .B(_0647_),
    .A_N(_0048_));
 sg13g2_o21ai_1 _1534_ (.B1(_0652_),
    .Y(_0653_),
    .A1(_0306_),
    .A2(_0651_));
 sg13g2_nand2b_1 _1535_ (.Y(_0654_),
    .B(_0650_),
    .A_N(_0653_));
 sg13g2_nor2_1 _1536_ (.A(_0619_),
    .B(_0622_),
    .Y(_0655_));
 sg13g2_nor2b_1 _1537_ (.A(_0621_),
    .B_N(_0623_),
    .Y(_0656_));
 sg13g2_o21ai_1 _1538_ (.B1(_0623_),
    .Y(_0657_),
    .A1(_0621_),
    .A2(_0643_));
 sg13g2_xnor2_1 _1539_ (.Y(_0658_),
    .A(_0655_),
    .B(_0657_));
 sg13g2_nor2_1 _1540_ (.A(_0308_),
    .B(_0658_),
    .Y(_0659_));
 sg13g2_a21oi_1 _1541_ (.A1(_0306_),
    .A2(_0651_),
    .Y(_0660_),
    .B1(_0659_));
 sg13g2_xnor2_1 _1542_ (.Y(_0661_),
    .A(_0643_),
    .B(_0656_));
 sg13g2_xnor2_1 _1543_ (.Y(_0662_),
    .A(_0638_),
    .B(_0639_));
 sg13g2_a22oi_1 _1544_ (.Y(_0663_),
    .B1(_0662_),
    .B2(_0331_),
    .A2(_0661_),
    .A1(_0313_));
 sg13g2_inv_1 _1545_ (.Y(_0664_),
    .A(_0663_));
 sg13g2_nor2_1 _1546_ (.A(_0331_),
    .B(_0662_),
    .Y(_0665_));
 sg13g2_xnor2_1 _1547_ (.Y(_0666_),
    .A(_0636_),
    .B(_0637_));
 sg13g2_nor2_1 _1548_ (.A(_0334_),
    .B(_0666_),
    .Y(_0667_));
 sg13g2_xnor2_1 _1549_ (.Y(_0668_),
    .A(\bitmap_yofs[0] ),
    .B(net249));
 sg13g2_xnor2_1 _1550_ (.Y(_0669_),
    .A(_0634_),
    .B(_0668_));
 sg13g2_a21oi_1 _1551_ (.A1(_0319_),
    .A2(_0669_),
    .Y(_0670_),
    .B1(_0667_));
 sg13g2_xnor2_1 _1552_ (.Y(_0671_),
    .A(_0632_),
    .B(_0633_));
 sg13g2_nor2_1 _1553_ (.A(_0316_),
    .B(_0671_),
    .Y(_0672_));
 sg13g2_xnor2_1 _1554_ (.Y(_0673_),
    .A(_0263_),
    .B(_0631_));
 sg13g2_nand2b_1 _1555_ (.Y(_0674_),
    .B(_0673_),
    .A_N(_0322_));
 sg13g2_and2_1 _1556_ (.A(_0316_),
    .B(_0671_),
    .X(_0675_));
 sg13g2_xnor2_1 _1557_ (.Y(_0676_),
    .A(_0322_),
    .B(_0673_));
 sg13g2_xor2_1 _1558_ (.B(_0671_),
    .A(_0316_),
    .X(_0677_));
 sg13g2_o21ai_1 _1559_ (.B1(_0266_),
    .Y(_0678_),
    .A1(net227),
    .A2(_0264_));
 sg13g2_nand3_1 _1560_ (.B(_0677_),
    .C(_0678_),
    .A(_0676_),
    .Y(_0679_));
 sg13g2_o21ai_1 _1561_ (.B1(_0679_),
    .Y(_0680_),
    .A1(_0674_),
    .A2(_0675_));
 sg13g2_nor2_1 _1562_ (.A(_0319_),
    .B(_0669_),
    .Y(_0681_));
 sg13g2_and4_1 _1563_ (.A(_0265_),
    .B(_0345_),
    .C(_0676_),
    .D(_0677_),
    .X(_0682_));
 sg13g2_nor2_1 _1564_ (.A(_0681_),
    .B(_0682_),
    .Y(_0683_));
 sg13g2_o21ai_1 _1565_ (.B1(_0683_),
    .Y(_0684_),
    .A1(_0672_),
    .A2(_0680_));
 sg13g2_a221oi_1 _1566_ (.B2(_0684_),
    .C1(_0665_),
    .B1(_0670_),
    .A1(_0334_),
    .Y(_0685_),
    .A2(_0666_));
 sg13g2_nor2_1 _1567_ (.A(_0313_),
    .B(_0661_),
    .Y(_0686_));
 sg13g2_a21oi_1 _1568_ (.A1(_0308_),
    .A2(_0658_),
    .Y(_0687_),
    .B1(_0686_));
 sg13g2_o21ai_1 _1569_ (.B1(_0687_),
    .Y(_0688_),
    .A1(_0664_),
    .A2(_0685_));
 sg13g2_a21o_1 _1570_ (.A2(_0688_),
    .A1(_0660_),
    .B1(_0654_),
    .X(_0689_));
 sg13g2_a21oi_1 _1571_ (.A1(_0649_),
    .A2(_0689_),
    .Y(_0003_),
    .B1(_0301_));
 sg13g2_nor2_1 _1572_ (.A(net287),
    .B(net98),
    .Y(_0690_));
 sg13g2_nor3_1 _1573_ (.A(net100),
    .B(net276),
    .C(_0410_),
    .Y(_0691_));
 sg13g2_nand4_1 _1574_ (.B(net259),
    .C(_0690_),
    .A(_0118_),
    .Y(_0692_),
    .D(_0691_));
 sg13g2_nand4_1 _1575_ (.B(net284),
    .C(net285),
    .A(net287),
    .Y(_0693_),
    .D(net276));
 sg13g2_o21ai_1 _1576_ (.B1(_0692_),
    .Y(_0694_),
    .A1(_0149_),
    .A2(_0693_));
 sg13g2_nor2_1 _1577_ (.A(net274),
    .B(_0694_),
    .Y(_0000_));
 sg13g2_nand2_1 _1578_ (.Y(_0695_),
    .A(net267),
    .B(\bitmap_yofs[0] ));
 sg13g2_nand4_1 _1579_ (.B(net265),
    .C(net267),
    .A(net264),
    .Y(_0696_),
    .D(\bitmap_yofs[0] ));
 sg13g2_a21oi_1 _1580_ (.A1(_0121_),
    .A2(_0122_),
    .Y(_0697_),
    .B1(_0696_));
 sg13g2_nor4_1 _1581_ (.A(net264),
    .B(net265),
    .C(net267),
    .D(\bitmap_yofs[0] ),
    .Y(_0698_));
 sg13g2_nor4_1 _1582_ (.A(net271),
    .B(\hvsync_gen.vpos[2] ),
    .C(net272),
    .D(net273),
    .Y(_0699_));
 sg13g2_a21oi_1 _1583_ (.A1(_0698_),
    .A2(_0699_),
    .Y(_0700_),
    .B1(\hvsync_gen.vpos[9] ));
 sg13g2_nand2b_1 _1584_ (.Y(_0701_),
    .B(_0700_),
    .A_N(\bitmap_yofs[4] ));
 sg13g2_o21ai_1 _1585_ (.B1(_0701_),
    .Y(_0001_),
    .A1(_0141_),
    .A2(_0697_));
 sg13g2_and2_1 _1586_ (.A(net287),
    .B(net98),
    .X(_0702_));
 sg13g2_nand3_1 _1587_ (.B(net285),
    .C(_0702_),
    .A(net284),
    .Y(_0703_));
 sg13g2_nor2b_2 _1588_ (.A(\bitmap_xofs[1] ),
    .B_N(net283),
    .Y(_0704_));
 sg13g2_nand2_1 _1589_ (.Y(_0705_),
    .A(net260),
    .B(_0704_));
 sg13g2_nor4_2 _1590_ (.A(net278),
    .B(_0143_),
    .C(_0703_),
    .Y(_0706_),
    .D(_0705_));
 sg13g2_or4_2 _1591_ (.A(net278),
    .B(_0143_),
    .C(_0703_),
    .D(_0705_),
    .X(_0707_));
 sg13g2_nor2b_2 _1592_ (.A(_0706_),
    .B_N(net288),
    .Y(_0708_));
 sg13g2_nand2_2 _1593_ (.Y(_0709_),
    .A(net288),
    .B(_0707_));
 sg13g2_nand4_1 _1594_ (.B(\hvsync_gen.vpos[2] ),
    .C(net272),
    .A(net271),
    .Y(_0710_),
    .D(net273));
 sg13g2_nor2_1 _1595_ (.A(_0695_),
    .B(_0710_),
    .Y(_0711_));
 sg13g2_nand4_1 _1596_ (.B(net265),
    .C(_0709_),
    .A(net264),
    .Y(_0712_),
    .D(_0711_));
 sg13g2_nand4_1 _1597_ (.B(\hvsync_gen.vpos[2] ),
    .C(\hvsync_gen.vpos[9] ),
    .A(net271),
    .Y(_0713_),
    .D(_0698_));
 sg13g2_or4_1 _1598_ (.A(net272),
    .B(net273),
    .C(\bitmap_yofs[4] ),
    .D(_0713_),
    .X(_0714_));
 sg13g2_o21ai_1 _1599_ (.B1(net288),
    .Y(_0715_),
    .A1(_0707_),
    .A2(_0714_));
 sg13g2_xnor2_1 _1600_ (.Y(_0716_),
    .A(\bitmap_yofs[4] ),
    .B(_0712_));
 sg13g2_nand2b_2 _1601_ (.Y(_0717_),
    .B(_0716_),
    .A_N(_0715_));
 sg13g2_inv_1 _1602_ (.Y(_0088_),
    .A(_0717_));
 sg13g2_and3_1 _1603_ (.X(_0718_),
    .A(net288),
    .B(_0706_),
    .C(_0714_));
 sg13g2_nand3_1 _1604_ (.B(_0706_),
    .C(_0714_),
    .A(net288),
    .Y(_0719_));
 sg13g2_nor3_1 _1605_ (.A(_0033_),
    .B(_0695_),
    .C(_0710_),
    .Y(_0720_));
 sg13g2_nor2b_1 _1606_ (.A(_0711_),
    .B_N(_0033_),
    .Y(_0721_));
 sg13g2_nor3_1 _1607_ (.A(_0719_),
    .B(_0720_),
    .C(_0721_),
    .Y(_0722_));
 sg13g2_a21oi_1 _1608_ (.A1(net265),
    .A2(_0708_),
    .Y(_0723_),
    .B1(_0722_));
 sg13g2_inv_1 _1609_ (.Y(_0086_),
    .A(net225));
 sg13g2_nor2_1 _1610_ (.A(net270),
    .B(_0710_),
    .Y(_0724_));
 sg13g2_xor2_1 _1611_ (.B(_0724_),
    .A(_0050_),
    .X(_0725_));
 sg13g2_nor2_1 _1612_ (.A(_0719_),
    .B(_0725_),
    .Y(_0726_));
 sg13g2_a21oi_2 _1613_ (.B1(_0726_),
    .Y(_0727_),
    .A2(_0708_),
    .A1(net267));
 sg13g2_inv_1 _1614_ (.Y(_0085_),
    .A(_0727_));
 sg13g2_xor2_1 _1615_ (.B(_0720_),
    .A(net97),
    .X(_0728_));
 sg13g2_nor2_1 _1616_ (.A(_0719_),
    .B(_0728_),
    .Y(_0729_));
 sg13g2_a21oi_1 _1617_ (.A1(net264),
    .A2(_0708_),
    .Y(_0730_),
    .B1(_0729_));
 sg13g2_inv_2 _1618_ (.Y(_0087_),
    .A(_0730_));
 sg13g2_nor2_1 _1619_ (.A(net218),
    .B(net223),
    .Y(_0731_));
 sg13g2_nor2_2 _1620_ (.A(net220),
    .B(net222),
    .Y(_0732_));
 sg13g2_nor3_1 _1621_ (.A(net220),
    .B(net218),
    .C(net223),
    .Y(_0733_));
 sg13g2_inv_1 _1622_ (.Y(_0734_),
    .A(_0733_));
 sg13g2_nor2_1 _1623_ (.A(net224),
    .B(_0727_),
    .Y(_0735_));
 sg13g2_nand2_2 _1624_ (.Y(_0736_),
    .A(net220),
    .B(net218));
 sg13g2_nand2_1 _1625_ (.Y(_0737_),
    .A(net223),
    .B(_0735_));
 sg13g2_a21oi_1 _1626_ (.A1(_0734_),
    .A2(_0737_),
    .Y(_0090_),
    .B1(net216));
 sg13g2_and2_1 _1627_ (.A(net270),
    .B(_0710_),
    .X(_0738_));
 sg13g2_nor3_1 _1628_ (.A(_0719_),
    .B(_0724_),
    .C(_0738_),
    .Y(_0739_));
 sg13g2_a21oi_2 _1629_ (.B1(_0739_),
    .Y(_0740_),
    .A2(net226),
    .A1(\bitmap_yofs[0] ));
 sg13g2_inv_2 _1630_ (.Y(_0084_),
    .A(_0740_));
 sg13g2_nand2_1 _1631_ (.Y(_0741_),
    .A(net224),
    .B(_0727_));
 sg13g2_nor2_1 _1632_ (.A(net218),
    .B(net221),
    .Y(_0742_));
 sg13g2_nand2_2 _1633_ (.Y(_0743_),
    .A(_0727_),
    .B(_0084_));
 sg13g2_o21ai_1 _1634_ (.B1(net222),
    .Y(_0744_),
    .A1(net220),
    .A2(_0743_));
 sg13g2_nand3b_1 _1635_ (.B(_0744_),
    .C(net217),
    .Y(_0745_),
    .A_N(_0732_));
 sg13g2_nand2b_1 _1636_ (.Y(_0027_),
    .B(_0745_),
    .A_N(_0090_));
 sg13g2_nand2_2 _1637_ (.Y(_0746_),
    .A(net224),
    .B(net221));
 sg13g2_nor2_2 _1638_ (.A(net218),
    .B(_0084_),
    .Y(_0747_));
 sg13g2_nor2_1 _1639_ (.A(net219),
    .B(_0746_),
    .Y(_0748_));
 sg13g2_nor2_1 _1640_ (.A(_0717_),
    .B(_0748_),
    .Y(_0749_));
 sg13g2_nand2_1 _1641_ (.Y(_0750_),
    .A(_0732_),
    .B(_0747_));
 sg13g2_o21ai_1 _1642_ (.B1(_0750_),
    .Y(_0028_),
    .A1(_0717_),
    .A2(_0748_));
 sg13g2_nor2_1 _1643_ (.A(net225),
    .B(net221),
    .Y(_0751_));
 sg13g2_nor2_1 _1644_ (.A(_0736_),
    .B(net221),
    .Y(_0752_));
 sg13g2_nor2_2 _1645_ (.A(net216),
    .B(_0087_),
    .Y(_0753_));
 sg13g2_nand2_1 _1646_ (.Y(_0754_),
    .A(_0752_),
    .B(_0753_));
 sg13g2_nand2_1 _1647_ (.Y(_0029_),
    .A(_0745_),
    .B(_0754_));
 sg13g2_nand2_1 _1648_ (.Y(_0755_),
    .A(net225),
    .B(net218));
 sg13g2_nor2_1 _1649_ (.A(_0727_),
    .B(_0084_),
    .Y(_0756_));
 sg13g2_nand2_2 _1650_ (.Y(_0757_),
    .A(net218),
    .B(net221));
 sg13g2_nor2_1 _1651_ (.A(net220),
    .B(_0757_),
    .Y(_0758_));
 sg13g2_nor2_1 _1652_ (.A(_0717_),
    .B(_0087_),
    .Y(_0759_));
 sg13g2_o21ai_1 _1653_ (.B1(net215),
    .Y(_0760_),
    .A1(_0752_),
    .A2(_0758_));
 sg13g2_nand2_1 _1654_ (.Y(_0761_),
    .A(net216),
    .B(_0732_));
 sg13g2_nand2_1 _1655_ (.Y(_0762_),
    .A(net216),
    .B(_0733_));
 sg13g2_nor2_2 _1656_ (.A(net224),
    .B(net218),
    .Y(_0763_));
 sg13g2_nor2_2 _1657_ (.A(net216),
    .B(net222),
    .Y(_0764_));
 sg13g2_nand2_1 _1658_ (.Y(_0765_),
    .A(_0763_),
    .B(_0764_));
 sg13g2_nand3_1 _1659_ (.B(_0762_),
    .C(_0765_),
    .A(_0760_),
    .Y(_0008_));
 sg13g2_nor2_1 _1660_ (.A(_0087_),
    .B(_0084_),
    .Y(_0766_));
 sg13g2_nand2b_1 _1661_ (.Y(_0767_),
    .B(_0766_),
    .A_N(_0763_));
 sg13g2_a21oi_1 _1662_ (.A1(_0732_),
    .A2(_0756_),
    .Y(_0768_),
    .B1(_0717_));
 sg13g2_nor2_1 _1663_ (.A(net222),
    .B(_0736_),
    .Y(_0769_));
 sg13g2_a221oi_1 _1664_ (.B2(_0766_),
    .C1(_0769_),
    .B1(_0735_),
    .A1(_0727_),
    .Y(_0770_),
    .A2(_0732_));
 sg13g2_a22oi_1 _1665_ (.Y(_0009_),
    .B1(_0770_),
    .B2(_0717_),
    .A2(_0768_),
    .A1(_0767_));
 sg13g2_nand2_1 _1666_ (.Y(_0771_),
    .A(_0731_),
    .B(_0746_));
 sg13g2_o21ai_1 _1667_ (.B1(_0771_),
    .Y(_0772_),
    .A1(_0737_),
    .A2(_0084_));
 sg13g2_nand2_1 _1668_ (.Y(_0773_),
    .A(_0717_),
    .B(_0772_));
 sg13g2_nand2_1 _1669_ (.Y(_0774_),
    .A(_0756_),
    .B(net215));
 sg13g2_nand3_1 _1670_ (.B(_0732_),
    .C(_0756_),
    .A(net217),
    .Y(_0775_));
 sg13g2_nand3_1 _1671_ (.B(_0774_),
    .C(_0775_),
    .A(_0773_),
    .Y(_0010_));
 sg13g2_and3_1 _1672_ (.X(_0776_),
    .A(net222),
    .B(_0741_),
    .C(_0746_));
 sg13g2_nand2_1 _1673_ (.Y(_0777_),
    .A(_0736_),
    .B(_0776_));
 sg13g2_a21oi_1 _1674_ (.A1(net222),
    .A2(_0752_),
    .Y(_0778_),
    .B1(net216));
 sg13g2_a22oi_1 _1675_ (.Y(_0011_),
    .B1(_0778_),
    .B2(_0750_),
    .A2(_0777_),
    .A1(_0768_));
 sg13g2_nand2_2 _1676_ (.Y(_0779_),
    .A(_0743_),
    .B(_0757_));
 sg13g2_inv_1 _1677_ (.Y(_0780_),
    .A(_0779_));
 sg13g2_nor3_1 _1678_ (.A(net216),
    .B(net224),
    .C(net222),
    .Y(_0781_));
 sg13g2_a22oi_1 _1679_ (.Y(_0782_),
    .B1(_0779_),
    .B2(_0781_),
    .A2(_0753_),
    .A1(_0747_));
 sg13g2_nand2_1 _1680_ (.Y(_0012_),
    .A(_0775_),
    .B(_0782_));
 sg13g2_nand2_1 _1681_ (.Y(_0783_),
    .A(_0755_),
    .B(_0766_));
 sg13g2_o21ai_1 _1682_ (.B1(_0783_),
    .Y(_0784_),
    .A1(_0751_),
    .A2(_0771_));
 sg13g2_nand2_1 _1683_ (.Y(_0785_),
    .A(_0717_),
    .B(_0784_));
 sg13g2_nand2_2 _1684_ (.Y(_0786_),
    .A(net220),
    .B(net221));
 sg13g2_nand3_1 _1685_ (.B(_0759_),
    .C(_0779_),
    .A(_0746_),
    .Y(_0787_));
 sg13g2_nand3_1 _1686_ (.B(_0785_),
    .C(_0787_),
    .A(_0775_),
    .Y(_0013_));
 sg13g2_xnor2_1 _1687_ (.Y(_0788_),
    .A(net224),
    .B(_0742_));
 sg13g2_nand3_1 _1688_ (.B(net215),
    .C(_0788_),
    .A(_0757_),
    .Y(_0789_));
 sg13g2_nand2_1 _1689_ (.Y(_0790_),
    .A(_0731_),
    .B(_0786_));
 sg13g2_nor3_1 _1690_ (.A(_0087_),
    .B(_0747_),
    .C(_0763_),
    .Y(_0791_));
 sg13g2_a21oi_1 _1691_ (.A1(_0731_),
    .A2(_0786_),
    .Y(_0792_),
    .B1(_0791_));
 sg13g2_o21ai_1 _1692_ (.B1(_0789_),
    .Y(_0014_),
    .A1(net217),
    .A2(_0792_));
 sg13g2_o21ai_1 _1693_ (.B1(_0789_),
    .Y(_0015_),
    .A1(_0751_),
    .A2(_0773_));
 sg13g2_nand3_1 _1694_ (.B(_0759_),
    .C(_0786_),
    .A(net219),
    .Y(_0793_));
 sg13g2_nand2_1 _1695_ (.Y(_0016_),
    .A(_0782_),
    .B(_0793_));
 sg13g2_nand2_1 _1696_ (.Y(_0794_),
    .A(net217),
    .B(_0750_));
 sg13g2_nor2_1 _1697_ (.A(_0776_),
    .B(_0794_),
    .Y(_0795_));
 sg13g2_a21oi_1 _1698_ (.A1(_0732_),
    .A2(_0740_),
    .Y(_0796_),
    .B1(net217));
 sg13g2_a21oi_1 _1699_ (.A1(_0783_),
    .A2(_0796_),
    .Y(_0017_),
    .B1(_0795_));
 sg13g2_nor2_1 _1700_ (.A(net224),
    .B(_0743_),
    .Y(_0797_));
 sg13g2_o21ai_1 _1701_ (.B1(net215),
    .Y(_0798_),
    .A1(_0758_),
    .A2(_0797_));
 sg13g2_and2_1 _1702_ (.A(_0754_),
    .B(_0798_),
    .X(_0799_));
 sg13g2_nand2_1 _1703_ (.Y(_0800_),
    .A(_0758_),
    .B(_0764_));
 sg13g2_nand2_1 _1704_ (.Y(_0018_),
    .A(_0799_),
    .B(_0800_));
 sg13g2_nor2_1 _1705_ (.A(net220),
    .B(_0779_),
    .Y(_0801_));
 sg13g2_nand2_1 _1706_ (.Y(_0802_),
    .A(_0753_),
    .B(_0801_));
 sg13g2_nand2_1 _1707_ (.Y(_0803_),
    .A(_0742_),
    .B(net215));
 sg13g2_nand2_1 _1708_ (.Y(_0019_),
    .A(_0802_),
    .B(_0803_));
 sg13g2_xnor2_1 _1709_ (.Y(_0804_),
    .A(net221),
    .B(_0769_));
 sg13g2_o21ai_1 _1710_ (.B1(_0798_),
    .Y(_0020_),
    .A1(net217),
    .A2(_0804_));
 sg13g2_o21ai_1 _1711_ (.B1(net215),
    .Y(_0805_),
    .A1(_0763_),
    .A2(_0801_));
 sg13g2_nand2b_1 _1712_ (.Y(_0806_),
    .B(_0786_),
    .A_N(_0744_));
 sg13g2_o21ai_1 _1713_ (.B1(_0806_),
    .Y(_0807_),
    .A1(net222),
    .A2(net221));
 sg13g2_o21ai_1 _1714_ (.B1(_0805_),
    .Y(_0021_),
    .A1(net216),
    .A2(_0807_));
 sg13g2_a22oi_1 _1715_ (.Y(_0022_),
    .B1(_0778_),
    .B2(_0790_),
    .A2(_0749_),
    .A1(_0737_));
 sg13g2_nor2_1 _1716_ (.A(_0753_),
    .B(_0776_),
    .Y(_0808_));
 sg13g2_nor2_1 _1717_ (.A(net224),
    .B(_0747_),
    .Y(_0809_));
 sg13g2_nor3_1 _1718_ (.A(_0748_),
    .B(_0808_),
    .C(_0809_),
    .Y(_0023_));
 sg13g2_nand2b_1 _1719_ (.Y(_0810_),
    .B(_0753_),
    .A_N(_0746_));
 sg13g2_o21ai_1 _1720_ (.B1(_0764_),
    .Y(_0811_),
    .A1(_0797_),
    .A2(_0801_));
 sg13g2_nand3_1 _1721_ (.B(_0810_),
    .C(_0811_),
    .A(_0799_),
    .Y(_0024_));
 sg13g2_nand3b_1 _1722_ (.B(_0779_),
    .C(_0753_),
    .Y(_0812_),
    .A_N(_0763_));
 sg13g2_nand3_1 _1723_ (.B(_0746_),
    .C(_0764_),
    .A(_0736_),
    .Y(_0813_));
 sg13g2_nand4_1 _1724_ (.B(_0798_),
    .C(_0812_),
    .A(_0762_),
    .Y(_0025_),
    .D(_0813_));
 sg13g2_nand4_1 _1725_ (.B(_0757_),
    .C(_0764_),
    .A(_0736_),
    .Y(_0814_),
    .D(_0786_));
 sg13g2_nand2_1 _1726_ (.Y(_0815_),
    .A(_0741_),
    .B(net215));
 sg13g2_nand3_1 _1727_ (.B(_0743_),
    .C(_0753_),
    .A(_0741_),
    .Y(_0816_));
 sg13g2_nand3_1 _1728_ (.B(_0815_),
    .C(_0816_),
    .A(_0814_),
    .Y(_0026_));
 sg13g2_nor2_2 _1729_ (.A(_0117_),
    .B(net283),
    .Y(_0817_));
 sg13g2_a221oi_1 _1730_ (.B2(\bitsTemp[2] ),
    .C1(net281),
    .B1(_0817_),
    .A1(\bitsTemp[4] ),
    .Y(_0818_),
    .A2(_0147_));
 sg13g2_a22oi_1 _1731_ (.Y(_0819_),
    .B1(_0704_),
    .B2(\bitsTemp[2] ),
    .A2(net259),
    .A1(\bitsTemp[3] ));
 sg13g2_a21oi_1 _1732_ (.A1(net281),
    .A2(_0819_),
    .Y(_0820_),
    .B1(_0818_));
 sg13g2_nand2_1 _1733_ (.Y(_0821_),
    .A(net281),
    .B(_0817_));
 sg13g2_a21oi_1 _1734_ (.A1(_0705_),
    .A2(_0821_),
    .Y(_0822_),
    .B1(_0138_));
 sg13g2_a21oi_1 _1735_ (.A1(\bitsTemp[12] ),
    .A2(net258),
    .Y(_0823_),
    .B1(net281));
 sg13g2_and2_1 _1736_ (.A(\bitsTemp[14] ),
    .B(_0704_),
    .X(_0824_));
 sg13g2_a221oi_1 _1737_ (.B2(\bitsTemp[13] ),
    .C1(_0824_),
    .B1(_0817_),
    .A1(\bitsTemp[15] ),
    .Y(_0825_),
    .A2(net259));
 sg13g2_a22oi_1 _1738_ (.Y(_0826_),
    .B1(_0817_),
    .B2(\bitsTemp[9] ),
    .A2(_0704_),
    .A1(\bitsTemp[10] ));
 sg13g2_a221oi_1 _1739_ (.B2(\bitsTemp[8] ),
    .C1(net260),
    .B1(net258),
    .A1(\bitsTemp[11] ),
    .Y(_0827_),
    .A2(_0144_));
 sg13g2_a221oi_1 _1740_ (.B2(_0827_),
    .C1(net278),
    .B1(_0826_),
    .A1(_0823_),
    .Y(_0828_),
    .A2(_0825_));
 sg13g2_o21ai_1 _1741_ (.B1(net278),
    .Y(_0829_),
    .A1(_0820_),
    .A2(_0822_));
 sg13g2_nand3b_1 _1742_ (.B(_0829_),
    .C(net276),
    .Y(_0830_),
    .A_N(_0828_));
 sg13g2_a22oi_1 _1743_ (.Y(_0831_),
    .B1(_0817_),
    .B2(\bitsTemp[21] ),
    .A2(net259),
    .A1(\bitsTemp[23] ));
 sg13g2_a22oi_1 _1744_ (.Y(_0832_),
    .B1(_0704_),
    .B2(\bitsTemp[22] ),
    .A2(net258),
    .A1(\bitsTemp[20] ));
 sg13g2_nand2_1 _1745_ (.Y(_0833_),
    .A(_0831_),
    .B(_0832_));
 sg13g2_nand3_1 _1746_ (.B(net260),
    .C(_0833_),
    .A(net278),
    .Y(_0834_));
 sg13g2_a22oi_1 _1747_ (.Y(_0835_),
    .B1(_0817_),
    .B2(\bitsTemp[17] ),
    .A2(net258),
    .A1(\bitsTemp[16] ));
 sg13g2_a22oi_1 _1748_ (.Y(_0836_),
    .B1(_0704_),
    .B2(\bitsTemp[18] ),
    .A2(net259),
    .A1(\bitsTemp[19] ));
 sg13g2_nand2_1 _1749_ (.Y(_0837_),
    .A(_0835_),
    .B(_0836_));
 sg13g2_nand3_1 _1750_ (.B(net282),
    .C(_0837_),
    .A(net278),
    .Y(_0838_));
 sg13g2_a22oi_1 _1751_ (.Y(_0839_),
    .B1(_0704_),
    .B2(\bitsTemp[30] ),
    .A2(net259),
    .A1(\bitsTemp[31] ));
 sg13g2_a221oi_1 _1752_ (.B2(\bitsTemp[29] ),
    .C1(net281),
    .B1(_0817_),
    .A1(\bitsTemp[28] ),
    .Y(_0840_),
    .A2(net258));
 sg13g2_a21oi_1 _1753_ (.A1(\bitsTemp[27] ),
    .A2(net259),
    .Y(_0841_),
    .B1(net260));
 sg13g2_nand2_1 _1754_ (.Y(_0842_),
    .A(\bitsTemp[25] ),
    .B(_0817_));
 sg13g2_a22oi_1 _1755_ (.Y(_0843_),
    .B1(_0704_),
    .B2(\bitsTemp[26] ),
    .A2(net258),
    .A1(\bitsTemp[24] ));
 sg13g2_nand3_1 _1756_ (.B(_0842_),
    .C(_0843_),
    .A(_0841_),
    .Y(_0844_));
 sg13g2_a21oi_1 _1757_ (.A1(_0839_),
    .A2(_0840_),
    .Y(_0845_),
    .B1(net278));
 sg13g2_a21oi_1 _1758_ (.A1(_0844_),
    .A2(_0845_),
    .Y(_0846_),
    .B1(net276));
 sg13g2_nand3_1 _1759_ (.B(_0838_),
    .C(_0846_),
    .A(_0834_),
    .Y(_0847_));
 sg13g2_nand4_1 _1760_ (.B(bmpOnV),
    .C(_0830_),
    .A(bmpOnH),
    .Y(_0848_),
    .D(_0847_));
 sg13g2_nand4_1 _1761_ (.B(net265),
    .C(net267),
    .A(net264),
    .Y(_0849_),
    .D(\bitmap_yofs[4] ));
 sg13g2_o21ai_1 _1762_ (.B1(net275),
    .Y(_0850_),
    .A1(net280),
    .A2(net277));
 sg13g2_and3_1 _1763_ (.X(_0851_),
    .A(_0124_),
    .B(_0849_),
    .C(_0850_));
 sg13g2_nand3_1 _1764_ (.B(test_h),
    .C(_0851_),
    .A(test_v),
    .Y(_0852_));
 sg13g2_xor2_1 _1765_ (.B(_0852_),
    .A(_0848_),
    .X(r));
 sg13g2_nand3_1 _1766_ (.B(test_g_v),
    .C(_0851_),
    .A(test_g_h),
    .Y(_0853_));
 sg13g2_xor2_1 _1767_ (.B(_0853_),
    .A(_0848_),
    .X(g));
 sg13g2_nand3_1 _1768_ (.B(test_b_v),
    .C(_0851_),
    .A(test_b_h),
    .Y(_0854_));
 sg13g2_xor2_1 _1769_ (.B(_0854_),
    .A(_0848_),
    .X(b));
 sg13g2_xnor2_1 _1770_ (.Y(_0855_),
    .A(_0067_),
    .B(net230));
 sg13g2_xnor2_1 _1771_ (.Y(_0056_),
    .A(net253),
    .B(_0855_));
 sg13g2_nor2_1 _1772_ (.A(_0127_),
    .B(net230),
    .Y(_0856_));
 sg13g2_xnor2_1 _1773_ (.Y(_0857_),
    .A(net250),
    .B(net230));
 sg13g2_a21oi_1 _1774_ (.A1(net230),
    .A2(_0186_),
    .Y(_0858_),
    .B1(net228));
 sg13g2_xor2_1 _1775_ (.B(_0858_),
    .A(_0857_),
    .X(_0057_));
 sg13g2_a21oi_1 _1776_ (.A1(_0857_),
    .A2(_0858_),
    .Y(_0859_),
    .B1(_0856_));
 sg13g2_xnor2_1 _1777_ (.Y(_0860_),
    .A(net247),
    .B(net230));
 sg13g2_xnor2_1 _1778_ (.Y(_0058_),
    .A(_0859_),
    .B(_0860_));
 sg13g2_xor2_1 _1779_ (.B(net229),
    .A(net246),
    .X(_0861_));
 sg13g2_a21oi_1 _1780_ (.A1(_0126_),
    .A2(net230),
    .Y(_0862_),
    .B1(_0859_));
 sg13g2_a21o_1 _1781_ (.A2(_0139_),
    .A1(net247),
    .B1(_0862_),
    .X(_0863_));
 sg13g2_nor2b_1 _1782_ (.A(_0861_),
    .B_N(_0863_),
    .Y(_0864_));
 sg13g2_xnor2_1 _1783_ (.Y(_0059_),
    .A(_0861_),
    .B(_0863_));
 sg13g2_a21oi_1 _1784_ (.A1(net246),
    .A2(_0139_),
    .Y(_0865_),
    .B1(_0864_));
 sg13g2_xnor2_1 _1785_ (.Y(_0866_),
    .A(net242),
    .B(v_offset_rev_flag));
 sg13g2_xnor2_1 _1786_ (.Y(_0060_),
    .A(_0865_),
    .B(_0866_));
 sg13g2_nor2b_1 _1787_ (.A(net230),
    .B_N(net238),
    .Y(_0867_));
 sg13g2_xnor2_1 _1788_ (.Y(_0868_),
    .A(net238),
    .B(v_offset_rev_flag));
 sg13g2_and2_1 _1789_ (.A(_0864_),
    .B(_0866_),
    .X(_0869_));
 sg13g2_nor2_1 _1790_ (.A(net229),
    .B(_0478_),
    .Y(_0870_));
 sg13g2_or2_1 _1791_ (.X(_0871_),
    .B(_0870_),
    .A(_0869_));
 sg13g2_xor2_1 _1792_ (.B(_0871_),
    .A(_0868_),
    .X(_0061_));
 sg13g2_xor2_1 _1793_ (.B(net229),
    .A(net236),
    .X(_0872_));
 sg13g2_inv_1 _1794_ (.Y(_0873_),
    .A(_0872_));
 sg13g2_a21oi_1 _1795_ (.A1(_0868_),
    .A2(_0871_),
    .Y(_0874_),
    .B1(_0867_));
 sg13g2_xnor2_1 _1796_ (.Y(_0062_),
    .A(_0873_),
    .B(_0874_));
 sg13g2_nor2b_1 _1797_ (.A(net229),
    .B_N(net232),
    .Y(_0875_));
 sg13g2_xnor2_1 _1798_ (.Y(_0876_),
    .A(net232),
    .B(net229));
 sg13g2_nand3_1 _1799_ (.B(_0869_),
    .C(_0873_),
    .A(_0868_),
    .Y(_0877_));
 sg13g2_o21ai_1 _1800_ (.B1(_0139_),
    .Y(_0878_),
    .A1(net236),
    .A2(net238));
 sg13g2_nand3b_1 _1801_ (.B(_0877_),
    .C(_0878_),
    .Y(_0879_),
    .A_N(_0870_));
 sg13g2_xor2_1 _1802_ (.B(_0879_),
    .A(_0876_),
    .X(_0063_));
 sg13g2_a21oi_1 _1803_ (.A1(_0876_),
    .A2(_0879_),
    .Y(_0880_),
    .B1(_0875_));
 sg13g2_xnor2_1 _1804_ (.Y(_0881_),
    .A(\v_offset[9] ),
    .B(net229));
 sg13g2_xnor2_1 _1805_ (.Y(_0064_),
    .A(_0880_),
    .B(_0881_));
 sg13g2_o21ai_1 _1806_ (.B1(_0803_),
    .Y(_0068_),
    .A1(_0761_),
    .A2(_0780_));
 sg13g2_nand2_1 _1807_ (.Y(_0069_),
    .A(_0762_),
    .B(_0803_));
 sg13g2_and2_1 _1808_ (.A(net76),
    .B(net226),
    .X(_0070_));
 sg13g2_nor3_1 _1809_ (.A(_0690_),
    .B(_0702_),
    .C(_0709_),
    .Y(_0071_));
 sg13g2_o21ai_1 _1810_ (.B1(net288),
    .Y(_0882_),
    .A1(net285),
    .A2(_0702_));
 sg13g2_a21oi_1 _1811_ (.A1(net285),
    .A2(_0702_),
    .Y(_0072_),
    .B1(_0882_));
 sg13g2_nor2b_1 _1812_ (.A(net79),
    .B_N(_0702_),
    .Y(_0883_));
 sg13g2_xnor2_1 _1813_ (.Y(_0884_),
    .A(net284),
    .B(_0883_));
 sg13g2_nor2_1 _1814_ (.A(_0709_),
    .B(net80),
    .Y(_0073_));
 sg13g2_xor2_1 _1815_ (.B(_0703_),
    .A(net283),
    .X(_0885_));
 sg13g2_nor2_1 _1816_ (.A(_0709_),
    .B(_0885_),
    .Y(_0074_));
 sg13g2_nor2_1 _1817_ (.A(_0043_),
    .B(_0703_),
    .Y(_0886_));
 sg13g2_xnor2_1 _1818_ (.Y(_0887_),
    .A(net92),
    .B(_0886_));
 sg13g2_nor2_1 _1819_ (.A(_0709_),
    .B(net93),
    .Y(_0075_));
 sg13g2_nor2_1 _1820_ (.A(_0148_),
    .B(_0703_),
    .Y(_0888_));
 sg13g2_xnor2_1 _1821_ (.Y(_0889_),
    .A(net281),
    .B(_0888_));
 sg13g2_nor2_1 _1822_ (.A(_0709_),
    .B(_0889_),
    .Y(_0076_));
 sg13g2_nor3_1 _1823_ (.A(net91),
    .B(_0148_),
    .C(_0703_),
    .Y(_0095_));
 sg13g2_o21ai_1 _1824_ (.B1(net226),
    .Y(_0096_),
    .A1(net279),
    .A2(_0095_));
 sg13g2_a21oi_1 _1825_ (.A1(net279),
    .A2(_0095_),
    .Y(_0077_),
    .B1(_0096_));
 sg13g2_nor2_1 _1826_ (.A(_0149_),
    .B(_0703_),
    .Y(_0097_));
 sg13g2_o21ai_1 _1827_ (.B1(net226),
    .Y(_0098_),
    .A1(net276),
    .A2(_0097_));
 sg13g2_a21oi_1 _1828_ (.A1(net276),
    .A2(_0097_),
    .Y(_0078_),
    .B1(_0098_));
 sg13g2_nor3_1 _1829_ (.A(net94),
    .B(_0149_),
    .C(_0703_),
    .Y(_0099_));
 sg13g2_o21ai_1 _1830_ (.B1(net226),
    .Y(_0100_),
    .A1(net275),
    .A2(_0099_));
 sg13g2_a21oi_1 _1831_ (.A1(net274),
    .A2(_0099_),
    .Y(_0079_),
    .B1(_0100_));
 sg13g2_a22oi_1 _1832_ (.Y(_0101_),
    .B1(_0718_),
    .B2(net77),
    .A2(net226),
    .A1(net273));
 sg13g2_inv_1 _1833_ (.Y(_0080_),
    .A(net78));
 sg13g2_nand2_1 _1834_ (.Y(_0102_),
    .A(net272),
    .B(net226));
 sg13g2_xnor2_1 _1835_ (.Y(_0103_),
    .A(net272),
    .B(net273));
 sg13g2_o21ai_1 _1836_ (.B1(_0102_),
    .Y(_0081_),
    .A1(_0719_),
    .A2(_0103_));
 sg13g2_nand3_1 _1837_ (.B(net273),
    .C(_0709_),
    .A(net272),
    .Y(_0104_));
 sg13g2_xnor2_1 _1838_ (.Y(_0105_),
    .A(_0122_),
    .B(_0104_));
 sg13g2_nor2_1 _1839_ (.A(_0715_),
    .B(_0105_),
    .Y(_0082_));
 sg13g2_nand2_1 _1840_ (.Y(_0106_),
    .A(net271),
    .B(net226));
 sg13g2_nand3_1 _1841_ (.B(net273),
    .C(_0137_),
    .A(net272),
    .Y(_0107_));
 sg13g2_xnor2_1 _1842_ (.Y(_0108_),
    .A(_0121_),
    .B(_0107_));
 sg13g2_o21ai_1 _1843_ (.B1(_0106_),
    .Y(_0083_),
    .A1(_0719_),
    .A2(_0108_));
 sg13g2_nor3_1 _1844_ (.A(_0049_),
    .B(_0696_),
    .C(_0710_),
    .Y(_0109_));
 sg13g2_o21ai_1 _1845_ (.B1(_0718_),
    .Y(_0110_),
    .A1(\hvsync_gen.vpos[9] ),
    .A2(_0109_));
 sg13g2_a21o_1 _1846_ (.A2(_0109_),
    .A1(\hvsync_gen.vpos[9] ),
    .B1(_0110_),
    .X(_0111_));
 sg13g2_o21ai_1 _1847_ (.B1(_0111_),
    .Y(_0089_),
    .A1(_0124_),
    .A2(_0709_));
 sg13g2_a221oi_1 _1848_ (.B2(_0087_),
    .C1(_0088_),
    .B1(_0743_),
    .A1(net220),
    .Y(_0091_),
    .A2(_0084_));
 sg13g2_nand3_1 _1849_ (.B(_0755_),
    .C(net215),
    .A(_0084_),
    .Y(_0112_));
 sg13g2_nand2_1 _1850_ (.Y(_0092_),
    .A(_0761_),
    .B(_0112_));
 sg13g2_nor2_1 _1851_ (.A(_0809_),
    .B(_0815_),
    .Y(_0093_));
 sg13g2_nand4_1 _1852_ (.B(_0214_),
    .C(_0241_),
    .A(_0152_),
    .Y(_0113_),
    .D(_0288_));
 sg13g2_nand4_1 _1853_ (.B(net228),
    .C(_0241_),
    .A(net236),
    .Y(_0114_),
    .D(_0350_));
 sg13g2_o21ai_1 _1854_ (.B1(net229),
    .Y(_0115_),
    .A1(_0481_),
    .A2(_0114_));
 sg13g2_nand2_1 _1855_ (.Y(_0094_),
    .A(_0113_),
    .B(_0115_));
 sg13g2_dfrbp_1 _1856_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net20),
    .D(_0068_),
    .Q_N(_0899_),
    .Q(\bitsTemp[3] ));
 sg13g2_dfrbp_1 _1857_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net21),
    .D(_0069_),
    .Q_N(_0900_),
    .Q(\bitsTemp[4] ));
 sg13g2_dfrbp_1 _1858_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net22),
    .D(_0027_),
    .Q_N(_0901_),
    .Q(\bitsTemp[8] ));
 sg13g2_dfrbp_1 _1859_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net23),
    .D(_0028_),
    .Q_N(_0902_),
    .Q(\bitsTemp[9] ));
 sg13g2_dfrbp_1 _1860_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net24),
    .D(_0029_),
    .Q_N(_0903_),
    .Q(\bitsTemp[10] ));
 sg13g2_dfrbp_1 _1861_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net25),
    .D(_0008_),
    .Q_N(_0904_),
    .Q(\bitsTemp[12] ));
 sg13g2_dfrbp_1 _1862_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net26),
    .D(_0009_),
    .Q_N(_0905_),
    .Q(\bitsTemp[13] ));
 sg13g2_dfrbp_1 _1863_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net27),
    .D(_0010_),
    .Q_N(_0906_),
    .Q(\bitsTemp[14] ));
 sg13g2_dfrbp_1 _1864_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net28),
    .D(_0011_),
    .Q_N(_0907_),
    .Q(\bitsTemp[15] ));
 sg13g2_dfrbp_1 _1865_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net29),
    .D(_0012_),
    .Q_N(_0908_),
    .Q(\bitsTemp[16] ));
 sg13g2_dfrbp_1 _1866_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net30),
    .D(_0013_),
    .Q_N(_0909_),
    .Q(\bitsTemp[17] ));
 sg13g2_dfrbp_1 _1867_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net31),
    .D(_0014_),
    .Q_N(_0910_),
    .Q(\bitsTemp[18] ));
 sg13g2_dfrbp_1 _1868_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net32),
    .D(_0015_),
    .Q_N(_0911_),
    .Q(\bitsTemp[19] ));
 sg13g2_dfrbp_1 _1869_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net33),
    .D(_0016_),
    .Q_N(_0912_),
    .Q(\bitsTemp[20] ));
 sg13g2_dfrbp_1 _1870_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net34),
    .D(_0017_),
    .Q_N(_0913_),
    .Q(\bitsTemp[22] ));
 sg13g2_dfrbp_1 _1871_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net35),
    .D(_0018_),
    .Q_N(_0914_),
    .Q(\bitsTemp[23] ));
 sg13g2_dfrbp_1 _1872_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net36),
    .D(_0019_),
    .Q_N(_0915_),
    .Q(\bitsTemp[24] ));
 sg13g2_dfrbp_1 _1873_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net37),
    .D(_0020_),
    .Q_N(_0916_),
    .Q(\bitsTemp[25] ));
 sg13g2_dfrbp_1 _1874_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net38),
    .D(_0021_),
    .Q_N(_0917_),
    .Q(\bitsTemp[26] ));
 sg13g2_dfrbp_1 _1875_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net39),
    .D(_0022_),
    .Q_N(_0918_),
    .Q(\bitsTemp[27] ));
 sg13g2_dfrbp_1 _1876_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net40),
    .D(_0023_),
    .Q_N(_0919_),
    .Q(\bitsTemp[28] ));
 sg13g2_dfrbp_1 _1877_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net41),
    .D(_0024_),
    .Q_N(_0920_),
    .Q(\bitsTemp[29] ));
 sg13g2_dfrbp_1 _1878_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net42),
    .D(_0025_),
    .Q_N(_0921_),
    .Q(\bitsTemp[30] ));
 sg13g2_dfrbp_1 _1879_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net43),
    .D(_0026_),
    .Q_N(_0922_),
    .Q(\bitsTemp[31] ));
 sg13g2_dfrbp_1 _1880_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net44),
    .D(_0001_),
    .Q_N(_0923_),
    .Q(bmpOnV));
 sg13g2_dfrbp_1 _1881_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net45),
    .D(_0000_),
    .Q_N(_0924_),
    .Q(bmpOnH));
 sg13g2_dfrbp_1 _1882_ (.CLK(net261),
    .RESET_B(net288),
    .D(_0067_),
    .Q_N(_0067_),
    .Q(\v_offset[0] ));
 sg13g2_dfrbp_1 _1883_ (.CLK(net261),
    .RESET_B(net289),
    .D(_0056_),
    .Q_N(_0925_),
    .Q(\v_offset[1] ));
 sg13g2_dfrbp_1 _1884_ (.CLK(net261),
    .RESET_B(net289),
    .D(_0057_),
    .Q_N(_0052_),
    .Q(\v_offset[2] ));
 sg13g2_dfrbp_1 _1885_ (.CLK(net261),
    .RESET_B(net288),
    .D(_0058_),
    .Q_N(_0055_),
    .Q(\v_offset[3] ));
 sg13g2_dfrbp_1 _1886_ (.CLK(net261),
    .RESET_B(net1),
    .D(_0059_),
    .Q_N(_0041_),
    .Q(\v_offset[4] ));
 sg13g2_dfrbp_1 _1887_ (.CLK(net261),
    .RESET_B(net1),
    .D(_0060_),
    .Q_N(_0035_),
    .Q(\v_offset[5] ));
 sg13g2_dfrbp_1 _1888_ (.CLK(net262),
    .RESET_B(net289),
    .D(_0061_),
    .Q_N(_0039_),
    .Q(\v_offset[6] ));
 sg13g2_dfrbp_1 _1889_ (.CLK(net262),
    .RESET_B(net289),
    .D(_0062_),
    .Q_N(_0038_),
    .Q(\v_offset[7] ));
 sg13g2_dfrbp_1 _1890_ (.CLK(net262),
    .RESET_B(net289),
    .D(_0063_),
    .Q_N(_0036_),
    .Q(\v_offset[8] ));
 sg13g2_dfrbp_1 _1891_ (.CLK(net261),
    .RESET_B(net289),
    .D(_0064_),
    .Q_N(_0048_),
    .Q(\v_offset[9] ));
 sg13g2_dfrbp_1 _1892_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net65),
    .D(_0070_),
    .Q_N(_0066_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 _1893_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net64),
    .D(_0071_),
    .Q_N(_0045_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _1894_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net63),
    .D(net90),
    .Q_N(_0044_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _1895_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net62),
    .D(_0073_),
    .Q_N(_0898_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _1896_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net61),
    .D(_0074_),
    .Q_N(_0043_),
    .Q(\bitmap_xofs[0] ));
 sg13g2_dfrbp_1 _1897_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net54),
    .D(_0075_),
    .Q_N(_0042_),
    .Q(\bitmap_xofs[1] ));
 sg13g2_dfrbp_1 _1898_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net53),
    .D(_0076_),
    .Q_N(_0040_),
    .Q(\bitmap_xofs[2] ));
 sg13g2_dfrbp_1 _1899_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net52),
    .D(_0077_),
    .Q_N(_0037_),
    .Q(\bitmap_xofs[3] ));
 sg13g2_dfrbp_1 _1900_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net51),
    .D(_0078_),
    .Q_N(_0046_),
    .Q(\bitmap_xofs[4] ));
 sg13g2_dfrbp_1 _1901_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net55),
    .D(net95),
    .Q_N(_0034_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _1902_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net56),
    .D(_0003_),
    .Q_N(_0926_),
    .Q(test_b_v));
 sg13g2_dfrbp_1 _1903_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net57),
    .D(_0002_),
    .Q_N(_0927_),
    .Q(test_b_h));
 sg13g2_dfrbp_1 _1904_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net58),
    .D(_0005_),
    .Q_N(_0928_),
    .Q(test_g_v));
 sg13g2_dfrbp_1 _1905_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net59),
    .D(_0004_),
    .Q_N(_0929_),
    .Q(test_g_h));
 sg13g2_dfrbp_1 _1906_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net60),
    .D(_0007_),
    .Q_N(_0930_),
    .Q(test_v));
 sg13g2_dfrbp_1 _1907_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net70),
    .D(_0006_),
    .Q_N(_0931_),
    .Q(test_h));
 sg13g2_dfrbp_1 _1908_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net50),
    .D(net82),
    .Q_N(_0897_),
    .Q(hsync));
 sg13g2_dfrbp_1 _1909_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net49),
    .D(_0080_),
    .Q_N(_0065_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _1910_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net47),
    .D(_0081_),
    .Q_N(_0054_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _1911_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net46),
    .D(_0082_),
    .Q_N(_0053_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _1912_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net18),
    .D(_0083_),
    .Q_N(_0896_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _1913_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net74),
    .D(_0084_),
    .Q_N(_0051_),
    .Q(\bitmap_yofs[0] ));
 sg13g2_dfrbp_1 _1914_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net72),
    .D(net219),
    .Q_N(_0050_),
    .Q(\bitmap_yofs[1] ));
 sg13g2_dfrbp_1 _1915_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net69),
    .D(_0086_),
    .Q_N(_0033_),
    .Q(\bitmap_yofs[2] ));
 sg13g2_dfrbp_1 _1916_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net67),
    .D(_0087_),
    .Q_N(_0032_),
    .Q(\bitmap_yofs[3] ));
 sg13g2_dfrbp_1 _1917_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net48),
    .D(_0088_),
    .Q_N(_0049_),
    .Q(\bitmap_yofs[4] ));
 sg13g2_dfrbp_1 _1918_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net75),
    .D(_0089_),
    .Q_N(_0047_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _1919_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net19),
    .D(net85),
    .Q_N(_0895_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 _1920_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net73),
    .D(_0090_),
    .Q_N(_0894_),
    .Q(\bitsTemp[11] ));
 sg13g2_dfrbp_1 _1921_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net71),
    .D(_0091_),
    .Q_N(_0893_),
    .Q(\bitsTemp[21] ));
 sg13g2_dfrbp_1 _1922_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net68),
    .D(_0092_),
    .Q_N(_0892_),
    .Q(\bitsTemp[2] ));
 sg13g2_dfrbp_1 _1923_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net66),
    .D(_0093_),
    .Q_N(_0891_),
    .Q(\bitsTemp[1] ));
 sg13g2_dfrbp_1 _1924_ (.CLK(net262),
    .RESET_B(net289),
    .D(_0094_),
    .Q_N(_0890_),
    .Q(v_offset_rev_flag));
 sg13g2_tiehi _1919__19 (.L_HI(net19));
 sg13g2_tiehi _1856__20 (.L_HI(net20));
 sg13g2_tiehi _1857__21 (.L_HI(net21));
 sg13g2_tiehi _1858__22 (.L_HI(net22));
 sg13g2_tiehi _1859__23 (.L_HI(net23));
 sg13g2_tiehi _1860__24 (.L_HI(net24));
 sg13g2_tiehi _1861__25 (.L_HI(net25));
 sg13g2_tiehi _1862__26 (.L_HI(net26));
 sg13g2_tiehi _1863__27 (.L_HI(net27));
 sg13g2_tiehi _1864__28 (.L_HI(net28));
 sg13g2_tiehi _1865__29 (.L_HI(net29));
 sg13g2_tiehi _1866__30 (.L_HI(net30));
 sg13g2_tiehi _1867__31 (.L_HI(net31));
 sg13g2_tiehi _1868__32 (.L_HI(net32));
 sg13g2_tiehi _1869__33 (.L_HI(net33));
 sg13g2_tiehi _1870__34 (.L_HI(net34));
 sg13g2_tiehi _1871__35 (.L_HI(net35));
 sg13g2_tiehi _1872__36 (.L_HI(net36));
 sg13g2_tiehi _1873__37 (.L_HI(net37));
 sg13g2_tiehi _1874__38 (.L_HI(net38));
 sg13g2_tiehi _1875__39 (.L_HI(net39));
 sg13g2_tiehi _1876__40 (.L_HI(net40));
 sg13g2_tiehi _1877__41 (.L_HI(net41));
 sg13g2_tiehi _1878__42 (.L_HI(net42));
 sg13g2_tiehi _1879__43 (.L_HI(net43));
 sg13g2_tiehi _1880__44 (.L_HI(net44));
 sg13g2_tiehi _1881__45 (.L_HI(net45));
 sg13g2_tiehi _1911__46 (.L_HI(net46));
 sg13g2_tiehi _1910__47 (.L_HI(net47));
 sg13g2_tiehi _1917__48 (.L_HI(net48));
 sg13g2_tiehi _1909__49 (.L_HI(net49));
 sg13g2_tiehi _1908__50 (.L_HI(net50));
 sg13g2_tiehi _1900__51 (.L_HI(net51));
 sg13g2_tiehi _1899__52 (.L_HI(net52));
 sg13g2_tiehi _1898__53 (.L_HI(net53));
 sg13g2_tiehi _1897__54 (.L_HI(net54));
 sg13g2_tiehi _1901__55 (.L_HI(net55));
 sg13g2_tiehi _1902__56 (.L_HI(net56));
 sg13g2_tiehi _1903__57 (.L_HI(net57));
 sg13g2_tiehi _1904__58 (.L_HI(net58));
 sg13g2_tiehi _1905__59 (.L_HI(net59));
 sg13g2_tiehi _1906__60 (.L_HI(net60));
 sg13g2_tiehi _1896__61 (.L_HI(net61));
 sg13g2_tiehi _1895__62 (.L_HI(net62));
 sg13g2_tiehi _1894__63 (.L_HI(net63));
 sg13g2_tiehi _1893__64 (.L_HI(net64));
 sg13g2_tiehi _1892__65 (.L_HI(net65));
 sg13g2_tiehi _1923__66 (.L_HI(net66));
 sg13g2_tiehi _1916__67 (.L_HI(net67));
 sg13g2_tiehi _1922__68 (.L_HI(net68));
 sg13g2_tiehi _1915__69 (.L_HI(net69));
 sg13g2_tiehi _1907__70 (.L_HI(net70));
 sg13g2_tiehi _1921__71 (.L_HI(net71));
 sg13g2_tiehi _1914__72 (.L_HI(net72));
 sg13g2_tiehi _1920__73 (.L_HI(net73));
 sg13g2_tiehi _1913__74 (.L_HI(net74));
 sg13g2_tiehi _1918__75 (.L_HI(net75));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_quarren42_demoscene_top_3 (.L_LO(net3));
 sg13g2_tielo tt_um_quarren42_demoscene_top_4 (.L_LO(net4));
 sg13g2_tielo tt_um_quarren42_demoscene_top_5 (.L_LO(net5));
 sg13g2_tielo tt_um_quarren42_demoscene_top_6 (.L_LO(net6));
 sg13g2_tielo tt_um_quarren42_demoscene_top_7 (.L_LO(net7));
 sg13g2_tielo tt_um_quarren42_demoscene_top_8 (.L_LO(net8));
 sg13g2_tielo tt_um_quarren42_demoscene_top_9 (.L_LO(net9));
 sg13g2_tielo tt_um_quarren42_demoscene_top_10 (.L_LO(net10));
 sg13g2_tielo tt_um_quarren42_demoscene_top_11 (.L_LO(net11));
 sg13g2_tielo tt_um_quarren42_demoscene_top_12 (.L_LO(net12));
 sg13g2_tielo tt_um_quarren42_demoscene_top_13 (.L_LO(net13));
 sg13g2_tielo tt_um_quarren42_demoscene_top_14 (.L_LO(net14));
 sg13g2_tielo tt_um_quarren42_demoscene_top_15 (.L_LO(net15));
 sg13g2_tielo tt_um_quarren42_demoscene_top_16 (.L_LO(net16));
 sg13g2_tielo tt_um_quarren42_demoscene_top_17 (.L_LO(net17));
 sg13g2_tiehi _1912__18 (.L_HI(net18));
 sg13g2_buf_1 _1999_ (.A(b),
    .X(uo_out[0]));
 sg13g2_buf_1 _2000_ (.A(g),
    .X(uo_out[1]));
 sg13g2_buf_1 _2001_ (.A(r),
    .X(uo_out[2]));
 sg13g2_buf_1 _2002_ (.A(net261),
    .X(uo_out[3]));
 sg13g2_buf_1 _2003_ (.A(b),
    .X(uo_out[4]));
 sg13g2_buf_1 _2004_ (.A(g),
    .X(uo_out[5]));
 sg13g2_buf_1 _2005_ (.A(r),
    .X(uo_out[6]));
 sg13g2_buf_1 _2006_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout215 (.A(_0759_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(net217),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_0088_),
    .X(net217));
 sg13g2_buf_4 fanout218 (.X(net218),
    .A(net219));
 sg13g2_buf_2 fanout219 (.A(_0085_),
    .X(net219));
 sg13g2_buf_4 fanout220 (.X(net220),
    .A(_0086_));
 sg13g2_buf_4 fanout221 (.X(net221),
    .A(_0740_));
 sg13g2_buf_2 fanout222 (.A(net223),
    .X(net222));
 sg13g2_buf_1 fanout223 (.A(_0730_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(net225),
    .X(net224));
 sg13g2_buf_1 fanout225 (.A(_0723_),
    .X(net225));
 sg13g2_buf_4 fanout226 (.X(net226),
    .A(_0708_));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(_0187_));
 sg13g2_buf_2 fanout228 (.A(_0152_),
    .X(net228));
 sg13g2_buf_4 fanout229 (.X(net229),
    .A(net230));
 sg13g2_buf_4 fanout230 (.X(net230),
    .A(v_offset_rev_flag));
 sg13g2_buf_2 fanout231 (.A(net232),
    .X(net231));
 sg13g2_buf_1 fanout232 (.A(net233),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(\v_offset[8] ),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(net236),
    .X(net234));
 sg13g2_buf_1 fanout235 (.A(net236),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(net237),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(\v_offset[7] ),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(net240),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(net240),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(\v_offset[6] ),
    .X(net240));
 sg13g2_buf_4 fanout241 (.X(net241),
    .A(net244));
 sg13g2_buf_2 fanout242 (.A(net244),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(net244),
    .X(net243));
 sg13g2_buf_1 fanout244 (.A(\v_offset[5] ),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(net246),
    .X(net245));
 sg13g2_buf_4 fanout246 (.X(net246),
    .A(\v_offset[4] ));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(net249));
 sg13g2_buf_2 fanout248 (.A(net249),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(\v_offset[3] ),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(net252),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(net252),
    .X(net251));
 sg13g2_buf_4 fanout252 (.X(net252),
    .A(\v_offset[2] ));
 sg13g2_buf_2 fanout253 (.A(net254),
    .X(net253));
 sg13g2_buf_1 fanout254 (.A(net255),
    .X(net254));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(\v_offset[1] ));
 sg13g2_buf_2 fanout256 (.A(net257),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(\v_offset[0] ),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_0147_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_0144_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_0118_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(\hvsync_gen.vsync ),
    .X(net261));
 sg13g2_buf_1 fanout262 (.A(\hvsync_gen.vsync ),
    .X(net262));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(net264));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(\bitmap_yofs[3] ));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(\bitmap_yofs[2] ));
 sg13g2_buf_2 fanout266 (.A(\bitmap_yofs[2] ),
    .X(net266));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(net83));
 sg13g2_buf_2 fanout268 (.A(\bitmap_yofs[1] ),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(net270),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_0051_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(net101),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(net99),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(\hvsync_gen.vpos[0] ),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(net275),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(\hvsync_gen.hpos[9] ),
    .X(net275));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(net88));
 sg13g2_buf_1 fanout277 (.A(\bitmap_xofs[4] ),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(net280),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(\bitmap_xofs[3] ),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(net96),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(\bitmap_xofs[2] ),
    .X(net282));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(net102));
 sg13g2_buf_2 fanout284 (.A(\hvsync_gen.hpos[3] ),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(net89),
    .X(net285));
 sg13g2_buf_1 fanout286 (.A(\hvsync_gen.hpos[2] ),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(\hvsync_gen.hpos[1] ),
    .X(net287));
 sg13g2_buf_4 fanout288 (.X(net288),
    .A(net289));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(net1));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_tielo tt_um_quarren42_demoscene_top_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0066_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0065_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0101_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0044_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0884_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0034_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0030_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold8 (.A(\bitmap_yofs[1] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0140_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0031_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0037_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0047_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold13 (.A(\bitmap_xofs[4] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold14 (.A(\hvsync_gen.hpos[2] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0072_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0040_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold17 (.A(\bitmap_xofs[1] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0887_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0046_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0079_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold21 (.A(\bitmap_xofs[2] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0032_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold23 (.A(\hvsync_gen.hpos[0] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold24 (.A(\hvsync_gen.vpos[1] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold25 (.A(\bitmap_xofs[3] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold26 (.A(\hvsync_gen.vpos[3] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold27 (.A(\bitmap_xofs[0] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold28 (.A(\bitmap_yofs[4] ),
    .X(net103));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_4 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_86 ();
 sg13g2_decap_8 FILLER_9_93 ();
 sg13g2_decap_8 FILLER_9_100 ();
 sg13g2_fill_1 FILLER_9_107 ();
 sg13g2_fill_2 FILLER_9_134 ();
 sg13g2_decap_4 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_170 ();
 sg13g2_decap_8 FILLER_9_177 ();
 sg13g2_decap_8 FILLER_9_184 ();
 sg13g2_decap_8 FILLER_9_191 ();
 sg13g2_decap_8 FILLER_9_198 ();
 sg13g2_decap_8 FILLER_9_205 ();
 sg13g2_decap_8 FILLER_9_212 ();
 sg13g2_decap_8 FILLER_9_219 ();
 sg13g2_decap_8 FILLER_9_226 ();
 sg13g2_decap_8 FILLER_9_233 ();
 sg13g2_decap_8 FILLER_9_240 ();
 sg13g2_decap_8 FILLER_9_247 ();
 sg13g2_decap_8 FILLER_9_254 ();
 sg13g2_decap_8 FILLER_9_261 ();
 sg13g2_decap_8 FILLER_9_268 ();
 sg13g2_decap_8 FILLER_9_275 ();
 sg13g2_decap_8 FILLER_9_282 ();
 sg13g2_decap_8 FILLER_9_289 ();
 sg13g2_decap_8 FILLER_9_296 ();
 sg13g2_decap_8 FILLER_9_303 ();
 sg13g2_decap_8 FILLER_9_310 ();
 sg13g2_decap_8 FILLER_9_317 ();
 sg13g2_decap_8 FILLER_9_324 ();
 sg13g2_decap_8 FILLER_9_331 ();
 sg13g2_decap_8 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_345 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_decap_8 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_fill_2 FILLER_10_28 ();
 sg13g2_fill_1 FILLER_10_34 ();
 sg13g2_decap_8 FILLER_10_41 ();
 sg13g2_decap_8 FILLER_10_48 ();
 sg13g2_fill_2 FILLER_10_55 ();
 sg13g2_fill_1 FILLER_10_57 ();
 sg13g2_fill_2 FILLER_10_68 ();
 sg13g2_fill_1 FILLER_10_70 ();
 sg13g2_decap_4 FILLER_10_75 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_4 FILLER_10_98 ();
 sg13g2_fill_2 FILLER_10_115 ();
 sg13g2_fill_1 FILLER_10_117 ();
 sg13g2_fill_2 FILLER_10_152 ();
 sg13g2_fill_1 FILLER_10_154 ();
 sg13g2_fill_2 FILLER_10_159 ();
 sg13g2_fill_1 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_188 ();
 sg13g2_decap_8 FILLER_10_195 ();
 sg13g2_decap_8 FILLER_10_202 ();
 sg13g2_decap_8 FILLER_10_209 ();
 sg13g2_decap_8 FILLER_10_216 ();
 sg13g2_decap_8 FILLER_10_223 ();
 sg13g2_decap_8 FILLER_10_230 ();
 sg13g2_decap_8 FILLER_10_237 ();
 sg13g2_decap_8 FILLER_10_244 ();
 sg13g2_decap_8 FILLER_10_251 ();
 sg13g2_decap_8 FILLER_10_258 ();
 sg13g2_decap_8 FILLER_10_265 ();
 sg13g2_decap_8 FILLER_10_272 ();
 sg13g2_decap_8 FILLER_10_279 ();
 sg13g2_decap_8 FILLER_10_286 ();
 sg13g2_decap_8 FILLER_10_293 ();
 sg13g2_decap_8 FILLER_10_300 ();
 sg13g2_decap_8 FILLER_10_307 ();
 sg13g2_decap_8 FILLER_10_314 ();
 sg13g2_decap_8 FILLER_10_321 ();
 sg13g2_decap_8 FILLER_10_328 ();
 sg13g2_decap_8 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_38 ();
 sg13g2_fill_2 FILLER_11_69 ();
 sg13g2_fill_2 FILLER_11_94 ();
 sg13g2_decap_4 FILLER_11_115 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_fill_2 FILLER_11_149 ();
 sg13g2_decap_8 FILLER_11_164 ();
 sg13g2_fill_2 FILLER_11_171 ();
 sg13g2_decap_8 FILLER_11_177 ();
 sg13g2_decap_8 FILLER_11_184 ();
 sg13g2_decap_8 FILLER_11_191 ();
 sg13g2_decap_8 FILLER_11_198 ();
 sg13g2_decap_8 FILLER_11_205 ();
 sg13g2_decap_8 FILLER_11_212 ();
 sg13g2_decap_8 FILLER_11_219 ();
 sg13g2_decap_8 FILLER_11_226 ();
 sg13g2_decap_8 FILLER_11_233 ();
 sg13g2_decap_8 FILLER_11_240 ();
 sg13g2_decap_8 FILLER_11_247 ();
 sg13g2_decap_8 FILLER_11_254 ();
 sg13g2_decap_8 FILLER_11_261 ();
 sg13g2_decap_8 FILLER_11_268 ();
 sg13g2_decap_8 FILLER_11_275 ();
 sg13g2_decap_8 FILLER_11_282 ();
 sg13g2_decap_8 FILLER_11_289 ();
 sg13g2_decap_8 FILLER_11_296 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_decap_8 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_317 ();
 sg13g2_decap_8 FILLER_11_324 ();
 sg13g2_decap_8 FILLER_11_331 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_decap_8 FILLER_11_345 ();
 sg13g2_decap_8 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_23 ();
 sg13g2_fill_2 FILLER_12_33 ();
 sg13g2_fill_2 FILLER_12_45 ();
 sg13g2_fill_1 FILLER_12_47 ();
 sg13g2_fill_2 FILLER_12_56 ();
 sg13g2_decap_4 FILLER_12_67 ();
 sg13g2_fill_1 FILLER_12_71 ();
 sg13g2_fill_1 FILLER_12_77 ();
 sg13g2_fill_1 FILLER_12_87 ();
 sg13g2_fill_2 FILLER_12_92 ();
 sg13g2_fill_1 FILLER_12_102 ();
 sg13g2_fill_2 FILLER_12_112 ();
 sg13g2_fill_1 FILLER_12_114 ();
 sg13g2_fill_1 FILLER_12_165 ();
 sg13g2_decap_8 FILLER_12_192 ();
 sg13g2_decap_8 FILLER_12_199 ();
 sg13g2_decap_8 FILLER_12_206 ();
 sg13g2_decap_8 FILLER_12_213 ();
 sg13g2_decap_8 FILLER_12_220 ();
 sg13g2_decap_8 FILLER_12_227 ();
 sg13g2_decap_8 FILLER_12_234 ();
 sg13g2_decap_8 FILLER_12_241 ();
 sg13g2_fill_1 FILLER_12_248 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_282 ();
 sg13g2_decap_8 FILLER_12_289 ();
 sg13g2_decap_8 FILLER_12_296 ();
 sg13g2_decap_8 FILLER_12_303 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_decap_8 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_338 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_2 ();
 sg13g2_fill_2 FILLER_13_17 ();
 sg13g2_fill_2 FILLER_13_51 ();
 sg13g2_fill_1 FILLER_13_53 ();
 sg13g2_fill_1 FILLER_13_60 ();
 sg13g2_fill_1 FILLER_13_79 ();
 sg13g2_fill_2 FILLER_13_87 ();
 sg13g2_fill_1 FILLER_13_89 ();
 sg13g2_fill_1 FILLER_13_134 ();
 sg13g2_decap_8 FILLER_13_158 ();
 sg13g2_fill_1 FILLER_13_165 ();
 sg13g2_fill_1 FILLER_13_198 ();
 sg13g2_decap_4 FILLER_13_203 ();
 sg13g2_decap_4 FILLER_13_211 ();
 sg13g2_decap_8 FILLER_13_223 ();
 sg13g2_decap_8 FILLER_13_230 ();
 sg13g2_fill_1 FILLER_13_237 ();
 sg13g2_fill_2 FILLER_13_247 ();
 sg13g2_fill_2 FILLER_13_257 ();
 sg13g2_fill_1 FILLER_13_259 ();
 sg13g2_decap_4 FILLER_13_264 ();
 sg13g2_fill_2 FILLER_13_278 ();
 sg13g2_fill_1 FILLER_13_280 ();
 sg13g2_fill_2 FILLER_13_307 ();
 sg13g2_fill_1 FILLER_13_309 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_2 FILLER_14_11 ();
 sg13g2_fill_2 FILLER_14_44 ();
 sg13g2_fill_2 FILLER_14_55 ();
 sg13g2_decap_4 FILLER_14_69 ();
 sg13g2_decap_4 FILLER_14_86 ();
 sg13g2_fill_2 FILLER_14_90 ();
 sg13g2_decap_8 FILLER_14_109 ();
 sg13g2_decap_4 FILLER_14_116 ();
 sg13g2_fill_1 FILLER_14_120 ();
 sg13g2_decap_8 FILLER_14_129 ();
 sg13g2_decap_8 FILLER_14_136 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_fill_2 FILLER_14_158 ();
 sg13g2_decap_4 FILLER_14_186 ();
 sg13g2_fill_1 FILLER_14_190 ();
 sg13g2_decap_4 FILLER_14_202 ();
 sg13g2_fill_2 FILLER_14_206 ();
 sg13g2_fill_2 FILLER_14_262 ();
 sg13g2_fill_1 FILLER_14_264 ();
 sg13g2_fill_2 FILLER_14_286 ();
 sg13g2_fill_1 FILLER_14_288 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_2 FILLER_14_316 ();
 sg13g2_fill_1 FILLER_14_318 ();
 sg13g2_fill_2 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_352 ();
 sg13g2_decap_8 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_366 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_27 ();
 sg13g2_fill_1 FILLER_15_32 ();
 sg13g2_decap_8 FILLER_15_37 ();
 sg13g2_decap_8 FILLER_15_44 ();
 sg13g2_decap_4 FILLER_15_51 ();
 sg13g2_decap_4 FILLER_15_59 ();
 sg13g2_decap_8 FILLER_15_93 ();
 sg13g2_fill_2 FILLER_15_100 ();
 sg13g2_decap_4 FILLER_15_107 ();
 sg13g2_decap_8 FILLER_15_163 ();
 sg13g2_fill_1 FILLER_15_170 ();
 sg13g2_fill_2 FILLER_15_180 ();
 sg13g2_fill_1 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_216 ();
 sg13g2_decap_8 FILLER_15_223 ();
 sg13g2_decap_4 FILLER_15_230 ();
 sg13g2_fill_2 FILLER_15_234 ();
 sg13g2_fill_2 FILLER_15_281 ();
 sg13g2_fill_2 FILLER_15_322 ();
 sg13g2_decap_4 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_11 ();
 sg13g2_fill_2 FILLER_16_16 ();
 sg13g2_fill_2 FILLER_16_70 ();
 sg13g2_fill_2 FILLER_16_87 ();
 sg13g2_fill_1 FILLER_16_89 ();
 sg13g2_decap_8 FILLER_16_116 ();
 sg13g2_decap_4 FILLER_16_127 ();
 sg13g2_fill_2 FILLER_16_131 ();
 sg13g2_fill_2 FILLER_16_188 ();
 sg13g2_fill_1 FILLER_16_258 ();
 sg13g2_fill_1 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_270 ();
 sg13g2_decap_4 FILLER_16_277 ();
 sg13g2_fill_1 FILLER_16_281 ();
 sg13g2_fill_2 FILLER_16_305 ();
 sg13g2_decap_4 FILLER_16_317 ();
 sg13g2_fill_2 FILLER_16_321 ();
 sg13g2_fill_1 FILLER_16_331 ();
 sg13g2_fill_2 FILLER_16_341 ();
 sg13g2_fill_1 FILLER_16_369 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_30 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_46 ();
 sg13g2_decap_8 FILLER_17_53 ();
 sg13g2_fill_2 FILLER_17_60 ();
 sg13g2_decap_4 FILLER_17_66 ();
 sg13g2_fill_2 FILLER_17_70 ();
 sg13g2_fill_1 FILLER_17_86 ();
 sg13g2_fill_1 FILLER_17_92 ();
 sg13g2_decap_4 FILLER_17_107 ();
 sg13g2_fill_1 FILLER_17_111 ();
 sg13g2_decap_8 FILLER_17_155 ();
 sg13g2_decap_4 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_166 ();
 sg13g2_fill_2 FILLER_17_181 ();
 sg13g2_decap_8 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_216 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_fill_1 FILLER_17_230 ();
 sg13g2_decap_8 FILLER_17_235 ();
 sg13g2_fill_2 FILLER_17_254 ();
 sg13g2_decap_4 FILLER_17_285 ();
 sg13g2_fill_1 FILLER_17_289 ();
 sg13g2_fill_2 FILLER_17_296 ();
 sg13g2_fill_1 FILLER_17_312 ();
 sg13g2_decap_4 FILLER_17_325 ();
 sg13g2_fill_2 FILLER_17_329 ();
 sg13g2_fill_1 FILLER_17_348 ();
 sg13g2_fill_2 FILLER_17_353 ();
 sg13g2_fill_1 FILLER_17_355 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_23 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_4 FILLER_18_124 ();
 sg13g2_fill_2 FILLER_18_128 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_fill_1 FILLER_18_156 ();
 sg13g2_decap_8 FILLER_18_187 ();
 sg13g2_decap_8 FILLER_18_194 ();
 sg13g2_decap_8 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_240 ();
 sg13g2_fill_2 FILLER_18_247 ();
 sg13g2_fill_1 FILLER_18_249 ();
 sg13g2_decap_4 FILLER_18_258 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_fill_2 FILLER_18_287 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_fill_1 FILLER_18_305 ();
 sg13g2_fill_1 FILLER_18_317 ();
 sg13g2_fill_2 FILLER_18_376 ();
 sg13g2_decap_4 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_fill_2 FILLER_19_55 ();
 sg13g2_decap_8 FILLER_19_61 ();
 sg13g2_decap_8 FILLER_19_68 ();
 sg13g2_fill_1 FILLER_19_75 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_2 FILLER_19_96 ();
 sg13g2_fill_1 FILLER_19_98 ();
 sg13g2_fill_1 FILLER_19_108 ();
 sg13g2_decap_8 FILLER_19_113 ();
 sg13g2_fill_2 FILLER_19_120 ();
 sg13g2_fill_1 FILLER_19_122 ();
 sg13g2_decap_8 FILLER_19_157 ();
 sg13g2_decap_4 FILLER_19_164 ();
 sg13g2_decap_8 FILLER_19_172 ();
 sg13g2_decap_4 FILLER_19_179 ();
 sg13g2_decap_4 FILLER_19_188 ();
 sg13g2_fill_1 FILLER_19_192 ();
 sg13g2_decap_8 FILLER_19_197 ();
 sg13g2_decap_8 FILLER_19_204 ();
 sg13g2_fill_2 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_213 ();
 sg13g2_decap_4 FILLER_19_256 ();
 sg13g2_fill_1 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_291 ();
 sg13g2_fill_1 FILLER_19_318 ();
 sg13g2_decap_8 FILLER_19_340 ();
 sg13g2_decap_4 FILLER_19_347 ();
 sg13g2_fill_1 FILLER_19_351 ();
 sg13g2_decap_4 FILLER_19_356 ();
 sg13g2_fill_1 FILLER_19_360 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_decap_4 FILLER_20_29 ();
 sg13g2_fill_2 FILLER_20_38 ();
 sg13g2_fill_1 FILLER_20_40 ();
 sg13g2_fill_2 FILLER_20_72 ();
 sg13g2_fill_2 FILLER_20_82 ();
 sg13g2_fill_2 FILLER_20_96 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_fill_2 FILLER_20_129 ();
 sg13g2_fill_1 FILLER_20_131 ();
 sg13g2_fill_2 FILLER_20_145 ();
 sg13g2_decap_4 FILLER_20_199 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_fill_1 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_235 ();
 sg13g2_fill_1 FILLER_20_237 ();
 sg13g2_decap_4 FILLER_20_242 ();
 sg13g2_fill_1 FILLER_20_246 ();
 sg13g2_decap_4 FILLER_20_252 ();
 sg13g2_fill_1 FILLER_20_256 ();
 sg13g2_decap_8 FILLER_20_265 ();
 sg13g2_decap_4 FILLER_20_272 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_fill_2 FILLER_20_295 ();
 sg13g2_fill_2 FILLER_20_306 ();
 sg13g2_fill_2 FILLER_20_331 ();
 sg13g2_fill_2 FILLER_20_354 ();
 sg13g2_decap_4 FILLER_20_386 ();
 sg13g2_fill_1 FILLER_20_390 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_18 ();
 sg13g2_decap_8 FILLER_21_25 ();
 sg13g2_decap_8 FILLER_21_32 ();
 sg13g2_fill_1 FILLER_21_39 ();
 sg13g2_fill_2 FILLER_21_44 ();
 sg13g2_decap_4 FILLER_21_51 ();
 sg13g2_fill_2 FILLER_21_55 ();
 sg13g2_fill_1 FILLER_21_60 ();
 sg13g2_fill_1 FILLER_21_88 ();
 sg13g2_fill_2 FILLER_21_94 ();
 sg13g2_decap_8 FILLER_21_100 ();
 sg13g2_fill_2 FILLER_21_107 ();
 sg13g2_fill_2 FILLER_21_128 ();
 sg13g2_fill_1 FILLER_21_130 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_fill_2 FILLER_21_167 ();
 sg13g2_fill_1 FILLER_21_169 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_decap_4 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_206 ();
 sg13g2_fill_1 FILLER_21_213 ();
 sg13g2_fill_1 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_245 ();
 sg13g2_fill_2 FILLER_21_255 ();
 sg13g2_decap_8 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_318 ();
 sg13g2_fill_2 FILLER_21_325 ();
 sg13g2_fill_1 FILLER_21_327 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_decap_4 FILLER_21_352 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_fill_2 FILLER_21_383 ();
 sg13g2_fill_1 FILLER_21_385 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_decap_8 FILLER_22_59 ();
 sg13g2_fill_1 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_89 ();
 sg13g2_decap_8 FILLER_22_96 ();
 sg13g2_fill_1 FILLER_22_103 ();
 sg13g2_decap_4 FILLER_22_110 ();
 sg13g2_fill_1 FILLER_22_114 ();
 sg13g2_fill_1 FILLER_22_150 ();
 sg13g2_fill_2 FILLER_22_163 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_fill_1 FILLER_22_203 ();
 sg13g2_decap_4 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_216 ();
 sg13g2_decap_4 FILLER_22_234 ();
 sg13g2_fill_2 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_257 ();
 sg13g2_decap_4 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_268 ();
 sg13g2_decap_4 FILLER_22_278 ();
 sg13g2_fill_2 FILLER_22_282 ();
 sg13g2_fill_2 FILLER_22_314 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_fill_1 FILLER_22_356 ();
 sg13g2_fill_1 FILLER_22_361 ();
 sg13g2_decap_4 FILLER_22_379 ();
 sg13g2_fill_2 FILLER_22_383 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_19 ();
 sg13g2_decap_8 FILLER_23_26 ();
 sg13g2_decap_8 FILLER_23_33 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_1 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_170 ();
 sg13g2_decap_4 FILLER_23_176 ();
 sg13g2_fill_1 FILLER_23_180 ();
 sg13g2_fill_2 FILLER_23_184 ();
 sg13g2_fill_1 FILLER_23_191 ();
 sg13g2_decap_8 FILLER_23_206 ();
 sg13g2_fill_1 FILLER_23_222 ();
 sg13g2_fill_1 FILLER_23_240 ();
 sg13g2_fill_2 FILLER_23_249 ();
 sg13g2_fill_1 FILLER_23_251 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_decap_4 FILLER_23_294 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_fill_1 FILLER_23_335 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_fill_2 FILLER_23_358 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_fill_2 FILLER_23_366 ();
 sg13g2_decap_4 FILLER_23_380 ();
 sg13g2_fill_1 FILLER_23_396 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_35 ();
 sg13g2_fill_1 FILLER_24_37 ();
 sg13g2_fill_2 FILLER_24_71 ();
 sg13g2_fill_1 FILLER_24_73 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_fill_2 FILLER_24_87 ();
 sg13g2_fill_1 FILLER_24_98 ();
 sg13g2_fill_2 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_139 ();
 sg13g2_fill_1 FILLER_24_169 ();
 sg13g2_fill_1 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_decap_4 FILLER_24_233 ();
 sg13g2_fill_2 FILLER_24_237 ();
 sg13g2_fill_1 FILLER_24_265 ();
 sg13g2_decap_8 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_fill_1 FILLER_24_285 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_fill_1 FILLER_24_305 ();
 sg13g2_decap_8 FILLER_24_309 ();
 sg13g2_decap_8 FILLER_24_316 ();
 sg13g2_fill_2 FILLER_24_341 ();
 sg13g2_decap_4 FILLER_24_356 ();
 sg13g2_decap_8 FILLER_24_365 ();
 sg13g2_fill_2 FILLER_24_372 ();
 sg13g2_fill_1 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_58 ();
 sg13g2_fill_1 FILLER_25_60 ();
 sg13g2_fill_1 FILLER_25_103 ();
 sg13g2_fill_2 FILLER_25_123 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_fill_2 FILLER_25_143 ();
 sg13g2_decap_8 FILLER_25_157 ();
 sg13g2_decap_4 FILLER_25_164 ();
 sg13g2_fill_1 FILLER_25_168 ();
 sg13g2_decap_4 FILLER_25_181 ();
 sg13g2_fill_1 FILLER_25_185 ();
 sg13g2_fill_1 FILLER_25_195 ();
 sg13g2_fill_2 FILLER_25_201 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_209 ();
 sg13g2_decap_4 FILLER_25_216 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_decap_8 FILLER_25_227 ();
 sg13g2_fill_2 FILLER_25_234 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_271 ();
 sg13g2_fill_1 FILLER_25_281 ();
 sg13g2_fill_2 FILLER_25_286 ();
 sg13g2_decap_4 FILLER_25_294 ();
 sg13g2_decap_4 FILLER_25_324 ();
 sg13g2_fill_1 FILLER_25_328 ();
 sg13g2_fill_2 FILLER_25_356 ();
 sg13g2_decap_4 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_fill_2 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_394 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_fill_1 FILLER_26_68 ();
 sg13g2_fill_2 FILLER_26_91 ();
 sg13g2_fill_1 FILLER_26_93 ();
 sg13g2_fill_2 FILLER_26_107 ();
 sg13g2_decap_4 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_fill_1 FILLER_26_142 ();
 sg13g2_decap_4 FILLER_26_167 ();
 sg13g2_fill_1 FILLER_26_171 ();
 sg13g2_fill_1 FILLER_26_193 ();
 sg13g2_decap_8 FILLER_26_248 ();
 sg13g2_decap_4 FILLER_26_255 ();
 sg13g2_fill_2 FILLER_26_259 ();
 sg13g2_fill_2 FILLER_26_290 ();
 sg13g2_fill_1 FILLER_26_292 ();
 sg13g2_decap_4 FILLER_26_317 ();
 sg13g2_decap_4 FILLER_26_329 ();
 sg13g2_fill_1 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_fill_2 FILLER_26_349 ();
 sg13g2_fill_1 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_fill_2 FILLER_26_377 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_49 ();
 sg13g2_fill_2 FILLER_27_57 ();
 sg13g2_fill_2 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_65 ();
 sg13g2_fill_1 FILLER_27_75 ();
 sg13g2_fill_2 FILLER_27_92 ();
 sg13g2_fill_1 FILLER_27_122 ();
 sg13g2_fill_2 FILLER_27_131 ();
 sg13g2_decap_4 FILLER_27_142 ();
 sg13g2_fill_2 FILLER_27_146 ();
 sg13g2_fill_2 FILLER_27_153 ();
 sg13g2_decap_8 FILLER_27_160 ();
 sg13g2_fill_1 FILLER_27_177 ();
 sg13g2_decap_4 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_186 ();
 sg13g2_decap_8 FILLER_27_197 ();
 sg13g2_fill_2 FILLER_27_204 ();
 sg13g2_fill_1 FILLER_27_206 ();
 sg13g2_fill_1 FILLER_27_212 ();
 sg13g2_decap_4 FILLER_27_218 ();
 sg13g2_fill_2 FILLER_27_222 ();
 sg13g2_decap_8 FILLER_27_229 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_decap_8 FILLER_27_279 ();
 sg13g2_fill_2 FILLER_27_286 ();
 sg13g2_fill_2 FILLER_27_313 ();
 sg13g2_fill_1 FILLER_27_315 ();
 sg13g2_fill_2 FILLER_27_324 ();
 sg13g2_decap_4 FILLER_27_350 ();
 sg13g2_decap_4 FILLER_27_378 ();
 sg13g2_fill_2 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_4 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_46 ();
 sg13g2_decap_4 FILLER_28_51 ();
 sg13g2_fill_1 FILLER_28_85 ();
 sg13g2_decap_8 FILLER_28_93 ();
 sg13g2_decap_4 FILLER_28_166 ();
 sg13g2_fill_1 FILLER_28_219 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_fill_2 FILLER_28_238 ();
 sg13g2_fill_1 FILLER_28_240 ();
 sg13g2_fill_2 FILLER_28_249 ();
 sg13g2_decap_8 FILLER_28_257 ();
 sg13g2_decap_4 FILLER_28_264 ();
 sg13g2_fill_2 FILLER_28_277 ();
 sg13g2_decap_8 FILLER_28_302 ();
 sg13g2_fill_2 FILLER_28_309 ();
 sg13g2_fill_1 FILLER_28_311 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_fill_2 FILLER_28_335 ();
 sg13g2_fill_1 FILLER_28_337 ();
 sg13g2_fill_2 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_348 ();
 sg13g2_decap_4 FILLER_28_361 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_110 ();
 sg13g2_decap_8 FILLER_29_117 ();
 sg13g2_fill_1 FILLER_29_132 ();
 sg13g2_decap_4 FILLER_29_141 ();
 sg13g2_fill_1 FILLER_29_145 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_4 FILLER_29_161 ();
 sg13g2_fill_2 FILLER_29_182 ();
 sg13g2_fill_1 FILLER_29_184 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_fill_2 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_219 ();
 sg13g2_decap_4 FILLER_29_239 ();
 sg13g2_fill_1 FILLER_29_243 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_decap_8 FILLER_29_272 ();
 sg13g2_decap_4 FILLER_29_279 ();
 sg13g2_fill_2 FILLER_29_288 ();
 sg13g2_fill_2 FILLER_29_326 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_fill_1 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_354 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_fill_2 FILLER_29_387 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_4 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_46 ();
 sg13g2_fill_1 FILLER_30_71 ();
 sg13g2_fill_2 FILLER_30_77 ();
 sg13g2_fill_1 FILLER_30_79 ();
 sg13g2_decap_8 FILLER_30_113 ();
 sg13g2_fill_2 FILLER_30_120 ();
 sg13g2_fill_2 FILLER_30_127 ();
 sg13g2_fill_1 FILLER_30_129 ();
 sg13g2_decap_8 FILLER_30_139 ();
 sg13g2_fill_2 FILLER_30_146 ();
 sg13g2_fill_2 FILLER_30_159 ();
 sg13g2_decap_8 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_fill_2 FILLER_30_193 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_fill_2 FILLER_30_210 ();
 sg13g2_fill_2 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_fill_2 FILLER_30_270 ();
 sg13g2_decap_4 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_281 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_4 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_341 ();
 sg13g2_decap_4 FILLER_30_358 ();
 sg13g2_decap_8 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_51 ();
 sg13g2_decap_4 FILLER_31_110 ();
 sg13g2_fill_2 FILLER_31_114 ();
 sg13g2_decap_4 FILLER_31_136 ();
 sg13g2_fill_2 FILLER_31_160 ();
 sg13g2_decap_8 FILLER_31_166 ();
 sg13g2_fill_1 FILLER_31_189 ();
 sg13g2_decap_4 FILLER_31_195 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_fill_2 FILLER_31_226 ();
 sg13g2_decap_8 FILLER_31_236 ();
 sg13g2_decap_4 FILLER_31_265 ();
 sg13g2_fill_2 FILLER_31_269 ();
 sg13g2_decap_4 FILLER_31_281 ();
 sg13g2_decap_8 FILLER_31_318 ();
 sg13g2_decap_4 FILLER_31_325 ();
 sg13g2_fill_2 FILLER_31_329 ();
 sg13g2_fill_2 FILLER_31_339 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_fill_2 FILLER_31_357 ();
 sg13g2_decap_4 FILLER_31_363 ();
 sg13g2_fill_2 FILLER_31_382 ();
 sg13g2_fill_1 FILLER_31_384 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_56 ();
 sg13g2_fill_2 FILLER_32_75 ();
 sg13g2_decap_4 FILLER_32_114 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_135 ();
 sg13g2_decap_4 FILLER_32_140 ();
 sg13g2_fill_2 FILLER_32_144 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_fill_2 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_190 ();
 sg13g2_decap_8 FILLER_32_197 ();
 sg13g2_fill_2 FILLER_32_204 ();
 sg13g2_fill_1 FILLER_32_206 ();
 sg13g2_fill_2 FILLER_32_215 ();
 sg13g2_fill_1 FILLER_32_217 ();
 sg13g2_fill_1 FILLER_32_226 ();
 sg13g2_fill_2 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_265 ();
 sg13g2_decap_8 FILLER_32_272 ();
 sg13g2_decap_8 FILLER_32_279 ();
 sg13g2_fill_2 FILLER_32_286 ();
 sg13g2_fill_1 FILLER_32_288 ();
 sg13g2_decap_4 FILLER_32_303 ();
 sg13g2_fill_2 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_322 ();
 sg13g2_fill_2 FILLER_32_335 ();
 sg13g2_decap_4 FILLER_32_358 ();
 sg13g2_fill_2 FILLER_32_362 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_4 FILLER_33_35 ();
 sg13g2_fill_2 FILLER_33_39 ();
 sg13g2_fill_2 FILLER_33_84 ();
 sg13g2_decap_4 FILLER_33_118 ();
 sg13g2_fill_2 FILLER_33_127 ();
 sg13g2_fill_2 FILLER_33_140 ();
 sg13g2_fill_1 FILLER_33_142 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_fill_1 FILLER_33_150 ();
 sg13g2_fill_2 FILLER_33_156 ();
 sg13g2_decap_4 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_194 ();
 sg13g2_fill_1 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_202 ();
 sg13g2_fill_2 FILLER_33_209 ();
 sg13g2_fill_1 FILLER_33_211 ();
 sg13g2_fill_2 FILLER_33_256 ();
 sg13g2_fill_1 FILLER_33_258 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_4 FILLER_33_336 ();
 sg13g2_fill_2 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_351 ();
 sg13g2_fill_1 FILLER_33_358 ();
 sg13g2_decap_8 FILLER_33_376 ();
 sg13g2_fill_2 FILLER_33_383 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_fill_2 FILLER_34_91 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_fill_1 FILLER_34_106 ();
 sg13g2_fill_1 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_128 ();
 sg13g2_fill_1 FILLER_34_130 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_fill_2 FILLER_34_168 ();
 sg13g2_fill_1 FILLER_34_170 ();
 sg13g2_decap_4 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_194 ();
 sg13g2_decap_8 FILLER_34_212 ();
 sg13g2_fill_2 FILLER_34_219 ();
 sg13g2_decap_8 FILLER_34_226 ();
 sg13g2_decap_4 FILLER_34_233 ();
 sg13g2_fill_2 FILLER_34_237 ();
 sg13g2_fill_1 FILLER_34_248 ();
 sg13g2_decap_8 FILLER_34_256 ();
 sg13g2_decap_8 FILLER_34_263 ();
 sg13g2_decap_8 FILLER_34_270 ();
 sg13g2_decap_8 FILLER_34_277 ();
 sg13g2_decap_8 FILLER_34_284 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_293 ();
 sg13g2_decap_4 FILLER_34_310 ();
 sg13g2_fill_2 FILLER_34_340 ();
 sg13g2_fill_1 FILLER_34_342 ();
 sg13g2_fill_1 FILLER_34_358 ();
 sg13g2_fill_2 FILLER_34_378 ();
 sg13g2_decap_4 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_114 ();
 sg13g2_decap_4 FILLER_35_133 ();
 sg13g2_fill_2 FILLER_35_137 ();
 sg13g2_fill_2 FILLER_35_149 ();
 sg13g2_decap_8 FILLER_35_180 ();
 sg13g2_decap_4 FILLER_35_187 ();
 sg13g2_fill_2 FILLER_35_232 ();
 sg13g2_fill_2 FILLER_35_289 ();
 sg13g2_fill_2 FILLER_35_296 ();
 sg13g2_fill_1 FILLER_35_298 ();
 sg13g2_decap_8 FILLER_35_330 ();
 sg13g2_fill_1 FILLER_35_337 ();
 sg13g2_decap_8 FILLER_35_352 ();
 sg13g2_fill_1 FILLER_35_359 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_63 ();
 sg13g2_decap_4 FILLER_36_88 ();
 sg13g2_fill_1 FILLER_36_92 ();
 sg13g2_fill_1 FILLER_36_102 ();
 sg13g2_fill_1 FILLER_36_115 ();
 sg13g2_decap_4 FILLER_36_124 ();
 sg13g2_fill_2 FILLER_36_140 ();
 sg13g2_decap_4 FILLER_36_168 ();
 sg13g2_fill_2 FILLER_36_193 ();
 sg13g2_decap_8 FILLER_36_215 ();
 sg13g2_fill_2 FILLER_36_222 ();
 sg13g2_decap_4 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_232 ();
 sg13g2_decap_4 FILLER_36_237 ();
 sg13g2_fill_1 FILLER_36_241 ();
 sg13g2_fill_2 FILLER_36_255 ();
 sg13g2_decap_4 FILLER_36_283 ();
 sg13g2_fill_2 FILLER_36_291 ();
 sg13g2_fill_1 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_302 ();
 sg13g2_fill_2 FILLER_36_316 ();
 sg13g2_decap_8 FILLER_36_328 ();
 sg13g2_decap_4 FILLER_36_335 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_fill_2 FILLER_36_350 ();
 sg13g2_fill_1 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_fill_1 FILLER_37_103 ();
 sg13g2_decap_8 FILLER_37_116 ();
 sg13g2_decap_8 FILLER_37_123 ();
 sg13g2_decap_4 FILLER_37_130 ();
 sg13g2_fill_1 FILLER_37_134 ();
 sg13g2_fill_2 FILLER_37_148 ();
 sg13g2_fill_2 FILLER_37_158 ();
 sg13g2_fill_2 FILLER_37_172 ();
 sg13g2_fill_1 FILLER_37_174 ();
 sg13g2_decap_8 FILLER_37_184 ();
 sg13g2_fill_2 FILLER_37_191 ();
 sg13g2_fill_1 FILLER_37_247 ();
 sg13g2_decap_8 FILLER_37_268 ();
 sg13g2_decap_8 FILLER_37_275 ();
 sg13g2_decap_8 FILLER_37_282 ();
 sg13g2_decap_8 FILLER_37_289 ();
 sg13g2_decap_4 FILLER_37_296 ();
 sg13g2_fill_2 FILLER_37_300 ();
 sg13g2_decap_4 FILLER_37_306 ();
 sg13g2_fill_1 FILLER_37_310 ();
 sg13g2_fill_2 FILLER_37_315 ();
 sg13g2_fill_1 FILLER_37_317 ();
 sg13g2_decap_4 FILLER_37_323 ();
 sg13g2_fill_1 FILLER_37_327 ();
 sg13g2_decap_8 FILLER_37_354 ();
 sg13g2_fill_2 FILLER_37_361 ();
 sg13g2_fill_1 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_fill_2 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_fill_2 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_150 ();
 sg13g2_fill_1 FILLER_38_181 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_4 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_223 ();
 sg13g2_fill_2 FILLER_38_230 ();
 sg13g2_fill_1 FILLER_38_232 ();
 sg13g2_decap_8 FILLER_38_237 ();
 sg13g2_decap_4 FILLER_38_244 ();
 sg13g2_fill_2 FILLER_38_248 ();
 sg13g2_decap_8 FILLER_38_272 ();
 sg13g2_decap_8 FILLER_38_279 ();
 sg13g2_decap_8 FILLER_38_286 ();
 sg13g2_decap_8 FILLER_38_293 ();
 sg13g2_decap_8 FILLER_38_326 ();
 sg13g2_decap_8 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_347 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_fill_1 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
endmodule

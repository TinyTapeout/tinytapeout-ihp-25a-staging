module tt_um_arandomdev_fir_engine_top (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire dac;
 wire \firEngine.adcDataValid ;
 wire \firEngine.adcData[0] ;
 wire \firEngine.adcData[1] ;
 wire \firEngine.adcData[2] ;
 wire \firEngine.adcData[3] ;
 wire \firEngine.adcData[4] ;
 wire \firEngine.adcData[5] ;
 wire \firEngine.adcData[6] ;
 wire \firEngine.adcData[7] ;
 wire \firEngine.clockConfig[0] ;
 wire \firEngine.clockConfig[1] ;
 wire \firEngine.clockConfig[2] ;
 wire \firEngine.clockConfig[3] ;
 wire \firEngine.configStore.serialOut ;
 wire \firEngine.firDataValid ;
 wire \firEngine.firInst.accQ[0] ;
 wire \firEngine.firInst.accQ[10] ;
 wire \firEngine.firInst.accQ[11] ;
 wire \firEngine.firInst.accQ[12] ;
 wire \firEngine.firInst.accQ[13] ;
 wire \firEngine.firInst.accQ[14] ;
 wire \firEngine.firInst.accQ[15] ;
 wire \firEngine.firInst.accQ[16] ;
 wire \firEngine.firInst.accQ[1] ;
 wire \firEngine.firInst.accQ[2] ;
 wire \firEngine.firInst.accQ[3] ;
 wire \firEngine.firInst.accQ[4] ;
 wire \firEngine.firInst.accQ[5] ;
 wire \firEngine.firInst.accQ[6] ;
 wire \firEngine.firInst.accQ[7] ;
 wire \firEngine.firInst.accQ[8] ;
 wire \firEngine.firInst.accQ[9] ;
 wire \firEngine.firInst.bit_cnt[0] ;
 wire \firEngine.firInst.bit_cnt[1] ;
 wire \firEngine.firInst.bit_cnt[2] ;
 wire \firEngine.firInst.coeffs[0][0] ;
 wire \firEngine.firInst.coeffs[0][1] ;
 wire \firEngine.firInst.coeffs[0][2] ;
 wire \firEngine.firInst.coeffs[0][3] ;
 wire \firEngine.firInst.coeffs[0][4] ;
 wire \firEngine.firInst.coeffs[0][5] ;
 wire \firEngine.firInst.coeffs[0][6] ;
 wire \firEngine.firInst.coeffs[0][7] ;
 wire \firEngine.firInst.coeffs[1][0] ;
 wire \firEngine.firInst.coeffs[1][1] ;
 wire \firEngine.firInst.coeffs[1][2] ;
 wire \firEngine.firInst.coeffs[1][3] ;
 wire \firEngine.firInst.coeffs[1][4] ;
 wire \firEngine.firInst.coeffs[1][5] ;
 wire \firEngine.firInst.coeffs[1][6] ;
 wire \firEngine.firInst.coeffs[1][7] ;
 wire \firEngine.firInst.coeffs[2][0] ;
 wire \firEngine.firInst.coeffs[2][1] ;
 wire \firEngine.firInst.coeffs[2][2] ;
 wire \firEngine.firInst.coeffs[2][3] ;
 wire \firEngine.firInst.coeffs[2][4] ;
 wire \firEngine.firInst.coeffs[2][5] ;
 wire \firEngine.firInst.coeffs[2][6] ;
 wire \firEngine.firInst.coeffs[2][7] ;
 wire \firEngine.firInst.coeffs[3][0] ;
 wire \firEngine.firInst.coeffs[3][1] ;
 wire \firEngine.firInst.coeffs[3][2] ;
 wire \firEngine.firInst.coeffs[3][3] ;
 wire \firEngine.firInst.coeffs[3][4] ;
 wire \firEngine.firInst.coeffs[3][5] ;
 wire \firEngine.firInst.coeffs[3][6] ;
 wire \firEngine.firInst.coeffs[3][7] ;
 wire \firEngine.firInst.coeffs[4][0] ;
 wire \firEngine.firInst.coeffs[4][1] ;
 wire \firEngine.firInst.coeffs[4][2] ;
 wire \firEngine.firInst.coeffs[4][3] ;
 wire \firEngine.firInst.coeffs[4][4] ;
 wire \firEngine.firInst.coeffs[4][5] ;
 wire \firEngine.firInst.coeffs[4][6] ;
 wire \firEngine.firInst.coeffs[4][7] ;
 wire \firEngine.firInst.coeffs[5][0] ;
 wire \firEngine.firInst.coeffs[5][1] ;
 wire \firEngine.firInst.coeffs[5][2] ;
 wire \firEngine.firInst.coeffs[5][3] ;
 wire \firEngine.firInst.coeffs[5][4] ;
 wire \firEngine.firInst.coeffs[5][5] ;
 wire \firEngine.firInst.coeffs[5][6] ;
 wire \firEngine.firInst.coeffs[5][7] ;
 wire \firEngine.firInst.sample_cnt[0] ;
 wire \firEngine.firInst.sample_cnt[1] ;
 wire \firEngine.firInst.sample_cnt[2] ;
 wire \firEngine.firInst.sample_cnt_en ;
 wire \firEngine.firInst.samples[0][0] ;
 wire \firEngine.firInst.samples[0][1] ;
 wire \firEngine.firInst.samples[0][2] ;
 wire \firEngine.firInst.samples[0][3] ;
 wire \firEngine.firInst.samples[0][4] ;
 wire \firEngine.firInst.samples[0][5] ;
 wire \firEngine.firInst.samples[0][6] ;
 wire \firEngine.firInst.samples[0][7] ;
 wire \firEngine.firInst.samples[10][0] ;
 wire \firEngine.firInst.samples[10][1] ;
 wire \firEngine.firInst.samples[10][2] ;
 wire \firEngine.firInst.samples[10][3] ;
 wire \firEngine.firInst.samples[10][4] ;
 wire \firEngine.firInst.samples[10][5] ;
 wire \firEngine.firInst.samples[10][6] ;
 wire \firEngine.firInst.samples[10][7] ;
 wire \firEngine.firInst.samples[1][0] ;
 wire \firEngine.firInst.samples[1][1] ;
 wire \firEngine.firInst.samples[1][2] ;
 wire \firEngine.firInst.samples[1][3] ;
 wire \firEngine.firInst.samples[1][4] ;
 wire \firEngine.firInst.samples[1][5] ;
 wire \firEngine.firInst.samples[1][6] ;
 wire \firEngine.firInst.samples[1][7] ;
 wire \firEngine.firInst.samples[2][0] ;
 wire \firEngine.firInst.samples[2][1] ;
 wire \firEngine.firInst.samples[2][2] ;
 wire \firEngine.firInst.samples[2][3] ;
 wire \firEngine.firInst.samples[2][4] ;
 wire \firEngine.firInst.samples[2][5] ;
 wire \firEngine.firInst.samples[2][6] ;
 wire \firEngine.firInst.samples[2][7] ;
 wire \firEngine.firInst.samples[3][0] ;
 wire \firEngine.firInst.samples[3][1] ;
 wire \firEngine.firInst.samples[3][2] ;
 wire \firEngine.firInst.samples[3][3] ;
 wire \firEngine.firInst.samples[3][4] ;
 wire \firEngine.firInst.samples[3][5] ;
 wire \firEngine.firInst.samples[3][6] ;
 wire \firEngine.firInst.samples[3][7] ;
 wire \firEngine.firInst.samples[4][0] ;
 wire \firEngine.firInst.samples[4][1] ;
 wire \firEngine.firInst.samples[4][2] ;
 wire \firEngine.firInst.samples[4][3] ;
 wire \firEngine.firInst.samples[4][4] ;
 wire \firEngine.firInst.samples[4][5] ;
 wire \firEngine.firInst.samples[4][6] ;
 wire \firEngine.firInst.samples[4][7] ;
 wire \firEngine.firInst.samples[5][0] ;
 wire \firEngine.firInst.samples[5][1] ;
 wire \firEngine.firInst.samples[5][2] ;
 wire \firEngine.firInst.samples[5][3] ;
 wire \firEngine.firInst.samples[5][4] ;
 wire \firEngine.firInst.samples[5][5] ;
 wire \firEngine.firInst.samples[5][6] ;
 wire \firEngine.firInst.samples[5][7] ;
 wire \firEngine.firInst.samples[6][0] ;
 wire \firEngine.firInst.samples[6][1] ;
 wire \firEngine.firInst.samples[6][2] ;
 wire \firEngine.firInst.samples[6][3] ;
 wire \firEngine.firInst.samples[6][4] ;
 wire \firEngine.firInst.samples[6][5] ;
 wire \firEngine.firInst.samples[6][6] ;
 wire \firEngine.firInst.samples[6][7] ;
 wire \firEngine.firInst.samples[7][0] ;
 wire \firEngine.firInst.samples[7][1] ;
 wire \firEngine.firInst.samples[7][2] ;
 wire \firEngine.firInst.samples[7][3] ;
 wire \firEngine.firInst.samples[7][4] ;
 wire \firEngine.firInst.samples[7][5] ;
 wire \firEngine.firInst.samples[7][6] ;
 wire \firEngine.firInst.samples[7][7] ;
 wire \firEngine.firInst.samples[8][0] ;
 wire \firEngine.firInst.samples[8][1] ;
 wire \firEngine.firInst.samples[8][2] ;
 wire \firEngine.firInst.samples[8][3] ;
 wire \firEngine.firInst.samples[8][4] ;
 wire \firEngine.firInst.samples[8][5] ;
 wire \firEngine.firInst.samples[8][6] ;
 wire \firEngine.firInst.samples[8][7] ;
 wire \firEngine.firInst.samples[9][0] ;
 wire \firEngine.firInst.samples[9][1] ;
 wire \firEngine.firInst.samples[9][2] ;
 wire \firEngine.firInst.samples[9][3] ;
 wire \firEngine.firInst.samples[9][4] ;
 wire \firEngine.firInst.samples[9][5] ;
 wire \firEngine.firInst.samples[9][6] ;
 wire \firEngine.firInst.samples[9][7] ;
 wire \firEngine.firInst.state[0] ;
 wire \firEngine.firInst.state[1] ;
 wire \firEngine.firInst.state[2] ;
 wire \firEngine.i2sController.adcQ ;
 wire \firEngine.i2sController.adcSynchronizer[0] ;
 wire \firEngine.i2sController.currentState[0] ;
 wire \firEngine.i2sController.currentState[1] ;
 wire \firEngine.i2sController.currentState[2] ;
 wire \firEngine.i2sController.dacDataQ[0] ;
 wire \firEngine.i2sController.dacDataQ[1] ;
 wire \firEngine.i2sController.dacDataQ[2] ;
 wire \firEngine.i2sController.dacDataQ[3] ;
 wire \firEngine.i2sController.dacDataQ[4] ;
 wire \firEngine.i2sController.dacDataQ[5] ;
 wire \firEngine.i2sController.dacDataQ[6] ;
 wire \firEngine.i2sController.dacDataQ[7] ;
 wire \firEngine.i2sController.lrck ;
 wire \firEngine.i2sController.lrckCounter[0] ;
 wire \firEngine.i2sController.lrckCounter[1] ;
 wire \firEngine.i2sController.lrckCounter[2] ;
 wire \firEngine.i2sController.lrckCounter[3] ;
 wire \firEngine.i2sController.lrckCounter[4] ;
 wire \firEngine.i2sController.mclk ;
 wire \firEngine.i2sController.mclkCounter[0] ;
 wire \firEngine.i2sController.mclkCounter[1] ;
 wire \firEngine.i2sController.mclkCounter[2] ;
 wire \firEngine.i2sController.mclkCounter[3] ;
 wire \firEngine.i2sController.nextState[0] ;
 wire \firEngine.i2sController.nextState[1] ;
 wire \firEngine.i2sController.sclk ;
 wire \firEngine.i2sController.sclkCounter ;
 wire \firEngine.spiSlave.cs ;
 wire \firEngine.spiSlave.csSynchronizer[0] ;
 wire \firEngine.spiSlave.mosi ;
 wire \firEngine.spiSlave.mosiSynchronizer[0] ;
 wire \firEngine.spiSlave.sclkSynchronizer[0] ;
 wire \firEngine.spiSlave.sclkSynchronizer[1] ;
 wire \firEngine.spiSlave.sclkSynchronizer[2] ;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire clknet_leaf_0_clk;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;

 sg13g2_inv_1 _1455_ (.Y(_0582_),
    .A(net239));
 sg13g2_inv_1 _1456_ (.Y(_0583_),
    .A(\firEngine.i2sController.mclk ));
 sg13g2_inv_1 _1457_ (.Y(_0584_),
    .A(net345));
 sg13g2_inv_1 _1458_ (.Y(_0585_),
    .A(net708));
 sg13g2_inv_1 _1459_ (.Y(_0586_),
    .A(\firEngine.i2sController.lrckCounter[0] ));
 sg13g2_inv_1 _1460_ (.Y(_0587_),
    .A(net297));
 sg13g2_inv_1 _1461_ (.Y(_0588_),
    .A(net256));
 sg13g2_inv_1 _1462_ (.Y(_0589_),
    .A(net279));
 sg13g2_inv_1 _1463_ (.Y(_0590_),
    .A(net247));
 sg13g2_inv_1 _1464_ (.Y(_0591_),
    .A(net263));
 sg13g2_inv_1 _1465_ (.Y(_0592_),
    .A(net277));
 sg13g2_inv_1 _1466_ (.Y(_0593_),
    .A(net258));
 sg13g2_inv_1 _1467_ (.Y(_0594_),
    .A(net267));
 sg13g2_inv_1 _1468_ (.Y(_0595_),
    .A(net254));
 sg13g2_inv_1 _1469_ (.Y(_0596_),
    .A(net291));
 sg13g2_inv_1 _1470_ (.Y(_0597_),
    .A(net293));
 sg13g2_inv_1 _1471_ (.Y(_0598_),
    .A(net251));
 sg13g2_inv_1 _1472_ (.Y(_0599_),
    .A(net249));
 sg13g2_inv_1 _1473_ (.Y(_0600_),
    .A(net269));
 sg13g2_inv_1 _1474_ (.Y(_0601_),
    .A(net282));
 sg13g2_inv_1 _1475_ (.Y(_0602_),
    .A(net261));
 sg13g2_inv_1 _1476_ (.Y(_0603_),
    .A(net374));
 sg13g2_inv_1 _1477_ (.Y(_0604_),
    .A(net550));
 sg13g2_inv_1 _1478_ (.Y(_0605_),
    .A(net314));
 sg13g2_inv_1 _1479_ (.Y(_0606_),
    .A(net298));
 sg13g2_inv_1 _1480_ (.Y(_0607_),
    .A(net364));
 sg13g2_inv_1 _1481_ (.Y(_0608_),
    .A(net405));
 sg13g2_inv_1 _1482_ (.Y(_0609_),
    .A(net610));
 sg13g2_inv_1 _1483_ (.Y(_0610_),
    .A(net670));
 sg13g2_inv_1 _1484_ (.Y(_0611_),
    .A(\firEngine.firInst.samples[4][0] ));
 sg13g2_inv_1 _1485_ (.Y(_0612_),
    .A(\firEngine.firInst.coeffs[0][7] ));
 sg13g2_inv_1 _1486_ (.Y(_0613_),
    .A(\firEngine.firInst.accQ[15] ));
 sg13g2_inv_1 _1487_ (.Y(_0614_),
    .A(\firEngine.firInst.accQ[14] ));
 sg13g2_inv_1 _1488_ (.Y(_0615_),
    .A(\firEngine.firInst.accQ[3] ));
 sg13g2_inv_1 _1489_ (.Y(_0616_),
    .A(net328));
 sg13g2_inv_1 _1490_ (.Y(_0617_),
    .A(net304));
 sg13g2_inv_1 _1491_ (.Y(_0618_),
    .A(net245));
 sg13g2_inv_1 _1492_ (.Y(_0619_),
    .A(net309));
 sg13g2_inv_1 _1493_ (.Y(_0620_),
    .A(net265));
 sg13g2_inv_1 _1494_ (.Y(_0621_),
    .A(net284));
 sg13g2_inv_1 _1495_ (.Y(_0622_),
    .A(net253));
 sg13g2_inv_1 _1496_ (.Y(_0623_),
    .A(net273));
 sg13g2_inv_1 _1497_ (.Y(_0624_),
    .A(net624));
 sg13g2_inv_1 _1498_ (.Y(_0625_),
    .A(net370));
 sg13g2_inv_1 _1499_ (.Y(_0626_),
    .A(\firEngine.clockConfig[0] ));
 sg13g2_inv_2 _1500_ (.Y(_0627_),
    .A(\firEngine.firInst.bit_cnt[2] ));
 sg13g2_inv_2 _1501_ (.Y(_0628_),
    .A(net557));
 sg13g2_inv_1 _1502_ (.Y(_0629_),
    .A(_0013_));
 sg13g2_inv_1 _1503_ (.Y(_0630_),
    .A(net275));
 sg13g2_inv_1 _1504_ (.Y(_0631_),
    .A(_0009_));
 sg13g2_inv_1 _1505_ (.Y(_0632_),
    .A(net283));
 sg13g2_inv_2 _1506_ (.Y(_0633_),
    .A(net590));
 sg13g2_inv_1 _1507_ (.Y(_0634_),
    .A(net678));
 sg13g2_inv_2 _1508_ (.Y(_0635_),
    .A(net307));
 sg13g2_inv_1 _1509_ (.Y(_0636_),
    .A(\firEngine.firInst.state[2] ));
 sg13g2_xnor2_1 _1510_ (.Y(_0637_),
    .A(\firEngine.clockConfig[1] ),
    .B(\firEngine.i2sController.mclkCounter[1] ));
 sg13g2_xnor2_1 _1511_ (.Y(_0638_),
    .A(\firEngine.clockConfig[0] ),
    .B(\firEngine.i2sController.mclkCounter[0] ));
 sg13g2_xnor2_1 _1512_ (.Y(_0639_),
    .A(\firEngine.clockConfig[3] ),
    .B(\firEngine.i2sController.mclkCounter[3] ));
 sg13g2_xnor2_1 _1513_ (.Y(_0640_),
    .A(\firEngine.clockConfig[2] ),
    .B(\firEngine.i2sController.mclkCounter[2] ));
 sg13g2_nand4_1 _1514_ (.B(_0638_),
    .C(_0639_),
    .A(_0637_),
    .Y(_0641_),
    .D(_0640_));
 sg13g2_nor2_1 _1515_ (.A(_0583_),
    .B(_0641_),
    .Y(_0642_));
 sg13g2_nand3_1 _1516_ (.B(\firEngine.i2sController.sclk ),
    .C(_0642_),
    .A(\firEngine.i2sController.sclkCounter ),
    .Y(_0643_));
 sg13g2_nor3_1 _1517_ (.A(_0585_),
    .B(_0586_),
    .C(_0643_),
    .Y(_0644_));
 sg13g2_and2_1 _1518_ (.A(net715),
    .B(_0644_),
    .X(_0645_));
 sg13g2_nand2_1 _1519_ (.Y(_0646_),
    .A(net705),
    .B(_0645_));
 sg13g2_nand4_1 _1520_ (.B(\firEngine.i2sController.lrckCounter[4] ),
    .C(\firEngine.i2sController.lrckCounter[3] ),
    .A(net294),
    .Y(_0647_),
    .D(_0645_));
 sg13g2_inv_1 _1521_ (.Y(_0648_),
    .A(net295));
 sg13g2_nor3_1 _1522_ (.A(\firEngine.i2sController.lrckCounter[2] ),
    .B(\firEngine.i2sController.lrckCounter[1] ),
    .C(_0586_),
    .Y(_0649_));
 sg13g2_nand3_1 _1523_ (.B(\firEngine.i2sController.lrckCounter[3] ),
    .C(_0649_),
    .A(net345),
    .Y(_0650_));
 sg13g2_a21oi_1 _1524_ (.A1(\firEngine.i2sController.currentState[0] ),
    .A2(net295),
    .Y(_0651_),
    .B1(net564));
 sg13g2_o21ai_1 _1525_ (.B1(_0651_),
    .Y(_0004_),
    .A1(_0634_),
    .A2(net346));
 sg13g2_nor2b_1 _1526_ (.A(_0011_),
    .B_N(\firEngine.firInst.sample_cnt[0] ),
    .Y(_0652_));
 sg13g2_nand2b_2 _1527_ (.Y(_0653_),
    .B(_0652_),
    .A_N(\firEngine.firInst.sample_cnt[1] ));
 sg13g2_inv_1 _1528_ (.Y(_0654_),
    .A(_0653_));
 sg13g2_a21oi_1 _1529_ (.A1(net280),
    .A2(\firEngine.firInst.sample_cnt[1] ),
    .Y(_0655_),
    .B1(_0654_));
 sg13g2_a21oi_1 _1530_ (.A1(\firEngine.firInst.bit_cnt[2] ),
    .A2(net556),
    .Y(_0656_),
    .B1(_0635_));
 sg13g2_a221oi_1 _1531_ (.B2(_0655_),
    .C1(_0656_),
    .B1(net683),
    .A1(net554),
    .Y(_0657_),
    .A2(net700));
 sg13g2_nor2_1 _1532_ (.A(net563),
    .B(net701),
    .Y(_0002_));
 sg13g2_a21oi_1 _1533_ (.A1(_0604_),
    .A2(\firEngine.firInst.state[0] ),
    .Y(_0658_),
    .B1(net421));
 sg13g2_nor3_2 _1534_ (.A(\firEngine.spiSlave.sclkSynchronizer[2] ),
    .B(_0632_),
    .C(net660),
    .Y(_0659_));
 sg13g2_or3_1 _1535_ (.A(\firEngine.spiSlave.sclkSynchronizer[2] ),
    .B(_0632_),
    .C(net720),
    .X(_0660_));
 sg13g2_nor3_1 _1536_ (.A(net563),
    .B(net422),
    .C(net511),
    .Y(_0003_));
 sg13g2_nand3_1 _1537_ (.B(net239),
    .C(_0642_),
    .A(\firEngine.i2sController.sclkCounter ),
    .Y(_0661_));
 sg13g2_inv_1 _1538_ (.Y(_0662_),
    .A(_0661_));
 sg13g2_a22oi_1 _1539_ (.Y(_0663_),
    .B1(_0661_),
    .B2(net664),
    .A2(_0648_),
    .A1(\firEngine.i2sController.currentState[0] ));
 sg13g2_nor2_1 _1540_ (.A(net564),
    .B(net665),
    .Y(\firEngine.i2sController.nextState[0] ));
 sg13g2_a22oi_1 _1541_ (.Y(_0664_),
    .B1(_0662_),
    .B2(net664),
    .A2(_0650_),
    .A1(net678));
 sg13g2_nor2_1 _1542_ (.A(net564),
    .B(net679),
    .Y(\firEngine.i2sController.nextState[1] ));
 sg13g2_nand2b_1 _1543_ (.Y(_0665_),
    .B(net683),
    .A_N(_0655_));
 sg13g2_o21ai_1 _1544_ (.B1(net593),
    .Y(_0666_),
    .A1(net422),
    .A2(_0659_));
 sg13g2_nand2b_1 _1545_ (.Y(_0001_),
    .B(net684),
    .A_N(_0666_));
 sg13g2_nor4_1 _1546_ (.A(_0627_),
    .B(_0628_),
    .C(net563),
    .D(_0635_),
    .Y(_0000_));
 sg13g2_and2_1 _1547_ (.A(net591),
    .B(net1),
    .X(_0032_));
 sg13g2_and2_1 _1548_ (.A(net592),
    .B(net235),
    .X(_0033_));
 sg13g2_a21oi_1 _1549_ (.A1(net324),
    .A2(_0659_),
    .Y(_0667_),
    .B1(net565));
 sg13g2_o21ai_1 _1550_ (.B1(net325),
    .Y(_0034_),
    .A1(_0626_),
    .A2(_0659_));
 sg13g2_a21oi_1 _1551_ (.A1(\firEngine.clockConfig[0] ),
    .A2(_0659_),
    .Y(_0668_),
    .B1(net565));
 sg13g2_o21ai_1 _1552_ (.B1(_0668_),
    .Y(_0035_),
    .A1(_0625_),
    .A2(_0659_));
 sg13g2_a21oi_1 _1553_ (.A1(net404),
    .A2(net511),
    .Y(_0669_),
    .B1(net565));
 sg13g2_o21ai_1 _1554_ (.B1(_0669_),
    .Y(_0036_),
    .A1(_0625_),
    .A2(net511));
 sg13g2_a21oi_1 _1555_ (.A1(net404),
    .A2(net661),
    .Y(_0670_),
    .B1(net565));
 sg13g2_o21ai_1 _1556_ (.B1(_0670_),
    .Y(_0037_),
    .A1(_0624_),
    .A2(net661));
 sg13g2_a21oi_1 _1557_ (.A1(\firEngine.configStore.serialOut ),
    .A2(net511),
    .Y(_0671_),
    .B1(net565));
 sg13g2_o21ai_1 _1558_ (.B1(_0671_),
    .Y(_0038_),
    .A1(_0624_),
    .A2(net511));
 sg13g2_nand2_1 _1559_ (.Y(_0672_),
    .A(net589),
    .B(_0641_));
 sg13g2_and3_1 _1560_ (.X(_0039_),
    .A(net589),
    .B(net234),
    .C(_0641_));
 sg13g2_and2_1 _1561_ (.A(\firEngine.i2sController.mclkCounter[0] ),
    .B(net318),
    .X(_0673_));
 sg13g2_nor2_1 _1562_ (.A(\firEngine.i2sController.mclkCounter[0] ),
    .B(net318),
    .Y(_0674_));
 sg13g2_nor3_1 _1563_ (.A(_0672_),
    .B(_0673_),
    .C(net319),
    .Y(_0040_));
 sg13g2_nand2_1 _1564_ (.Y(_0675_),
    .A(\firEngine.i2sController.mclkCounter[2] ),
    .B(_0673_));
 sg13g2_xnor2_1 _1565_ (.Y(_0676_),
    .A(net419),
    .B(_0673_));
 sg13g2_nor2_1 _1566_ (.A(_0672_),
    .B(net420),
    .Y(_0041_));
 sg13g2_xor2_1 _1567_ (.B(_0675_),
    .A(net380),
    .X(_0677_));
 sg13g2_nor2_1 _1568_ (.A(_0672_),
    .B(net381),
    .Y(_0042_));
 sg13g2_and2_1 _1569_ (.A(net592),
    .B(net3),
    .X(_0043_));
 sg13g2_and2_1 _1570_ (.A(net592),
    .B(net237),
    .X(_0044_));
 sg13g2_nor2_1 _1571_ (.A(_0632_),
    .B(net565),
    .Y(_0045_));
 sg13g2_and2_1 _1572_ (.A(net592),
    .B(net2),
    .X(_0046_));
 sg13g2_and2_1 _1573_ (.A(net592),
    .B(net236),
    .X(_0047_));
 sg13g2_a21oi_1 _1574_ (.A1(net560),
    .A2(_0653_),
    .Y(_0678_),
    .B1(net547));
 sg13g2_a21o_1 _1575_ (.A2(_0653_),
    .A1(net560),
    .B1(net547),
    .X(_0679_));
 sg13g2_o21ai_1 _1576_ (.B1(net571),
    .Y(_0680_),
    .A1(\firEngine.firInst.samples[10][0] ),
    .A2(net463));
 sg13g2_a21oi_1 _1577_ (.A1(_0623_),
    .A2(net463),
    .Y(_0048_),
    .B1(_0680_));
 sg13g2_o21ai_1 _1578_ (.B1(net572),
    .Y(_0681_),
    .A1(net260),
    .A2(net461));
 sg13g2_a21oi_1 _1579_ (.A1(_0622_),
    .A2(net461),
    .Y(_0049_),
    .B1(_0681_));
 sg13g2_o21ai_1 _1580_ (.B1(net566),
    .Y(_0682_),
    .A1(net286),
    .A2(net461));
 sg13g2_a21oi_1 _1581_ (.A1(_0621_),
    .A2(net461),
    .Y(_0050_),
    .B1(_0682_));
 sg13g2_o21ai_1 _1582_ (.B1(net566),
    .Y(_0683_),
    .A1(\firEngine.firInst.samples[10][3] ),
    .A2(net462));
 sg13g2_a21oi_1 _1583_ (.A1(_0620_),
    .A2(net462),
    .Y(_0051_),
    .B1(_0683_));
 sg13g2_o21ai_1 _1584_ (.B1(net574),
    .Y(_0684_),
    .A1(\firEngine.firInst.samples[10][4] ),
    .A2(net467));
 sg13g2_a21oi_1 _1585_ (.A1(_0619_),
    .A2(net467),
    .Y(_0052_),
    .B1(_0684_));
 sg13g2_o21ai_1 _1586_ (.B1(net569),
    .Y(_0685_),
    .A1(\firEngine.firInst.samples[10][5] ),
    .A2(net466));
 sg13g2_a21oi_1 _1587_ (.A1(_0618_),
    .A2(net466),
    .Y(_0053_),
    .B1(_0685_));
 sg13g2_o21ai_1 _1588_ (.B1(net574),
    .Y(_0686_),
    .A1(net311),
    .A2(net478));
 sg13g2_a21oi_1 _1589_ (.A1(_0617_),
    .A2(net466),
    .Y(_0054_),
    .B1(_0686_));
 sg13g2_o21ai_1 _1590_ (.B1(net568),
    .Y(_0687_),
    .A1(\firEngine.firInst.samples[10][7] ),
    .A2(net466));
 sg13g2_a21oi_1 _1591_ (.A1(_0616_),
    .A2(net466),
    .Y(_0055_),
    .B1(_0687_));
 sg13g2_o21ai_1 _1592_ (.B1(net571),
    .Y(_0688_),
    .A1(net282),
    .A2(net482));
 sg13g2_a21oi_1 _1593_ (.A1(_0623_),
    .A2(net481),
    .Y(_0056_),
    .B1(_0688_));
 sg13g2_o21ai_1 _1594_ (.B1(net566),
    .Y(_0689_),
    .A1(net249),
    .A2(net481));
 sg13g2_a21oi_1 _1595_ (.A1(_0622_),
    .A2(net481),
    .Y(_0057_),
    .B1(_0689_));
 sg13g2_o21ai_1 _1596_ (.B1(net566),
    .Y(_0690_),
    .A1(\firEngine.firInst.samples[8][2] ),
    .A2(net479));
 sg13g2_a21oi_1 _1597_ (.A1(_0621_),
    .A2(net479),
    .Y(_0058_),
    .B1(_0690_));
 sg13g2_o21ai_1 _1598_ (.B1(net567),
    .Y(_0691_),
    .A1(net254),
    .A2(net480));
 sg13g2_a21oi_1 _1599_ (.A1(_0620_),
    .A2(net480),
    .Y(_0059_),
    .B1(_0691_));
 sg13g2_o21ai_1 _1600_ (.B1(net568),
    .Y(_0692_),
    .A1(net258),
    .A2(net483));
 sg13g2_a21oi_1 _1601_ (.A1(_0619_),
    .A2(net483),
    .Y(_0060_),
    .B1(_0692_));
 sg13g2_o21ai_1 _1602_ (.B1(net569),
    .Y(_0693_),
    .A1(net263),
    .A2(net484));
 sg13g2_a21oi_1 _1603_ (.A1(_0618_),
    .A2(net485),
    .Y(_0061_),
    .B1(_0693_));
 sg13g2_o21ai_1 _1604_ (.B1(net578),
    .Y(_0694_),
    .A1(net279),
    .A2(net485));
 sg13g2_a21oi_1 _1605_ (.A1(_0617_),
    .A2(net485),
    .Y(_0062_),
    .B1(_0694_));
 sg13g2_o21ai_1 _1606_ (.B1(net570),
    .Y(_0695_),
    .A1(net297),
    .A2(net484));
 sg13g2_a21oi_1 _1607_ (.A1(_0616_),
    .A2(net484),
    .Y(_0063_),
    .B1(_0695_));
 sg13g2_a21oi_1 _1608_ (.A1(net558),
    .A2(_0629_),
    .Y(_0696_),
    .B1(net556));
 sg13g2_o21ai_1 _1609_ (.B1(_0696_),
    .Y(_0697_),
    .A1(net558),
    .A2(_0012_));
 sg13g2_mux2_1 _1610_ (.A0(_0014_),
    .A1(_0015_),
    .S(net558),
    .X(_0698_));
 sg13g2_a21oi_1 _1611_ (.A1(net556),
    .A2(_0698_),
    .Y(_0699_),
    .B1(\firEngine.firInst.bit_cnt[2] ));
 sg13g2_nor2b_1 _1612_ (.A(_0017_),
    .B_N(net559),
    .Y(_0700_));
 sg13g2_o21ai_1 _1613_ (.B1(_0628_),
    .Y(_0701_),
    .A1(net559),
    .A2(_0016_));
 sg13g2_mux2_1 _1614_ (.A0(_0018_),
    .A1(_0019_),
    .S(net559),
    .X(_0702_));
 sg13g2_a21oi_1 _1615_ (.A1(net557),
    .A2(_0702_),
    .Y(_0703_),
    .B1(_0627_));
 sg13g2_o21ai_1 _1616_ (.B1(_0703_),
    .Y(_0704_),
    .A1(_0700_),
    .A2(_0701_));
 sg13g2_a21oi_1 _1617_ (.A1(_0697_),
    .A2(_0699_),
    .Y(_0705_),
    .B1(_0653_));
 sg13g2_mux2_1 _1618_ (.A0(\firEngine.firInst.samples[0][4] ),
    .A1(\firEngine.firInst.samples[0][5] ),
    .S(net558),
    .X(_0706_));
 sg13g2_nand2_1 _1619_ (.Y(_0707_),
    .A(_0628_),
    .B(_0706_));
 sg13g2_mux2_1 _1620_ (.A0(\firEngine.firInst.samples[0][6] ),
    .A1(\firEngine.firInst.samples[0][7] ),
    .S(net558),
    .X(_0708_));
 sg13g2_a21oi_1 _1621_ (.A1(net556),
    .A2(_0708_),
    .Y(_0709_),
    .B1(_0627_));
 sg13g2_mux4_1 _1622_ (.S0(net558),
    .A0(\firEngine.firInst.samples[0][0] ),
    .A1(\firEngine.firInst.samples[0][1] ),
    .A2(\firEngine.firInst.samples[0][2] ),
    .A3(\firEngine.firInst.samples[0][3] ),
    .S1(net556),
    .X(_0710_));
 sg13g2_nor2_1 _1623_ (.A(\firEngine.firInst.bit_cnt[2] ),
    .B(_0710_),
    .Y(_0711_));
 sg13g2_a21oi_2 _1624_ (.B1(_0711_),
    .Y(_0712_),
    .A2(_0709_),
    .A1(_0707_));
 sg13g2_mux2_1 _1625_ (.A0(\firEngine.firInst.samples[10][4] ),
    .A1(\firEngine.firInst.samples[10][5] ),
    .S(net558),
    .X(_0713_));
 sg13g2_nand2_1 _1626_ (.Y(_0714_),
    .A(_0628_),
    .B(_0713_));
 sg13g2_mux2_1 _1627_ (.A0(\firEngine.firInst.samples[10][6] ),
    .A1(\firEngine.firInst.samples[10][7] ),
    .S(net559),
    .X(_0715_));
 sg13g2_a21oi_1 _1628_ (.A1(net556),
    .A2(_0715_),
    .Y(_0716_),
    .B1(_0627_));
 sg13g2_mux4_1 _1629_ (.S0(net558),
    .A0(\firEngine.firInst.samples[10][0] ),
    .A1(\firEngine.firInst.samples[10][1] ),
    .A2(\firEngine.firInst.samples[10][2] ),
    .A3(\firEngine.firInst.samples[10][3] ),
    .S1(net556),
    .X(_0717_));
 sg13g2_nor2_1 _1630_ (.A(\firEngine.firInst.bit_cnt[2] ),
    .B(_0717_),
    .Y(_0718_));
 sg13g2_a21oi_2 _1631_ (.B1(_0718_),
    .Y(_0719_),
    .A2(_0716_),
    .A1(_0714_));
 sg13g2_xnor2_1 _1632_ (.Y(_0720_),
    .A(_0712_),
    .B(_0719_));
 sg13g2_a22oi_1 _1633_ (.Y(_0721_),
    .B1(_0720_),
    .B2(_0653_),
    .A2(_0705_),
    .A1(_0704_));
 sg13g2_xnor2_1 _1634_ (.Y(_0722_),
    .A(\firEngine.configStore.serialOut ),
    .B(_0712_));
 sg13g2_and3_1 _1635_ (.X(_0723_),
    .A(_0653_),
    .B(_0719_),
    .C(_0722_));
 sg13g2_nor2_2 _1636_ (.A(_0721_),
    .B(_0723_),
    .Y(_0724_));
 sg13g2_or2_2 _1637_ (.X(_0725_),
    .B(_0723_),
    .A(_0721_));
 sg13g2_nand4_1 _1638_ (.B(_0719_),
    .C(_0720_),
    .A(_0653_),
    .Y(_0726_),
    .D(_0722_));
 sg13g2_nand2_2 _1639_ (.Y(_0727_),
    .A(net559),
    .B(net557));
 sg13g2_nor2_1 _1640_ (.A(net717),
    .B(_0727_),
    .Y(_0728_));
 sg13g2_or2_2 _1641_ (.X(_0729_),
    .B(_0727_),
    .A(_0010_));
 sg13g2_nor2_1 _1642_ (.A(_0726_),
    .B(_0729_),
    .Y(_0730_));
 sg13g2_nand2b_1 _1643_ (.Y(_0731_),
    .B(net492),
    .A_N(net460));
 sg13g2_xnor2_1 _1644_ (.Y(_0732_),
    .A(_0630_),
    .B(net460));
 sg13g2_xnor2_1 _1645_ (.Y(_0733_),
    .A(_0029_),
    .B(net460));
 sg13g2_nand2_1 _1646_ (.Y(_0734_),
    .A(_0631_),
    .B(_0733_));
 sg13g2_xnor2_1 _1647_ (.Y(_0735_),
    .A(net559),
    .B(net557));
 sg13g2_inv_1 _1648_ (.Y(_0736_),
    .A(_0735_));
 sg13g2_mux2_2 _1649_ (.A0(_0736_),
    .A1(net556),
    .S(net460),
    .X(_0737_));
 sg13g2_mux2_1 _1650_ (.A0(_0735_),
    .A1(_0628_),
    .S(net460),
    .X(_0738_));
 sg13g2_nand3_1 _1651_ (.B(_0733_),
    .C(net453),
    .A(_0631_),
    .Y(_0739_));
 sg13g2_xnor2_1 _1652_ (.Y(_0740_),
    .A(_0627_),
    .B(_0727_));
 sg13g2_inv_1 _1653_ (.Y(_0741_),
    .A(_0740_));
 sg13g2_nand2b_1 _1654_ (.Y(_0742_),
    .B(_0740_),
    .A_N(net460));
 sg13g2_nand2_1 _1655_ (.Y(_0743_),
    .A(_0627_),
    .B(net460));
 sg13g2_mux2_1 _1656_ (.A0(_0741_),
    .A1(\firEngine.firInst.bit_cnt[2] ),
    .S(net460),
    .X(_0744_));
 sg13g2_nand2_1 _1657_ (.Y(_0745_),
    .A(_0742_),
    .B(_0743_));
 sg13g2_nor4_2 _1658_ (.A(_0009_),
    .B(_0732_),
    .C(_0737_),
    .Y(_0746_),
    .D(net452));
 sg13g2_and2_1 _1659_ (.A(net454),
    .B(_0746_),
    .X(_0747_));
 sg13g2_nand2_1 _1660_ (.Y(_0748_),
    .A(net454),
    .B(_0746_));
 sg13g2_nor2_2 _1661_ (.A(net458),
    .B(_0748_),
    .Y(_0749_));
 sg13g2_nand2_1 _1662_ (.Y(_0750_),
    .A(_0008_),
    .B(_0749_));
 sg13g2_nor2_1 _1663_ (.A(net560),
    .B(net307),
    .Y(_0751_));
 sg13g2_or2_1 _1664_ (.X(_0752_),
    .B(\firEngine.firInst.state[1] ),
    .A(net560));
 sg13g2_xor2_1 _1665_ (.B(_0749_),
    .A(_0008_),
    .X(_0753_));
 sg13g2_nor2_1 _1666_ (.A(net554),
    .B(net563),
    .Y(_0754_));
 sg13g2_nand2_1 _1667_ (.Y(_0755_),
    .A(net537),
    .B(net593));
 sg13g2_o21ai_1 _1668_ (.B1(net530),
    .Y(_0756_),
    .A1(net366),
    .A2(net531));
 sg13g2_a21oi_1 _1669_ (.A1(net531),
    .A2(_0753_),
    .Y(_0064_),
    .B1(_0756_));
 sg13g2_xor2_1 _1670_ (.B(_0726_),
    .A(net559),
    .X(_0757_));
 sg13g2_mux2_1 _1671_ (.A0(_0009_),
    .A1(_0022_),
    .S(_0757_),
    .X(_0758_));
 sg13g2_nor3_1 _1672_ (.A(_0737_),
    .B(net452),
    .C(_0758_),
    .Y(_0759_));
 sg13g2_nor4_2 _1673_ (.A(net457),
    .B(_0737_),
    .C(net452),
    .Y(_0760_),
    .D(_0758_));
 sg13g2_or4_1 _1674_ (.A(net456),
    .B(_0737_),
    .C(net452),
    .D(_0758_),
    .X(_0761_));
 sg13g2_nor2_1 _1675_ (.A(_0739_),
    .B(_0761_),
    .Y(_0762_));
 sg13g2_nand2b_1 _1676_ (.Y(_0763_),
    .B(_0760_),
    .A_N(_0739_));
 sg13g2_nand2_1 _1677_ (.Y(_0764_),
    .A(_0721_),
    .B(_0723_));
 sg13g2_inv_1 _1678_ (.Y(_0765_),
    .A(net450));
 sg13g2_a21oi_1 _1679_ (.A1(_0748_),
    .A2(_0761_),
    .Y(_0766_),
    .B1(net451));
 sg13g2_o21ai_1 _1680_ (.B1(net448),
    .Y(_0767_),
    .A1(_0747_),
    .A2(_0760_));
 sg13g2_nor2_1 _1681_ (.A(net458),
    .B(_0761_),
    .Y(_0768_));
 sg13g2_nand3_1 _1682_ (.B(_0760_),
    .C(net451),
    .A(_0725_),
    .Y(_0769_));
 sg13g2_o21ai_1 _1683_ (.B1(_0769_),
    .Y(_0770_),
    .A1(_0762_),
    .A2(_0767_));
 sg13g2_a221oi_1 _1684_ (.B2(net451),
    .C1(_0749_),
    .B1(_0768_),
    .A1(_0763_),
    .Y(_0771_),
    .A2(_0766_));
 sg13g2_xnor2_1 _1685_ (.Y(_0772_),
    .A(_0749_),
    .B(_0770_));
 sg13g2_and2_1 _1686_ (.A(\firEngine.firInst.accQ[1] ),
    .B(_0772_),
    .X(_0773_));
 sg13g2_xor2_1 _1687_ (.B(_0772_),
    .A(\firEngine.firInst.accQ[1] ),
    .X(_0774_));
 sg13g2_xnor2_1 _1688_ (.Y(_0775_),
    .A(_0750_),
    .B(_0774_));
 sg13g2_o21ai_1 _1689_ (.B1(net530),
    .Y(_0776_),
    .A1(net658),
    .A2(net531));
 sg13g2_a21oi_1 _1690_ (.A1(net531),
    .A2(_0775_),
    .Y(_0065_),
    .B1(_0776_));
 sg13g2_a21oi_2 _1691_ (.B1(_0773_),
    .Y(_0777_),
    .A2(_0774_),
    .A1(_0750_));
 sg13g2_mux2_1 _1692_ (.A0(_0022_),
    .A1(_0023_),
    .S(_0757_),
    .X(_0778_));
 sg13g2_a21oi_1 _1693_ (.A1(_0631_),
    .A2(_0733_),
    .Y(_0779_),
    .B1(net453));
 sg13g2_a221oi_1 _1694_ (.B2(net453),
    .C1(_0779_),
    .B1(_0778_),
    .A1(_0742_),
    .Y(_0780_),
    .A2(_0743_));
 sg13g2_and2_1 _1695_ (.A(net454),
    .B(_0780_),
    .X(_0781_));
 sg13g2_nand2_1 _1696_ (.Y(_0782_),
    .A(net455),
    .B(_0780_));
 sg13g2_nand3_1 _1697_ (.B(net454),
    .C(_0780_),
    .A(_0725_),
    .Y(_0783_));
 sg13g2_mux2_1 _1698_ (.A0(_0781_),
    .A1(_0783_),
    .S(_0767_),
    .X(_0784_));
 sg13g2_nand2_1 _1699_ (.Y(_0785_),
    .A(_0771_),
    .B(_0784_));
 sg13g2_xnor2_1 _1700_ (.Y(_0786_),
    .A(_0771_),
    .B(_0784_));
 sg13g2_nand2_1 _1701_ (.Y(_0787_),
    .A(\firEngine.firInst.accQ[2] ),
    .B(_0786_));
 sg13g2_nor2_1 _1702_ (.A(\firEngine.firInst.accQ[2] ),
    .B(_0786_),
    .Y(_0788_));
 sg13g2_xor2_1 _1703_ (.B(_0786_),
    .A(net671),
    .X(_0789_));
 sg13g2_xor2_1 _1704_ (.B(_0789_),
    .A(_0777_),
    .X(_0790_));
 sg13g2_o21ai_1 _1705_ (.B1(net530),
    .Y(_0791_),
    .A1(net671),
    .A2(net531));
 sg13g2_a21oi_1 _1706_ (.A1(net531),
    .A2(_0790_),
    .Y(_0066_),
    .B1(_0791_));
 sg13g2_o21ai_1 _1707_ (.B1(_0787_),
    .Y(_0792_),
    .A1(_0777_),
    .A2(_0788_));
 sg13g2_mux4_1 _1708_ (.S0(_0757_),
    .A0(_0009_),
    .A1(_0022_),
    .A2(_0023_),
    .A3(_0024_),
    .S1(net453),
    .X(_0793_));
 sg13g2_nor2_1 _1709_ (.A(net452),
    .B(_0793_),
    .Y(_0794_));
 sg13g2_nor3_2 _1710_ (.A(net456),
    .B(net452),
    .C(_0793_),
    .Y(_0795_));
 sg13g2_a21oi_1 _1711_ (.A1(_0771_),
    .A2(_0784_),
    .Y(_0796_),
    .B1(net451));
 sg13g2_or2_1 _1712_ (.X(_0797_),
    .B(_0796_),
    .A(_0795_));
 sg13g2_a21oi_1 _1713_ (.A1(_0795_),
    .A2(_0796_),
    .Y(_0798_),
    .B1(net458));
 sg13g2_a21oi_1 _1714_ (.A1(_0771_),
    .A2(_0784_),
    .Y(_0799_),
    .B1(net492));
 sg13g2_nand3_1 _1715_ (.B(_0798_),
    .C(_0799_),
    .A(_0797_),
    .Y(_0800_));
 sg13g2_a21o_1 _1716_ (.A2(_0798_),
    .A1(_0797_),
    .B1(_0799_),
    .X(_0801_));
 sg13g2_a21oi_1 _1717_ (.A1(_0800_),
    .A2(_0801_),
    .Y(_0802_),
    .B1(_0615_));
 sg13g2_nand3_1 _1718_ (.B(_0800_),
    .C(_0801_),
    .A(_0615_),
    .Y(_0803_));
 sg13g2_nor2b_1 _1719_ (.A(_0802_),
    .B_N(_0803_),
    .Y(_0804_));
 sg13g2_xnor2_1 _1720_ (.Y(_0805_),
    .A(_0792_),
    .B(_0804_));
 sg13g2_o21ai_1 _1721_ (.B1(net530),
    .Y(_0806_),
    .A1(net338),
    .A2(net532));
 sg13g2_a21oi_1 _1722_ (.A1(net532),
    .A2(_0805_),
    .Y(_0067_),
    .B1(_0806_));
 sg13g2_a21oi_2 _1723_ (.B1(_0802_),
    .Y(_0807_),
    .A2(_0803_),
    .A1(_0792_));
 sg13g2_mux2_1 _1724_ (.A0(_0024_),
    .A1(_0025_),
    .S(_0757_),
    .X(_0808_));
 sg13g2_mux4_1 _1725_ (.S0(_0757_),
    .A0(_0022_),
    .A1(_0023_),
    .A2(_0024_),
    .A3(_0025_),
    .S1(net453),
    .X(_0809_));
 sg13g2_mux2_1 _1726_ (.A0(_0739_),
    .A1(_0809_),
    .S(_0745_),
    .X(_0810_));
 sg13g2_nor2_1 _1727_ (.A(net457),
    .B(_0810_),
    .Y(_0811_));
 sg13g2_nand2b_1 _1728_ (.Y(_0812_),
    .B(net455),
    .A_N(_0810_));
 sg13g2_nor3_2 _1729_ (.A(_0747_),
    .B(_0760_),
    .C(_0795_),
    .Y(_0813_));
 sg13g2_a21oi_1 _1730_ (.A1(_0782_),
    .A2(_0813_),
    .Y(_0814_),
    .B1(net451));
 sg13g2_or2_1 _1731_ (.X(_0815_),
    .B(_0814_),
    .A(_0811_));
 sg13g2_a21oi_1 _1732_ (.A1(_0811_),
    .A2(_0814_),
    .Y(_0816_),
    .B1(_0724_));
 sg13g2_nand2_1 _1733_ (.Y(_0817_),
    .A(_0815_),
    .B(_0816_));
 sg13g2_a21oi_1 _1734_ (.A1(_0725_),
    .A2(_0795_),
    .Y(_0818_),
    .B1(_0785_));
 sg13g2_nor2_1 _1735_ (.A(net493),
    .B(_0818_),
    .Y(_0819_));
 sg13g2_xor2_1 _1736_ (.B(_0819_),
    .A(_0817_),
    .X(_0820_));
 sg13g2_nand2_1 _1737_ (.Y(_0821_),
    .A(\firEngine.firInst.accQ[4] ),
    .B(_0820_));
 sg13g2_xnor2_1 _1738_ (.Y(_0822_),
    .A(net646),
    .B(_0820_));
 sg13g2_xnor2_1 _1739_ (.Y(_0823_),
    .A(_0807_),
    .B(_0822_));
 sg13g2_o21ai_1 _1740_ (.B1(net530),
    .Y(_0824_),
    .A1(net646),
    .A2(net531));
 sg13g2_a21oi_1 _1741_ (.A1(net531),
    .A2(_0823_),
    .Y(_0068_),
    .B1(_0824_));
 sg13g2_o21ai_1 _1742_ (.B1(_0821_),
    .Y(_0825_),
    .A1(_0807_),
    .A2(_0822_));
 sg13g2_mux2_1 _1743_ (.A0(_0025_),
    .A1(_0026_),
    .S(_0757_),
    .X(_0826_));
 sg13g2_mux4_1 _1744_ (.S0(_0757_),
    .A0(_0023_),
    .A1(_0024_),
    .A2(_0025_),
    .A3(_0026_),
    .S1(net453),
    .X(_0827_));
 sg13g2_nor2_1 _1745_ (.A(net452),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_nor3_1 _1746_ (.A(_0737_),
    .B(net449),
    .C(_0758_),
    .Y(_0829_));
 sg13g2_o21ai_1 _1747_ (.B1(net454),
    .Y(_0830_),
    .A1(_0828_),
    .A2(_0829_));
 sg13g2_inv_1 _1748_ (.Y(_0831_),
    .A(_0830_));
 sg13g2_nand3_1 _1749_ (.B(_0812_),
    .C(_0813_),
    .A(_0782_),
    .Y(_0832_));
 sg13g2_nand3_1 _1750_ (.B(_0831_),
    .C(_0832_),
    .A(_0765_),
    .Y(_0833_));
 sg13g2_a21o_1 _1751_ (.A2(_0832_),
    .A1(net448),
    .B1(_0831_),
    .X(_0834_));
 sg13g2_nand3_1 _1752_ (.B(_0833_),
    .C(_0834_),
    .A(_0725_),
    .Y(_0835_));
 sg13g2_a221oi_1 _1753_ (.B2(_0816_),
    .C1(_0785_),
    .B1(_0815_),
    .A1(_0725_),
    .Y(_0836_),
    .A2(_0795_));
 sg13g2_nor2_1 _1754_ (.A(net493),
    .B(_0836_),
    .Y(_0837_));
 sg13g2_xor2_1 _1755_ (.B(_0837_),
    .A(_0835_),
    .X(_0838_));
 sg13g2_and2_1 _1756_ (.A(\firEngine.firInst.accQ[5] ),
    .B(_0838_),
    .X(_0839_));
 sg13g2_or2_1 _1757_ (.X(_0840_),
    .B(_0838_),
    .A(\firEngine.firInst.accQ[5] ));
 sg13g2_nand2b_1 _1758_ (.Y(_0841_),
    .B(_0840_),
    .A_N(_0839_));
 sg13g2_xor2_1 _1759_ (.B(_0841_),
    .A(_0825_),
    .X(_0842_));
 sg13g2_o21ai_1 _1760_ (.B1(_0754_),
    .Y(_0843_),
    .A1(net655),
    .A2(_0752_));
 sg13g2_a21oi_1 _1761_ (.A1(net536),
    .A2(_0842_),
    .Y(_0069_),
    .B1(net656));
 sg13g2_a21oi_2 _1762_ (.B1(_0839_),
    .Y(_0844_),
    .A2(_0840_),
    .A1(_0825_));
 sg13g2_mux2_1 _1763_ (.A0(_0026_),
    .A1(_0027_),
    .S(_0757_),
    .X(_0845_));
 sg13g2_mux2_1 _1764_ (.A0(_0808_),
    .A1(_0845_),
    .S(net453),
    .X(_0846_));
 sg13g2_mux4_1 _1765_ (.S0(net453),
    .A0(_0734_),
    .A1(_0778_),
    .A2(_0808_),
    .A3(_0845_),
    .S1(net449),
    .X(_0847_));
 sg13g2_nand2b_2 _1766_ (.Y(_0848_),
    .B(net455),
    .A_N(_0847_));
 sg13g2_inv_1 _1767_ (.Y(_0849_),
    .A(_0848_));
 sg13g2_and4_1 _1768_ (.A(_0782_),
    .B(_0812_),
    .C(_0813_),
    .D(_0830_),
    .X(_0850_));
 sg13g2_nand4_1 _1769_ (.B(_0812_),
    .C(_0813_),
    .A(_0782_),
    .Y(_0851_),
    .D(_0830_));
 sg13g2_nor3_1 _1770_ (.A(net450),
    .B(_0848_),
    .C(_0850_),
    .Y(_0852_));
 sg13g2_a21oi_1 _1771_ (.A1(net448),
    .A2(_0851_),
    .Y(_0853_),
    .B1(_0849_));
 sg13g2_nor3_2 _1772_ (.A(net458),
    .B(_0852_),
    .C(_0853_),
    .Y(_0854_));
 sg13g2_a21oi_2 _1773_ (.B1(net493),
    .Y(_0855_),
    .A2(_0836_),
    .A1(_0835_));
 sg13g2_xor2_1 _1774_ (.B(_0855_),
    .A(_0854_),
    .X(_0856_));
 sg13g2_nand2b_1 _1775_ (.Y(_0857_),
    .B(\firEngine.firInst.accQ[6] ),
    .A_N(_0856_));
 sg13g2_xor2_1 _1776_ (.B(_0856_),
    .A(net626),
    .X(_0858_));
 sg13g2_xnor2_1 _1777_ (.Y(_0859_),
    .A(_0844_),
    .B(_0858_));
 sg13g2_o21ai_1 _1778_ (.B1(net529),
    .Y(_0860_),
    .A1(net626),
    .A2(net536));
 sg13g2_a21oi_1 _1779_ (.A1(net536),
    .A2(_0859_),
    .Y(_0070_),
    .B1(_0860_));
 sg13g2_o21ai_1 _1780_ (.B1(_0857_),
    .Y(_0861_),
    .A1(_0844_),
    .A2(_0858_));
 sg13g2_mux2_1 _1781_ (.A0(_0027_),
    .A1(_0028_),
    .S(_0733_),
    .X(_0862_));
 sg13g2_mux2_1 _1782_ (.A0(_0826_),
    .A1(_0862_),
    .S(_0738_),
    .X(_0863_));
 sg13g2_mux2_2 _1783_ (.A0(_0793_),
    .A1(_0863_),
    .S(net449),
    .X(_0864_));
 sg13g2_inv_1 _1784_ (.Y(_0865_),
    .A(_0864_));
 sg13g2_nor2_1 _1785_ (.A(net457),
    .B(_0864_),
    .Y(_0866_));
 sg13g2_nor2_1 _1786_ (.A(net450),
    .B(_0848_),
    .Y(_0867_));
 sg13g2_a21oi_2 _1787_ (.B1(net451),
    .Y(_0868_),
    .A2(_0850_),
    .A1(_0848_));
 sg13g2_a221oi_1 _1788_ (.B2(_0731_),
    .C1(_0867_),
    .B1(_0865_),
    .A1(net448),
    .Y(_0869_),
    .A2(_0851_));
 sg13g2_a21o_1 _1789_ (.A2(_0868_),
    .A1(_0866_),
    .B1(_0724_),
    .X(_0870_));
 sg13g2_nor2_1 _1790_ (.A(_0869_),
    .B(_0870_),
    .Y(_0871_));
 sg13g2_and2_1 _1791_ (.A(_0729_),
    .B(_0854_),
    .X(_0872_));
 sg13g2_nor2_1 _1792_ (.A(_0855_),
    .B(_0872_),
    .Y(_0873_));
 sg13g2_xor2_1 _1793_ (.B(_0873_),
    .A(_0871_),
    .X(_0874_));
 sg13g2_and2_1 _1794_ (.A(\firEngine.firInst.accQ[7] ),
    .B(_0874_),
    .X(_0875_));
 sg13g2_or2_1 _1795_ (.X(_0876_),
    .B(_0874_),
    .A(\firEngine.firInst.accQ[7] ));
 sg13g2_nor2b_1 _1796_ (.A(_0875_),
    .B_N(_0876_),
    .Y(_0877_));
 sg13g2_xnor2_1 _1797_ (.Y(_0878_),
    .A(_0861_),
    .B(_0877_));
 sg13g2_o21ai_1 _1798_ (.B1(net530),
    .Y(_0879_),
    .A1(net704),
    .A2(net536));
 sg13g2_a21oi_1 _1799_ (.A1(net536),
    .A2(_0878_),
    .Y(_0071_),
    .B1(_0879_));
 sg13g2_a21oi_1 _1800_ (.A1(_0861_),
    .A2(_0876_),
    .Y(_0880_),
    .B1(_0875_));
 sg13g2_a21o_1 _1801_ (.A2(_0876_),
    .A1(_0861_),
    .B1(_0875_),
    .X(_0881_));
 sg13g2_nor3_1 _1802_ (.A(net493),
    .B(_0869_),
    .C(_0870_),
    .Y(_0882_));
 sg13g2_nor3_1 _1803_ (.A(_0855_),
    .B(_0872_),
    .C(_0882_),
    .Y(_0883_));
 sg13g2_nor3_1 _1804_ (.A(net457),
    .B(net450),
    .C(_0864_),
    .Y(_0884_));
 sg13g2_mux2_1 _1805_ (.A0(_0612_),
    .A1(_0845_),
    .S(_0737_),
    .X(_0885_));
 sg13g2_mux2_1 _1806_ (.A0(_0809_),
    .A1(_0885_),
    .S(net449),
    .X(_0886_));
 sg13g2_nor2_1 _1807_ (.A(net454),
    .B(_0746_),
    .Y(_0887_));
 sg13g2_a21o_2 _1808_ (.A2(_0886_),
    .A1(net455),
    .B1(_0887_),
    .X(_0888_));
 sg13g2_o21ai_1 _1809_ (.B1(_0888_),
    .Y(_0889_),
    .A1(_0868_),
    .A2(_0884_));
 sg13g2_or4_1 _1810_ (.A(_0724_),
    .B(_0868_),
    .C(_0884_),
    .D(_0888_),
    .X(_0890_));
 sg13g2_nand2_1 _1811_ (.Y(_0891_),
    .A(_0889_),
    .B(_0890_));
 sg13g2_xor2_1 _1812_ (.B(_0891_),
    .A(_0883_),
    .X(_0892_));
 sg13g2_nand2_1 _1813_ (.Y(_0893_),
    .A(\firEngine.firInst.accQ[8] ),
    .B(_0892_));
 sg13g2_xnor2_1 _1814_ (.Y(_0894_),
    .A(\firEngine.firInst.accQ[8] ),
    .B(_0892_));
 sg13g2_xnor2_1 _1815_ (.Y(_0895_),
    .A(_0880_),
    .B(_0894_));
 sg13g2_o21ai_1 _1816_ (.B1(net530),
    .Y(_0896_),
    .A1(net713),
    .A2(net536));
 sg13g2_a21oi_1 _1817_ (.A1(net536),
    .A2(_0895_),
    .Y(_0072_),
    .B1(_0896_));
 sg13g2_a21oi_1 _1818_ (.A1(_0889_),
    .A2(_0890_),
    .Y(_0897_),
    .B1(net492));
 sg13g2_or4_1 _1819_ (.A(_0855_),
    .B(_0872_),
    .C(_0882_),
    .D(_0897_),
    .X(_0898_));
 sg13g2_nor2_1 _1820_ (.A(net450),
    .B(_0888_),
    .Y(_0899_));
 sg13g2_a21oi_1 _1821_ (.A1(_0869_),
    .A2(_0888_),
    .Y(_0900_),
    .B1(net450));
 sg13g2_mux2_1 _1822_ (.A0(_0612_),
    .A1(_0862_),
    .S(_0737_),
    .X(_0901_));
 sg13g2_nand2_1 _1823_ (.Y(_0902_),
    .A(_0744_),
    .B(_0827_));
 sg13g2_a21oi_1 _1824_ (.A1(net449),
    .A2(_0901_),
    .Y(_0903_),
    .B1(net456));
 sg13g2_a22oi_1 _1825_ (.Y(_0904_),
    .B1(_0902_),
    .B2(_0903_),
    .A2(_0759_),
    .A1(net456));
 sg13g2_nor2_1 _1826_ (.A(net458),
    .B(_0904_),
    .Y(_0905_));
 sg13g2_mux2_1 _1827_ (.A0(_0905_),
    .A1(_0904_),
    .S(_0900_),
    .X(_0906_));
 sg13g2_xnor2_1 _1828_ (.Y(_0907_),
    .A(_0898_),
    .B(_0906_));
 sg13g2_nor2_1 _1829_ (.A(\firEngine.firInst.accQ[9] ),
    .B(_0907_),
    .Y(_0908_));
 sg13g2_nand2_1 _1830_ (.Y(_0909_),
    .A(\firEngine.firInst.accQ[9] ),
    .B(_0907_));
 sg13g2_nand2b_1 _1831_ (.Y(_0910_),
    .B(_0909_),
    .A_N(_0908_));
 sg13g2_o21ai_1 _1832_ (.B1(_0893_),
    .Y(_0911_),
    .A1(_0880_),
    .A2(_0894_));
 sg13g2_nor2_1 _1833_ (.A(_0910_),
    .B(_0911_),
    .Y(_0912_));
 sg13g2_nand2_1 _1834_ (.Y(_0913_),
    .A(_0910_),
    .B(_0911_));
 sg13g2_nor2_1 _1835_ (.A(_0751_),
    .B(_0912_),
    .Y(_0914_));
 sg13g2_o21ai_1 _1836_ (.B1(net529),
    .Y(_0915_),
    .A1(net703),
    .A2(net534));
 sg13g2_a21oi_1 _1837_ (.A1(_0913_),
    .A2(_0914_),
    .Y(_0073_),
    .B1(_0915_));
 sg13g2_nand2_1 _1838_ (.Y(_0916_),
    .A(_0729_),
    .B(_0906_));
 sg13g2_nor2b_1 _1839_ (.A(_0898_),
    .B_N(_0916_),
    .Y(_0917_));
 sg13g2_nand2_1 _1840_ (.Y(_0918_),
    .A(net452),
    .B(_0846_));
 sg13g2_a21oi_1 _1841_ (.A1(_0028_),
    .A2(_0745_),
    .Y(_0919_),
    .B1(net456));
 sg13g2_a22oi_1 _1842_ (.Y(_0920_),
    .B1(_0918_),
    .B2(_0919_),
    .A2(_0780_),
    .A1(net456));
 sg13g2_nor2_1 _1843_ (.A(net451),
    .B(_0904_),
    .Y(_0921_));
 sg13g2_nor4_1 _1844_ (.A(_0868_),
    .B(_0884_),
    .C(_0899_),
    .D(_0921_),
    .Y(_0922_));
 sg13g2_nor2_1 _1845_ (.A(net458),
    .B(_0920_),
    .Y(_0923_));
 sg13g2_mux2_1 _1846_ (.A0(_0920_),
    .A1(_0923_),
    .S(_0922_),
    .X(_0924_));
 sg13g2_xor2_1 _1847_ (.B(_0924_),
    .A(_0917_),
    .X(_0925_));
 sg13g2_nand2_1 _1848_ (.Y(_0926_),
    .A(\firEngine.firInst.accQ[10] ),
    .B(_0925_));
 sg13g2_nor2_1 _1849_ (.A(\firEngine.firInst.accQ[10] ),
    .B(_0925_),
    .Y(_0927_));
 sg13g2_xor2_1 _1850_ (.B(_0925_),
    .A(\firEngine.firInst.accQ[10] ),
    .X(_0928_));
 sg13g2_nor2_1 _1851_ (.A(_0894_),
    .B(_0910_),
    .Y(_0929_));
 sg13g2_o21ai_1 _1852_ (.B1(_0909_),
    .Y(_0930_),
    .A1(_0893_),
    .A2(_0908_));
 sg13g2_a21oi_1 _1853_ (.A1(_0881_),
    .A2(_0929_),
    .Y(_0931_),
    .B1(_0930_));
 sg13g2_xor2_1 _1854_ (.B(_0931_),
    .A(_0928_),
    .X(_0932_));
 sg13g2_o21ai_1 _1855_ (.B1(net529),
    .Y(_0933_),
    .A1(net712),
    .A2(net534));
 sg13g2_a21oi_1 _1856_ (.A1(net534),
    .A2(_0932_),
    .Y(_0074_),
    .B1(_0933_));
 sg13g2_nand2_1 _1857_ (.Y(_0934_),
    .A(_0729_),
    .B(_0924_));
 sg13g2_nand3b_1 _1858_ (.B(_0916_),
    .C(_0934_),
    .Y(_0935_),
    .A_N(_0898_));
 sg13g2_nand2_1 _1859_ (.Y(_0936_),
    .A(_0744_),
    .B(_0863_));
 sg13g2_a22oi_1 _1860_ (.Y(_0937_),
    .B1(_0919_),
    .B2(_0936_),
    .A2(_0794_),
    .A1(net456));
 sg13g2_and4_1 _1861_ (.A(_0869_),
    .B(_0888_),
    .C(_0904_),
    .D(_0920_),
    .X(_0938_));
 sg13g2_nand3b_1 _1862_ (.B(_0937_),
    .C(net448),
    .Y(_0939_),
    .A_N(_0938_));
 sg13g2_nor2_1 _1863_ (.A(net458),
    .B(_0937_),
    .Y(_0940_));
 sg13g2_o21ai_1 _1864_ (.B1(_0940_),
    .Y(_0941_),
    .A1(net450),
    .A2(_0938_));
 sg13g2_and2_1 _1865_ (.A(_0939_),
    .B(_0941_),
    .X(_0942_));
 sg13g2_xnor2_1 _1866_ (.Y(_0943_),
    .A(_0935_),
    .B(_0942_));
 sg13g2_nand2b_1 _1867_ (.Y(_0944_),
    .B(_0943_),
    .A_N(\firEngine.firInst.accQ[11] ));
 sg13g2_nand2b_1 _1868_ (.Y(_0945_),
    .B(\firEngine.firInst.accQ[11] ),
    .A_N(_0943_));
 sg13g2_nand2_1 _1869_ (.Y(_0946_),
    .A(_0944_),
    .B(_0945_));
 sg13g2_o21ai_1 _1870_ (.B1(_0926_),
    .Y(_0947_),
    .A1(_0927_),
    .A2(_0931_));
 sg13g2_xor2_1 _1871_ (.B(_0947_),
    .A(_0946_),
    .X(_0948_));
 sg13g2_o21ai_1 _1872_ (.B1(net529),
    .Y(_0949_),
    .A1(net697),
    .A2(net533));
 sg13g2_a21oi_1 _1873_ (.A1(net534),
    .A2(_0948_),
    .Y(_0075_),
    .B1(_0949_));
 sg13g2_nand2_1 _1874_ (.Y(_0950_),
    .A(_0926_),
    .B(_0945_));
 sg13g2_a21o_1 _1875_ (.A2(_0950_),
    .A1(_0944_),
    .B1(_0930_),
    .X(_0951_));
 sg13g2_a21o_1 _1876_ (.A2(_0929_),
    .A1(_0881_),
    .B1(_0951_),
    .X(_0952_));
 sg13g2_nand2_1 _1877_ (.Y(_0953_),
    .A(_0927_),
    .B(_0945_));
 sg13g2_nand3_1 _1878_ (.B(_0952_),
    .C(_0953_),
    .A(_0944_),
    .Y(_0954_));
 sg13g2_nor2_1 _1879_ (.A(net492),
    .B(_0942_),
    .Y(_0955_));
 sg13g2_or2_1 _1880_ (.X(_0956_),
    .B(_0955_),
    .A(_0935_));
 sg13g2_nand2_1 _1881_ (.Y(_0957_),
    .A(_0730_),
    .B(_0810_));
 sg13g2_a21oi_1 _1882_ (.A1(\firEngine.firInst.coeffs[0][7] ),
    .A2(net449),
    .Y(_0958_),
    .B1(net456));
 sg13g2_o21ai_1 _1883_ (.B1(_0958_),
    .Y(_0959_),
    .A1(net449),
    .A2(_0885_));
 sg13g2_nand2_1 _1884_ (.Y(_0960_),
    .A(_0957_),
    .B(_0959_));
 sg13g2_a21oi_1 _1885_ (.A1(_0937_),
    .A2(_0938_),
    .Y(_0961_),
    .B1(net450));
 sg13g2_nor3_1 _1886_ (.A(net458),
    .B(_0960_),
    .C(_0961_),
    .Y(_0962_));
 sg13g2_a21o_1 _1887_ (.A2(_0961_),
    .A1(_0960_),
    .B1(_0962_),
    .X(_0963_));
 sg13g2_xnor2_1 _1888_ (.Y(_0964_),
    .A(_0956_),
    .B(_0963_));
 sg13g2_nand2_1 _1889_ (.Y(_0965_),
    .A(\firEngine.firInst.accQ[12] ),
    .B(_0964_));
 sg13g2_xnor2_1 _1890_ (.Y(_0966_),
    .A(\firEngine.firInst.accQ[12] ),
    .B(_0964_));
 sg13g2_xnor2_1 _1891_ (.Y(_0967_),
    .A(_0954_),
    .B(_0966_));
 sg13g2_o21ai_1 _1892_ (.B1(net529),
    .Y(_0968_),
    .A1(net694),
    .A2(net533));
 sg13g2_a21oi_1 _1893_ (.A1(net533),
    .A2(_0967_),
    .Y(_0076_),
    .B1(_0968_));
 sg13g2_a21oi_1 _1894_ (.A1(_0729_),
    .A2(_0963_),
    .Y(_0969_),
    .B1(_0956_));
 sg13g2_nand3_1 _1895_ (.B(_0938_),
    .C(_0960_),
    .A(_0937_),
    .Y(_0970_));
 sg13g2_nand2_1 _1896_ (.Y(_0971_),
    .A(net448),
    .B(_0970_));
 sg13g2_nor3_1 _1897_ (.A(net454),
    .B(_0828_),
    .C(_0829_),
    .Y(_0972_));
 sg13g2_o21ai_1 _1898_ (.B1(_0958_),
    .Y(_0973_),
    .A1(net449),
    .A2(_0901_));
 sg13g2_nor2b_2 _1899_ (.A(_0972_),
    .B_N(_0973_),
    .Y(_0974_));
 sg13g2_nand2_1 _1900_ (.Y(_0975_),
    .A(_0725_),
    .B(_0974_));
 sg13g2_mux2_1 _1901_ (.A0(_0974_),
    .A1(_0975_),
    .S(_0971_),
    .X(_0976_));
 sg13g2_xnor2_1 _1902_ (.Y(_0977_),
    .A(_0969_),
    .B(_0976_));
 sg13g2_nor2_1 _1903_ (.A(\firEngine.firInst.accQ[13] ),
    .B(_0977_),
    .Y(_0978_));
 sg13g2_xor2_1 _1904_ (.B(_0977_),
    .A(\firEngine.firInst.accQ[13] ),
    .X(_0979_));
 sg13g2_o21ai_1 _1905_ (.B1(_0965_),
    .Y(_0980_),
    .A1(_0954_),
    .A2(_0966_));
 sg13g2_xnor2_1 _1906_ (.Y(_0981_),
    .A(_0979_),
    .B(_0980_));
 sg13g2_o21ai_1 _1907_ (.B1(net529),
    .Y(_0982_),
    .A1(net714),
    .A2(net533));
 sg13g2_a21oi_1 _1908_ (.A1(net533),
    .A2(_0981_),
    .Y(_0077_),
    .B1(_0982_));
 sg13g2_nor2b_1 _1909_ (.A(_0966_),
    .B_N(_0979_),
    .Y(_0983_));
 sg13g2_nand4_1 _1910_ (.B(_0952_),
    .C(_0953_),
    .A(_0944_),
    .Y(_0984_),
    .D(_0983_));
 sg13g2_nor2_1 _1911_ (.A(_0965_),
    .B(_0978_),
    .Y(_0985_));
 sg13g2_a21oi_2 _1912_ (.B1(_0985_),
    .Y(_0986_),
    .A2(_0977_),
    .A1(\firEngine.firInst.accQ[13] ));
 sg13g2_and2_1 _1913_ (.A(_0028_),
    .B(net454),
    .X(_0987_));
 sg13g2_a21o_1 _1914_ (.A2(_0847_),
    .A1(net457),
    .B1(_0987_),
    .X(_0988_));
 sg13g2_o21ai_1 _1915_ (.B1(net448),
    .Y(_0989_),
    .A1(_0970_),
    .A2(_0974_));
 sg13g2_nand2_1 _1916_ (.Y(_0990_),
    .A(_0988_),
    .B(_0989_));
 sg13g2_o21ai_1 _1917_ (.B1(_0725_),
    .Y(_0991_),
    .A1(_0988_),
    .A2(_0989_));
 sg13g2_nor2b_1 _1918_ (.A(_0991_),
    .B_N(_0990_),
    .Y(_0992_));
 sg13g2_inv_1 _1919_ (.Y(_0993_),
    .A(_0992_));
 sg13g2_nor2_1 _1920_ (.A(net492),
    .B(_0976_),
    .Y(_0994_));
 sg13g2_nor2b_1 _1921_ (.A(_0994_),
    .B_N(_0969_),
    .Y(_0995_));
 sg13g2_xnor2_1 _1922_ (.Y(_0996_),
    .A(_0992_),
    .B(_0995_));
 sg13g2_xnor2_1 _1923_ (.Y(_0997_),
    .A(_0021_),
    .B(_0996_));
 sg13g2_and3_1 _1924_ (.X(_0998_),
    .A(_0984_),
    .B(_0986_),
    .C(_0997_));
 sg13g2_a21oi_1 _1925_ (.A1(_0984_),
    .A2(_0986_),
    .Y(_0999_),
    .B1(_0997_));
 sg13g2_or2_1 _1926_ (.X(_1000_),
    .B(_0999_),
    .A(_0998_));
 sg13g2_o21ai_1 _1927_ (.B1(net529),
    .Y(_1001_),
    .A1(net642),
    .A2(net533));
 sg13g2_a21oi_1 _1928_ (.A1(net533),
    .A2(_1000_),
    .Y(_0078_),
    .B1(_1001_));
 sg13g2_nand2b_1 _1929_ (.Y(_1002_),
    .B(\firEngine.firInst.accQ[14] ),
    .A_N(_0996_));
 sg13g2_nor2b_1 _1930_ (.A(_0999_),
    .B_N(_1002_),
    .Y(_1003_));
 sg13g2_a21oi_1 _1931_ (.A1(_0993_),
    .A2(_0995_),
    .Y(_1004_),
    .B1(net492));
 sg13g2_nand2_1 _1932_ (.Y(_1005_),
    .A(net448),
    .B(_0990_));
 sg13g2_a21o_1 _1933_ (.A2(_0864_),
    .A1(net457),
    .B1(_0987_),
    .X(_1006_));
 sg13g2_o21ai_1 _1934_ (.B1(_0725_),
    .Y(_1007_),
    .A1(_1005_),
    .A2(_1006_));
 sg13g2_a21oi_1 _1935_ (.A1(_1005_),
    .A2(_1006_),
    .Y(_1008_),
    .B1(_1007_));
 sg13g2_xnor2_1 _1936_ (.Y(_1009_),
    .A(_1004_),
    .B(_1008_));
 sg13g2_or2_1 _1937_ (.X(_1010_),
    .B(_1009_),
    .A(_0020_));
 sg13g2_nand2_1 _1938_ (.Y(_1011_),
    .A(_0020_),
    .B(_1009_));
 sg13g2_xor2_1 _1939_ (.B(_1009_),
    .A(_0020_),
    .X(_1012_));
 sg13g2_xnor2_1 _1940_ (.Y(_1013_),
    .A(_1003_),
    .B(_1012_));
 sg13g2_o21ai_1 _1941_ (.B1(net529),
    .Y(_1014_),
    .A1(net672),
    .A2(net533));
 sg13g2_a21oi_1 _1942_ (.A1(net535),
    .A2(_1013_),
    .Y(_0079_),
    .B1(_1014_));
 sg13g2_nand2_1 _1943_ (.Y(_1015_),
    .A(net398),
    .B(_0751_));
 sg13g2_a221oi_1 _1944_ (.B2(_1011_),
    .C1(_0997_),
    .B1(_1010_),
    .A1(_0984_),
    .Y(_1016_),
    .A2(_0986_));
 sg13g2_nand2_1 _1945_ (.Y(_1017_),
    .A(\firEngine.firInst.accQ[15] ),
    .B(_1009_));
 sg13g2_o21ai_1 _1946_ (.B1(_1017_),
    .Y(_1018_),
    .A1(_1002_),
    .A2(_1012_));
 sg13g2_a21o_1 _1947_ (.A2(_0886_),
    .A1(net457),
    .B1(_0987_),
    .X(_1019_));
 sg13g2_a21oi_1 _1948_ (.A1(_0989_),
    .A2(_1019_),
    .Y(_1020_),
    .B1(_1007_));
 sg13g2_xor2_1 _1949_ (.B(_1020_),
    .A(\firEngine.firInst.accQ[16] ),
    .X(_1021_));
 sg13g2_xnor2_1 _1950_ (.Y(_1022_),
    .A(_1004_),
    .B(_1021_));
 sg13g2_o21ai_1 _1951_ (.B1(_1022_),
    .Y(_1023_),
    .A1(_1016_),
    .A2(_1018_));
 sg13g2_or3_1 _1952_ (.A(_1016_),
    .B(_1018_),
    .C(_1022_),
    .X(_1024_));
 sg13g2_nand3_1 _1953_ (.B(_1023_),
    .C(_1024_),
    .A(net535),
    .Y(_1025_));
 sg13g2_a21oi_1 _1954_ (.A1(_1015_),
    .A2(_1025_),
    .Y(_0080_),
    .B1(_0755_));
 sg13g2_nand2_1 _1955_ (.Y(_1026_),
    .A(\firEngine.firInst.state[2] ),
    .B(_0659_));
 sg13g2_nand3_1 _1956_ (.B(_0635_),
    .C(_1026_),
    .A(net593),
    .Y(_1027_));
 sg13g2_nand2_1 _1957_ (.Y(_1028_),
    .A(net565),
    .B(net271));
 sg13g2_o21ai_1 _1958_ (.B1(_1028_),
    .Y(_0081_),
    .A1(_0665_),
    .A2(_1027_));
 sg13g2_a21oi_1 _1959_ (.A1(_0635_),
    .A2(_0636_),
    .Y(_1029_),
    .B1(\firEngine.firInst.sample_cnt_en ));
 sg13g2_inv_1 _1960_ (.Y(_1030_),
    .A(_1029_));
 sg13g2_o21ai_1 _1961_ (.B1(net593),
    .Y(_1031_),
    .A1(net330),
    .A2(net560));
 sg13g2_a21oi_1 _1962_ (.A1(net330),
    .A2(_1030_),
    .Y(_0082_),
    .B1(_1031_));
 sg13g2_nand2_1 _1963_ (.Y(_1032_),
    .A(net608),
    .B(net330));
 sg13g2_a22oi_1 _1964_ (.Y(_1033_),
    .B1(_1032_),
    .B2(net560),
    .A2(_1029_),
    .A1(net608));
 sg13g2_o21ai_1 _1965_ (.B1(net593),
    .Y(_1034_),
    .A1(net608),
    .A2(net330));
 sg13g2_nor2_1 _1966_ (.A(net609),
    .B(_1034_),
    .Y(_0083_));
 sg13g2_o21ai_1 _1967_ (.B1(net560),
    .Y(_1035_),
    .A1(_0011_),
    .A2(_1032_));
 sg13g2_a21oi_1 _1968_ (.A1(_0011_),
    .A2(_1032_),
    .Y(_1036_),
    .B1(_1035_));
 sg13g2_a21oi_1 _1969_ (.A1(net280),
    .A2(_1029_),
    .Y(_1037_),
    .B1(_1036_));
 sg13g2_nor2_1 _1970_ (.A(net563),
    .B(net281),
    .Y(_0084_));
 sg13g2_nand2_1 _1971_ (.Y(_1038_),
    .A(net560),
    .B(net1));
 sg13g2_nand2b_1 _1972_ (.Y(_1039_),
    .B(net524),
    .A_N(net438));
 sg13g2_o21ai_1 _1973_ (.B1(_1039_),
    .Y(_1040_),
    .A1(net662),
    .A2(net524));
 sg13g2_o21ai_1 _1974_ (.B1(net584),
    .Y(_1041_),
    .A1(net711),
    .A2(net509));
 sg13g2_a21oi_1 _1975_ (.A1(net509),
    .A2(_1040_),
    .Y(_0085_),
    .B1(_1041_));
 sg13g2_nand2b_1 _1976_ (.Y(_1042_),
    .B(net522),
    .A_N(\firEngine.firInst.coeffs[0][1] ));
 sg13g2_o21ai_1 _1977_ (.B1(_1042_),
    .Y(_1043_),
    .A1(\firEngine.firInst.coeffs[1][1] ),
    .A2(net522));
 sg13g2_o21ai_1 _1978_ (.B1(net578),
    .Y(_1044_),
    .A1(net438),
    .A2(net509));
 sg13g2_a21oi_1 _1979_ (.A1(net497),
    .A2(_1043_),
    .Y(_0086_),
    .B1(_1044_));
 sg13g2_nand2b_1 _1980_ (.Y(_1045_),
    .B(net515),
    .A_N(net396));
 sg13g2_o21ai_1 _1981_ (.B1(_1045_),
    .Y(_1046_),
    .A1(net432),
    .A2(net515));
 sg13g2_o21ai_1 _1982_ (.B1(net583),
    .Y(_1047_),
    .A1(net643),
    .A2(net497));
 sg13g2_a21oi_1 _1983_ (.A1(net497),
    .A2(_1046_),
    .Y(_0087_),
    .B1(_1047_));
 sg13g2_nand2b_1 _1984_ (.Y(_1048_),
    .B(net513),
    .A_N(\firEngine.firInst.coeffs[0][3] ));
 sg13g2_o21ai_1 _1985_ (.B1(_1048_),
    .Y(_1049_),
    .A1(net354),
    .A2(net514));
 sg13g2_o21ai_1 _1986_ (.B1(net577),
    .Y(_1050_),
    .A1(net396),
    .A2(net495));
 sg13g2_a21oi_1 _1987_ (.A1(net496),
    .A2(_1049_),
    .Y(_0088_),
    .B1(_1050_));
 sg13g2_nand2b_1 _1988_ (.Y(_1051_),
    .B(net520),
    .A_N(\firEngine.firInst.coeffs[0][4] ));
 sg13g2_o21ai_1 _1989_ (.B1(_1051_),
    .Y(_1052_),
    .A1(\firEngine.firInst.coeffs[1][4] ),
    .A2(net520));
 sg13g2_o21ai_1 _1990_ (.B1(net579),
    .Y(_1053_),
    .A1(net615),
    .A2(net501));
 sg13g2_a21oi_1 _1991_ (.A1(net501),
    .A2(_1052_),
    .Y(_0089_),
    .B1(_1053_));
 sg13g2_nand2b_1 _1992_ (.Y(_1054_),
    .B(net526),
    .A_N(net650));
 sg13g2_o21ai_1 _1993_ (.B1(_1054_),
    .Y(_1055_),
    .A1(net352),
    .A2(net520));
 sg13g2_o21ai_1 _1994_ (.B1(net580),
    .Y(_1056_),
    .A1(net676),
    .A2(net506));
 sg13g2_a21oi_1 _1995_ (.A1(net506),
    .A2(_1055_),
    .Y(_0090_),
    .B1(_1056_));
 sg13g2_nand2b_1 _1996_ (.Y(_1057_),
    .B(net527),
    .A_N(net638));
 sg13g2_o21ai_1 _1997_ (.B1(_1057_),
    .Y(_0237_),
    .A1(\firEngine.firInst.coeffs[1][6] ),
    .A2(net527));
 sg13g2_o21ai_1 _1998_ (.B1(net580),
    .Y(_0238_),
    .A1(net650),
    .A2(net507));
 sg13g2_a21oi_1 _1999_ (.A1(net507),
    .A2(_0237_),
    .Y(_0091_),
    .B1(_0238_));
 sg13g2_nand2_1 _2000_ (.Y(_0239_),
    .A(_0612_),
    .B(net524));
 sg13g2_o21ai_1 _2001_ (.B1(_0239_),
    .Y(_0240_),
    .A1(\firEngine.firInst.coeffs[1][7] ),
    .A2(net524));
 sg13g2_o21ai_1 _2002_ (.B1(net584),
    .Y(_0241_),
    .A1(net638),
    .A2(net507));
 sg13g2_a21oi_1 _2003_ (.A1(net507),
    .A2(_0240_),
    .Y(_0092_),
    .B1(_0241_));
 sg13g2_nand2b_1 _2004_ (.Y(_0242_),
    .B(net522),
    .A_N(net662));
 sg13g2_o21ai_1 _2005_ (.B1(_0242_),
    .Y(_0243_),
    .A1(net699),
    .A2(net522));
 sg13g2_o21ai_1 _2006_ (.B1(net585),
    .Y(_0244_),
    .A1(net707),
    .A2(net509));
 sg13g2_a21oi_1 _2007_ (.A1(net509),
    .A2(_0243_),
    .Y(_0093_),
    .B1(_0244_));
 sg13g2_nand2b_1 _2008_ (.Y(_0245_),
    .B(net516),
    .A_N(\firEngine.firInst.coeffs[1][1] ));
 sg13g2_o21ai_1 _2009_ (.B1(_0245_),
    .Y(_0246_),
    .A1(\firEngine.firInst.coeffs[2][1] ),
    .A2(net516));
 sg13g2_o21ai_1 _2010_ (.B1(net578),
    .Y(_0247_),
    .A1(net662),
    .A2(net498));
 sg13g2_a21oi_1 _2011_ (.A1(net499),
    .A2(_0246_),
    .Y(_0094_),
    .B1(_0247_));
 sg13g2_nand2b_1 _2012_ (.Y(_0248_),
    .B(net514),
    .A_N(net432));
 sg13g2_o21ai_1 _2013_ (.B1(_0248_),
    .Y(_0249_),
    .A1(net657),
    .A2(net512));
 sg13g2_o21ai_1 _2014_ (.B1(net577),
    .Y(_0250_),
    .A1(net698),
    .A2(net495));
 sg13g2_a21oi_1 _2015_ (.A1(net495),
    .A2(_0249_),
    .Y(_0095_),
    .B1(_0250_));
 sg13g2_nand2b_1 _2016_ (.Y(_0251_),
    .B(net513),
    .A_N(net354));
 sg13g2_o21ai_1 _2017_ (.B1(_0251_),
    .Y(_0252_),
    .A1(\firEngine.firInst.coeffs[2][3] ),
    .A2(net513));
 sg13g2_o21ai_1 _2018_ (.B1(net576),
    .Y(_0253_),
    .A1(net432),
    .A2(net494));
 sg13g2_a21oi_1 _2019_ (.A1(net500),
    .A2(_0252_),
    .Y(_0096_),
    .B1(_0253_));
 sg13g2_nand2b_1 _2020_ (.Y(_0254_),
    .B(net517),
    .A_N(\firEngine.firInst.coeffs[1][4] ));
 sg13g2_o21ai_1 _2021_ (.B1(_0254_),
    .Y(_0255_),
    .A1(\firEngine.firInst.coeffs[2][4] ),
    .A2(net517));
 sg13g2_o21ai_1 _2022_ (.B1(net579),
    .Y(_0256_),
    .A1(net354),
    .A2(net500));
 sg13g2_a21oi_1 _2023_ (.A1(net500),
    .A2(_0255_),
    .Y(_0097_),
    .B1(_0256_));
 sg13g2_nand2b_1 _2024_ (.Y(_0257_),
    .B(net520),
    .A_N(net352));
 sg13g2_o21ai_1 _2025_ (.B1(_0257_),
    .Y(_0258_),
    .A1(net617),
    .A2(net519));
 sg13g2_o21ai_1 _2026_ (.B1(net579),
    .Y(_0259_),
    .A1(net627),
    .A2(net503));
 sg13g2_a21oi_1 _2027_ (.A1(net505),
    .A2(_0258_),
    .Y(_0098_),
    .B1(_0259_));
 sg13g2_nand2b_1 _2028_ (.Y(_0260_),
    .B(net525),
    .A_N(\firEngine.firInst.coeffs[1][6] ));
 sg13g2_o21ai_1 _2029_ (.B1(_0260_),
    .Y(_0261_),
    .A1(\firEngine.firInst.coeffs[2][6] ),
    .A2(net525));
 sg13g2_o21ai_1 _2030_ (.B1(net580),
    .Y(_0262_),
    .A1(net352),
    .A2(net504));
 sg13g2_a21oi_1 _2031_ (.A1(net504),
    .A2(_0261_),
    .Y(_0099_),
    .B1(_0262_));
 sg13g2_nand2b_1 _2032_ (.Y(_0263_),
    .B(net526),
    .A_N(\firEngine.firInst.coeffs[1][7] ));
 sg13g2_o21ai_1 _2033_ (.B1(_0263_),
    .Y(_0264_),
    .A1(\firEngine.firInst.coeffs[2][7] ),
    .A2(net526));
 sg13g2_o21ai_1 _2034_ (.B1(net584),
    .Y(_0265_),
    .A1(net652),
    .A2(net508));
 sg13g2_a21oi_1 _2035_ (.A1(net507),
    .A2(_0264_),
    .Y(_0100_),
    .B1(_0265_));
 sg13g2_nand2b_1 _2036_ (.Y(_0266_),
    .B(net522),
    .A_N(\firEngine.firInst.coeffs[2][0] ));
 sg13g2_o21ai_1 _2037_ (.B1(_0266_),
    .Y(_0267_),
    .A1(net680),
    .A2(net522));
 sg13g2_o21ai_1 _2038_ (.B1(net580),
    .Y(_0268_),
    .A1(\firEngine.firInst.coeffs[1][7] ),
    .A2(net507));
 sg13g2_a21oi_1 _2039_ (.A1(net498),
    .A2(net681),
    .Y(_0101_),
    .B1(_0268_));
 sg13g2_nand2b_1 _2040_ (.Y(_0269_),
    .B(net515),
    .A_N(net693));
 sg13g2_o21ai_1 _2041_ (.B1(_0269_),
    .Y(_0270_),
    .A1(net634),
    .A2(net515));
 sg13g2_o21ai_1 _2042_ (.B1(net578),
    .Y(_0271_),
    .A1(net699),
    .A2(net497));
 sg13g2_a21oi_1 _2043_ (.A1(net497),
    .A2(_0270_),
    .Y(_0102_),
    .B1(_0271_));
 sg13g2_nand2b_1 _2044_ (.Y(_0272_),
    .B(net512),
    .A_N(net657));
 sg13g2_o21ai_1 _2045_ (.B1(_0272_),
    .Y(_0273_),
    .A1(net385),
    .A2(net512));
 sg13g2_o21ai_1 _2046_ (.B1(net576),
    .Y(_0274_),
    .A1(net693),
    .A2(net495));
 sg13g2_a21oi_1 _2047_ (.A1(net494),
    .A2(_0273_),
    .Y(_0103_),
    .B1(_0274_));
 sg13g2_nand2b_1 _2048_ (.Y(_0275_),
    .B(net517),
    .A_N(net434));
 sg13g2_o21ai_1 _2049_ (.B1(_0275_),
    .Y(_0276_),
    .A1(net372),
    .A2(net513));
 sg13g2_o21ai_1 _2050_ (.B1(net576),
    .Y(_0277_),
    .A1(net657),
    .A2(net496));
 sg13g2_a21oi_1 _2051_ (.A1(net500),
    .A2(_0276_),
    .Y(_0104_),
    .B1(_0277_));
 sg13g2_nand2b_1 _2052_ (.Y(_0278_),
    .B(net518),
    .A_N(\firEngine.firInst.coeffs[2][4] ));
 sg13g2_o21ai_1 _2053_ (.B1(_0278_),
    .Y(_0279_),
    .A1(\firEngine.firInst.coeffs[3][4] ),
    .A2(net518));
 sg13g2_o21ai_1 _2054_ (.B1(net579),
    .Y(_0280_),
    .A1(net434),
    .A2(net501));
 sg13g2_a21oi_1 _2055_ (.A1(net502),
    .A2(_0279_),
    .Y(_0105_),
    .B1(_0280_));
 sg13g2_nand2b_1 _2056_ (.Y(_0281_),
    .B(net519),
    .A_N(net617));
 sg13g2_o21ai_1 _2057_ (.B1(_0281_),
    .Y(_0282_),
    .A1(net644),
    .A2(net519));
 sg13g2_o21ai_1 _2058_ (.B1(net582),
    .Y(_0283_),
    .A1(net654),
    .A2(net503));
 sg13g2_a21oi_1 _2059_ (.A1(net502),
    .A2(_0282_),
    .Y(_0106_),
    .B1(_0283_));
 sg13g2_nand2b_1 _2060_ (.Y(_0284_),
    .B(net525),
    .A_N(net362));
 sg13g2_o21ai_1 _2061_ (.B1(_0284_),
    .Y(_0285_),
    .A1(net596),
    .A2(net525));
 sg13g2_o21ai_1 _2062_ (.B1(net581),
    .Y(_0286_),
    .A1(net617),
    .A2(net505));
 sg13g2_a21oi_1 _2063_ (.A1(net504),
    .A2(_0285_),
    .Y(_0107_),
    .B1(_0286_));
 sg13g2_nand2b_1 _2064_ (.Y(_0287_),
    .B(net526),
    .A_N(\firEngine.firInst.coeffs[2][7] ));
 sg13g2_o21ai_1 _2065_ (.B1(_0287_),
    .Y(_0288_),
    .A1(\firEngine.firInst.coeffs[3][7] ),
    .A2(net526));
 sg13g2_o21ai_1 _2066_ (.B1(net581),
    .Y(_0289_),
    .A1(net362),
    .A2(net504));
 sg13g2_a21oi_1 _2067_ (.A1(net504),
    .A2(_0288_),
    .Y(_0108_),
    .B1(_0289_));
 sg13g2_nand2b_1 _2068_ (.Y(_0290_),
    .B(net523),
    .A_N(\firEngine.firInst.coeffs[3][0] ));
 sg13g2_o21ai_1 _2069_ (.B1(_0290_),
    .Y(_0291_),
    .A1(\firEngine.firInst.coeffs[4][0] ),
    .A2(net523));
 sg13g2_o21ai_1 _2070_ (.B1(net580),
    .Y(_0292_),
    .A1(net674),
    .A2(net506));
 sg13g2_a21oi_1 _2071_ (.A1(net506),
    .A2(_0291_),
    .Y(_0109_),
    .B1(_0292_));
 sg13g2_nand2b_1 _2072_ (.Y(_0293_),
    .B(net514),
    .A_N(net634));
 sg13g2_o21ai_1 _2073_ (.B1(_0293_),
    .Y(_0294_),
    .A1(net647),
    .A2(net515));
 sg13g2_o21ai_1 _2074_ (.B1(net578),
    .Y(_0295_),
    .A1(net680),
    .A2(net497));
 sg13g2_a21oi_1 _2075_ (.A1(net495),
    .A2(_0294_),
    .Y(_0110_),
    .B1(_0295_));
 sg13g2_nand2b_1 _2076_ (.Y(_0296_),
    .B(net512),
    .A_N(net385));
 sg13g2_o21ai_1 _2077_ (.B1(_0296_),
    .Y(_0297_),
    .A1(net598),
    .A2(net512));
 sg13g2_o21ai_1 _2078_ (.B1(net576),
    .Y(_0298_),
    .A1(net634),
    .A2(net494));
 sg13g2_a21oi_1 _2079_ (.A1(net494),
    .A2(_0297_),
    .Y(_0111_),
    .B1(_0298_));
 sg13g2_nand2b_1 _2080_ (.Y(_0299_),
    .B(net517),
    .A_N(net372));
 sg13g2_o21ai_1 _2081_ (.B1(_0299_),
    .Y(_0300_),
    .A1(net350),
    .A2(net513));
 sg13g2_o21ai_1 _2082_ (.B1(net576),
    .Y(_0301_),
    .A1(net385),
    .A2(net494));
 sg13g2_a21oi_1 _2083_ (.A1(net500),
    .A2(_0300_),
    .Y(_0112_),
    .B1(_0301_));
 sg13g2_nand2b_1 _2084_ (.Y(_0302_),
    .B(net518),
    .A_N(\firEngine.firInst.coeffs[3][4] ));
 sg13g2_o21ai_1 _2085_ (.B1(_0302_),
    .Y(_0303_),
    .A1(\firEngine.firInst.coeffs[4][4] ),
    .A2(net517));
 sg13g2_o21ai_1 _2086_ (.B1(net579),
    .Y(_0304_),
    .A1(net372),
    .A2(net501));
 sg13g2_a21oi_1 _2087_ (.A1(net502),
    .A2(_0303_),
    .Y(_0113_),
    .B1(_0304_));
 sg13g2_nand2b_1 _2088_ (.Y(_0305_),
    .B(net519),
    .A_N(net644));
 sg13g2_o21ai_1 _2089_ (.B1(_0305_),
    .Y(_0306_),
    .A1(\firEngine.firInst.coeffs[4][5] ),
    .A2(net519));
 sg13g2_o21ai_1 _2090_ (.B1(net582),
    .Y(_0307_),
    .A1(net688),
    .A2(net502));
 sg13g2_a21oi_1 _2091_ (.A1(net502),
    .A2(_0306_),
    .Y(_0114_),
    .B1(_0307_));
 sg13g2_nand2b_1 _2092_ (.Y(_0308_),
    .B(net525),
    .A_N(net596));
 sg13g2_o21ai_1 _2093_ (.B1(_0308_),
    .Y(_0309_),
    .A1(\firEngine.firInst.coeffs[4][6] ),
    .A2(net525));
 sg13g2_o21ai_1 _2094_ (.B1(net581),
    .Y(_0310_),
    .A1(net644),
    .A2(net505));
 sg13g2_a21oi_1 _2095_ (.A1(net504),
    .A2(_0309_),
    .Y(_0115_),
    .B1(_0310_));
 sg13g2_nand2b_1 _2096_ (.Y(_0311_),
    .B(net525),
    .A_N(\firEngine.firInst.coeffs[3][7] ));
 sg13g2_o21ai_1 _2097_ (.B1(_0311_),
    .Y(_0312_),
    .A1(\firEngine.firInst.coeffs[4][7] ),
    .A2(net525));
 sg13g2_o21ai_1 _2098_ (.B1(net581),
    .Y(_0313_),
    .A1(net596),
    .A2(net504));
 sg13g2_a21oi_1 _2099_ (.A1(net508),
    .A2(_0312_),
    .Y(_0116_),
    .B1(_0313_));
 sg13g2_nand2b_1 _2100_ (.Y(_0314_),
    .B(net523),
    .A_N(\firEngine.firInst.coeffs[4][0] ));
 sg13g2_o21ai_1 _2101_ (.B1(_0314_),
    .Y(_0315_),
    .A1(net677),
    .A2(net523));
 sg13g2_o21ai_1 _2102_ (.B1(net580),
    .Y(_0316_),
    .A1(net686),
    .A2(net506));
 sg13g2_a21oi_1 _2103_ (.A1(net506),
    .A2(_0315_),
    .Y(_0117_),
    .B1(_0316_));
 sg13g2_nand2b_1 _2104_ (.Y(_0317_),
    .B(net515),
    .A_N(net647));
 sg13g2_o21ai_1 _2105_ (.B1(_0317_),
    .Y(_0318_),
    .A1(net640),
    .A2(net515));
 sg13g2_o21ai_1 _2106_ (.B1(net578),
    .Y(_0319_),
    .A1(net706),
    .A2(net497));
 sg13g2_a21oi_1 _2107_ (.A1(net497),
    .A2(_0318_),
    .Y(_0118_),
    .B1(_0319_));
 sg13g2_nand2b_1 _2108_ (.Y(_0320_),
    .B(net512),
    .A_N(net598));
 sg13g2_o21ai_1 _2109_ (.B1(_0320_),
    .Y(_0321_),
    .A1(net399),
    .A2(net512));
 sg13g2_o21ai_1 _2110_ (.B1(net576),
    .Y(_0322_),
    .A1(net647),
    .A2(net495));
 sg13g2_a21oi_1 _2111_ (.A1(net494),
    .A2(_0321_),
    .Y(_0119_),
    .B1(_0322_));
 sg13g2_nand2b_1 _2112_ (.Y(_0323_),
    .B(net513),
    .A_N(net350));
 sg13g2_o21ai_1 _2113_ (.B1(_0323_),
    .Y(_0324_),
    .A1(net356),
    .A2(net513));
 sg13g2_o21ai_1 _2114_ (.B1(net576),
    .Y(_0325_),
    .A1(net598),
    .A2(net494));
 sg13g2_a21oi_1 _2115_ (.A1(net500),
    .A2(_0324_),
    .Y(_0120_),
    .B1(_0325_));
 sg13g2_nand2b_1 _2116_ (.Y(_0326_),
    .B(net518),
    .A_N(\firEngine.firInst.coeffs[4][4] ));
 sg13g2_o21ai_1 _2117_ (.B1(_0326_),
    .Y(_0327_),
    .A1(\firEngine.firInst.coeffs[5][4] ),
    .A2(net517));
 sg13g2_o21ai_1 _2118_ (.B1(net579),
    .Y(_0328_),
    .A1(net350),
    .A2(net501));
 sg13g2_a21oi_1 _2119_ (.A1(net502),
    .A2(_0327_),
    .Y(_0121_),
    .B1(_0328_));
 sg13g2_nand2b_1 _2120_ (.Y(_0329_),
    .B(net519),
    .A_N(\firEngine.firInst.coeffs[4][5] ));
 sg13g2_o21ai_1 _2121_ (.B1(_0329_),
    .Y(_0330_),
    .A1(\firEngine.firInst.coeffs[5][5] ),
    .A2(net519));
 sg13g2_o21ai_1 _2122_ (.B1(net582),
    .Y(_0331_),
    .A1(net620),
    .A2(net503));
 sg13g2_a21oi_1 _2123_ (.A1(net502),
    .A2(_0330_),
    .Y(_0122_),
    .B1(_0331_));
 sg13g2_nand2b_1 _2124_ (.Y(_0332_),
    .B(net526),
    .A_N(\firEngine.firInst.coeffs[4][6] ));
 sg13g2_o21ai_1 _2125_ (.B1(_0332_),
    .Y(_0333_),
    .A1(net447),
    .A2(net526));
 sg13g2_o21ai_1 _2126_ (.B1(net580),
    .Y(_0334_),
    .A1(net690),
    .A2(net505));
 sg13g2_a21oi_1 _2127_ (.A1(net504),
    .A2(_0333_),
    .Y(_0123_),
    .B1(_0334_));
 sg13g2_nand2b_1 _2128_ (.Y(_0335_),
    .B(net527),
    .A_N(\firEngine.firInst.coeffs[4][7] ));
 sg13g2_o21ai_1 _2129_ (.B1(_0335_),
    .Y(_0336_),
    .A1(net631),
    .A2(net527));
 sg13g2_o21ai_1 _2130_ (.B1(net584),
    .Y(_0337_),
    .A1(\firEngine.firInst.coeffs[4][6] ),
    .A2(net508));
 sg13g2_a21oi_1 _2131_ (.A1(net508),
    .A2(net632),
    .Y(_0124_),
    .B1(_0337_));
 sg13g2_nand2b_1 _2132_ (.Y(_0338_),
    .B(net522),
    .A_N(\firEngine.firInst.coeffs[5][0] ));
 sg13g2_o21ai_1 _2133_ (.B1(_0338_),
    .Y(_0339_),
    .A1(net438),
    .A2(net522));
 sg13g2_o21ai_1 _2134_ (.B1(net584),
    .Y(_0340_),
    .A1(net668),
    .A2(net507));
 sg13g2_a21oi_1 _2135_ (.A1(net507),
    .A2(_0339_),
    .Y(_0125_),
    .B1(_0340_));
 sg13g2_nand2b_1 _2136_ (.Y(_0341_),
    .B(net516),
    .A_N(net640));
 sg13g2_o21ai_1 _2137_ (.B1(_0341_),
    .Y(_0342_),
    .A1(net643),
    .A2(net515));
 sg13g2_o21ai_1 _2138_ (.B1(net578),
    .Y(_0343_),
    .A1(net677),
    .A2(net498));
 sg13g2_a21oi_1 _2139_ (.A1(net498),
    .A2(_0342_),
    .Y(_0126_),
    .B1(_0343_));
 sg13g2_nand2b_1 _2140_ (.Y(_0344_),
    .B(net514),
    .A_N(net399));
 sg13g2_o21ai_1 _2141_ (.B1(_0344_),
    .Y(_0345_),
    .A1(net396),
    .A2(net512));
 sg13g2_o21ai_1 _2142_ (.B1(net577),
    .Y(_0346_),
    .A1(net640),
    .A2(net495));
 sg13g2_a21oi_1 _2143_ (.A1(net495),
    .A2(_0345_),
    .Y(_0127_),
    .B1(_0346_));
 sg13g2_nand2b_1 _2144_ (.Y(_0347_),
    .B(net513),
    .A_N(net356));
 sg13g2_o21ai_1 _2145_ (.B1(_0347_),
    .Y(_0348_),
    .A1(\firEngine.firInst.coeffs[0][3] ),
    .A2(net514));
 sg13g2_o21ai_1 _2146_ (.B1(net576),
    .Y(_0349_),
    .A1(net399),
    .A2(net494));
 sg13g2_a21oi_1 _2147_ (.A1(net500),
    .A2(_0348_),
    .Y(_0128_),
    .B1(_0349_));
 sg13g2_nand2b_1 _2148_ (.Y(_0350_),
    .B(net517),
    .A_N(\firEngine.firInst.coeffs[5][4] ));
 sg13g2_o21ai_1 _2149_ (.B1(_0350_),
    .Y(_0351_),
    .A1(\firEngine.firInst.coeffs[0][4] ),
    .A2(net517));
 sg13g2_o21ai_1 _2150_ (.B1(net579),
    .Y(_0352_),
    .A1(net356),
    .A2(net500));
 sg13g2_a21oi_1 _2151_ (.A1(net501),
    .A2(_0351_),
    .Y(_0129_),
    .B1(_0352_));
 sg13g2_nand2b_1 _2152_ (.Y(_0353_),
    .B(net519),
    .A_N(net692));
 sg13g2_o21ai_1 _2153_ (.B1(_0353_),
    .Y(_0354_),
    .A1(net650),
    .A2(net520));
 sg13g2_o21ai_1 _2154_ (.B1(net579),
    .Y(_0355_),
    .A1(net702),
    .A2(net502));
 sg13g2_a21oi_1 _2155_ (.A1(net505),
    .A2(_0354_),
    .Y(_0130_),
    .B1(_0355_));
 sg13g2_nand2b_1 _2156_ (.Y(_0356_),
    .B(net527),
    .A_N(net447));
 sg13g2_o21ai_1 _2157_ (.B1(_0356_),
    .Y(_0357_),
    .A1(net638),
    .A2(net528));
 sg13g2_o21ai_1 _2158_ (.B1(net580),
    .Y(_0358_),
    .A1(net692),
    .A2(net505));
 sg13g2_a21oi_1 _2159_ (.A1(net508),
    .A2(_0357_),
    .Y(_0131_),
    .B1(_0358_));
 sg13g2_nand2b_1 _2160_ (.Y(_0359_),
    .B(net527),
    .A_N(\firEngine.firInst.coeffs[5][7] ));
 sg13g2_o21ai_1 _2161_ (.B1(_0359_),
    .Y(_0360_),
    .A1(\firEngine.firInst.coeffs[0][7] ),
    .A2(net527));
 sg13g2_o21ai_1 _2162_ (.B1(net584),
    .Y(_0361_),
    .A1(net447),
    .A2(net508));
 sg13g2_a21oi_1 _2163_ (.A1(net508),
    .A2(_0360_),
    .Y(_0132_),
    .B1(_0361_));
 sg13g2_nor2b_1 _2164_ (.A(net551),
    .B_N(net401),
    .Y(_0362_));
 sg13g2_a21oi_1 _2165_ (.A1(net445),
    .A2(net552),
    .Y(_0363_),
    .B1(_0362_));
 sg13g2_o21ai_1 _2166_ (.B1(net587),
    .Y(_0364_),
    .A1(\firEngine.firInst.samples[0][0] ),
    .A2(net471));
 sg13g2_a21oi_1 _2167_ (.A1(net471),
    .A2(_0363_),
    .Y(_0133_),
    .B1(_0364_));
 sg13g2_nor2b_1 _2168_ (.A(net551),
    .B_N(\firEngine.firInst.samples[1][1] ),
    .Y(_0365_));
 sg13g2_a21oi_1 _2169_ (.A1(net287),
    .A2(net551),
    .Y(_0366_),
    .B1(_0365_));
 sg13g2_o21ai_1 _2170_ (.B1(net587),
    .Y(_0367_),
    .A1(net390),
    .A2(net471));
 sg13g2_a21oi_1 _2171_ (.A1(net471),
    .A2(_0366_),
    .Y(_0134_),
    .B1(_0367_));
 sg13g2_nor2b_1 _2172_ (.A(net549),
    .B_N(\firEngine.firInst.samples[1][2] ),
    .Y(_0368_));
 sg13g2_a21oi_1 _2173_ (.A1(net327),
    .A2(net549),
    .Y(_0369_),
    .B1(_0368_));
 sg13g2_o21ai_1 _2174_ (.B1(net586),
    .Y(_0370_),
    .A1(net410),
    .A2(net468));
 sg13g2_a21oi_1 _2175_ (.A1(net472),
    .A2(_0369_),
    .Y(_0135_),
    .B1(_0370_));
 sg13g2_nor2b_1 _2176_ (.A(net541),
    .B_N(net636),
    .Y(_0371_));
 sg13g2_a21oi_1 _2177_ (.A1(net305),
    .A2(net548),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_o21ai_1 _2178_ (.B1(net572),
    .Y(_0373_),
    .A1(net641),
    .A2(net469));
 sg13g2_a21oi_1 _2179_ (.A1(net469),
    .A2(_0372_),
    .Y(_0136_),
    .B1(_0373_));
 sg13g2_nor2b_1 _2180_ (.A(net550),
    .B_N(net395),
    .Y(_0374_));
 sg13g2_a21oi_1 _2181_ (.A1(net302),
    .A2(net550),
    .Y(_0375_),
    .B1(_0374_));
 sg13g2_o21ai_1 _2182_ (.B1(net588),
    .Y(_0376_),
    .A1(net388),
    .A2(net476));
 sg13g2_a21oi_1 _2183_ (.A1(net473),
    .A2(_0375_),
    .Y(_0137_),
    .B1(_0376_));
 sg13g2_nor2b_1 _2184_ (.A(net542),
    .B_N(net444),
    .Y(_0377_));
 sg13g2_a21oi_1 _2185_ (.A1(net337),
    .A2(net542),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_o21ai_1 _2186_ (.B1(net574),
    .Y(_0379_),
    .A1(net340),
    .A2(net475));
 sg13g2_a21oi_1 _2187_ (.A1(net475),
    .A2(_0378_),
    .Y(_0138_),
    .B1(_0379_));
 sg13g2_nor2b_1 _2188_ (.A(net554),
    .B_N(\firEngine.firInst.samples[1][6] ),
    .Y(_0380_));
 sg13g2_a21oi_1 _2189_ (.A1(net289),
    .A2(net554),
    .Y(_0381_),
    .B1(_0380_));
 sg13g2_o21ai_1 _2190_ (.B1(net588),
    .Y(_0382_),
    .A1(net312),
    .A2(net477));
 sg13g2_a21oi_1 _2191_ (.A1(net476),
    .A2(_0381_),
    .Y(_0139_),
    .B1(_0382_));
 sg13g2_nor2b_1 _2192_ (.A(net553),
    .B_N(\firEngine.firInst.samples[1][7] ),
    .Y(_0383_));
 sg13g2_a21oi_1 _2193_ (.A1(net241),
    .A2(net553),
    .Y(_0384_),
    .B1(_0383_));
 sg13g2_o21ai_1 _2194_ (.B1(net588),
    .Y(_0385_),
    .A1(net316),
    .A2(net476));
 sg13g2_a21oi_1 _2195_ (.A1(net476),
    .A2(_0384_),
    .Y(_0140_),
    .B1(_0385_));
 sg13g2_nor2b_1 _2196_ (.A(net551),
    .B_N(\firEngine.firInst.samples[2][0] ),
    .Y(_0386_));
 sg13g2_a21oi_1 _2197_ (.A1(net551),
    .A2(\firEngine.firInst.samples[0][0] ),
    .Y(_0387_),
    .B1(_0386_));
 sg13g2_o21ai_1 _2198_ (.B1(net587),
    .Y(_0388_),
    .A1(net401),
    .A2(net470));
 sg13g2_a21oi_1 _2199_ (.A1(net470),
    .A2(_0387_),
    .Y(_0141_),
    .B1(_0388_));
 sg13g2_nor2b_1 _2200_ (.A(net549),
    .B_N(net613),
    .Y(_0389_));
 sg13g2_a21oi_1 _2201_ (.A1(net551),
    .A2(net390),
    .Y(_0390_),
    .B1(_0389_));
 sg13g2_o21ai_1 _2202_ (.B1(net587),
    .Y(_0391_),
    .A1(net604),
    .A2(net470));
 sg13g2_a21oi_1 _2203_ (.A1(net470),
    .A2(_0390_),
    .Y(_0142_),
    .B1(_0391_));
 sg13g2_nor2b_1 _2204_ (.A(net548),
    .B_N(net602),
    .Y(_0392_));
 sg13g2_a21oi_1 _2205_ (.A1(net548),
    .A2(net410),
    .Y(_0393_),
    .B1(_0392_));
 sg13g2_o21ai_1 _2206_ (.B1(net586),
    .Y(_0394_),
    .A1(net635),
    .A2(net468));
 sg13g2_a21oi_1 _2207_ (.A1(net468),
    .A2(_0393_),
    .Y(_0143_),
    .B1(_0394_));
 sg13g2_nor2b_1 _2208_ (.A(net540),
    .B_N(net622),
    .Y(_0395_));
 sg13g2_a21oi_1 _2209_ (.A1(net541),
    .A2(\firEngine.firInst.samples[0][3] ),
    .Y(_0396_),
    .B1(_0395_));
 sg13g2_o21ai_1 _2210_ (.B1(net573),
    .Y(_0397_),
    .A1(net636),
    .A2(net468));
 sg13g2_a21oi_1 _2211_ (.A1(net468),
    .A2(_0396_),
    .Y(_0144_),
    .B1(_0397_));
 sg13g2_nor2b_1 _2212_ (.A(net550),
    .B_N(net386),
    .Y(_0398_));
 sg13g2_a21oi_1 _2213_ (.A1(net550),
    .A2(net388),
    .Y(_0399_),
    .B1(_0398_));
 sg13g2_o21ai_1 _2214_ (.B1(net586),
    .Y(_0400_),
    .A1(net395),
    .A2(net473));
 sg13g2_a21oi_1 _2215_ (.A1(net473),
    .A2(_0399_),
    .Y(_0145_),
    .B1(_0400_));
 sg13g2_nor2b_1 _2216_ (.A(net542),
    .B_N(net442),
    .Y(_0401_));
 sg13g2_a21oi_1 _2217_ (.A1(net542),
    .A2(net340),
    .Y(_0402_),
    .B1(_0401_));
 sg13g2_o21ai_1 _2218_ (.B1(net572),
    .Y(_0403_),
    .A1(net444),
    .A2(net464));
 sg13g2_a21oi_1 _2219_ (.A1(net464),
    .A2(_0402_),
    .Y(_0146_),
    .B1(_0403_));
 sg13g2_nor2b_1 _2220_ (.A(net553),
    .B_N(net403),
    .Y(_0404_));
 sg13g2_a21oi_1 _2221_ (.A1(net553),
    .A2(net312),
    .Y(_0405_),
    .B1(_0404_));
 sg13g2_o21ai_1 _2222_ (.B1(net588),
    .Y(_0406_),
    .A1(net630),
    .A2(net477));
 sg13g2_a21oi_1 _2223_ (.A1(net475),
    .A2(_0405_),
    .Y(_0147_),
    .B1(_0406_));
 sg13g2_nor2b_1 _2224_ (.A(net553),
    .B_N(net412),
    .Y(_0407_));
 sg13g2_a21oi_1 _2225_ (.A1(net553),
    .A2(net316),
    .Y(_0408_),
    .B1(_0407_));
 sg13g2_o21ai_1 _2226_ (.B1(net588),
    .Y(_0409_),
    .A1(net407),
    .A2(net477));
 sg13g2_a21oi_1 _2227_ (.A1(net477),
    .A2(_0408_),
    .Y(_0148_),
    .B1(_0409_));
 sg13g2_nor2b_1 _2228_ (.A(net549),
    .B_N(net618),
    .Y(_0410_));
 sg13g2_a21oi_1 _2229_ (.A1(net551),
    .A2(net401),
    .Y(_0411_),
    .B1(_0410_));
 sg13g2_o21ai_1 _2230_ (.B1(net587),
    .Y(_0412_),
    .A1(net629),
    .A2(net470));
 sg13g2_a21oi_1 _2231_ (.A1(net470),
    .A2(_0411_),
    .Y(_0149_),
    .B1(_0412_));
 sg13g2_nor2b_1 _2232_ (.A(net549),
    .B_N(\firEngine.firInst.samples[3][1] ),
    .Y(_0413_));
 sg13g2_a21oi_1 _2233_ (.A1(net551),
    .A2(net604),
    .Y(_0414_),
    .B1(_0413_));
 sg13g2_o21ai_1 _2234_ (.B1(net587),
    .Y(_0415_),
    .A1(\firEngine.firInst.samples[2][1] ),
    .A2(net470));
 sg13g2_a21oi_1 _2235_ (.A1(net470),
    .A2(net605),
    .Y(_0150_),
    .B1(_0415_));
 sg13g2_nor2b_1 _2236_ (.A(net548),
    .B_N(net599),
    .Y(_0416_));
 sg13g2_a21oi_1 _2237_ (.A1(net548),
    .A2(\firEngine.firInst.samples[1][2] ),
    .Y(_0417_),
    .B1(_0416_));
 sg13g2_o21ai_1 _2238_ (.B1(net586),
    .Y(_0418_),
    .A1(net602),
    .A2(net469));
 sg13g2_a21oi_1 _2239_ (.A1(net469),
    .A2(_0417_),
    .Y(_0151_),
    .B1(_0418_));
 sg13g2_nor2b_1 _2240_ (.A(net540),
    .B_N(\firEngine.firInst.samples[3][3] ),
    .Y(_0419_));
 sg13g2_a21oi_1 _2241_ (.A1(net540),
    .A2(\firEngine.firInst.samples[1][3] ),
    .Y(_0420_),
    .B1(_0419_));
 sg13g2_o21ai_1 _2242_ (.B1(net572),
    .Y(_0421_),
    .A1(net622),
    .A2(net468));
 sg13g2_a21oi_1 _2243_ (.A1(net468),
    .A2(_0420_),
    .Y(_0152_),
    .B1(_0421_));
 sg13g2_nor2b_1 _2244_ (.A(net552),
    .B_N(\firEngine.firInst.samples[3][4] ),
    .Y(_0422_));
 sg13g2_a21oi_1 _2245_ (.A1(net552),
    .A2(\firEngine.firInst.samples[1][4] ),
    .Y(_0423_),
    .B1(_0422_));
 sg13g2_o21ai_1 _2246_ (.B1(net587),
    .Y(_0424_),
    .A1(net386),
    .A2(net474));
 sg13g2_a21oi_1 _2247_ (.A1(net474),
    .A2(_0423_),
    .Y(_0153_),
    .B1(_0424_));
 sg13g2_nor2b_1 _2248_ (.A(net539),
    .B_N(net428),
    .Y(_0425_));
 sg13g2_a21oi_1 _2249_ (.A1(net539),
    .A2(\firEngine.firInst.samples[1][5] ),
    .Y(_0426_),
    .B1(_0425_));
 sg13g2_o21ai_1 _2250_ (.B1(net572),
    .Y(_0427_),
    .A1(net442),
    .A2(net463));
 sg13g2_a21oi_1 _2251_ (.A1(net464),
    .A2(_0426_),
    .Y(_0154_),
    .B1(_0427_));
 sg13g2_nor2b_1 _2252_ (.A(net547),
    .B_N(net344),
    .Y(_0428_));
 sg13g2_a21oi_1 _2253_ (.A1(net553),
    .A2(net630),
    .Y(_0429_),
    .B1(_0428_));
 sg13g2_o21ai_1 _2254_ (.B1(net588),
    .Y(_0430_),
    .A1(net403),
    .A2(net475));
 sg13g2_a21oi_1 _2255_ (.A1(net475),
    .A2(_0429_),
    .Y(_0155_),
    .B1(_0430_));
 sg13g2_nor2b_1 _2256_ (.A(net546),
    .B_N(\firEngine.firInst.samples[3][7] ),
    .Y(_0431_));
 sg13g2_a21oi_1 _2257_ (.A1(net553),
    .A2(net407),
    .Y(_0432_),
    .B1(_0431_));
 sg13g2_o21ai_1 _2258_ (.B1(net588),
    .Y(_0433_),
    .A1(\firEngine.firInst.samples[2][7] ),
    .A2(net476));
 sg13g2_a21oi_1 _2259_ (.A1(net476),
    .A2(net408),
    .Y(_0156_),
    .B1(_0433_));
 sg13g2_nor2_1 _2260_ (.A(net549),
    .B(_0611_),
    .Y(_0434_));
 sg13g2_a21oi_1 _2261_ (.A1(net549),
    .A2(\firEngine.firInst.samples[2][0] ),
    .Y(_0435_),
    .B1(_0434_));
 sg13g2_o21ai_1 _2262_ (.B1(net586),
    .Y(_0436_),
    .A1(net618),
    .A2(net472));
 sg13g2_a21oi_1 _2263_ (.A1(net472),
    .A2(_0435_),
    .Y(_0157_),
    .B1(_0436_));
 sg13g2_nor2_1 _2264_ (.A(net548),
    .B(_0610_),
    .Y(_0437_));
 sg13g2_a21oi_1 _2265_ (.A1(net549),
    .A2(net613),
    .Y(_0438_),
    .B1(_0437_));
 sg13g2_o21ai_1 _2266_ (.B1(net586),
    .Y(_0439_),
    .A1(net666),
    .A2(net472));
 sg13g2_a21oi_1 _2267_ (.A1(net472),
    .A2(_0438_),
    .Y(_0158_),
    .B1(_0439_));
 sg13g2_nor2_1 _2268_ (.A(net541),
    .B(_0609_),
    .Y(_0440_));
 sg13g2_a21oi_1 _2269_ (.A1(net541),
    .A2(net602),
    .Y(_0441_),
    .B1(_0440_));
 sg13g2_o21ai_1 _2270_ (.B1(net586),
    .Y(_0442_),
    .A1(net599),
    .A2(net469));
 sg13g2_a21oi_1 _2271_ (.A1(net468),
    .A2(_0441_),
    .Y(_0159_),
    .B1(_0442_));
 sg13g2_nor2_1 _2272_ (.A(net540),
    .B(_0608_),
    .Y(_0443_));
 sg13g2_a21oi_1 _2273_ (.A1(net540),
    .A2(net622),
    .Y(_0444_),
    .B1(_0443_));
 sg13g2_o21ai_1 _2274_ (.B1(net573),
    .Y(_0445_),
    .A1(net628),
    .A2(net463));
 sg13g2_a21oi_1 _2275_ (.A1(net463),
    .A2(_0444_),
    .Y(_0160_),
    .B1(_0445_));
 sg13g2_nor2_1 _2276_ (.A(net542),
    .B(_0607_),
    .Y(_0446_));
 sg13g2_a21oi_1 _2277_ (.A1(net550),
    .A2(net386),
    .Y(_0447_),
    .B1(_0446_));
 sg13g2_o21ai_1 _2278_ (.B1(net586),
    .Y(_0448_),
    .A1(net607),
    .A2(net469));
 sg13g2_a21oi_1 _2279_ (.A1(net469),
    .A2(_0447_),
    .Y(_0161_),
    .B1(_0448_));
 sg13g2_nor2_1 _2280_ (.A(net543),
    .B(_0606_),
    .Y(_0449_));
 sg13g2_a21oi_1 _2281_ (.A1(net543),
    .A2(\firEngine.firInst.samples[2][5] ),
    .Y(_0450_),
    .B1(_0449_));
 sg13g2_o21ai_1 _2282_ (.B1(net571),
    .Y(_0451_),
    .A1(net428),
    .A2(net463));
 sg13g2_a21oi_1 _2283_ (.A1(net464),
    .A2(_0450_),
    .Y(_0162_),
    .B1(_0451_));
 sg13g2_nor2_1 _2284_ (.A(net546),
    .B(_0605_),
    .Y(_0452_));
 sg13g2_a21oi_1 _2285_ (.A1(net546),
    .A2(net403),
    .Y(_0453_),
    .B1(_0452_));
 sg13g2_o21ai_1 _2286_ (.B1(net574),
    .Y(_0454_),
    .A1(net344),
    .A2(net475));
 sg13g2_a21oi_1 _2287_ (.A1(net475),
    .A2(_0453_),
    .Y(_0163_),
    .B1(_0454_));
 sg13g2_nor2_1 _2288_ (.A(_0603_),
    .B(net546),
    .Y(_0455_));
 sg13g2_a21oi_1 _2289_ (.A1(net546),
    .A2(net412),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_o21ai_1 _2290_ (.B1(net575),
    .Y(_0457_),
    .A1(net601),
    .A2(net476));
 sg13g2_a21oi_1 _2291_ (.A1(net475),
    .A2(_0456_),
    .Y(_0164_),
    .B1(_0457_));
 sg13g2_nand2_1 _2292_ (.Y(_0458_),
    .A(net537),
    .B(net648));
 sg13g2_a21oi_1 _2293_ (.A1(net548),
    .A2(net618),
    .Y(_0459_),
    .B1(net488));
 sg13g2_a221oi_1 _2294_ (.B2(_0459_),
    .C1(net562),
    .B1(_0458_),
    .A1(_0611_),
    .Y(_0165_),
    .A2(net488));
 sg13g2_nand2_1 _2295_ (.Y(_0460_),
    .A(net537),
    .B(net390));
 sg13g2_a21oi_1 _2296_ (.A1(net548),
    .A2(net666),
    .Y(_0461_),
    .B1(net488));
 sg13g2_a221oi_1 _2297_ (.B2(_0461_),
    .C1(net562),
    .B1(_0460_),
    .A1(_0610_),
    .Y(_0166_),
    .A2(net488));
 sg13g2_nand2_1 _2298_ (.Y(_0462_),
    .A(net537),
    .B(net410));
 sg13g2_a21oi_1 _2299_ (.A1(net541),
    .A2(net599),
    .Y(_0463_),
    .B1(net488));
 sg13g2_a221oi_1 _2300_ (.B2(_0463_),
    .C1(net561),
    .B1(_0462_),
    .A1(_0609_),
    .Y(_0167_),
    .A2(net487));
 sg13g2_nand2_1 _2301_ (.Y(_0464_),
    .A(net537),
    .B(\firEngine.firInst.samples[0][3] ));
 sg13g2_a21oi_1 _2302_ (.A1(net540),
    .A2(\firEngine.firInst.samples[3][3] ),
    .Y(_0465_),
    .B1(net487));
 sg13g2_a221oi_1 _2303_ (.B2(_0465_),
    .C1(net561),
    .B1(_0464_),
    .A1(_0608_),
    .Y(_0168_),
    .A2(net487));
 sg13g2_nand2_1 _2304_ (.Y(_0466_),
    .A(net537),
    .B(net388));
 sg13g2_a21oi_1 _2305_ (.A1(net542),
    .A2(\firEngine.firInst.samples[3][4] ),
    .Y(_0467_),
    .B1(net487));
 sg13g2_a221oi_1 _2306_ (.B2(_0467_),
    .C1(net561),
    .B1(_0466_),
    .A1(_0607_),
    .Y(_0169_),
    .A2(net489));
 sg13g2_nand2_1 _2307_ (.Y(_0468_),
    .A(net537),
    .B(net340));
 sg13g2_a21oi_1 _2308_ (.A1(net539),
    .A2(\firEngine.firInst.samples[3][5] ),
    .Y(_0469_),
    .B1(net487));
 sg13g2_a221oi_1 _2309_ (.B2(_0469_),
    .C1(net561),
    .B1(_0468_),
    .A1(_0606_),
    .Y(_0170_),
    .A2(net489));
 sg13g2_nand2_1 _2310_ (.Y(_0470_),
    .A(_0604_),
    .B(net312));
 sg13g2_a21oi_1 _2311_ (.A1(net546),
    .A2(net344),
    .Y(_0471_),
    .B1(net489));
 sg13g2_a221oi_1 _2312_ (.B2(_0471_),
    .C1(net561),
    .B1(_0470_),
    .A1(_0605_),
    .Y(_0171_),
    .A2(net489));
 sg13g2_nand2_1 _2313_ (.Y(_0472_),
    .A(net537),
    .B(net316));
 sg13g2_a21oi_1 _2314_ (.A1(net546),
    .A2(net601),
    .Y(_0473_),
    .B1(net489));
 sg13g2_a221oi_1 _2315_ (.B2(_0473_),
    .C1(net561),
    .B1(_0472_),
    .A1(_0603_),
    .Y(_0172_),
    .A2(net489));
 sg13g2_o21ai_1 _2316_ (.B1(net573),
    .Y(_0474_),
    .A1(net540),
    .A2(net368));
 sg13g2_a21oi_1 _2317_ (.A1(net541),
    .A2(_0611_),
    .Y(_0173_),
    .B1(_0474_));
 sg13g2_o21ai_1 _2318_ (.B1(net573),
    .Y(_0475_),
    .A1(net538),
    .A2(net426));
 sg13g2_a21oi_1 _2319_ (.A1(net540),
    .A2(_0610_),
    .Y(_0174_),
    .B1(_0475_));
 sg13g2_o21ai_1 _2320_ (.B1(net572),
    .Y(_0476_),
    .A1(net538),
    .A2(net332));
 sg13g2_a21oi_1 _2321_ (.A1(net538),
    .A2(_0609_),
    .Y(_0175_),
    .B1(_0476_));
 sg13g2_o21ai_1 _2322_ (.B1(net572),
    .Y(_0477_),
    .A1(net538),
    .A2(net358));
 sg13g2_a21oi_1 _2323_ (.A1(net539),
    .A2(_0608_),
    .Y(_0176_),
    .B1(_0477_));
 sg13g2_o21ai_1 _2324_ (.B1(net575),
    .Y(_0478_),
    .A1(net544),
    .A2(\firEngine.firInst.samples[5][4] ));
 sg13g2_a21oi_1 _2325_ (.A1(net546),
    .A2(_0607_),
    .Y(_0177_),
    .B1(_0478_));
 sg13g2_o21ai_1 _2326_ (.B1(net574),
    .Y(_0479_),
    .A1(net544),
    .A2(\firEngine.firInst.samples[5][5] ));
 sg13g2_a21oi_1 _2327_ (.A1(net545),
    .A2(_0606_),
    .Y(_0178_),
    .B1(_0479_));
 sg13g2_o21ai_1 _2328_ (.B1(net574),
    .Y(_0480_),
    .A1(net545),
    .A2(\firEngine.firInst.samples[5][6] ));
 sg13g2_a21oi_1 _2329_ (.A1(net544),
    .A2(_0605_),
    .Y(_0179_),
    .B1(_0480_));
 sg13g2_o21ai_1 _2330_ (.B1(net574),
    .Y(_0481_),
    .A1(\firEngine.firInst.samples[5][7] ),
    .A2(net545));
 sg13g2_a21oi_1 _2331_ (.A1(_0603_),
    .A2(net544),
    .Y(_0180_),
    .B1(_0481_));
 sg13g2_nor2b_1 _2332_ (.A(net539),
    .B_N(\firEngine.firInst.samples[10][0] ),
    .Y(_0482_));
 sg13g2_a21oi_1 _2333_ (.A1(net539),
    .A2(\firEngine.firInst.samples[5][0] ),
    .Y(_0483_),
    .B1(_0482_));
 sg13g2_o21ai_1 _2334_ (.B1(net571),
    .Y(_0484_),
    .A1(net342),
    .A2(net463));
 sg13g2_a21oi_1 _2335_ (.A1(net463),
    .A2(_0483_),
    .Y(_0181_),
    .B1(_0484_));
 sg13g2_nor2b_1 _2336_ (.A(net538),
    .B_N(net260),
    .Y(_0485_));
 sg13g2_a21oi_1 _2337_ (.A1(net538),
    .A2(\firEngine.firInst.samples[5][1] ),
    .Y(_0486_),
    .B1(_0485_));
 sg13g2_o21ai_1 _2338_ (.B1(net571),
    .Y(_0487_),
    .A1(net415),
    .A2(net461));
 sg13g2_a21oi_1 _2339_ (.A1(net461),
    .A2(_0486_),
    .Y(_0182_),
    .B1(_0487_));
 sg13g2_nor2b_1 _2340_ (.A(net538),
    .B_N(net286),
    .Y(_0488_));
 sg13g2_a21oi_1 _2341_ (.A1(net538),
    .A2(net332),
    .Y(_0489_),
    .B1(_0488_));
 sg13g2_o21ai_1 _2342_ (.B1(net566),
    .Y(_0490_),
    .A1(net614),
    .A2(net461));
 sg13g2_a21oi_1 _2343_ (.A1(net461),
    .A2(_0489_),
    .Y(_0183_),
    .B1(_0490_));
 sg13g2_nor2b_1 _2344_ (.A(net539),
    .B_N(\firEngine.firInst.samples[10][3] ),
    .Y(_0491_));
 sg13g2_a21oi_1 _2345_ (.A1(net543),
    .A2(net358),
    .Y(_0492_),
    .B1(_0491_));
 sg13g2_o21ai_1 _2346_ (.B1(net567),
    .Y(_0493_),
    .A1(net360),
    .A2(net462));
 sg13g2_a21oi_1 _2347_ (.A1(net462),
    .A2(_0492_),
    .Y(_0184_),
    .B1(_0493_));
 sg13g2_nor2b_1 _2348_ (.A(net544),
    .B_N(\firEngine.firInst.samples[10][4] ),
    .Y(_0494_));
 sg13g2_a21oi_1 _2349_ (.A1(net544),
    .A2(\firEngine.firInst.samples[5][4] ),
    .Y(_0495_),
    .B1(_0494_));
 sg13g2_o21ai_1 _2350_ (.B1(net574),
    .Y(_0496_),
    .A1(net413),
    .A2(net467));
 sg13g2_a21oi_1 _2351_ (.A1(net467),
    .A2(_0495_),
    .Y(_0185_),
    .B1(_0496_));
 sg13g2_nor2b_1 _2352_ (.A(net544),
    .B_N(\firEngine.firInst.samples[10][5] ),
    .Y(_0497_));
 sg13g2_a21oi_1 _2353_ (.A1(net544),
    .A2(\firEngine.firInst.samples[5][5] ),
    .Y(_0498_),
    .B1(_0497_));
 sg13g2_o21ai_1 _2354_ (.B1(net568),
    .Y(_0499_),
    .A1(net348),
    .A2(net467));
 sg13g2_a21oi_1 _2355_ (.A1(net467),
    .A2(_0498_),
    .Y(_0186_),
    .B1(_0499_));
 sg13g2_nor2b_1 _2356_ (.A(net545),
    .B_N(net311),
    .Y(_0500_));
 sg13g2_a21oi_1 _2357_ (.A1(net545),
    .A2(\firEngine.firInst.samples[5][6] ),
    .Y(_0501_),
    .B1(_0500_));
 sg13g2_o21ai_1 _2358_ (.B1(net569),
    .Y(_0502_),
    .A1(net376),
    .A2(net466));
 sg13g2_a21oi_1 _2359_ (.A1(net467),
    .A2(_0501_),
    .Y(_0187_),
    .B1(_0502_));
 sg13g2_nor2b_1 _2360_ (.A(net545),
    .B_N(\firEngine.firInst.samples[10][7] ),
    .Y(_0503_));
 sg13g2_a21oi_1 _2361_ (.A1(\firEngine.firInst.samples[5][7] ),
    .A2(net545),
    .Y(_0504_),
    .B1(_0503_));
 sg13g2_o21ai_1 _2362_ (.B1(net568),
    .Y(_0505_),
    .A1(net430),
    .A2(net466));
 sg13g2_a21oi_1 _2363_ (.A1(net466),
    .A2(_0504_),
    .Y(_0188_),
    .B1(_0505_));
 sg13g2_o21ai_1 _2364_ (.B1(net571),
    .Y(_0506_),
    .A1(\firEngine.firInst.samples[6][0] ),
    .A2(net487));
 sg13g2_a21oi_1 _2365_ (.A1(_0602_),
    .A2(net487),
    .Y(_0189_),
    .B1(_0506_));
 sg13g2_o21ai_1 _2366_ (.B1(net571),
    .Y(_0507_),
    .A1(\firEngine.firInst.samples[6][1] ),
    .A2(net481));
 sg13g2_a21oi_1 _2367_ (.A1(_0600_),
    .A2(net481),
    .Y(_0190_),
    .B1(_0507_));
 sg13g2_o21ai_1 _2368_ (.B1(net566),
    .Y(_0508_),
    .A1(\firEngine.firInst.samples[6][2] ),
    .A2(net479));
 sg13g2_a21oi_1 _2369_ (.A1(_0598_),
    .A2(net479),
    .Y(_0191_),
    .B1(_0508_));
 sg13g2_o21ai_1 _2370_ (.B1(net567),
    .Y(_0509_),
    .A1(\firEngine.firInst.samples[6][3] ),
    .A2(net479));
 sg13g2_a21oi_1 _2371_ (.A1(_0596_),
    .A2(net479),
    .Y(_0192_),
    .B1(_0509_));
 sg13g2_o21ai_1 _2372_ (.B1(net568),
    .Y(_0510_),
    .A1(\firEngine.firInst.samples[6][4] ),
    .A2(net490));
 sg13g2_a21oi_1 _2373_ (.A1(_0594_),
    .A2(net483),
    .Y(_0193_),
    .B1(_0510_));
 sg13g2_o21ai_1 _2374_ (.B1(net568),
    .Y(_0511_),
    .A1(\firEngine.firInst.samples[6][5] ),
    .A2(net486));
 sg13g2_a21oi_1 _2375_ (.A1(_0592_),
    .A2(net483),
    .Y(_0194_),
    .B1(_0511_));
 sg13g2_o21ai_1 _2376_ (.B1(net569),
    .Y(_0512_),
    .A1(\firEngine.firInst.samples[6][6] ),
    .A2(net485));
 sg13g2_a21oi_1 _2377_ (.A1(_0590_),
    .A2(net485),
    .Y(_0195_),
    .B1(_0512_));
 sg13g2_o21ai_1 _2378_ (.B1(net568),
    .Y(_0513_),
    .A1(\firEngine.firInst.samples[6][7] ),
    .A2(net485));
 sg13g2_a21oi_1 _2379_ (.A1(_0588_),
    .A2(net484),
    .Y(_0196_),
    .B1(_0513_));
 sg13g2_o21ai_1 _2380_ (.B1(net571),
    .Y(_0514_),
    .A1(net261),
    .A2(net487));
 sg13g2_a21oi_1 _2381_ (.A1(_0601_),
    .A2(net481),
    .Y(_0197_),
    .B1(_0514_));
 sg13g2_o21ai_1 _2382_ (.B1(net566),
    .Y(_0515_),
    .A1(\firEngine.firInst.samples[7][1] ),
    .A2(net481));
 sg13g2_a21oi_1 _2383_ (.A1(_0599_),
    .A2(net481),
    .Y(_0198_),
    .B1(_0515_));
 sg13g2_o21ai_1 _2384_ (.B1(net566),
    .Y(_0516_),
    .A1(net251),
    .A2(net479));
 sg13g2_a21oi_1 _2385_ (.A1(_0597_),
    .A2(net479),
    .Y(_0199_),
    .B1(_0516_));
 sg13g2_o21ai_1 _2386_ (.B1(net567),
    .Y(_0517_),
    .A1(\firEngine.firInst.samples[7][3] ),
    .A2(net480));
 sg13g2_a21oi_1 _2387_ (.A1(_0595_),
    .A2(net480),
    .Y(_0200_),
    .B1(_0517_));
 sg13g2_o21ai_1 _2388_ (.B1(net568),
    .Y(_0518_),
    .A1(\firEngine.firInst.samples[7][4] ),
    .A2(net483));
 sg13g2_a21oi_1 _2389_ (.A1(_0593_),
    .A2(net483),
    .Y(_0201_),
    .B1(_0518_));
 sg13g2_o21ai_1 _2390_ (.B1(net570),
    .Y(_0519_),
    .A1(\firEngine.firInst.samples[7][5] ),
    .A2(net483));
 sg13g2_a21oi_1 _2391_ (.A1(_0591_),
    .A2(net483),
    .Y(_0202_),
    .B1(_0519_));
 sg13g2_o21ai_1 _2392_ (.B1(net578),
    .Y(_0520_),
    .A1(net247),
    .A2(net484));
 sg13g2_a21oi_1 _2393_ (.A1(_0589_),
    .A2(net484),
    .Y(_0203_),
    .B1(_0520_));
 sg13g2_o21ai_1 _2394_ (.B1(net570),
    .Y(_0521_),
    .A1(net256),
    .A2(net484));
 sg13g2_a21oi_1 _2395_ (.A1(_0587_),
    .A2(net484),
    .Y(_0204_),
    .B1(_0521_));
 sg13g2_o21ai_1 _2396_ (.B1(net589),
    .Y(_0522_),
    .A1(net321),
    .A2(_0643_));
 sg13g2_a21oi_1 _2397_ (.A1(_0586_),
    .A2(_0643_),
    .Y(_0205_),
    .B1(net322));
 sg13g2_and2_1 _2398_ (.A(_0585_),
    .B(_0643_),
    .X(_0523_));
 sg13g2_o21ai_1 _2399_ (.B1(net589),
    .Y(_0524_),
    .A1(net708),
    .A2(\firEngine.i2sController.lrckCounter[0] ));
 sg13g2_nor3_1 _2400_ (.A(_0644_),
    .B(_0523_),
    .C(net709),
    .Y(_0206_));
 sg13g2_o21ai_1 _2401_ (.B1(net589),
    .Y(_0525_),
    .A1(net715),
    .A2(_0644_));
 sg13g2_nor2_1 _2402_ (.A(_0645_),
    .B(_0525_),
    .Y(_0207_));
 sg13g2_o21ai_1 _2403_ (.B1(net590),
    .Y(_0526_),
    .A1(net705),
    .A2(_0645_));
 sg13g2_nor2b_1 _2404_ (.A(_0526_),
    .B_N(_0646_),
    .Y(_0208_));
 sg13g2_xnor2_1 _2405_ (.Y(_0527_),
    .A(_0584_),
    .B(_0646_));
 sg13g2_nor2_1 _2406_ (.A(net564),
    .B(_0527_),
    .Y(_0209_));
 sg13g2_o21ai_1 _2407_ (.B1(\firEngine.firInst.accQ[16] ),
    .Y(_0528_),
    .A1(_0613_),
    .A2(_0614_));
 sg13g2_nor2_1 _2408_ (.A(\firEngine.i2sController.currentState[0] ),
    .B(\firEngine.i2sController.currentState[2] ),
    .Y(_0529_));
 sg13g2_nor2b_1 _2409_ (.A(_0529_),
    .B_N(net271),
    .Y(_0530_));
 sg13g2_nor2_1 _2410_ (.A(\firEngine.firInst.accQ[15] ),
    .B(\firEngine.firInst.accQ[14] ),
    .Y(_0531_));
 sg13g2_o21ai_1 _2411_ (.B1(net491),
    .Y(_0532_),
    .A1(\firEngine.firInst.accQ[16] ),
    .A2(_0531_));
 sg13g2_a21oi_1 _2412_ (.A1(\firEngine.firInst.accQ[7] ),
    .A2(_0528_),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_o21ai_1 _2413_ (.B1(net591),
    .Y(_0534_),
    .A1(net392),
    .A2(_0530_));
 sg13g2_nor2_1 _2414_ (.A(_0533_),
    .B(net393),
    .Y(_0210_));
 sg13g2_a21oi_1 _2415_ (.A1(\firEngine.firInst.accQ[8] ),
    .A2(_0528_),
    .Y(_0535_),
    .B1(_0532_));
 sg13g2_o21ai_1 _2416_ (.B1(net591),
    .Y(_0536_),
    .A1(net436),
    .A2(net491));
 sg13g2_nor2_1 _2417_ (.A(_0535_),
    .B(_0536_),
    .Y(_0211_));
 sg13g2_a21oi_1 _2418_ (.A1(\firEngine.firInst.accQ[9] ),
    .A2(_0528_),
    .Y(_0537_),
    .B1(_0532_));
 sg13g2_o21ai_1 _2419_ (.B1(net591),
    .Y(_0538_),
    .A1(net417),
    .A2(net491));
 sg13g2_nor2_1 _2420_ (.A(_0537_),
    .B(_0538_),
    .Y(_0212_));
 sg13g2_a21oi_1 _2421_ (.A1(\firEngine.firInst.accQ[10] ),
    .A2(_0528_),
    .Y(_0539_),
    .B1(_0532_));
 sg13g2_o21ai_1 _2422_ (.B1(net591),
    .Y(_0540_),
    .A1(net378),
    .A2(net491));
 sg13g2_nor2_1 _2423_ (.A(_0539_),
    .B(_0540_),
    .Y(_0213_));
 sg13g2_a21oi_1 _2424_ (.A1(\firEngine.firInst.accQ[11] ),
    .A2(_0528_),
    .Y(_0541_),
    .B1(_0532_));
 sg13g2_o21ai_1 _2425_ (.B1(net591),
    .Y(_0542_),
    .A1(net440),
    .A2(net491));
 sg13g2_nor2_1 _2426_ (.A(_0541_),
    .B(_0542_),
    .Y(_0214_));
 sg13g2_a21oi_1 _2427_ (.A1(\firEngine.firInst.accQ[12] ),
    .A2(_0528_),
    .Y(_0543_),
    .B1(_0532_));
 sg13g2_o21ai_1 _2428_ (.B1(net591),
    .Y(_0544_),
    .A1(net424),
    .A2(net491));
 sg13g2_nor2_1 _2429_ (.A(_0543_),
    .B(_0544_),
    .Y(_0215_));
 sg13g2_a21oi_1 _2430_ (.A1(\firEngine.firInst.accQ[13] ),
    .A2(_0528_),
    .Y(_0545_),
    .B1(_0532_));
 sg13g2_o21ai_1 _2431_ (.B1(net591),
    .Y(_0546_),
    .A1(net611),
    .A2(net491));
 sg13g2_nor2_1 _2432_ (.A(_0545_),
    .B(_0546_),
    .Y(_0216_));
 sg13g2_nor2b_1 _2433_ (.A(net491),
    .B_N(\firEngine.i2sController.dacDataQ[7] ),
    .Y(_0547_));
 sg13g2_a21oi_1 _2434_ (.A1(net695),
    .A2(_0528_),
    .Y(_0548_),
    .B1(_0532_));
 sg13g2_nor2_1 _2435_ (.A(_0547_),
    .B(_0548_),
    .Y(_0549_));
 sg13g2_nor2_1 _2436_ (.A(net565),
    .B(net696),
    .Y(_0217_));
 sg13g2_a21oi_1 _2437_ (.A1(\firEngine.i2sController.currentState[1] ),
    .A2(_0643_),
    .Y(_0550_),
    .B1(\firEngine.i2sController.currentState[2] ));
 sg13g2_xor2_1 _2438_ (.B(\firEngine.i2sController.lrckCounter[0] ),
    .A(\firEngine.i2sController.lrckCounter[1] ),
    .X(_0551_));
 sg13g2_xnor2_1 _2439_ (.Y(_0552_),
    .A(_0030_),
    .B(_0551_));
 sg13g2_mux4_1 _2440_ (.S0(\firEngine.i2sController.lrckCounter[0] ),
    .A0(\firEngine.i2sController.dacDataQ[7] ),
    .A1(\firEngine.i2sController.dacDataQ[6] ),
    .A2(\firEngine.i2sController.dacDataQ[5] ),
    .A3(\firEngine.i2sController.dacDataQ[4] ),
    .S1(_0552_),
    .X(_0553_));
 sg13g2_mux4_1 _2441_ (.S0(\firEngine.i2sController.lrckCounter[0] ),
    .A0(\firEngine.i2sController.dacDataQ[3] ),
    .A1(\firEngine.i2sController.dacDataQ[2] ),
    .A2(\firEngine.i2sController.dacDataQ[1] ),
    .A3(\firEngine.i2sController.dacDataQ[0] ),
    .S1(_0552_),
    .X(_0554_));
 sg13g2_nor2b_1 _2442_ (.A(_0554_),
    .B_N(\firEngine.i2sController.lrckCounter[2] ),
    .Y(_0555_));
 sg13g2_nand2_1 _2443_ (.Y(_0556_),
    .A(_0584_),
    .B(\firEngine.i2sController.currentState[1] ));
 sg13g2_nor3_1 _2444_ (.A(\firEngine.i2sController.lrckCounter[3] ),
    .B(_0555_),
    .C(_0556_),
    .Y(_0557_));
 sg13g2_o21ai_1 _2445_ (.B1(_0557_),
    .Y(_0558_),
    .A1(\firEngine.i2sController.lrckCounter[2] ),
    .A2(_0553_));
 sg13g2_o21ai_1 _2446_ (.B1(net590),
    .Y(_0559_),
    .A1(net382),
    .A2(_0550_));
 sg13g2_a21oi_1 _2447_ (.A1(_0550_),
    .A2(_0558_),
    .Y(_0218_),
    .B1(net383));
 sg13g2_nor3_1 _2448_ (.A(\firEngine.i2sController.lrckCounter[2] ),
    .B(\firEngine.i2sController.lrckCounter[1] ),
    .C(\firEngine.i2sController.lrckCounter[0] ),
    .Y(_0560_));
 sg13g2_nor2b_1 _2449_ (.A(_0560_),
    .B_N(\firEngine.i2sController.lrckCounter[3] ),
    .Y(_0561_));
 sg13g2_nor3_1 _2450_ (.A(_0661_),
    .B(_0556_),
    .C(_0561_),
    .Y(_0562_));
 sg13g2_a21oi_2 _2451_ (.B1(net459),
    .Y(_0563_),
    .A2(net719),
    .A1(_0634_));
 sg13g2_a22oi_1 _2452_ (.Y(_0564_),
    .B1(_0563_),
    .B2(\firEngine.adcData[0] ),
    .A2(net459),
    .A1(net300));
 sg13g2_nor2_1 _2453_ (.A(net564),
    .B(net301),
    .Y(_0219_));
 sg13g2_a22oi_1 _2454_ (.Y(_0565_),
    .B1(_0563_),
    .B2(net287),
    .A2(_0562_),
    .A1(\firEngine.adcData[0] ));
 sg13g2_nor2_1 _2455_ (.A(net564),
    .B(net288),
    .Y(_0220_));
 sg13g2_a22oi_1 _2456_ (.Y(_0566_),
    .B1(_0563_),
    .B2(net327),
    .A2(net459),
    .A1(net287));
 sg13g2_nor2_1 _2457_ (.A(net564),
    .B(_0566_),
    .Y(_0221_));
 sg13g2_a22oi_1 _2458_ (.Y(_0567_),
    .B1(_0563_),
    .B2(net305),
    .A2(net459),
    .A1(\firEngine.adcData[2] ));
 sg13g2_nor2_1 _2459_ (.A(net562),
    .B(net306),
    .Y(_0222_));
 sg13g2_a22oi_1 _2460_ (.Y(_0568_),
    .B1(_0563_),
    .B2(net302),
    .A2(net459),
    .A1(\firEngine.adcData[3] ));
 sg13g2_nor2_1 _2461_ (.A(net561),
    .B(net303),
    .Y(_0223_));
 sg13g2_a22oi_1 _2462_ (.Y(_0569_),
    .B1(_0563_),
    .B2(net337),
    .A2(net459),
    .A1(net302));
 sg13g2_nor2_1 _2463_ (.A(net561),
    .B(_0569_),
    .Y(_0224_));
 sg13g2_a22oi_1 _2464_ (.Y(_0570_),
    .B1(_0563_),
    .B2(net289),
    .A2(net459),
    .A1(\firEngine.adcData[5] ));
 sg13g2_nor2_1 _2465_ (.A(net562),
    .B(net290),
    .Y(_0225_));
 sg13g2_a22oi_1 _2466_ (.Y(_0571_),
    .B1(_0563_),
    .B2(net241),
    .A2(net459),
    .A1(\firEngine.adcData[6] ));
 sg13g2_nor2_1 _2467_ (.A(net562),
    .B(net242),
    .Y(_0226_));
 sg13g2_nand2_1 _2468_ (.Y(_0572_),
    .A(net584),
    .B(net532));
 sg13g2_nor3_1 _2469_ (.A(_0630_),
    .B(net492),
    .C(_0572_),
    .Y(_0227_));
 sg13g2_nor2_1 _2470_ (.A(_0735_),
    .B(_0572_),
    .Y(_0228_));
 sg13g2_nor3_1 _2471_ (.A(net492),
    .B(_0740_),
    .C(_0572_),
    .Y(_0229_));
 sg13g2_or2_1 _2472_ (.X(_0573_),
    .B(\firEngine.i2sController.currentState[1] ),
    .A(\firEngine.i2sController.currentState[0] ));
 sg13g2_and3_1 _2473_ (.X(_0574_),
    .A(net589),
    .B(net716),
    .C(_0634_));
 sg13g2_and4_1 _2474_ (.A(net589),
    .B(_0663_),
    .C(_0664_),
    .D(_0573_),
    .X(_0575_));
 sg13g2_nor2_1 _2475_ (.A(net552),
    .B(_0575_),
    .Y(_0576_));
 sg13g2_nor2_1 _2476_ (.A(_0574_),
    .B(_0576_),
    .Y(_0230_));
 sg13g2_o21ai_1 _2477_ (.B1(net590),
    .Y(_0577_),
    .A1(net243),
    .A2(_0641_));
 sg13g2_a21oi_1 _2478_ (.A1(_0583_),
    .A2(_0641_),
    .Y(_0231_),
    .B1(_0577_));
 sg13g2_o21ai_1 _2479_ (.B1(\firEngine.i2sController.lrck ),
    .Y(_0578_),
    .A1(_0584_),
    .A2(_0646_));
 sg13g2_a21oi_1 _2480_ (.A1(net295),
    .A2(_0578_),
    .Y(_0232_),
    .B1(net564));
 sg13g2_nor3_2 _2481_ (.A(net334),
    .B(_0583_),
    .C(_0641_),
    .Y(_0579_));
 sg13g2_o21ai_1 _2482_ (.B1(net590),
    .Y(_0580_),
    .A1(\firEngine.i2sController.sclk ),
    .A2(_0579_));
 sg13g2_a21oi_1 _2483_ (.A1(_0582_),
    .A2(_0579_),
    .Y(_0233_),
    .B1(_0580_));
 sg13g2_and2_1 _2484_ (.A(net589),
    .B(net4),
    .X(_0234_));
 sg13g2_and2_1 _2485_ (.A(net590),
    .B(net238),
    .X(_0235_));
 sg13g2_o21ai_1 _2486_ (.B1(net590),
    .Y(_0581_),
    .A1(\firEngine.i2sController.sclkCounter ),
    .A2(_0642_));
 sg13g2_nor2_1 _2487_ (.A(net335),
    .B(_0581_),
    .Y(_0236_));
 sg13g2_dfrbp_1 _2488_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net17),
    .D(net685),
    .Q_N(_1237_),
    .Q(\firEngine.firInst.state[0] ));
 sg13g2_dfrbp_1 _2489_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net18),
    .D(_0002_),
    .Q_N(_1238_),
    .Q(\firEngine.firInst.state[1] ));
 sg13g2_dfrbp_1 _2490_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net19),
    .D(net423),
    .Q_N(_1239_),
    .Q(\firEngine.firInst.state[2] ));
 sg13g2_dfrbp_1 _2491_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net20),
    .D(net308),
    .Q_N(_1240_),
    .Q(\firEngine.firInst.sample_cnt_en ));
 sg13g2_dfrbp_1 _2492_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net21),
    .D(net347),
    .Q_N(_1241_),
    .Q(\firEngine.i2sController.currentState[0] ));
 sg13g2_dfrbp_1 _2493_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net123),
    .D(\firEngine.i2sController.nextState[1] ),
    .Q_N(_1242_),
    .Q(\firEngine.i2sController.currentState[1] ));
 sg13g2_dfrbp_1 _2494_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net16),
    .D(\firEngine.i2sController.nextState[0] ),
    .Q_N(_1236_),
    .Q(\firEngine.i2sController.currentState[2] ));
 sg13g2_dfrbp_1 _2495_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net128),
    .D(_0032_),
    .Q_N(_1235_),
    .Q(\firEngine.spiSlave.csSynchronizer[0] ));
 sg13g2_dfrbp_1 _2496_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net127),
    .D(_0033_),
    .Q_N(_1234_),
    .Q(\firEngine.spiSlave.cs ));
 sg13g2_dfrbp_1 _2497_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net126),
    .D(net326),
    .Q_N(_1233_),
    .Q(\firEngine.clockConfig[0] ));
 sg13g2_dfrbp_1 _2498_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net124),
    .D(net371),
    .Q_N(_1232_),
    .Q(\firEngine.clockConfig[1] ));
 sg13g2_dfrbp_1 _2499_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net122),
    .D(_0036_),
    .Q_N(_1231_),
    .Q(\firEngine.clockConfig[2] ));
 sg13g2_dfrbp_1 _2500_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net120),
    .D(_0037_),
    .Q_N(_1230_),
    .Q(\firEngine.clockConfig[3] ));
 sg13g2_dfrbp_1 _2501_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net118),
    .D(net625),
    .Q_N(_1229_),
    .Q(\firEngine.configStore.serialOut ));
 sg13g2_dfrbp_1 _2502_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net116),
    .D(_0039_),
    .Q_N(_0031_),
    .Q(\firEngine.i2sController.mclkCounter[0] ));
 sg13g2_dfrbp_1 _2503_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net115),
    .D(net320),
    .Q_N(_1228_),
    .Q(\firEngine.i2sController.mclkCounter[1] ));
 sg13g2_dfrbp_1 _2504_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net114),
    .D(_0041_),
    .Q_N(_1227_),
    .Q(\firEngine.i2sController.mclkCounter[2] ));
 sg13g2_dfrbp_1 _2505_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net113),
    .D(_0042_),
    .Q_N(_1226_),
    .Q(\firEngine.i2sController.mclkCounter[3] ));
 sg13g2_dfrbp_1 _2506_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net112),
    .D(_0043_),
    .Q_N(_1225_),
    .Q(\firEngine.spiSlave.sclkSynchronizer[0] ));
 sg13g2_dfrbp_1 _2507_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net111),
    .D(_0044_),
    .Q_N(_1224_),
    .Q(\firEngine.spiSlave.sclkSynchronizer[1] ));
 sg13g2_dfrbp_1 _2508_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net110),
    .D(_0045_),
    .Q_N(_1223_),
    .Q(\firEngine.spiSlave.sclkSynchronizer[2] ));
 sg13g2_dfrbp_1 _2509_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net109),
    .D(_0046_),
    .Q_N(_1222_),
    .Q(\firEngine.spiSlave.mosiSynchronizer[0] ));
 sg13g2_dfrbp_1 _2510_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net108),
    .D(_0047_),
    .Q_N(_1221_),
    .Q(\firEngine.spiSlave.mosi ));
 sg13g2_dfrbp_1 _2511_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net107),
    .D(net274),
    .Q_N(_1220_),
    .Q(\firEngine.firInst.samples[10][0] ));
 sg13g2_dfrbp_1 _2512_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net105),
    .D(_0049_),
    .Q_N(_1219_),
    .Q(\firEngine.firInst.samples[10][1] ));
 sg13g2_dfrbp_1 _2513_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net103),
    .D(_0050_),
    .Q_N(_1218_),
    .Q(\firEngine.firInst.samples[10][2] ));
 sg13g2_dfrbp_1 _2514_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net101),
    .D(net266),
    .Q_N(_1217_),
    .Q(\firEngine.firInst.samples[10][3] ));
 sg13g2_dfrbp_1 _2515_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net99),
    .D(net310),
    .Q_N(_1216_),
    .Q(\firEngine.firInst.samples[10][4] ));
 sg13g2_dfrbp_1 _2516_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net97),
    .D(net246),
    .Q_N(_1215_),
    .Q(\firEngine.firInst.samples[10][5] ));
 sg13g2_dfrbp_1 _2517_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net95),
    .D(_0054_),
    .Q_N(_1214_),
    .Q(\firEngine.firInst.samples[10][6] ));
 sg13g2_dfrbp_1 _2518_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net93),
    .D(net329),
    .Q_N(_1213_),
    .Q(\firEngine.firInst.samples[10][7] ));
 sg13g2_dfrbp_1 _2519_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net91),
    .D(_0056_),
    .Q_N(_1212_),
    .Q(\firEngine.firInst.samples[9][0] ));
 sg13g2_dfrbp_1 _2520_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net89),
    .D(_0057_),
    .Q_N(_1211_),
    .Q(\firEngine.firInst.samples[9][1] ));
 sg13g2_dfrbp_1 _2521_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net87),
    .D(net285),
    .Q_N(_1210_),
    .Q(\firEngine.firInst.samples[9][2] ));
 sg13g2_dfrbp_1 _2522_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net85),
    .D(_0059_),
    .Q_N(_1209_),
    .Q(\firEngine.firInst.samples[9][3] ));
 sg13g2_dfrbp_1 _2523_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net83),
    .D(_0060_),
    .Q_N(_1208_),
    .Q(\firEngine.firInst.samples[9][4] ));
 sg13g2_dfrbp_1 _2524_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net81),
    .D(_0061_),
    .Q_N(_1207_),
    .Q(\firEngine.firInst.samples[9][5] ));
 sg13g2_dfrbp_1 _2525_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net79),
    .D(_0062_),
    .Q_N(_1206_),
    .Q(\firEngine.firInst.samples[9][6] ));
 sg13g2_dfrbp_1 _2526_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net77),
    .D(_0063_),
    .Q_N(_1205_),
    .Q(\firEngine.firInst.samples[9][7] ));
 sg13g2_dfrbp_1 _2527_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net75),
    .D(net367),
    .Q_N(_0008_),
    .Q(\firEngine.firInst.accQ[0] ));
 sg13g2_dfrbp_1 _2528_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net73),
    .D(net659),
    .Q_N(_1204_),
    .Q(\firEngine.firInst.accQ[1] ));
 sg13g2_dfrbp_1 _2529_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net71),
    .D(_0066_),
    .Q_N(_1203_),
    .Q(\firEngine.firInst.accQ[2] ));
 sg13g2_dfrbp_1 _2530_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net69),
    .D(net339),
    .Q_N(_1202_),
    .Q(\firEngine.firInst.accQ[3] ));
 sg13g2_dfrbp_1 _2531_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net67),
    .D(_0068_),
    .Q_N(_1201_),
    .Q(\firEngine.firInst.accQ[4] ));
 sg13g2_dfrbp_1 _2532_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net65),
    .D(_0069_),
    .Q_N(_1200_),
    .Q(\firEngine.firInst.accQ[5] ));
 sg13g2_dfrbp_1 _2533_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net63),
    .D(_0070_),
    .Q_N(_1199_),
    .Q(\firEngine.firInst.accQ[6] ));
 sg13g2_dfrbp_1 _2534_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net61),
    .D(_0071_),
    .Q_N(_1198_),
    .Q(\firEngine.firInst.accQ[7] ));
 sg13g2_dfrbp_1 _2535_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net59),
    .D(_0072_),
    .Q_N(_1197_),
    .Q(\firEngine.firInst.accQ[8] ));
 sg13g2_dfrbp_1 _2536_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net57),
    .D(_0073_),
    .Q_N(_1196_),
    .Q(\firEngine.firInst.accQ[9] ));
 sg13g2_dfrbp_1 _2537_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net55),
    .D(_0074_),
    .Q_N(_1195_),
    .Q(\firEngine.firInst.accQ[10] ));
 sg13g2_dfrbp_1 _2538_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net53),
    .D(_0075_),
    .Q_N(_1194_),
    .Q(\firEngine.firInst.accQ[11] ));
 sg13g2_dfrbp_1 _2539_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net51),
    .D(_0076_),
    .Q_N(_1193_),
    .Q(\firEngine.firInst.accQ[12] ));
 sg13g2_dfrbp_1 _2540_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net49),
    .D(_0077_),
    .Q_N(_1192_),
    .Q(\firEngine.firInst.accQ[13] ));
 sg13g2_dfrbp_1 _2541_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net47),
    .D(_0078_),
    .Q_N(_0021_),
    .Q(\firEngine.firInst.accQ[14] ));
 sg13g2_dfrbp_1 _2542_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net45),
    .D(net673),
    .Q_N(_0020_),
    .Q(\firEngine.firInst.accQ[15] ));
 sg13g2_dfrbp_1 _2543_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net43),
    .D(_0080_),
    .Q_N(_1191_),
    .Q(\firEngine.firInst.accQ[16] ));
 sg13g2_dfrbp_1 _2544_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net41),
    .D(net272),
    .Q_N(_1190_),
    .Q(\firEngine.firDataValid ));
 sg13g2_dfrbp_1 _2545_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net40),
    .D(net331),
    .Q_N(_1189_),
    .Q(\firEngine.firInst.sample_cnt[0] ));
 sg13g2_dfrbp_1 _2546_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net38),
    .D(_0083_),
    .Q_N(_1188_),
    .Q(\firEngine.firInst.sample_cnt[1] ));
 sg13g2_dfrbp_1 _2547_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net36),
    .D(_0084_),
    .Q_N(_0011_),
    .Q(\firEngine.firInst.sample_cnt[2] ));
 sg13g2_dfrbp_1 _2548_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net34),
    .D(_0085_),
    .Q_N(_0009_),
    .Q(\firEngine.firInst.coeffs[0][0] ));
 sg13g2_dfrbp_1 _2549_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net32),
    .D(net439),
    .Q_N(_0022_),
    .Q(\firEngine.firInst.coeffs[0][1] ));
 sg13g2_dfrbp_1 _2550_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net30),
    .D(_0087_),
    .Q_N(_0023_),
    .Q(\firEngine.firInst.coeffs[0][2] ));
 sg13g2_dfrbp_1 _2551_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net28),
    .D(net397),
    .Q_N(_0024_),
    .Q(\firEngine.firInst.coeffs[0][3] ));
 sg13g2_dfrbp_1 _2552_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net26),
    .D(net616),
    .Q_N(_0025_),
    .Q(\firEngine.firInst.coeffs[0][4] ));
 sg13g2_dfrbp_1 _2553_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net24),
    .D(_0090_),
    .Q_N(_0026_),
    .Q(\firEngine.firInst.coeffs[0][5] ));
 sg13g2_dfrbp_1 _2554_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net22),
    .D(net651),
    .Q_N(_0027_),
    .Q(\firEngine.firInst.coeffs[0][6] ));
 sg13g2_dfrbp_1 _2555_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net226),
    .D(net639),
    .Q_N(_0028_),
    .Q(\firEngine.firInst.coeffs[0][7] ));
 sg13g2_dfrbp_1 _2556_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net224),
    .D(_0093_),
    .Q_N(_1187_),
    .Q(\firEngine.firInst.coeffs[1][0] ));
 sg13g2_dfrbp_1 _2557_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net222),
    .D(net663),
    .Q_N(_1186_),
    .Q(\firEngine.firInst.coeffs[1][1] ));
 sg13g2_dfrbp_1 _2558_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net220),
    .D(_0095_),
    .Q_N(_1185_),
    .Q(\firEngine.firInst.coeffs[1][2] ));
 sg13g2_dfrbp_1 _2559_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net218),
    .D(net433),
    .Q_N(_1184_),
    .Q(\firEngine.firInst.coeffs[1][3] ));
 sg13g2_dfrbp_1 _2560_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net216),
    .D(net355),
    .Q_N(_1183_),
    .Q(\firEngine.firInst.coeffs[1][4] ));
 sg13g2_dfrbp_1 _2561_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net214),
    .D(_0098_),
    .Q_N(_1182_),
    .Q(\firEngine.firInst.coeffs[1][5] ));
 sg13g2_dfrbp_1 _2562_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net212),
    .D(net353),
    .Q_N(_1181_),
    .Q(\firEngine.firInst.coeffs[1][6] ));
 sg13g2_dfrbp_1 _2563_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net210),
    .D(net653),
    .Q_N(_1180_),
    .Q(\firEngine.firInst.coeffs[1][7] ));
 sg13g2_dfrbp_1 _2564_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net208),
    .D(net682),
    .Q_N(_1179_),
    .Q(\firEngine.firInst.coeffs[2][0] ));
 sg13g2_dfrbp_1 _2565_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net206),
    .D(_0102_),
    .Q_N(_1178_),
    .Q(\firEngine.firInst.coeffs[2][1] ));
 sg13g2_dfrbp_1 _2566_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net204),
    .D(_0103_),
    .Q_N(_1177_),
    .Q(\firEngine.firInst.coeffs[2][2] ));
 sg13g2_dfrbp_1 _2567_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net202),
    .D(_0104_),
    .Q_N(_1176_),
    .Q(\firEngine.firInst.coeffs[2][3] ));
 sg13g2_dfrbp_1 _2568_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net200),
    .D(net435),
    .Q_N(_1175_),
    .Q(\firEngine.firInst.coeffs[2][4] ));
 sg13g2_dfrbp_1 _2569_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net198),
    .D(_0106_),
    .Q_N(_1174_),
    .Q(\firEngine.firInst.coeffs[2][5] ));
 sg13g2_dfrbp_1 _2570_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net196),
    .D(_0107_),
    .Q_N(_1173_),
    .Q(\firEngine.firInst.coeffs[2][6] ));
 sg13g2_dfrbp_1 _2571_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net194),
    .D(net363),
    .Q_N(_1172_),
    .Q(\firEngine.firInst.coeffs[2][7] ));
 sg13g2_dfrbp_1 _2572_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net192),
    .D(net675),
    .Q_N(_1171_),
    .Q(\firEngine.firInst.coeffs[3][0] ));
 sg13g2_dfrbp_1 _2573_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net190),
    .D(_0110_),
    .Q_N(_1170_),
    .Q(\firEngine.firInst.coeffs[3][1] ));
 sg13g2_dfrbp_1 _2574_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net188),
    .D(_0111_),
    .Q_N(_1169_),
    .Q(\firEngine.firInst.coeffs[3][2] ));
 sg13g2_dfrbp_1 _2575_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net186),
    .D(_0112_),
    .Q_N(_1168_),
    .Q(\firEngine.firInst.coeffs[3][3] ));
 sg13g2_dfrbp_1 _2576_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net184),
    .D(net373),
    .Q_N(_1167_),
    .Q(\firEngine.firInst.coeffs[3][4] ));
 sg13g2_dfrbp_1 _2577_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net182),
    .D(net689),
    .Q_N(_1166_),
    .Q(\firEngine.firInst.coeffs[3][5] ));
 sg13g2_dfrbp_1 _2578_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net180),
    .D(net645),
    .Q_N(_1165_),
    .Q(\firEngine.firInst.coeffs[3][6] ));
 sg13g2_dfrbp_1 _2579_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net178),
    .D(net597),
    .Q_N(_1164_),
    .Q(\firEngine.firInst.coeffs[3][7] ));
 sg13g2_dfrbp_1 _2580_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net176),
    .D(net687),
    .Q_N(_1163_),
    .Q(\firEngine.firInst.coeffs[4][0] ));
 sg13g2_dfrbp_1 _2581_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net174),
    .D(_0118_),
    .Q_N(_1162_),
    .Q(\firEngine.firInst.coeffs[4][1] ));
 sg13g2_dfrbp_1 _2582_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net172),
    .D(_0119_),
    .Q_N(_1161_),
    .Q(\firEngine.firInst.coeffs[4][2] ));
 sg13g2_dfrbp_1 _2583_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net170),
    .D(_0120_),
    .Q_N(_1160_),
    .Q(\firEngine.firInst.coeffs[4][3] ));
 sg13g2_dfrbp_1 _2584_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net168),
    .D(net351),
    .Q_N(_1159_),
    .Q(\firEngine.firInst.coeffs[4][4] ));
 sg13g2_dfrbp_1 _2585_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net166),
    .D(net621),
    .Q_N(_1158_),
    .Q(\firEngine.firInst.coeffs[4][5] ));
 sg13g2_dfrbp_1 _2586_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net164),
    .D(net691),
    .Q_N(_1157_),
    .Q(\firEngine.firInst.coeffs[4][6] ));
 sg13g2_dfrbp_1 _2587_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net162),
    .D(net633),
    .Q_N(_1156_),
    .Q(\firEngine.firInst.coeffs[4][7] ));
 sg13g2_dfrbp_1 _2588_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net160),
    .D(net669),
    .Q_N(_1155_),
    .Q(\firEngine.firInst.coeffs[5][0] ));
 sg13g2_dfrbp_1 _2589_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net158),
    .D(_0126_),
    .Q_N(_1154_),
    .Q(\firEngine.firInst.coeffs[5][1] ));
 sg13g2_dfrbp_1 _2590_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net156),
    .D(_0127_),
    .Q_N(_1153_),
    .Q(\firEngine.firInst.coeffs[5][2] ));
 sg13g2_dfrbp_1 _2591_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net154),
    .D(net400),
    .Q_N(_1152_),
    .Q(\firEngine.firInst.coeffs[5][3] ));
 sg13g2_dfrbp_1 _2592_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net152),
    .D(net357),
    .Q_N(_1151_),
    .Q(\firEngine.firInst.coeffs[5][4] ));
 sg13g2_dfrbp_1 _2593_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net150),
    .D(_0130_),
    .Q_N(_1150_),
    .Q(\firEngine.firInst.coeffs[5][5] ));
 sg13g2_dfrbp_1 _2594_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net148),
    .D(_0131_),
    .Q_N(_1149_),
    .Q(\firEngine.firInst.coeffs[5][6] ));
 sg13g2_dfrbp_1 _2595_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net146),
    .D(net595),
    .Q_N(_1148_),
    .Q(\firEngine.firInst.coeffs[5][7] ));
 sg13g2_dfrbp_1 _2596_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net144),
    .D(net446),
    .Q_N(_1147_),
    .Q(\firEngine.firInst.samples[0][0] ));
 sg13g2_dfrbp_1 _2597_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net142),
    .D(net391),
    .Q_N(_1146_),
    .Q(\firEngine.firInst.samples[0][1] ));
 sg13g2_dfrbp_1 _2598_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net140),
    .D(net411),
    .Q_N(_1145_),
    .Q(\firEngine.firInst.samples[0][2] ));
 sg13g2_dfrbp_1 _2599_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net138),
    .D(_0136_),
    .Q_N(_1144_),
    .Q(\firEngine.firInst.samples[0][3] ));
 sg13g2_dfrbp_1 _2600_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net136),
    .D(_0137_),
    .Q_N(_1143_),
    .Q(\firEngine.firInst.samples[0][4] ));
 sg13g2_dfrbp_1 _2601_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net134),
    .D(_0138_),
    .Q_N(_1142_),
    .Q(\firEngine.firInst.samples[0][5] ));
 sg13g2_dfrbp_1 _2602_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net132),
    .D(net313),
    .Q_N(_1141_),
    .Q(\firEngine.firInst.samples[0][6] ));
 sg13g2_dfrbp_1 _2603_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net130),
    .D(net317),
    .Q_N(_1140_),
    .Q(\firEngine.firInst.samples[0][7] ));
 sg13g2_dfrbp_1 _2604_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net125),
    .D(net402),
    .Q_N(_1139_),
    .Q(\firEngine.firInst.samples[1][0] ));
 sg13g2_dfrbp_1 _2605_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net121),
    .D(_0142_),
    .Q_N(_1138_),
    .Q(\firEngine.firInst.samples[1][1] ));
 sg13g2_dfrbp_1 _2606_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net117),
    .D(_0143_),
    .Q_N(_1137_),
    .Q(\firEngine.firInst.samples[1][2] ));
 sg13g2_dfrbp_1 _2607_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net104),
    .D(net637),
    .Q_N(_1136_),
    .Q(\firEngine.firInst.samples[1][3] ));
 sg13g2_dfrbp_1 _2608_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net100),
    .D(_0145_),
    .Q_N(_1135_),
    .Q(\firEngine.firInst.samples[1][4] ));
 sg13g2_dfrbp_1 _2609_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net96),
    .D(_0146_),
    .Q_N(_1134_),
    .Q(\firEngine.firInst.samples[1][5] ));
 sg13g2_dfrbp_1 _2610_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net92),
    .D(_0147_),
    .Q_N(_1133_),
    .Q(\firEngine.firInst.samples[1][6] ));
 sg13g2_dfrbp_1 _2611_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net88),
    .D(_0148_),
    .Q_N(_1132_),
    .Q(\firEngine.firInst.samples[1][7] ));
 sg13g2_dfrbp_1 _2612_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net84),
    .D(_0149_),
    .Q_N(_1131_),
    .Q(\firEngine.firInst.samples[2][0] ));
 sg13g2_dfrbp_1 _2613_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net80),
    .D(net606),
    .Q_N(_1130_),
    .Q(\firEngine.firInst.samples[2][1] ));
 sg13g2_dfrbp_1 _2614_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net76),
    .D(net603),
    .Q_N(_1129_),
    .Q(\firEngine.firInst.samples[2][2] ));
 sg13g2_dfrbp_1 _2615_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net72),
    .D(net623),
    .Q_N(_1128_),
    .Q(\firEngine.firInst.samples[2][3] ));
 sg13g2_dfrbp_1 _2616_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net68),
    .D(net387),
    .Q_N(_1127_),
    .Q(\firEngine.firInst.samples[2][4] ));
 sg13g2_dfrbp_1 _2617_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net64),
    .D(net443),
    .Q_N(_1126_),
    .Q(\firEngine.firInst.samples[2][5] ));
 sg13g2_dfrbp_1 _2618_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net60),
    .D(_0155_),
    .Q_N(_1125_),
    .Q(\firEngine.firInst.samples[2][6] ));
 sg13g2_dfrbp_1 _2619_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net56),
    .D(net409),
    .Q_N(_1124_),
    .Q(\firEngine.firInst.samples[2][7] ));
 sg13g2_dfrbp_1 _2620_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net52),
    .D(net619),
    .Q_N(_1123_),
    .Q(\firEngine.firInst.samples[3][0] ));
 sg13g2_dfrbp_1 _2621_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net48),
    .D(net667),
    .Q_N(_1122_),
    .Q(\firEngine.firInst.samples[3][1] ));
 sg13g2_dfrbp_1 _2622_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net44),
    .D(_0159_),
    .Q_N(_1121_),
    .Q(\firEngine.firInst.samples[3][2] ));
 sg13g2_dfrbp_1 _2623_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net39),
    .D(_0160_),
    .Q_N(_1120_),
    .Q(\firEngine.firInst.samples[3][3] ));
 sg13g2_dfrbp_1 _2624_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net35),
    .D(_0161_),
    .Q_N(_1119_),
    .Q(\firEngine.firInst.samples[3][4] ));
 sg13g2_dfrbp_1 _2625_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net31),
    .D(net429),
    .Q_N(_1118_),
    .Q(\firEngine.firInst.samples[3][5] ));
 sg13g2_dfrbp_1 _2626_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net27),
    .D(_0163_),
    .Q_N(_1117_),
    .Q(\firEngine.firInst.samples[3][6] ));
 sg13g2_dfrbp_1 _2627_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net23),
    .D(_0164_),
    .Q_N(_1116_),
    .Q(\firEngine.firInst.samples[3][7] ));
 sg13g2_dfrbp_1 _2628_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net225),
    .D(net649),
    .Q_N(_1115_),
    .Q(\firEngine.firInst.samples[4][0] ));
 sg13g2_dfrbp_1 _2629_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net221),
    .D(_0166_),
    .Q_N(_1114_),
    .Q(\firEngine.firInst.samples[4][1] ));
 sg13g2_dfrbp_1 _2630_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net217),
    .D(net600),
    .Q_N(_1113_),
    .Q(\firEngine.firInst.samples[4][2] ));
 sg13g2_dfrbp_1 _2631_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net213),
    .D(net406),
    .Q_N(_1112_),
    .Q(\firEngine.firInst.samples[4][3] ));
 sg13g2_dfrbp_1 _2632_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net209),
    .D(net389),
    .Q_N(_1111_),
    .Q(\firEngine.firInst.samples[4][4] ));
 sg13g2_dfrbp_1 _2633_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net205),
    .D(net341),
    .Q_N(_1110_),
    .Q(\firEngine.firInst.samples[4][5] ));
 sg13g2_dfrbp_1 _2634_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net201),
    .D(_0171_),
    .Q_N(_1109_),
    .Q(\firEngine.firInst.samples[4][6] ));
 sg13g2_dfrbp_1 _2635_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net197),
    .D(_0172_),
    .Q_N(_1108_),
    .Q(\firEngine.firInst.samples[4][7] ));
 sg13g2_dfrbp_1 _2636_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net193),
    .D(net369),
    .Q_N(_0012_),
    .Q(\firEngine.firInst.samples[5][0] ));
 sg13g2_dfrbp_1 _2637_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net189),
    .D(net427),
    .Q_N(_0013_),
    .Q(\firEngine.firInst.samples[5][1] ));
 sg13g2_dfrbp_1 _2638_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net185),
    .D(net333),
    .Q_N(_0014_),
    .Q(\firEngine.firInst.samples[5][2] ));
 sg13g2_dfrbp_1 _2639_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net181),
    .D(net359),
    .Q_N(_0015_),
    .Q(\firEngine.firInst.samples[5][3] ));
 sg13g2_dfrbp_1 _2640_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net177),
    .D(net365),
    .Q_N(_0016_),
    .Q(\firEngine.firInst.samples[5][4] ));
 sg13g2_dfrbp_1 _2641_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net173),
    .D(net299),
    .Q_N(_0017_),
    .Q(\firEngine.firInst.samples[5][5] ));
 sg13g2_dfrbp_1 _2642_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net169),
    .D(net315),
    .Q_N(_0018_),
    .Q(\firEngine.firInst.samples[5][6] ));
 sg13g2_dfrbp_1 _2643_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net165),
    .D(net375),
    .Q_N(_0019_),
    .Q(\firEngine.firInst.samples[5][7] ));
 sg13g2_dfrbp_1 _2644_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net161),
    .D(net343),
    .Q_N(_1107_),
    .Q(\firEngine.firInst.samples[6][0] ));
 sg13g2_dfrbp_1 _2645_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net157),
    .D(net416),
    .Q_N(_1106_),
    .Q(\firEngine.firInst.samples[6][1] ));
 sg13g2_dfrbp_1 _2646_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net153),
    .D(_0183_),
    .Q_N(_1105_),
    .Q(\firEngine.firInst.samples[6][2] ));
 sg13g2_dfrbp_1 _2647_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net149),
    .D(net361),
    .Q_N(_1104_),
    .Q(\firEngine.firInst.samples[6][3] ));
 sg13g2_dfrbp_1 _2648_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net145),
    .D(net414),
    .Q_N(_1103_),
    .Q(\firEngine.firInst.samples[6][4] ));
 sg13g2_dfrbp_1 _2649_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net141),
    .D(net349),
    .Q_N(_1102_),
    .Q(\firEngine.firInst.samples[6][5] ));
 sg13g2_dfrbp_1 _2650_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net137),
    .D(net377),
    .Q_N(_1101_),
    .Q(\firEngine.firInst.samples[6][6] ));
 sg13g2_dfrbp_1 _2651_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net133),
    .D(net431),
    .Q_N(_1100_),
    .Q(\firEngine.firInst.samples[6][7] ));
 sg13g2_dfrbp_1 _2652_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net129),
    .D(net262),
    .Q_N(_1099_),
    .Q(\firEngine.firInst.samples[7][0] ));
 sg13g2_dfrbp_1 _2653_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net119),
    .D(net270),
    .Q_N(_1098_),
    .Q(\firEngine.firInst.samples[7][1] ));
 sg13g2_dfrbp_1 _2654_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net102),
    .D(net252),
    .Q_N(_1097_),
    .Q(\firEngine.firInst.samples[7][2] ));
 sg13g2_dfrbp_1 _2655_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net94),
    .D(net292),
    .Q_N(_1096_),
    .Q(\firEngine.firInst.samples[7][3] ));
 sg13g2_dfrbp_1 _2656_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net86),
    .D(net268),
    .Q_N(_1095_),
    .Q(\firEngine.firInst.samples[7][4] ));
 sg13g2_dfrbp_1 _2657_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net78),
    .D(net278),
    .Q_N(_1094_),
    .Q(\firEngine.firInst.samples[7][5] ));
 sg13g2_dfrbp_1 _2658_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net70),
    .D(net248),
    .Q_N(_1093_),
    .Q(\firEngine.firInst.samples[7][6] ));
 sg13g2_dfrbp_1 _2659_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net62),
    .D(net257),
    .Q_N(_1092_),
    .Q(\firEngine.firInst.samples[7][7] ));
 sg13g2_dfrbp_1 _2660_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net54),
    .D(_0197_),
    .Q_N(_1091_),
    .Q(\firEngine.firInst.samples[8][0] ));
 sg13g2_dfrbp_1 _2661_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net46),
    .D(net250),
    .Q_N(_1090_),
    .Q(\firEngine.firInst.samples[8][1] ));
 sg13g2_dfrbp_1 _2662_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net37),
    .D(_0199_),
    .Q_N(_1089_),
    .Q(\firEngine.firInst.samples[8][2] ));
 sg13g2_dfrbp_1 _2663_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net29),
    .D(net255),
    .Q_N(_1088_),
    .Q(\firEngine.firInst.samples[8][3] ));
 sg13g2_dfrbp_1 _2664_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net15),
    .D(net259),
    .Q_N(_1087_),
    .Q(\firEngine.firInst.samples[8][4] ));
 sg13g2_dfrbp_1 _2665_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net219),
    .D(net264),
    .Q_N(_1086_),
    .Q(\firEngine.firInst.samples[8][5] ));
 sg13g2_dfrbp_1 _2666_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net211),
    .D(_0203_),
    .Q_N(_1085_),
    .Q(\firEngine.firInst.samples[8][6] ));
 sg13g2_dfrbp_1 _2667_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net203),
    .D(_0204_),
    .Q_N(_1084_),
    .Q(\firEngine.firInst.samples[8][7] ));
 sg13g2_dfrbp_1 _2668_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net195),
    .D(net323),
    .Q_N(_0030_),
    .Q(\firEngine.i2sController.lrckCounter[0] ));
 sg13g2_dfrbp_1 _2669_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net187),
    .D(net710),
    .Q_N(_1083_),
    .Q(\firEngine.i2sController.lrckCounter[1] ));
 sg13g2_dfrbp_1 _2670_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net179),
    .D(_0207_),
    .Q_N(_1082_),
    .Q(\firEngine.i2sController.lrckCounter[2] ));
 sg13g2_dfrbp_1 _2671_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net171),
    .D(_0208_),
    .Q_N(_1081_),
    .Q(\firEngine.i2sController.lrckCounter[3] ));
 sg13g2_dfrbp_1 _2672_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net163),
    .D(_0209_),
    .Q_N(_1080_),
    .Q(\firEngine.i2sController.lrckCounter[4] ));
 sg13g2_dfrbp_1 _2673_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net155),
    .D(net394),
    .Q_N(_1079_),
    .Q(\firEngine.i2sController.dacDataQ[0] ));
 sg13g2_dfrbp_1 _2674_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net147),
    .D(net437),
    .Q_N(_1078_),
    .Q(\firEngine.i2sController.dacDataQ[1] ));
 sg13g2_dfrbp_1 _2675_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net139),
    .D(net418),
    .Q_N(_1077_),
    .Q(\firEngine.i2sController.dacDataQ[2] ));
 sg13g2_dfrbp_1 _2676_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net131),
    .D(net379),
    .Q_N(_1076_),
    .Q(\firEngine.i2sController.dacDataQ[3] ));
 sg13g2_dfrbp_1 _2677_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net106),
    .D(net441),
    .Q_N(_1075_),
    .Q(\firEngine.i2sController.dacDataQ[4] ));
 sg13g2_dfrbp_1 _2678_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net90),
    .D(net425),
    .Q_N(_1074_),
    .Q(\firEngine.i2sController.dacDataQ[5] ));
 sg13g2_dfrbp_1 _2679_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net74),
    .D(net612),
    .Q_N(_1073_),
    .Q(\firEngine.i2sController.dacDataQ[6] ));
 sg13g2_dfrbp_1 _2680_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net58),
    .D(_0217_),
    .Q_N(_1072_),
    .Q(\firEngine.i2sController.dacDataQ[7] ));
 sg13g2_dfrbp_1 _2681_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net42),
    .D(net384),
    .Q_N(_1071_),
    .Q(dac));
 sg13g2_dfrbp_1 _2682_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net25),
    .D(_0219_),
    .Q_N(_1070_),
    .Q(\firEngine.adcData[0] ));
 sg13g2_dfrbp_1 _2683_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net215),
    .D(_0220_),
    .Q_N(_1069_),
    .Q(\firEngine.adcData[1] ));
 sg13g2_dfrbp_1 _2684_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net199),
    .D(_0221_),
    .Q_N(_1068_),
    .Q(\firEngine.adcData[2] ));
 sg13g2_dfrbp_1 _2685_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net183),
    .D(_0222_),
    .Q_N(_1067_),
    .Q(\firEngine.adcData[3] ));
 sg13g2_dfrbp_1 _2686_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net167),
    .D(_0223_),
    .Q_N(_1066_),
    .Q(\firEngine.adcData[4] ));
 sg13g2_dfrbp_1 _2687_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net151),
    .D(_0224_),
    .Q_N(_1065_),
    .Q(\firEngine.adcData[5] ));
 sg13g2_dfrbp_1 _2688_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net135),
    .D(_0225_),
    .Q_N(_1064_),
    .Q(\firEngine.adcData[6] ));
 sg13g2_dfrbp_1 _2689_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net98),
    .D(_0226_),
    .Q_N(_1063_),
    .Q(\firEngine.adcData[7] ));
 sg13g2_dfrbp_1 _2690_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net66),
    .D(net276),
    .Q_N(_0029_),
    .Q(\firEngine.firInst.bit_cnt[0] ));
 sg13g2_dfrbp_1 _2691_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net50),
    .D(_0228_),
    .Q_N(_1062_),
    .Q(\firEngine.firInst.bit_cnt[1] ));
 sg13g2_dfrbp_1 _2692_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net33),
    .D(_0229_),
    .Q_N(_0010_),
    .Q(\firEngine.firInst.bit_cnt[2] ));
 sg13g2_dfrbp_1 _2693_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net223),
    .D(_0230_),
    .Q_N(_1061_),
    .Q(\firEngine.adcDataValid ));
 sg13g2_dfrbp_1 _2694_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net207),
    .D(net244),
    .Q_N(_0007_),
    .Q(\firEngine.i2sController.mclk ));
 sg13g2_dfrbp_1 _2695_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net175),
    .D(net296),
    .Q_N(_0005_),
    .Q(\firEngine.i2sController.lrck ));
 sg13g2_dfrbp_1 _2696_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net143),
    .D(net240),
    .Q_N(_0006_),
    .Q(\firEngine.i2sController.sclk ));
 sg13g2_dfrbp_1 _2697_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net82),
    .D(_0234_),
    .Q_N(_1060_),
    .Q(\firEngine.i2sController.adcSynchronizer[0] ));
 sg13g2_dfrbp_1 _2698_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net191),
    .D(_0235_),
    .Q_N(_1059_),
    .Q(\firEngine.i2sController.adcQ ));
 sg13g2_dfrbp_1 _2699_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net159),
    .D(net336),
    .Q_N(_1058_),
    .Q(\firEngine.i2sController.sclkCounter ));
 sg13g2_tiehi _2494__16 (.L_HI(net16));
 sg13g2_tiehi _2488__17 (.L_HI(net17));
 sg13g2_tiehi _2489__18 (.L_HI(net18));
 sg13g2_tiehi _2490__19 (.L_HI(net19));
 sg13g2_tiehi _2491__20 (.L_HI(net20));
 sg13g2_tiehi _2492__21 (.L_HI(net21));
 sg13g2_tiehi _2554__22 (.L_HI(net22));
 sg13g2_tiehi _2627__23 (.L_HI(net23));
 sg13g2_tiehi _2553__24 (.L_HI(net24));
 sg13g2_tiehi _2682__25 (.L_HI(net25));
 sg13g2_tiehi _2552__26 (.L_HI(net26));
 sg13g2_tiehi _2626__27 (.L_HI(net27));
 sg13g2_tiehi _2551__28 (.L_HI(net28));
 sg13g2_tiehi _2663__29 (.L_HI(net29));
 sg13g2_tiehi _2550__30 (.L_HI(net30));
 sg13g2_tiehi _2625__31 (.L_HI(net31));
 sg13g2_tiehi _2549__32 (.L_HI(net32));
 sg13g2_tiehi _2692__33 (.L_HI(net33));
 sg13g2_tiehi _2548__34 (.L_HI(net34));
 sg13g2_tiehi _2624__35 (.L_HI(net35));
 sg13g2_tiehi _2547__36 (.L_HI(net36));
 sg13g2_tiehi _2662__37 (.L_HI(net37));
 sg13g2_tiehi _2546__38 (.L_HI(net38));
 sg13g2_tiehi _2623__39 (.L_HI(net39));
 sg13g2_tiehi _2545__40 (.L_HI(net40));
 sg13g2_tiehi _2544__41 (.L_HI(net41));
 sg13g2_tiehi _2681__42 (.L_HI(net42));
 sg13g2_tiehi _2543__43 (.L_HI(net43));
 sg13g2_tiehi _2622__44 (.L_HI(net44));
 sg13g2_tiehi _2542__45 (.L_HI(net45));
 sg13g2_tiehi _2661__46 (.L_HI(net46));
 sg13g2_tiehi _2541__47 (.L_HI(net47));
 sg13g2_tiehi _2621__48 (.L_HI(net48));
 sg13g2_tiehi _2540__49 (.L_HI(net49));
 sg13g2_tiehi _2691__50 (.L_HI(net50));
 sg13g2_tiehi _2539__51 (.L_HI(net51));
 sg13g2_tiehi _2620__52 (.L_HI(net52));
 sg13g2_tiehi _2538__53 (.L_HI(net53));
 sg13g2_tiehi _2660__54 (.L_HI(net54));
 sg13g2_tiehi _2537__55 (.L_HI(net55));
 sg13g2_tiehi _2619__56 (.L_HI(net56));
 sg13g2_tiehi _2536__57 (.L_HI(net57));
 sg13g2_tiehi _2680__58 (.L_HI(net58));
 sg13g2_tiehi _2535__59 (.L_HI(net59));
 sg13g2_tiehi _2618__60 (.L_HI(net60));
 sg13g2_tiehi _2534__61 (.L_HI(net61));
 sg13g2_tiehi _2659__62 (.L_HI(net62));
 sg13g2_tiehi _2533__63 (.L_HI(net63));
 sg13g2_tiehi _2617__64 (.L_HI(net64));
 sg13g2_tiehi _2532__65 (.L_HI(net65));
 sg13g2_tiehi _2690__66 (.L_HI(net66));
 sg13g2_tiehi _2531__67 (.L_HI(net67));
 sg13g2_tiehi _2616__68 (.L_HI(net68));
 sg13g2_tiehi _2530__69 (.L_HI(net69));
 sg13g2_tiehi _2658__70 (.L_HI(net70));
 sg13g2_tiehi _2529__71 (.L_HI(net71));
 sg13g2_tiehi _2615__72 (.L_HI(net72));
 sg13g2_tiehi _2528__73 (.L_HI(net73));
 sg13g2_tiehi _2679__74 (.L_HI(net74));
 sg13g2_tiehi _2527__75 (.L_HI(net75));
 sg13g2_tiehi _2614__76 (.L_HI(net76));
 sg13g2_tiehi _2526__77 (.L_HI(net77));
 sg13g2_tiehi _2657__78 (.L_HI(net78));
 sg13g2_tiehi _2525__79 (.L_HI(net79));
 sg13g2_tiehi _2613__80 (.L_HI(net80));
 sg13g2_tiehi _2524__81 (.L_HI(net81));
 sg13g2_tiehi _2697__82 (.L_HI(net82));
 sg13g2_tiehi _2523__83 (.L_HI(net83));
 sg13g2_tiehi _2612__84 (.L_HI(net84));
 sg13g2_tiehi _2522__85 (.L_HI(net85));
 sg13g2_tiehi _2656__86 (.L_HI(net86));
 sg13g2_tiehi _2521__87 (.L_HI(net87));
 sg13g2_tiehi _2611__88 (.L_HI(net88));
 sg13g2_tiehi _2520__89 (.L_HI(net89));
 sg13g2_tiehi _2678__90 (.L_HI(net90));
 sg13g2_tiehi _2519__91 (.L_HI(net91));
 sg13g2_tiehi _2610__92 (.L_HI(net92));
 sg13g2_tiehi _2518__93 (.L_HI(net93));
 sg13g2_tiehi _2655__94 (.L_HI(net94));
 sg13g2_tiehi _2517__95 (.L_HI(net95));
 sg13g2_tiehi _2609__96 (.L_HI(net96));
 sg13g2_tiehi _2516__97 (.L_HI(net97));
 sg13g2_tiehi _2689__98 (.L_HI(net98));
 sg13g2_tiehi _2515__99 (.L_HI(net99));
 sg13g2_tiehi _2608__100 (.L_HI(net100));
 sg13g2_tiehi _2514__101 (.L_HI(net101));
 sg13g2_tiehi _2654__102 (.L_HI(net102));
 sg13g2_tiehi _2513__103 (.L_HI(net103));
 sg13g2_tiehi _2607__104 (.L_HI(net104));
 sg13g2_tiehi _2512__105 (.L_HI(net105));
 sg13g2_tiehi _2677__106 (.L_HI(net106));
 sg13g2_tiehi _2511__107 (.L_HI(net107));
 sg13g2_tiehi _2510__108 (.L_HI(net108));
 sg13g2_tiehi _2509__109 (.L_HI(net109));
 sg13g2_tiehi _2508__110 (.L_HI(net110));
 sg13g2_tiehi _2507__111 (.L_HI(net111));
 sg13g2_tiehi _2506__112 (.L_HI(net112));
 sg13g2_tiehi _2505__113 (.L_HI(net113));
 sg13g2_tiehi _2504__114 (.L_HI(net114));
 sg13g2_tiehi _2503__115 (.L_HI(net115));
 sg13g2_tiehi _2502__116 (.L_HI(net116));
 sg13g2_tiehi _2606__117 (.L_HI(net117));
 sg13g2_tiehi _2501__118 (.L_HI(net118));
 sg13g2_tiehi _2653__119 (.L_HI(net119));
 sg13g2_tiehi _2500__120 (.L_HI(net120));
 sg13g2_tiehi _2605__121 (.L_HI(net121));
 sg13g2_tiehi _2499__122 (.L_HI(net122));
 sg13g2_tiehi _2493__123 (.L_HI(net123));
 sg13g2_tiehi _2498__124 (.L_HI(net124));
 sg13g2_tiehi _2604__125 (.L_HI(net125));
 sg13g2_tiehi _2497__126 (.L_HI(net126));
 sg13g2_tiehi _2496__127 (.L_HI(net127));
 sg13g2_tiehi _2495__128 (.L_HI(net128));
 sg13g2_tiehi _2652__129 (.L_HI(net129));
 sg13g2_tiehi _2603__130 (.L_HI(net130));
 sg13g2_tiehi _2676__131 (.L_HI(net131));
 sg13g2_tiehi _2602__132 (.L_HI(net132));
 sg13g2_tiehi _2651__133 (.L_HI(net133));
 sg13g2_tiehi _2601__134 (.L_HI(net134));
 sg13g2_tiehi _2688__135 (.L_HI(net135));
 sg13g2_tiehi _2600__136 (.L_HI(net136));
 sg13g2_tiehi _2650__137 (.L_HI(net137));
 sg13g2_tiehi _2599__138 (.L_HI(net138));
 sg13g2_tiehi _2675__139 (.L_HI(net139));
 sg13g2_tiehi _2598__140 (.L_HI(net140));
 sg13g2_tiehi _2649__141 (.L_HI(net141));
 sg13g2_tiehi _2597__142 (.L_HI(net142));
 sg13g2_tiehi _2696__143 (.L_HI(net143));
 sg13g2_tiehi _2596__144 (.L_HI(net144));
 sg13g2_tiehi _2648__145 (.L_HI(net145));
 sg13g2_tiehi _2595__146 (.L_HI(net146));
 sg13g2_tiehi _2674__147 (.L_HI(net147));
 sg13g2_tiehi _2594__148 (.L_HI(net148));
 sg13g2_tiehi _2647__149 (.L_HI(net149));
 sg13g2_tiehi _2593__150 (.L_HI(net150));
 sg13g2_tiehi _2687__151 (.L_HI(net151));
 sg13g2_tiehi _2592__152 (.L_HI(net152));
 sg13g2_tiehi _2646__153 (.L_HI(net153));
 sg13g2_tiehi _2591__154 (.L_HI(net154));
 sg13g2_tiehi _2673__155 (.L_HI(net155));
 sg13g2_tiehi _2590__156 (.L_HI(net156));
 sg13g2_tiehi _2645__157 (.L_HI(net157));
 sg13g2_tiehi _2589__158 (.L_HI(net158));
 sg13g2_tiehi _2699__159 (.L_HI(net159));
 sg13g2_tiehi _2588__160 (.L_HI(net160));
 sg13g2_tiehi _2644__161 (.L_HI(net161));
 sg13g2_tiehi _2587__162 (.L_HI(net162));
 sg13g2_tiehi _2672__163 (.L_HI(net163));
 sg13g2_tiehi _2586__164 (.L_HI(net164));
 sg13g2_tiehi _2643__165 (.L_HI(net165));
 sg13g2_tiehi _2585__166 (.L_HI(net166));
 sg13g2_tiehi _2686__167 (.L_HI(net167));
 sg13g2_tiehi _2584__168 (.L_HI(net168));
 sg13g2_tiehi _2642__169 (.L_HI(net169));
 sg13g2_tiehi _2583__170 (.L_HI(net170));
 sg13g2_tiehi _2671__171 (.L_HI(net171));
 sg13g2_tiehi _2582__172 (.L_HI(net172));
 sg13g2_tiehi _2641__173 (.L_HI(net173));
 sg13g2_tiehi _2581__174 (.L_HI(net174));
 sg13g2_tiehi _2695__175 (.L_HI(net175));
 sg13g2_tiehi _2580__176 (.L_HI(net176));
 sg13g2_tiehi _2640__177 (.L_HI(net177));
 sg13g2_tiehi _2579__178 (.L_HI(net178));
 sg13g2_tiehi _2670__179 (.L_HI(net179));
 sg13g2_tiehi _2578__180 (.L_HI(net180));
 sg13g2_tiehi _2639__181 (.L_HI(net181));
 sg13g2_tiehi _2577__182 (.L_HI(net182));
 sg13g2_tiehi _2685__183 (.L_HI(net183));
 sg13g2_tiehi _2576__184 (.L_HI(net184));
 sg13g2_tiehi _2638__185 (.L_HI(net185));
 sg13g2_tiehi _2575__186 (.L_HI(net186));
 sg13g2_tiehi _2669__187 (.L_HI(net187));
 sg13g2_tiehi _2574__188 (.L_HI(net188));
 sg13g2_tiehi _2637__189 (.L_HI(net189));
 sg13g2_tiehi _2573__190 (.L_HI(net190));
 sg13g2_tiehi _2698__191 (.L_HI(net191));
 sg13g2_tiehi _2572__192 (.L_HI(net192));
 sg13g2_tiehi _2636__193 (.L_HI(net193));
 sg13g2_tiehi _2571__194 (.L_HI(net194));
 sg13g2_tiehi _2668__195 (.L_HI(net195));
 sg13g2_tiehi _2570__196 (.L_HI(net196));
 sg13g2_tiehi _2635__197 (.L_HI(net197));
 sg13g2_tiehi _2569__198 (.L_HI(net198));
 sg13g2_tiehi _2684__199 (.L_HI(net199));
 sg13g2_tiehi _2568__200 (.L_HI(net200));
 sg13g2_tiehi _2634__201 (.L_HI(net201));
 sg13g2_tiehi _2567__202 (.L_HI(net202));
 sg13g2_tiehi _2667__203 (.L_HI(net203));
 sg13g2_tiehi _2566__204 (.L_HI(net204));
 sg13g2_tiehi _2633__205 (.L_HI(net205));
 sg13g2_tiehi _2565__206 (.L_HI(net206));
 sg13g2_tiehi _2694__207 (.L_HI(net207));
 sg13g2_tiehi _2564__208 (.L_HI(net208));
 sg13g2_tiehi _2632__209 (.L_HI(net209));
 sg13g2_tiehi _2563__210 (.L_HI(net210));
 sg13g2_tiehi _2666__211 (.L_HI(net211));
 sg13g2_tiehi _2562__212 (.L_HI(net212));
 sg13g2_tiehi _2631__213 (.L_HI(net213));
 sg13g2_tiehi _2561__214 (.L_HI(net214));
 sg13g2_tiehi _2683__215 (.L_HI(net215));
 sg13g2_tiehi _2560__216 (.L_HI(net216));
 sg13g2_tiehi _2630__217 (.L_HI(net217));
 sg13g2_tiehi _2559__218 (.L_HI(net218));
 sg13g2_tiehi _2665__219 (.L_HI(net219));
 sg13g2_tiehi _2558__220 (.L_HI(net220));
 sg13g2_tiehi _2629__221 (.L_HI(net221));
 sg13g2_tiehi _2557__222 (.L_HI(net222));
 sg13g2_tiehi _2693__223 (.L_HI(net223));
 sg13g2_tiehi _2556__224 (.L_HI(net224));
 sg13g2_tiehi _2628__225 (.L_HI(net225));
 sg13g2_tiehi _2555__226 (.L_HI(net226));
 sg13g2_tiehi tt_um_arandomdev_fir_engine_top_227 (.L_HI(net227));
 sg13g2_tiehi tt_um_arandomdev_fir_engine_top_228 (.L_HI(net228));
 sg13g2_tiehi tt_um_arandomdev_fir_engine_top_229 (.L_HI(net229));
 sg13g2_tiehi tt_um_arandomdev_fir_engine_top_230 (.L_HI(net230));
 sg13g2_tiehi tt_um_arandomdev_fir_engine_top_231 (.L_HI(net231));
 sg13g2_tiehi tt_um_arandomdev_fir_engine_top_232 (.L_HI(net232));
 sg13g2_tiehi tt_um_arandomdev_fir_engine_top_233 (.L_HI(net233));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_arandomdev_fir_engine_top_6 (.L_LO(net6));
 sg13g2_tielo tt_um_arandomdev_fir_engine_top_7 (.L_LO(net7));
 sg13g2_tielo tt_um_arandomdev_fir_engine_top_8 (.L_LO(net8));
 sg13g2_tielo tt_um_arandomdev_fir_engine_top_9 (.L_LO(net9));
 sg13g2_tielo tt_um_arandomdev_fir_engine_top_10 (.L_LO(net10));
 sg13g2_tielo tt_um_arandomdev_fir_engine_top_11 (.L_LO(net11));
 sg13g2_tielo tt_um_arandomdev_fir_engine_top_12 (.L_LO(net12));
 sg13g2_tielo tt_um_arandomdev_fir_engine_top_13 (.L_LO(net13));
 sg13g2_tielo tt_um_arandomdev_fir_engine_top_14 (.L_LO(net14));
 sg13g2_tiehi _2664__15 (.L_HI(net15));
 sg13g2_buf_1 _2929_ (.A(\firEngine.i2sController.mclk ),
    .X(uio_out[0]));
 sg13g2_buf_1 _2930_ (.A(\firEngine.i2sController.lrck ),
    .X(uio_out[1]));
 sg13g2_buf_1 _2931_ (.A(\firEngine.i2sController.sclk ),
    .X(uio_out[2]));
 sg13g2_buf_1 _2932_ (.A(dac),
    .X(uio_out[3]));
 sg13g2_buf_1 _2933_ (.A(\firEngine.i2sController.mclk ),
    .X(uio_out[4]));
 sg13g2_buf_1 _2934_ (.A(\firEngine.i2sController.lrck ),
    .X(uio_out[5]));
 sg13g2_buf_1 _2935_ (.A(\firEngine.i2sController.sclk ),
    .X(uio_out[6]));
 sg13g2_buf_2 fanout448 (.A(_0765_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_0745_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(net451),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_0764_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_0744_),
    .X(net452));
 sg13g2_buf_4 fanout453 (.X(net453),
    .A(_0738_));
 sg13g2_buf_2 fanout454 (.A(_0731_),
    .X(net454));
 sg13g2_buf_1 fanout455 (.A(_0731_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(net457),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_0730_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_0724_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_0562_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_0726_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(net465),
    .X(net461));
 sg13g2_buf_1 fanout462 (.A(net465),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(net465),
    .X(net463));
 sg13g2_buf_1 fanout464 (.A(net465),
    .X(net464));
 sg13g2_buf_1 fanout465 (.A(net478),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(net467),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(net478),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(net469),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(net474),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(net472),
    .X(net470));
 sg13g2_buf_1 fanout471 (.A(net472),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(net473),
    .X(net472));
 sg13g2_buf_1 fanout473 (.A(net474),
    .X(net473));
 sg13g2_buf_1 fanout474 (.A(net478),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(net476),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(net478),
    .X(net476));
 sg13g2_buf_1 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_0679_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(net482),
    .X(net479));
 sg13g2_buf_1 fanout480 (.A(net482),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(net482),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(net490),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(net486),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(net486),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_1 fanout486 (.A(net490),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(net489),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(net489),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(net490),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_0678_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_0530_),
    .X(net491));
 sg13g2_buf_4 fanout492 (.X(net492),
    .A(_0728_));
 sg13g2_buf_2 fanout493 (.A(_0728_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(net496),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(net496),
    .X(net495));
 sg13g2_buf_1 fanout496 (.A(net499),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(net499),
    .X(net497));
 sg13g2_buf_1 fanout498 (.A(net499),
    .X(net498));
 sg13g2_buf_1 fanout499 (.A(net510),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(net501),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(net503),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(net503),
    .X(net502));
 sg13g2_buf_1 fanout503 (.A(net510),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(net505),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(net506),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(net510),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(net509),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_1 fanout510 (.A(net511),
    .X(net510));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(_0660_));
 sg13g2_buf_2 fanout512 (.A(net514),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(net514),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(net521),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(net516),
    .X(net515));
 sg13g2_buf_1 fanout516 (.A(net521),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(net521),
    .X(net517));
 sg13g2_buf_1 fanout518 (.A(net521),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(net520),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(net521),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(net528),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(net524),
    .X(net522));
 sg13g2_buf_1 fanout523 (.A(net524),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(net528),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(net526),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(net527),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_1038_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(net530),
    .X(net529));
 sg13g2_buf_4 fanout530 (.X(net530),
    .A(_0754_));
 sg13g2_buf_2 fanout531 (.A(net532),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_0752_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(net535),
    .X(net533));
 sg13g2_buf_1 fanout534 (.A(net535),
    .X(net534));
 sg13g2_buf_1 fanout535 (.A(net536),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_0752_),
    .X(net536));
 sg13g2_buf_4 fanout537 (.X(net537),
    .A(_0604_));
 sg13g2_buf_2 fanout538 (.A(net539),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(net543),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(net541),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(net542),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(net543),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(net555),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(net545),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net555),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(net547),
    .X(net546));
 sg13g2_buf_1 fanout547 (.A(net555),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net550),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(net550),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(net552),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(net555),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(\firEngine.adcDataValid ),
    .X(net555));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(\firEngine.firInst.bit_cnt[1] ));
 sg13g2_buf_2 fanout557 (.A(net718),
    .X(net557));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(\firEngine.firInst.bit_cnt[0] ));
 sg13g2_buf_2 fanout559 (.A(\firEngine.firInst.bit_cnt[0] ),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(\firEngine.firInst.sample_cnt_en ),
    .X(net560));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(net563));
 sg13g2_buf_2 fanout562 (.A(net563),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_0633_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_0633_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_0633_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(net567),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(net585),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(net570),
    .X(net568));
 sg13g2_buf_1 fanout569 (.A(net570),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(net585),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(net575),
    .X(net572));
 sg13g2_buf_1 fanout573 (.A(net575),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net575),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(net585),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(net577),
    .X(net576));
 sg13g2_buf_1 fanout577 (.A(net583),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(net583),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(net582),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(net582),
    .X(net580));
 sg13g2_buf_1 fanout581 (.A(net582),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(net583),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(net584),
    .X(net583));
 sg13g2_buf_4 fanout584 (.X(net584),
    .A(net585));
 sg13g2_buf_2 fanout585 (.A(net594),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(net587),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net588),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(net594),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(net594));
 sg13g2_buf_2 fanout591 (.A(net593),
    .X(net591));
 sg13g2_buf_1 fanout592 (.A(net593),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(net594),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(rst_n),
    .X(net594));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[7]),
    .X(net4));
 sg13g2_tielo tt_um_arandomdev_fir_engine_top_5 (.L_LO(net5));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_8 clkload3 (.A(clknet_leaf_27_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_leaf_28_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_24_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_17_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_18_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_16_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0031_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold2 (.A(\firEngine.spiSlave.csSynchronizer[0] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold3 (.A(\firEngine.spiSlave.mosiSynchronizer[0] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold4 (.A(\firEngine.spiSlave.sclkSynchronizer[0] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold5 (.A(\firEngine.i2sController.adcSynchronizer[0] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0006_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0233_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold8 (.A(\firEngine.adcData[7] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0571_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0007_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0231_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold12 (.A(\firEngine.firInst.samples[9][5] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0053_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold14 (.A(\firEngine.firInst.samples[7][6] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0195_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold16 (.A(\firEngine.firInst.samples[8][1] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0198_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold18 (.A(\firEngine.firInst.samples[7][2] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0191_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold20 (.A(\firEngine.firInst.samples[9][1] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold21 (.A(\firEngine.firInst.samples[8][3] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0200_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold23 (.A(\firEngine.firInst.samples[7][7] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0196_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold25 (.A(\firEngine.firInst.samples[8][4] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0201_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold27 (.A(\firEngine.firInst.samples[10][1] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold28 (.A(\firEngine.firInst.samples[7][0] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0189_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold30 (.A(\firEngine.firInst.samples[8][5] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0202_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold32 (.A(\firEngine.firInst.samples[9][3] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0051_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold34 (.A(\firEngine.firInst.samples[7][4] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0193_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold36 (.A(\firEngine.firInst.samples[7][1] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0190_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold38 (.A(\firEngine.firDataValid ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0081_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold40 (.A(\firEngine.firInst.samples[9][0] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0048_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0029_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0227_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold44 (.A(\firEngine.firInst.samples[7][5] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0194_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold46 (.A(\firEngine.firInst.samples[8][6] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold47 (.A(\firEngine.firInst.sample_cnt[2] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold48 (.A(_1037_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold49 (.A(\firEngine.firInst.samples[8][0] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold50 (.A(\firEngine.spiSlave.sclkSynchronizer[1] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold51 (.A(\firEngine.firInst.samples[9][2] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0058_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold53 (.A(\firEngine.firInst.samples[10][2] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold54 (.A(\firEngine.adcData[1] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0565_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold56 (.A(\firEngine.adcData[6] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0570_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold58 (.A(\firEngine.firInst.samples[7][3] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0192_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold60 (.A(\firEngine.firInst.samples[8][2] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0005_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0647_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0232_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold64 (.A(\firEngine.firInst.samples[8][7] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold65 (.A(\firEngine.firInst.samples[4][5] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0178_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold67 (.A(\firEngine.i2sController.adcQ ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0564_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold69 (.A(\firEngine.adcData[4] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0568_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold71 (.A(\firEngine.firInst.samples[9][6] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold72 (.A(\firEngine.adcData[3] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0567_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold74 (.A(\firEngine.firInst.state[1] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0000_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold76 (.A(\firEngine.firInst.samples[9][4] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0052_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold78 (.A(\firEngine.firInst.samples[10][6] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold79 (.A(\firEngine.firInst.samples[0][6] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0139_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold81 (.A(\firEngine.firInst.samples[4][6] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0179_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold83 (.A(\firEngine.firInst.samples[0][7] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0140_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold85 (.A(\firEngine.i2sController.mclkCounter[1] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0674_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0040_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0030_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0522_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0205_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold91 (.A(\firEngine.spiSlave.mosi ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0667_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0034_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold94 (.A(\firEngine.adcData[2] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold95 (.A(\firEngine.firInst.samples[9][7] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0055_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold97 (.A(\firEngine.firInst.sample_cnt[0] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0082_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold99 (.A(\firEngine.firInst.samples[5][2] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0175_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold101 (.A(_1058_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0579_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0236_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold104 (.A(\firEngine.adcData[5] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold105 (.A(\firEngine.firInst.accQ[3] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0067_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold107 (.A(\firEngine.firInst.samples[0][5] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0170_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold109 (.A(\firEngine.firInst.samples[6][0] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0181_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold111 (.A(\firEngine.firInst.samples[3][6] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold112 (.A(\firEngine.i2sController.lrckCounter[4] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0650_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0004_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold115 (.A(\firEngine.firInst.samples[6][5] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0186_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold117 (.A(\firEngine.firInst.coeffs[4][3] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0121_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold119 (.A(\firEngine.firInst.coeffs[1][5] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0099_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold121 (.A(\firEngine.firInst.coeffs[1][3] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0097_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold123 (.A(\firEngine.firInst.coeffs[5][3] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0129_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold125 (.A(\firEngine.firInst.samples[5][3] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0176_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold127 (.A(\firEngine.firInst.samples[6][3] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0184_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold129 (.A(\firEngine.firInst.coeffs[2][6] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0108_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold131 (.A(\firEngine.firInst.samples[4][4] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0177_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold133 (.A(\firEngine.firInst.accQ[0] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0064_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold135 (.A(\firEngine.firInst.samples[5][0] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0173_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold137 (.A(\firEngine.clockConfig[1] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0035_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold139 (.A(\firEngine.firInst.coeffs[3][3] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0113_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold141 (.A(\firEngine.firInst.samples[4][7] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0180_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold143 (.A(\firEngine.firInst.samples[6][6] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0187_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold145 (.A(\firEngine.i2sController.dacDataQ[3] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0213_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold147 (.A(\firEngine.i2sController.mclkCounter[3] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0677_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold149 (.A(dac),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0559_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0218_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold152 (.A(\firEngine.firInst.coeffs[3][2] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold153 (.A(\firEngine.firInst.samples[2][4] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0153_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold155 (.A(\firEngine.firInst.samples[0][4] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0169_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold157 (.A(\firEngine.firInst.samples[0][1] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0134_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold159 (.A(\firEngine.i2sController.dacDataQ[0] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0534_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0210_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold162 (.A(\firEngine.firInst.samples[1][4] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold163 (.A(\firEngine.firInst.coeffs[0][2] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0088_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold165 (.A(\firEngine.firInst.accQ[16] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold166 (.A(\firEngine.firInst.coeffs[5][2] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0128_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold168 (.A(\firEngine.firInst.samples[1][0] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0141_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold170 (.A(\firEngine.firInst.samples[2][6] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold171 (.A(\firEngine.clockConfig[2] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold172 (.A(\firEngine.firInst.samples[4][3] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0168_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold174 (.A(\firEngine.firInst.samples[1][7] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0432_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0156_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold177 (.A(\firEngine.firInst.samples[0][2] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0135_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold179 (.A(\firEngine.firInst.samples[2][7] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold180 (.A(\firEngine.firInst.samples[6][4] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0185_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold182 (.A(\firEngine.firInst.samples[6][1] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0182_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold184 (.A(\firEngine.i2sController.dacDataQ[2] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0212_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold186 (.A(\firEngine.i2sController.mclkCounter[2] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0676_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold188 (.A(\firEngine.firInst.state[2] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0658_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0003_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold191 (.A(\firEngine.i2sController.dacDataQ[5] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0215_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold193 (.A(\firEngine.firInst.samples[5][1] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0174_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold195 (.A(\firEngine.firInst.samples[3][5] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0162_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold197 (.A(\firEngine.firInst.samples[6][7] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0188_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold199 (.A(\firEngine.firInst.coeffs[1][2] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0096_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold201 (.A(\firEngine.firInst.coeffs[2][3] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0105_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold203 (.A(\firEngine.i2sController.dacDataQ[1] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0211_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold205 (.A(\firEngine.firInst.coeffs[0][0] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0086_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold207 (.A(\firEngine.i2sController.dacDataQ[4] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0214_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold209 (.A(\firEngine.firInst.samples[2][5] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0154_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold211 (.A(\firEngine.firInst.samples[1][5] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold212 (.A(\firEngine.adcData[0] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0133_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold214 (.A(\firEngine.firInst.coeffs[5][6] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0132_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold216 (.A(\firEngine.firInst.coeffs[3][6] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0116_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold218 (.A(\firEngine.firInst.coeffs[4][2] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold219 (.A(\firEngine.firInst.samples[3][2] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0167_),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold221 (.A(\firEngine.firInst.samples[3][7] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold222 (.A(\firEngine.firInst.samples[2][2] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0151_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold224 (.A(\firEngine.firInst.samples[1][1] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0414_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0150_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold227 (.A(\firEngine.firInst.samples[3][4] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold228 (.A(\firEngine.firInst.sample_cnt[1] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold229 (.A(_1033_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold230 (.A(\firEngine.firInst.samples[4][2] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold231 (.A(\firEngine.i2sController.dacDataQ[6] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0216_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold233 (.A(\firEngine.firInst.samples[2][1] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold234 (.A(\firEngine.firInst.samples[6][2] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold235 (.A(\firEngine.firInst.coeffs[0][3] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0089_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold237 (.A(\firEngine.firInst.coeffs[2][5] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold238 (.A(\firEngine.firInst.samples[3][0] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0157_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold240 (.A(\firEngine.firInst.coeffs[4][4] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0122_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold242 (.A(\firEngine.firInst.samples[2][3] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0152_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold244 (.A(\firEngine.clockConfig[3] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0038_),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold246 (.A(\firEngine.firInst.accQ[6] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold247 (.A(\firEngine.firInst.coeffs[1][4] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold248 (.A(\firEngine.firInst.samples[3][3] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold249 (.A(\firEngine.firInst.samples[2][0] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold250 (.A(\firEngine.firInst.samples[1][6] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold251 (.A(\firEngine.firInst.coeffs[5][7] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0336_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0124_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold254 (.A(\firEngine.firInst.coeffs[3][1] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold255 (.A(\firEngine.firInst.samples[1][2] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold256 (.A(\firEngine.firInst.samples[1][3] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0144_),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold258 (.A(\firEngine.firInst.coeffs[0][6] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0092_),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold260 (.A(\firEngine.firInst.coeffs[5][1] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold261 (.A(\firEngine.firInst.samples[0][3] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold262 (.A(\firEngine.firInst.accQ[14] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold263 (.A(\firEngine.firInst.coeffs[0][1] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold264 (.A(\firEngine.firInst.coeffs[3][5] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0115_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold266 (.A(\firEngine.firInst.accQ[4] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold267 (.A(\firEngine.firInst.coeffs[4][1] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold268 (.A(\firEngine.firInst.samples[0][0] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0165_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold270 (.A(\firEngine.firInst.coeffs[0][5] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0091_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold272 (.A(\firEngine.firInst.coeffs[1][6] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0100_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold274 (.A(\firEngine.firInst.coeffs[2][4] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold275 (.A(\firEngine.firInst.accQ[5] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0843_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold277 (.A(\firEngine.firInst.coeffs[2][2] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold278 (.A(\firEngine.firInst.accQ[1] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0065_),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold280 (.A(\firEngine.spiSlave.cs ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0659_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold282 (.A(\firEngine.firInst.coeffs[1][0] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0094_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold284 (.A(\firEngine.i2sController.currentState[2] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0663_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold286 (.A(\firEngine.firInst.samples[3][1] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0158_),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold288 (.A(\firEngine.firInst.coeffs[4][7] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0125_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold290 (.A(\firEngine.firInst.samples[4][1] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold291 (.A(\firEngine.firInst.accQ[2] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold292 (.A(\firEngine.firInst.accQ[15] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0079_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold294 (.A(\firEngine.firInst.coeffs[2][7] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0109_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold296 (.A(\firEngine.firInst.coeffs[0][4] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold297 (.A(\firEngine.firInst.coeffs[5][0] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold298 (.A(\firEngine.i2sController.currentState[1] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0664_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold300 (.A(\firEngine.firInst.coeffs[3][0] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0267_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0101_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold303 (.A(\firEngine.firInst.sample_cnt_en ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0665_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0001_),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold306 (.A(\firEngine.firInst.coeffs[3][7] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0117_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold308 (.A(\firEngine.firInst.coeffs[3][4] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0114_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold310 (.A(\firEngine.firInst.coeffs[4][5] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0123_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold312 (.A(\firEngine.firInst.coeffs[5][5] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold313 (.A(\firEngine.firInst.coeffs[2][1] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold314 (.A(\firEngine.firInst.accQ[12] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0021_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0549_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold317 (.A(\firEngine.firInst.accQ[11] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold318 (.A(\firEngine.firInst.coeffs[1][1] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold319 (.A(\firEngine.firInst.coeffs[2][0] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold320 (.A(\firEngine.firInst.state[0] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0657_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold322 (.A(\firEngine.firInst.coeffs[5][4] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold323 (.A(\firEngine.firInst.accQ[9] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold324 (.A(\firEngine.firInst.accQ[7] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold325 (.A(\firEngine.i2sController.lrckCounter[3] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold326 (.A(\firEngine.firInst.coeffs[4][0] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold327 (.A(\firEngine.firInst.coeffs[0][7] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold328 (.A(\firEngine.i2sController.lrckCounter[1] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0524_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0206_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold331 (.A(\firEngine.configStore.serialOut ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold332 (.A(\firEngine.firInst.accQ[10] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold333 (.A(\firEngine.firInst.accQ[8] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold334 (.A(\firEngine.firInst.accQ[13] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold335 (.A(\firEngine.i2sController.lrckCounter[2] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold336 (.A(\firEngine.i2sController.currentState[0] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0010_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold338 (.A(\firEngine.firInst.bit_cnt[1] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold339 (.A(\firEngine.i2sController.currentState[2] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold340 (.A(\firEngine.spiSlave.cs ),
    .X(net720));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(rst_n));
 sg13g2_antennanp ANTENNA_4 (.A(rst_n));
 sg13g2_antennanp ANTENNA_5 (.A(rst_n));
 sg13g2_antennanp ANTENNA_6 (.A(rst_n));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_4 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_310 ();
 sg13g2_decap_8 FILLER_3_317 ();
 sg13g2_decap_8 FILLER_3_324 ();
 sg13g2_decap_8 FILLER_3_331 ();
 sg13g2_decap_8 FILLER_3_338 ();
 sg13g2_decap_8 FILLER_3_345 ();
 sg13g2_decap_8 FILLER_3_352 ();
 sg13g2_decap_8 FILLER_3_359 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_decap_8 FILLER_3_373 ();
 sg13g2_decap_8 FILLER_3_380 ();
 sg13g2_decap_8 FILLER_3_387 ();
 sg13g2_decap_8 FILLER_3_394 ();
 sg13g2_decap_8 FILLER_3_401 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_fill_2 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_decap_8 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_338 ();
 sg13g2_decap_8 FILLER_4_345 ();
 sg13g2_decap_8 FILLER_4_352 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_4 FILLER_5_259 ();
 sg13g2_fill_1 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_268 ();
 sg13g2_decap_8 FILLER_5_275 ();
 sg13g2_fill_2 FILLER_5_282 ();
 sg13g2_fill_1 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_fill_1 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_346 ();
 sg13g2_decap_8 FILLER_6_353 ();
 sg13g2_decap_8 FILLER_6_360 ();
 sg13g2_decap_8 FILLER_6_367 ();
 sg13g2_decap_8 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_381 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_decap_8 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_fill_2 FILLER_7_276 ();
 sg13g2_fill_1 FILLER_7_278 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_fill_2 FILLER_8_252 ();
 sg13g2_fill_1 FILLER_8_254 ();
 sg13g2_fill_2 FILLER_8_279 ();
 sg13g2_fill_1 FILLER_8_300 ();
 sg13g2_fill_2 FILLER_8_324 ();
 sg13g2_decap_8 FILLER_8_352 ();
 sg13g2_decap_8 FILLER_8_359 ();
 sg13g2_decap_8 FILLER_8_366 ();
 sg13g2_decap_8 FILLER_8_373 ();
 sg13g2_decap_8 FILLER_8_380 ();
 sg13g2_decap_8 FILLER_8_387 ();
 sg13g2_decap_8 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_4 FILLER_9_231 ();
 sg13g2_fill_2 FILLER_9_235 ();
 sg13g2_decap_4 FILLER_9_277 ();
 sg13g2_fill_1 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_fill_2 FILLER_10_245 ();
 sg13g2_fill_1 FILLER_10_247 ();
 sg13g2_decap_4 FILLER_10_252 ();
 sg13g2_fill_2 FILLER_10_256 ();
 sg13g2_decap_4 FILLER_10_268 ();
 sg13g2_fill_2 FILLER_10_272 ();
 sg13g2_fill_2 FILLER_10_338 ();
 sg13g2_fill_1 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_fill_2 FILLER_11_245 ();
 sg13g2_fill_1 FILLER_11_247 ();
 sg13g2_decap_4 FILLER_11_279 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_4 FILLER_12_231 ();
 sg13g2_fill_2 FILLER_12_235 ();
 sg13g2_fill_1 FILLER_12_277 ();
 sg13g2_fill_1 FILLER_12_321 ();
 sg13g2_fill_2 FILLER_12_327 ();
 sg13g2_fill_1 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_370 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_4 FILLER_13_238 ();
 sg13g2_fill_1 FILLER_13_242 ();
 sg13g2_fill_2 FILLER_13_256 ();
 sg13g2_fill_1 FILLER_13_258 ();
 sg13g2_fill_2 FILLER_13_279 ();
 sg13g2_fill_1 FILLER_13_281 ();
 sg13g2_fill_1 FILLER_13_313 ();
 sg13g2_fill_2 FILLER_13_348 ();
 sg13g2_fill_1 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_372 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_4 FILLER_14_262 ();
 sg13g2_fill_1 FILLER_14_266 ();
 sg13g2_fill_1 FILLER_14_287 ();
 sg13g2_fill_2 FILLER_14_329 ();
 sg13g2_fill_1 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_fill_2 FILLER_15_210 ();
 sg13g2_fill_1 FILLER_15_212 ();
 sg13g2_fill_2 FILLER_15_220 ();
 sg13g2_fill_2 FILLER_15_231 ();
 sg13g2_fill_1 FILLER_15_233 ();
 sg13g2_decap_4 FILLER_15_260 ();
 sg13g2_fill_1 FILLER_15_264 ();
 sg13g2_decap_4 FILLER_15_280 ();
 sg13g2_decap_4 FILLER_15_302 ();
 sg13g2_fill_2 FILLER_15_306 ();
 sg13g2_fill_2 FILLER_15_326 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_4 FILLER_16_196 ();
 sg13g2_fill_2 FILLER_16_200 ();
 sg13g2_fill_1 FILLER_16_233 ();
 sg13g2_fill_2 FILLER_16_323 ();
 sg13g2_fill_1 FILLER_16_334 ();
 sg13g2_fill_2 FILLER_16_340 ();
 sg13g2_fill_1 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_4 FILLER_17_147 ();
 sg13g2_fill_2 FILLER_17_151 ();
 sg13g2_decap_8 FILLER_17_160 ();
 sg13g2_decap_4 FILLER_17_167 ();
 sg13g2_fill_1 FILLER_17_171 ();
 sg13g2_decap_4 FILLER_17_176 ();
 sg13g2_fill_1 FILLER_17_180 ();
 sg13g2_fill_2 FILLER_17_252 ();
 sg13g2_decap_4 FILLER_17_274 ();
 sg13g2_fill_1 FILLER_17_305 ();
 sg13g2_fill_2 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_327 ();
 sg13g2_fill_2 FILLER_17_334 ();
 sg13g2_fill_1 FILLER_17_336 ();
 sg13g2_decap_4 FILLER_17_361 ();
 sg13g2_fill_1 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_4 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_137 ();
 sg13g2_decap_4 FILLER_18_142 ();
 sg13g2_fill_1 FILLER_18_146 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_fill_2 FILLER_18_172 ();
 sg13g2_fill_1 FILLER_18_200 ();
 sg13g2_fill_2 FILLER_18_235 ();
 sg13g2_fill_2 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_265 ();
 sg13g2_fill_2 FILLER_18_286 ();
 sg13g2_fill_1 FILLER_18_288 ();
 sg13g2_fill_1 FILLER_18_322 ();
 sg13g2_fill_1 FILLER_18_328 ();
 sg13g2_fill_1 FILLER_18_344 ();
 sg13g2_decap_8 FILLER_18_370 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_4 FILLER_19_105 ();
 sg13g2_fill_2 FILLER_19_109 ();
 sg13g2_fill_2 FILLER_19_241 ();
 sg13g2_fill_2 FILLER_19_256 ();
 sg13g2_fill_1 FILLER_19_258 ();
 sg13g2_fill_2 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_270 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_fill_2 FILLER_20_112 ();
 sg13g2_fill_2 FILLER_20_154 ();
 sg13g2_fill_2 FILLER_20_230 ();
 sg13g2_fill_1 FILLER_20_232 ();
 sg13g2_decap_8 FILLER_20_236 ();
 sg13g2_decap_8 FILLER_20_243 ();
 sg13g2_fill_2 FILLER_20_250 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_fill_2 FILLER_20_272 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_4 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_fill_2 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_220 ();
 sg13g2_fill_2 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_317 ();
 sg13g2_fill_2 FILLER_21_356 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_fill_1 FILLER_22_105 ();
 sg13g2_fill_2 FILLER_22_176 ();
 sg13g2_fill_1 FILLER_22_311 ();
 sg13g2_fill_2 FILLER_22_351 ();
 sg13g2_fill_2 FILLER_22_367 ();
 sg13g2_fill_1 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_122 ();
 sg13g2_fill_1 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_197 ();
 sg13g2_fill_1 FILLER_23_260 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_312 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_fill_1 FILLER_23_358 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_119 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_1 FILLER_24_129 ();
 sg13g2_fill_2 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_208 ();
 sg13g2_fill_1 FILLER_24_214 ();
 sg13g2_fill_2 FILLER_24_260 ();
 sg13g2_fill_1 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_fill_1 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_4 FILLER_25_84 ();
 sg13g2_fill_1 FILLER_25_88 ();
 sg13g2_decap_8 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_162 ();
 sg13g2_fill_2 FILLER_25_171 ();
 sg13g2_fill_1 FILLER_25_186 ();
 sg13g2_fill_2 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_204 ();
 sg13g2_decap_4 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_229 ();
 sg13g2_fill_2 FILLER_25_308 ();
 sg13g2_fill_2 FILLER_25_356 ();
 sg13g2_fill_1 FILLER_25_358 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_fill_1 FILLER_26_165 ();
 sg13g2_fill_2 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_225 ();
 sg13g2_fill_1 FILLER_26_227 ();
 sg13g2_fill_2 FILLER_26_254 ();
 sg13g2_fill_1 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_318 ();
 sg13g2_decap_8 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_4 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_126 ();
 sg13g2_fill_2 FILLER_27_142 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_fill_2 FILLER_28_84 ();
 sg13g2_fill_1 FILLER_28_86 ();
 sg13g2_fill_2 FILLER_28_126 ();
 sg13g2_fill_2 FILLER_28_143 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_decap_4 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_172 ();
 sg13g2_fill_2 FILLER_28_200 ();
 sg13g2_fill_1 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_decap_4 FILLER_28_254 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_fill_2 FILLER_28_320 ();
 sg13g2_fill_2 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_348 ();
 sg13g2_decap_8 FILLER_28_372 ();
 sg13g2_decap_8 FILLER_28_379 ();
 sg13g2_decap_8 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_fill_1 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_115 ();
 sg13g2_fill_1 FILLER_29_117 ();
 sg13g2_fill_1 FILLER_29_131 ();
 sg13g2_fill_2 FILLER_29_160 ();
 sg13g2_decap_4 FILLER_29_167 ();
 sg13g2_fill_2 FILLER_29_171 ();
 sg13g2_fill_2 FILLER_29_195 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_fill_1 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_214 ();
 sg13g2_fill_2 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_226 ();
 sg13g2_decap_8 FILLER_29_249 ();
 sg13g2_decap_4 FILLER_29_256 ();
 sg13g2_fill_2 FILLER_29_260 ();
 sg13g2_decap_4 FILLER_29_267 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_fill_1 FILLER_29_296 ();
 sg13g2_fill_2 FILLER_29_328 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_fill_2 FILLER_29_345 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_4 FILLER_30_84 ();
 sg13g2_fill_1 FILLER_30_88 ();
 sg13g2_fill_1 FILLER_30_172 ();
 sg13g2_decap_4 FILLER_30_183 ();
 sg13g2_fill_1 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_312 ();
 sg13g2_fill_2 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_320 ();
 sg13g2_decap_8 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_4 FILLER_31_126 ();
 sg13g2_fill_2 FILLER_31_209 ();
 sg13g2_fill_2 FILLER_31_251 ();
 sg13g2_decap_4 FILLER_31_284 ();
 sg13g2_decap_4 FILLER_31_309 ();
 sg13g2_fill_2 FILLER_31_316 ();
 sg13g2_fill_1 FILLER_31_318 ();
 sg13g2_fill_2 FILLER_31_344 ();
 sg13g2_decap_8 FILLER_31_374 ();
 sg13g2_decap_8 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_4 FILLER_32_84 ();
 sg13g2_fill_1 FILLER_32_114 ();
 sg13g2_fill_1 FILLER_32_138 ();
 sg13g2_fill_1 FILLER_32_179 ();
 sg13g2_decap_4 FILLER_32_216 ();
 sg13g2_fill_1 FILLER_32_225 ();
 sg13g2_fill_2 FILLER_32_252 ();
 sg13g2_fill_1 FILLER_32_254 ();
 sg13g2_decap_4 FILLER_32_276 ();
 sg13g2_fill_2 FILLER_32_280 ();
 sg13g2_decap_4 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_91 ();
 sg13g2_decap_4 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_191 ();
 sg13g2_fill_2 FILLER_33_201 ();
 sg13g2_fill_1 FILLER_33_213 ();
 sg13g2_fill_2 FILLER_33_224 ();
 sg13g2_decap_4 FILLER_33_230 ();
 sg13g2_decap_8 FILLER_33_247 ();
 sg13g2_decap_8 FILLER_33_254 ();
 sg13g2_decap_8 FILLER_33_261 ();
 sg13g2_fill_2 FILLER_33_268 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_decap_4 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_4 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_95 ();
 sg13g2_decap_4 FILLER_34_149 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_4 FILLER_34_172 ();
 sg13g2_decap_8 FILLER_34_181 ();
 sg13g2_decap_8 FILLER_34_207 ();
 sg13g2_decap_4 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_218 ();
 sg13g2_decap_4 FILLER_34_224 ();
 sg13g2_fill_1 FILLER_34_228 ();
 sg13g2_fill_2 FILLER_34_237 ();
 sg13g2_fill_1 FILLER_34_239 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_252 ();
 sg13g2_fill_1 FILLER_34_254 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_4 FILLER_34_297 ();
 sg13g2_fill_1 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_338 ();
 sg13g2_decap_8 FILLER_34_348 ();
 sg13g2_decap_8 FILLER_34_355 ();
 sg13g2_decap_8 FILLER_34_362 ();
 sg13g2_decap_8 FILLER_34_369 ();
 sg13g2_decap_8 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_34_383 ();
 sg13g2_decap_8 FILLER_34_390 ();
 sg13g2_decap_8 FILLER_34_397 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_4 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_132 ();
 sg13g2_fill_1 FILLER_35_134 ();
 sg13g2_fill_2 FILLER_35_150 ();
 sg13g2_fill_2 FILLER_35_188 ();
 sg13g2_fill_1 FILLER_35_190 ();
 sg13g2_fill_1 FILLER_35_210 ();
 sg13g2_fill_2 FILLER_35_231 ();
 sg13g2_fill_1 FILLER_35_233 ();
 sg13g2_fill_2 FILLER_35_278 ();
 sg13g2_fill_2 FILLER_35_298 ();
 sg13g2_fill_1 FILLER_35_300 ();
 sg13g2_fill_2 FILLER_35_321 ();
 sg13g2_decap_8 FILLER_35_327 ();
 sg13g2_decap_8 FILLER_35_334 ();
 sg13g2_decap_8 FILLER_35_341 ();
 sg13g2_decap_4 FILLER_35_348 ();
 sg13g2_decap_8 FILLER_35_370 ();
 sg13g2_decap_8 FILLER_35_377 ();
 sg13g2_decap_8 FILLER_35_384 ();
 sg13g2_decap_8 FILLER_35_391 ();
 sg13g2_decap_8 FILLER_35_398 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_117 ();
 sg13g2_decap_4 FILLER_36_185 ();
 sg13g2_fill_2 FILLER_36_241 ();
 sg13g2_fill_1 FILLER_36_243 ();
 sg13g2_fill_2 FILLER_36_252 ();
 sg13g2_fill_1 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_283 ();
 sg13g2_decap_8 FILLER_36_295 ();
 sg13g2_decap_8 FILLER_36_302 ();
 sg13g2_decap_8 FILLER_36_318 ();
 sg13g2_decap_8 FILLER_36_325 ();
 sg13g2_decap_8 FILLER_36_332 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_1 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_377 ();
 sg13g2_decap_8 FILLER_36_384 ();
 sg13g2_decap_8 FILLER_36_391 ();
 sg13g2_decap_8 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_4 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_207 ();
 sg13g2_decap_4 FILLER_37_253 ();
 sg13g2_fill_2 FILLER_37_266 ();
 sg13g2_fill_1 FILLER_37_268 ();
 sg13g2_decap_4 FILLER_37_288 ();
 sg13g2_fill_1 FILLER_37_306 ();
 sg13g2_fill_2 FILLER_37_317 ();
 sg13g2_decap_8 FILLER_37_327 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_fill_1 FILLER_38_98 ();
 sg13g2_fill_2 FILLER_38_193 ();
 sg13g2_fill_2 FILLER_38_241 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_fill_2 FILLER_38_254 ();
 sg13g2_fill_2 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_305 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_1 FILLER_38_334 ();
 sg13g2_fill_1 FILLER_38_340 ();
 sg13g2_fill_2 FILLER_38_350 ();
 sg13g2_fill_1 FILLER_38_352 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_fill_1 FILLER_39_98 ();
 sg13g2_fill_1 FILLER_39_112 ();
 sg13g2_fill_1 FILLER_39_182 ();
 sg13g2_decap_4 FILLER_39_214 ();
 sg13g2_fill_2 FILLER_39_218 ();
 sg13g2_fill_2 FILLER_39_239 ();
 sg13g2_fill_1 FILLER_39_241 ();
 sg13g2_decap_4 FILLER_39_245 ();
 sg13g2_fill_1 FILLER_39_342 ();
 sg13g2_decap_8 FILLER_39_365 ();
 sg13g2_decap_8 FILLER_39_372 ();
 sg13g2_decap_8 FILLER_39_379 ();
 sg13g2_decap_8 FILLER_39_386 ();
 sg13g2_decap_8 FILLER_39_393 ();
 sg13g2_decap_8 FILLER_39_400 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_fill_2 FILLER_40_91 ();
 sg13g2_fill_2 FILLER_40_119 ();
 sg13g2_fill_2 FILLER_40_143 ();
 sg13g2_fill_1 FILLER_40_169 ();
 sg13g2_decap_8 FILLER_40_190 ();
 sg13g2_decap_4 FILLER_40_206 ();
 sg13g2_fill_1 FILLER_40_210 ();
 sg13g2_fill_2 FILLER_40_219 ();
 sg13g2_decap_4 FILLER_40_224 ();
 sg13g2_fill_2 FILLER_40_237 ();
 sg13g2_fill_2 FILLER_40_271 ();
 sg13g2_fill_1 FILLER_40_273 ();
 sg13g2_fill_1 FILLER_40_284 ();
 sg13g2_fill_2 FILLER_40_327 ();
 sg13g2_fill_2 FILLER_40_358 ();
 sg13g2_fill_1 FILLER_40_360 ();
 sg13g2_decap_8 FILLER_40_373 ();
 sg13g2_decap_8 FILLER_40_380 ();
 sg13g2_decap_8 FILLER_40_387 ();
 sg13g2_decap_8 FILLER_40_394 ();
 sg13g2_decap_8 FILLER_40_401 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_fill_2 FILLER_41_98 ();
 sg13g2_fill_1 FILLER_41_100 ();
 sg13g2_fill_2 FILLER_41_129 ();
 sg13g2_fill_1 FILLER_41_131 ();
 sg13g2_fill_1 FILLER_41_146 ();
 sg13g2_decap_4 FILLER_41_178 ();
 sg13g2_fill_1 FILLER_41_201 ();
 sg13g2_fill_2 FILLER_41_228 ();
 sg13g2_fill_1 FILLER_41_238 ();
 sg13g2_fill_2 FILLER_41_287 ();
 sg13g2_fill_2 FILLER_41_294 ();
 sg13g2_fill_1 FILLER_41_296 ();
 sg13g2_fill_2 FILLER_41_327 ();
 sg13g2_decap_4 FILLER_41_347 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_fill_2 FILLER_42_91 ();
 sg13g2_fill_2 FILLER_42_119 ();
 sg13g2_fill_2 FILLER_42_161 ();
 sg13g2_fill_2 FILLER_42_167 ();
 sg13g2_decap_8 FILLER_42_199 ();
 sg13g2_fill_2 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_254 ();
 sg13g2_fill_2 FILLER_42_261 ();
 sg13g2_decap_8 FILLER_42_271 ();
 sg13g2_fill_1 FILLER_42_278 ();
 sg13g2_fill_2 FILLER_42_283 ();
 sg13g2_decap_8 FILLER_42_289 ();
 sg13g2_decap_8 FILLER_42_296 ();
 sg13g2_decap_4 FILLER_42_303 ();
 sg13g2_decap_4 FILLER_42_315 ();
 sg13g2_fill_1 FILLER_42_319 ();
 sg13g2_decap_4 FILLER_42_339 ();
 sg13g2_fill_2 FILLER_42_351 ();
 sg13g2_fill_1 FILLER_42_353 ();
 sg13g2_fill_2 FILLER_42_373 ();
 sg13g2_fill_1 FILLER_42_375 ();
 sg13g2_decap_8 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_fill_2 FILLER_43_91 ();
 sg13g2_fill_1 FILLER_43_93 ();
 sg13g2_fill_1 FILLER_43_113 ();
 sg13g2_decap_8 FILLER_43_159 ();
 sg13g2_decap_8 FILLER_43_166 ();
 sg13g2_decap_4 FILLER_43_191 ();
 sg13g2_fill_1 FILLER_43_195 ();
 sg13g2_fill_1 FILLER_43_209 ();
 sg13g2_fill_2 FILLER_43_220 ();
 sg13g2_fill_1 FILLER_43_235 ();
 sg13g2_fill_2 FILLER_43_258 ();
 sg13g2_fill_2 FILLER_43_276 ();
 sg13g2_fill_1 FILLER_43_278 ();
 sg13g2_decap_8 FILLER_43_293 ();
 sg13g2_decap_4 FILLER_43_304 ();
 sg13g2_fill_1 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_313 ();
 sg13g2_decap_8 FILLER_43_320 ();
 sg13g2_fill_1 FILLER_43_327 ();
 sg13g2_fill_1 FILLER_43_333 ();
 sg13g2_decap_8 FILLER_43_358 ();
 sg13g2_decap_8 FILLER_43_365 ();
 sg13g2_fill_1 FILLER_43_372 ();
 sg13g2_decap_8 FILLER_43_377 ();
 sg13g2_decap_8 FILLER_43_384 ();
 sg13g2_decap_8 FILLER_43_391 ();
 sg13g2_decap_8 FILLER_43_398 ();
 sg13g2_decap_4 FILLER_43_405 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_fill_2 FILLER_44_91 ();
 sg13g2_fill_1 FILLER_44_93 ();
 sg13g2_fill_2 FILLER_44_141 ();
 sg13g2_fill_2 FILLER_44_161 ();
 sg13g2_fill_2 FILLER_44_184 ();
 sg13g2_fill_1 FILLER_44_186 ();
 sg13g2_decap_4 FILLER_44_200 ();
 sg13g2_fill_1 FILLER_44_204 ();
 sg13g2_fill_1 FILLER_44_219 ();
 sg13g2_fill_2 FILLER_44_225 ();
 sg13g2_fill_1 FILLER_44_227 ();
 sg13g2_fill_1 FILLER_44_256 ();
 sg13g2_decap_8 FILLER_44_327 ();
 sg13g2_decap_8 FILLER_44_334 ();
 sg13g2_fill_2 FILLER_44_341 ();
 sg13g2_fill_1 FILLER_44_343 ();
 sg13g2_decap_8 FILLER_44_369 ();
 sg13g2_decap_8 FILLER_44_376 ();
 sg13g2_decap_8 FILLER_44_383 ();
 sg13g2_decap_8 FILLER_44_390 ();
 sg13g2_decap_8 FILLER_44_397 ();
 sg13g2_decap_4 FILLER_44_404 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_4 FILLER_45_98 ();
 sg13g2_decap_4 FILLER_45_115 ();
 sg13g2_fill_2 FILLER_45_208 ();
 sg13g2_fill_1 FILLER_45_210 ();
 sg13g2_fill_2 FILLER_45_215 ();
 sg13g2_fill_2 FILLER_45_273 ();
 sg13g2_fill_1 FILLER_45_275 ();
 sg13g2_fill_1 FILLER_45_284 ();
 sg13g2_decap_8 FILLER_45_290 ();
 sg13g2_decap_4 FILLER_45_297 ();
 sg13g2_fill_2 FILLER_45_305 ();
 sg13g2_fill_2 FILLER_45_315 ();
 sg13g2_fill_2 FILLER_45_322 ();
 sg13g2_fill_1 FILLER_45_330 ();
 sg13g2_fill_2 FILLER_45_346 ();
 sg13g2_decap_8 FILLER_45_387 ();
 sg13g2_decap_8 FILLER_45_394 ();
 sg13g2_decap_8 FILLER_45_401 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_fill_2 FILLER_46_91 ();
 sg13g2_fill_1 FILLER_46_93 ();
 sg13g2_fill_1 FILLER_46_130 ();
 sg13g2_fill_2 FILLER_46_136 ();
 sg13g2_fill_1 FILLER_46_138 ();
 sg13g2_fill_2 FILLER_46_198 ();
 sg13g2_fill_2 FILLER_46_226 ();
 sg13g2_decap_4 FILLER_46_238 ();
 sg13g2_fill_1 FILLER_46_242 ();
 sg13g2_fill_2 FILLER_46_272 ();
 sg13g2_decap_4 FILLER_46_292 ();
 sg13g2_fill_1 FILLER_46_296 ();
 sg13g2_decap_4 FILLER_46_304 ();
 sg13g2_fill_2 FILLER_46_308 ();
 sg13g2_fill_1 FILLER_46_339 ();
 sg13g2_fill_2 FILLER_46_348 ();
 sg13g2_fill_1 FILLER_46_350 ();
 sg13g2_fill_2 FILLER_46_359 ();
 sg13g2_fill_1 FILLER_46_361 ();
 sg13g2_fill_1 FILLER_46_376 ();
 sg13g2_decap_8 FILLER_46_386 ();
 sg13g2_decap_8 FILLER_46_393 ();
 sg13g2_decap_8 FILLER_46_400 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_fill_2 FILLER_47_91 ();
 sg13g2_fill_2 FILLER_47_124 ();
 sg13g2_fill_1 FILLER_47_214 ();
 sg13g2_decap_8 FILLER_47_241 ();
 sg13g2_decap_4 FILLER_47_248 ();
 sg13g2_decap_8 FILLER_47_261 ();
 sg13g2_decap_8 FILLER_47_268 ();
 sg13g2_decap_8 FILLER_47_275 ();
 sg13g2_decap_4 FILLER_47_282 ();
 sg13g2_fill_1 FILLER_47_286 ();
 sg13g2_fill_1 FILLER_47_295 ();
 sg13g2_fill_1 FILLER_47_310 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_fill_2 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_fill_2 FILLER_47_406 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_4 FILLER_48_98 ();
 sg13g2_decap_4 FILLER_48_111 ();
 sg13g2_fill_2 FILLER_48_130 ();
 sg13g2_fill_1 FILLER_48_142 ();
 sg13g2_decap_4 FILLER_48_166 ();
 sg13g2_fill_1 FILLER_48_170 ();
 sg13g2_fill_2 FILLER_48_180 ();
 sg13g2_fill_1 FILLER_48_197 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_fill_2 FILLER_48_217 ();
 sg13g2_fill_1 FILLER_48_219 ();
 sg13g2_fill_2 FILLER_48_225 ();
 sg13g2_decap_8 FILLER_48_234 ();
 sg13g2_fill_2 FILLER_48_241 ();
 sg13g2_fill_1 FILLER_48_243 ();
 sg13g2_fill_2 FILLER_48_257 ();
 sg13g2_fill_2 FILLER_48_280 ();
 sg13g2_fill_2 FILLER_48_287 ();
 sg13g2_fill_1 FILLER_48_289 ();
 sg13g2_fill_2 FILLER_48_310 ();
 sg13g2_fill_1 FILLER_48_312 ();
 sg13g2_fill_2 FILLER_48_317 ();
 sg13g2_decap_4 FILLER_48_343 ();
 sg13g2_fill_1 FILLER_48_347 ();
 sg13g2_decap_8 FILLER_48_373 ();
 sg13g2_decap_8 FILLER_48_380 ();
 sg13g2_decap_8 FILLER_48_387 ();
 sg13g2_decap_8 FILLER_48_394 ();
 sg13g2_decap_8 FILLER_48_401 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_179 ();
 sg13g2_decap_8 FILLER_49_195 ();
 sg13g2_fill_2 FILLER_49_202 ();
 sg13g2_fill_1 FILLER_49_204 ();
 sg13g2_fill_2 FILLER_49_213 ();
 sg13g2_fill_1 FILLER_49_289 ();
 sg13g2_fill_1 FILLER_49_313 ();
 sg13g2_decap_4 FILLER_49_345 ();
 sg13g2_decap_8 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_decap_4 FILLER_49_403 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_fill_2 FILLER_50_91 ();
 sg13g2_fill_2 FILLER_50_119 ();
 sg13g2_fill_2 FILLER_50_148 ();
 sg13g2_fill_1 FILLER_50_181 ();
 sg13g2_fill_2 FILLER_50_291 ();
 sg13g2_fill_2 FILLER_50_305 ();
 sg13g2_fill_1 FILLER_50_307 ();
 sg13g2_fill_2 FILLER_50_316 ();
 sg13g2_decap_8 FILLER_50_340 ();
 sg13g2_decap_8 FILLER_50_347 ();
 sg13g2_decap_8 FILLER_50_354 ();
 sg13g2_decap_4 FILLER_50_361 ();
 sg13g2_decap_8 FILLER_50_369 ();
 sg13g2_decap_8 FILLER_50_376 ();
 sg13g2_decap_8 FILLER_50_383 ();
 sg13g2_decap_8 FILLER_50_390 ();
 sg13g2_decap_8 FILLER_50_397 ();
 sg13g2_decap_4 FILLER_50_404 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_4 FILLER_51_91 ();
 sg13g2_fill_1 FILLER_51_95 ();
 sg13g2_fill_2 FILLER_51_150 ();
 sg13g2_fill_1 FILLER_51_152 ();
 sg13g2_fill_1 FILLER_51_167 ();
 sg13g2_fill_1 FILLER_51_182 ();
 sg13g2_fill_2 FILLER_51_240 ();
 sg13g2_fill_1 FILLER_51_242 ();
 sg13g2_fill_2 FILLER_51_248 ();
 sg13g2_fill_2 FILLER_51_270 ();
 sg13g2_fill_1 FILLER_51_272 ();
 sg13g2_fill_1 FILLER_51_310 ();
 sg13g2_fill_2 FILLER_51_334 ();
 sg13g2_fill_1 FILLER_51_345 ();
 sg13g2_decap_8 FILLER_51_361 ();
 sg13g2_decap_8 FILLER_51_368 ();
 sg13g2_decap_8 FILLER_51_375 ();
 sg13g2_decap_8 FILLER_51_382 ();
 sg13g2_decap_8 FILLER_51_389 ();
 sg13g2_decap_8 FILLER_51_396 ();
 sg13g2_decap_4 FILLER_51_403 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_fill_2 FILLER_52_112 ();
 sg13g2_fill_2 FILLER_52_133 ();
 sg13g2_fill_1 FILLER_52_135 ();
 sg13g2_fill_2 FILLER_52_172 ();
 sg13g2_fill_1 FILLER_52_184 ();
 sg13g2_fill_2 FILLER_52_216 ();
 sg13g2_fill_1 FILLER_52_218 ();
 sg13g2_fill_1 FILLER_52_228 ();
 sg13g2_fill_1 FILLER_52_242 ();
 sg13g2_fill_2 FILLER_52_252 ();
 sg13g2_fill_1 FILLER_52_254 ();
 sg13g2_fill_1 FILLER_52_278 ();
 sg13g2_decap_4 FILLER_52_288 ();
 sg13g2_fill_2 FILLER_52_292 ();
 sg13g2_fill_2 FILLER_52_301 ();
 sg13g2_fill_1 FILLER_52_308 ();
 sg13g2_fill_2 FILLER_52_333 ();
 sg13g2_fill_1 FILLER_52_335 ();
 sg13g2_fill_1 FILLER_52_352 ();
 sg13g2_decap_8 FILLER_52_381 ();
 sg13g2_decap_8 FILLER_52_388 ();
 sg13g2_decap_8 FILLER_52_395 ();
 sg13g2_decap_8 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_fill_1 FILLER_53_139 ();
 sg13g2_fill_1 FILLER_53_195 ();
 sg13g2_fill_1 FILLER_53_205 ();
 sg13g2_fill_2 FILLER_53_236 ();
 sg13g2_fill_1 FILLER_53_238 ();
 sg13g2_fill_2 FILLER_53_243 ();
 sg13g2_fill_1 FILLER_53_258 ();
 sg13g2_fill_2 FILLER_53_269 ();
 sg13g2_fill_2 FILLER_53_280 ();
 sg13g2_fill_1 FILLER_53_282 ();
 sg13g2_decap_8 FILLER_53_298 ();
 sg13g2_decap_4 FILLER_53_305 ();
 sg13g2_fill_2 FILLER_53_309 ();
 sg13g2_fill_1 FILLER_53_319 ();
 sg13g2_fill_2 FILLER_53_337 ();
 sg13g2_decap_8 FILLER_53_373 ();
 sg13g2_decap_8 FILLER_53_380 ();
 sg13g2_decap_8 FILLER_53_387 ();
 sg13g2_decap_8 FILLER_53_394 ();
 sg13g2_decap_8 FILLER_53_401 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_fill_2 FILLER_54_91 ();
 sg13g2_fill_2 FILLER_54_119 ();
 sg13g2_fill_1 FILLER_54_121 ();
 sg13g2_fill_1 FILLER_54_147 ();
 sg13g2_fill_2 FILLER_54_153 ();
 sg13g2_fill_2 FILLER_54_184 ();
 sg13g2_fill_1 FILLER_54_217 ();
 sg13g2_fill_2 FILLER_54_223 ();
 sg13g2_fill_1 FILLER_54_225 ();
 sg13g2_decap_8 FILLER_54_311 ();
 sg13g2_fill_2 FILLER_54_318 ();
 sg13g2_decap_8 FILLER_54_341 ();
 sg13g2_decap_8 FILLER_54_369 ();
 sg13g2_decap_8 FILLER_54_376 ();
 sg13g2_decap_8 FILLER_54_383 ();
 sg13g2_decap_8 FILLER_54_390 ();
 sg13g2_decap_8 FILLER_54_397 ();
 sg13g2_decap_4 FILLER_54_404 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_fill_1 FILLER_55_130 ();
 sg13g2_fill_1 FILLER_55_292 ();
 sg13g2_fill_2 FILLER_55_309 ();
 sg13g2_fill_2 FILLER_55_331 ();
 sg13g2_decap_4 FILLER_55_337 ();
 sg13g2_decap_8 FILLER_55_359 ();
 sg13g2_decap_8 FILLER_55_366 ();
 sg13g2_decap_8 FILLER_55_373 ();
 sg13g2_decap_8 FILLER_55_380 ();
 sg13g2_decap_8 FILLER_55_387 ();
 sg13g2_decap_8 FILLER_55_394 ();
 sg13g2_decap_8 FILLER_55_401 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_4 FILLER_56_91 ();
 sg13g2_fill_1 FILLER_56_95 ();
 sg13g2_fill_2 FILLER_56_145 ();
 sg13g2_fill_2 FILLER_56_178 ();
 sg13g2_fill_2 FILLER_56_259 ();
 sg13g2_fill_1 FILLER_56_296 ();
 sg13g2_fill_2 FILLER_56_315 ();
 sg13g2_decap_8 FILLER_56_333 ();
 sg13g2_fill_2 FILLER_56_340 ();
 sg13g2_fill_1 FILLER_56_342 ();
 sg13g2_decap_8 FILLER_56_356 ();
 sg13g2_decap_8 FILLER_56_363 ();
 sg13g2_decap_8 FILLER_56_370 ();
 sg13g2_decap_8 FILLER_56_377 ();
 sg13g2_decap_8 FILLER_56_384 ();
 sg13g2_decap_8 FILLER_56_391 ();
 sg13g2_decap_8 FILLER_56_398 ();
 sg13g2_decap_4 FILLER_56_405 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_fill_2 FILLER_57_98 ();
 sg13g2_fill_2 FILLER_57_117 ();
 sg13g2_fill_2 FILLER_57_138 ();
 sg13g2_fill_1 FILLER_57_140 ();
 sg13g2_fill_2 FILLER_57_229 ();
 sg13g2_fill_1 FILLER_57_231 ();
 sg13g2_fill_1 FILLER_57_272 ();
 sg13g2_decap_8 FILLER_57_297 ();
 sg13g2_decap_8 FILLER_57_304 ();
 sg13g2_decap_4 FILLER_57_311 ();
 sg13g2_fill_1 FILLER_57_315 ();
 sg13g2_decap_8 FILLER_57_321 ();
 sg13g2_decap_8 FILLER_57_328 ();
 sg13g2_fill_2 FILLER_57_335 ();
 sg13g2_decap_8 FILLER_57_368 ();
 sg13g2_decap_8 FILLER_57_375 ();
 sg13g2_decap_8 FILLER_57_382 ();
 sg13g2_decap_8 FILLER_57_389 ();
 sg13g2_decap_8 FILLER_57_396 ();
 sg13g2_decap_4 FILLER_57_403 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_fill_2 FILLER_58_105 ();
 sg13g2_fill_2 FILLER_58_127 ();
 sg13g2_fill_2 FILLER_58_214 ();
 sg13g2_fill_1 FILLER_58_216 ();
 sg13g2_fill_1 FILLER_58_221 ();
 sg13g2_fill_1 FILLER_58_279 ();
 sg13g2_fill_2 FILLER_58_290 ();
 sg13g2_fill_1 FILLER_58_292 ();
 sg13g2_decap_8 FILLER_58_309 ();
 sg13g2_decap_4 FILLER_58_316 ();
 sg13g2_fill_1 FILLER_58_320 ();
 sg13g2_fill_2 FILLER_58_329 ();
 sg13g2_fill_2 FILLER_58_335 ();
 sg13g2_decap_4 FILLER_58_342 ();
 sg13g2_decap_8 FILLER_58_367 ();
 sg13g2_decap_8 FILLER_58_374 ();
 sg13g2_decap_8 FILLER_58_381 ();
 sg13g2_decap_8 FILLER_58_388 ();
 sg13g2_decap_8 FILLER_58_395 ();
 sg13g2_decap_8 FILLER_58_402 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_4 FILLER_59_91 ();
 sg13g2_fill_2 FILLER_59_95 ();
 sg13g2_fill_2 FILLER_59_123 ();
 sg13g2_fill_1 FILLER_59_125 ();
 sg13g2_fill_2 FILLER_59_135 ();
 sg13g2_decap_8 FILLER_59_211 ();
 sg13g2_fill_1 FILLER_59_218 ();
 sg13g2_fill_2 FILLER_59_259 ();
 sg13g2_fill_1 FILLER_59_313 ();
 sg13g2_fill_2 FILLER_59_339 ();
 sg13g2_fill_1 FILLER_59_341 ();
 sg13g2_decap_8 FILLER_59_352 ();
 sg13g2_decap_8 FILLER_59_359 ();
 sg13g2_decap_8 FILLER_59_366 ();
 sg13g2_decap_8 FILLER_59_373 ();
 sg13g2_decap_8 FILLER_59_380 ();
 sg13g2_decap_8 FILLER_59_387 ();
 sg13g2_decap_8 FILLER_59_394 ();
 sg13g2_decap_8 FILLER_59_401 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_4 FILLER_60_84 ();
 sg13g2_fill_1 FILLER_60_88 ();
 sg13g2_fill_2 FILLER_60_112 ();
 sg13g2_fill_1 FILLER_60_173 ();
 sg13g2_fill_2 FILLER_60_183 ();
 sg13g2_decap_8 FILLER_60_194 ();
 sg13g2_fill_2 FILLER_60_201 ();
 sg13g2_fill_1 FILLER_60_203 ();
 sg13g2_fill_1 FILLER_60_213 ();
 sg13g2_fill_2 FILLER_60_219 ();
 sg13g2_fill_1 FILLER_60_234 ();
 sg13g2_fill_2 FILLER_60_301 ();
 sg13g2_fill_1 FILLER_60_303 ();
 sg13g2_fill_2 FILLER_60_340 ();
 sg13g2_fill_1 FILLER_60_342 ();
 sg13g2_decap_4 FILLER_60_348 ();
 sg13g2_fill_2 FILLER_60_352 ();
 sg13g2_decap_8 FILLER_60_359 ();
 sg13g2_decap_8 FILLER_60_366 ();
 sg13g2_decap_8 FILLER_60_373 ();
 sg13g2_decap_8 FILLER_60_380 ();
 sg13g2_decap_8 FILLER_60_387 ();
 sg13g2_decap_8 FILLER_60_394 ();
 sg13g2_decap_8 FILLER_60_401 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_4 FILLER_61_91 ();
 sg13g2_fill_2 FILLER_61_95 ();
 sg13g2_fill_1 FILLER_61_133 ();
 sg13g2_fill_2 FILLER_61_148 ();
 sg13g2_fill_1 FILLER_61_176 ();
 sg13g2_fill_2 FILLER_61_182 ();
 sg13g2_fill_1 FILLER_61_184 ();
 sg13g2_fill_1 FILLER_61_229 ();
 sg13g2_fill_2 FILLER_61_244 ();
 sg13g2_fill_2 FILLER_61_310 ();
 sg13g2_fill_2 FILLER_61_326 ();
 sg13g2_fill_2 FILLER_61_354 ();
 sg13g2_decap_8 FILLER_61_365 ();
 sg13g2_decap_8 FILLER_61_372 ();
 sg13g2_decap_8 FILLER_61_379 ();
 sg13g2_decap_8 FILLER_61_386 ();
 sg13g2_decap_8 FILLER_61_393 ();
 sg13g2_decap_8 FILLER_61_400 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_4 FILLER_62_98 ();
 sg13g2_fill_2 FILLER_62_119 ();
 sg13g2_fill_1 FILLER_62_121 ();
 sg13g2_fill_2 FILLER_62_132 ();
 sg13g2_fill_1 FILLER_62_165 ();
 sg13g2_fill_2 FILLER_62_170 ();
 sg13g2_fill_1 FILLER_62_172 ();
 sg13g2_fill_2 FILLER_62_187 ();
 sg13g2_fill_2 FILLER_62_196 ();
 sg13g2_fill_1 FILLER_62_207 ();
 sg13g2_decap_4 FILLER_62_221 ();
 sg13g2_fill_1 FILLER_62_225 ();
 sg13g2_fill_2 FILLER_62_252 ();
 sg13g2_fill_1 FILLER_62_254 ();
 sg13g2_fill_2 FILLER_62_316 ();
 sg13g2_fill_2 FILLER_62_328 ();
 sg13g2_fill_1 FILLER_62_330 ();
 sg13g2_decap_8 FILLER_62_381 ();
 sg13g2_decap_8 FILLER_62_388 ();
 sg13g2_decap_8 FILLER_62_395 ();
 sg13g2_decap_8 FILLER_62_402 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_fill_1 FILLER_63_160 ();
 sg13g2_decap_8 FILLER_63_226 ();
 sg13g2_decap_4 FILLER_63_233 ();
 sg13g2_decap_8 FILLER_63_241 ();
 sg13g2_decap_4 FILLER_63_248 ();
 sg13g2_fill_2 FILLER_63_252 ();
 sg13g2_fill_2 FILLER_63_306 ();
 sg13g2_fill_1 FILLER_63_308 ();
 sg13g2_fill_2 FILLER_63_318 ();
 sg13g2_fill_2 FILLER_63_332 ();
 sg13g2_fill_1 FILLER_63_334 ();
 sg13g2_decap_8 FILLER_63_370 ();
 sg13g2_decap_8 FILLER_63_377 ();
 sg13g2_decap_8 FILLER_63_384 ();
 sg13g2_decap_8 FILLER_63_391 ();
 sg13g2_decap_8 FILLER_63_398 ();
 sg13g2_decap_4 FILLER_63_405 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_fill_2 FILLER_64_98 ();
 sg13g2_fill_1 FILLER_64_152 ();
 sg13g2_fill_2 FILLER_64_235 ();
 sg13g2_fill_1 FILLER_64_237 ();
 sg13g2_fill_2 FILLER_64_246 ();
 sg13g2_fill_2 FILLER_64_293 ();
 sg13g2_decap_8 FILLER_64_359 ();
 sg13g2_decap_8 FILLER_64_366 ();
 sg13g2_decap_8 FILLER_64_373 ();
 sg13g2_decap_8 FILLER_64_380 ();
 sg13g2_decap_8 FILLER_64_387 ();
 sg13g2_decap_8 FILLER_64_394 ();
 sg13g2_decap_8 FILLER_64_401 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_4 FILLER_65_105 ();
 sg13g2_fill_2 FILLER_65_139 ();
 sg13g2_fill_1 FILLER_65_141 ();
 sg13g2_fill_1 FILLER_65_229 ();
 sg13g2_fill_1 FILLER_65_256 ();
 sg13g2_fill_1 FILLER_65_295 ();
 sg13g2_decap_8 FILLER_65_356 ();
 sg13g2_decap_8 FILLER_65_363 ();
 sg13g2_decap_8 FILLER_65_370 ();
 sg13g2_decap_8 FILLER_65_377 ();
 sg13g2_decap_8 FILLER_65_384 ();
 sg13g2_decap_8 FILLER_65_391 ();
 sg13g2_decap_8 FILLER_65_398 ();
 sg13g2_decap_4 FILLER_65_405 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_4 FILLER_66_112 ();
 sg13g2_fill_1 FILLER_66_129 ();
 sg13g2_fill_1 FILLER_66_205 ();
 sg13g2_fill_2 FILLER_66_261 ();
 sg13g2_fill_1 FILLER_66_263 ();
 sg13g2_fill_2 FILLER_66_295 ();
 sg13g2_fill_1 FILLER_66_297 ();
 sg13g2_fill_2 FILLER_66_324 ();
 sg13g2_decap_8 FILLER_66_352 ();
 sg13g2_decap_8 FILLER_66_359 ();
 sg13g2_decap_8 FILLER_66_366 ();
 sg13g2_decap_8 FILLER_66_373 ();
 sg13g2_decap_8 FILLER_66_380 ();
 sg13g2_decap_8 FILLER_66_387 ();
 sg13g2_decap_8 FILLER_66_394 ();
 sg13g2_decap_8 FILLER_66_401 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_4 FILLER_67_119 ();
 sg13g2_fill_2 FILLER_67_123 ();
 sg13g2_fill_1 FILLER_67_130 ();
 sg13g2_fill_1 FILLER_67_144 ();
 sg13g2_fill_2 FILLER_67_204 ();
 sg13g2_fill_1 FILLER_67_260 ();
 sg13g2_fill_1 FILLER_67_270 ();
 sg13g2_fill_2 FILLER_67_293 ();
 sg13g2_fill_1 FILLER_67_305 ();
 sg13g2_fill_2 FILLER_67_341 ();
 sg13g2_fill_1 FILLER_67_343 ();
 sg13g2_decap_8 FILLER_67_353 ();
 sg13g2_decap_8 FILLER_67_360 ();
 sg13g2_decap_8 FILLER_67_367 ();
 sg13g2_decap_8 FILLER_67_374 ();
 sg13g2_decap_8 FILLER_67_381 ();
 sg13g2_decap_8 FILLER_67_388 ();
 sg13g2_decap_8 FILLER_67_395 ();
 sg13g2_decap_8 FILLER_67_402 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_4 FILLER_68_119 ();
 sg13g2_fill_2 FILLER_68_123 ();
 sg13g2_fill_1 FILLER_68_154 ();
 sg13g2_fill_1 FILLER_68_164 ();
 sg13g2_fill_1 FILLER_68_191 ();
 sg13g2_fill_1 FILLER_68_221 ();
 sg13g2_fill_2 FILLER_68_252 ();
 sg13g2_fill_1 FILLER_68_289 ();
 sg13g2_fill_2 FILLER_68_299 ();
 sg13g2_fill_1 FILLER_68_310 ();
 sg13g2_fill_2 FILLER_68_324 ();
 sg13g2_decap_8 FILLER_68_344 ();
 sg13g2_decap_8 FILLER_68_351 ();
 sg13g2_decap_8 FILLER_68_358 ();
 sg13g2_decap_8 FILLER_68_365 ();
 sg13g2_decap_8 FILLER_68_372 ();
 sg13g2_decap_8 FILLER_68_379 ();
 sg13g2_decap_8 FILLER_68_386 ();
 sg13g2_decap_8 FILLER_68_393 ();
 sg13g2_decap_8 FILLER_68_400 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_4 FILLER_69_126 ();
 sg13g2_fill_1 FILLER_69_166 ();
 sg13g2_fill_1 FILLER_69_180 ();
 sg13g2_fill_1 FILLER_69_206 ();
 sg13g2_decap_8 FILLER_69_346 ();
 sg13g2_decap_8 FILLER_69_353 ();
 sg13g2_decap_8 FILLER_69_360 ();
 sg13g2_decap_8 FILLER_69_367 ();
 sg13g2_decap_8 FILLER_69_374 ();
 sg13g2_decap_8 FILLER_69_381 ();
 sg13g2_decap_8 FILLER_69_388 ();
 sg13g2_decap_8 FILLER_69_395 ();
 sg13g2_decap_8 FILLER_69_402 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_4 FILLER_70_133 ();
 sg13g2_fill_1 FILLER_70_137 ();
 sg13g2_fill_1 FILLER_70_155 ();
 sg13g2_fill_2 FILLER_70_183 ();
 sg13g2_fill_2 FILLER_70_199 ();
 sg13g2_fill_1 FILLER_70_224 ();
 sg13g2_fill_2 FILLER_70_274 ();
 sg13g2_decap_8 FILLER_70_332 ();
 sg13g2_decap_8 FILLER_70_339 ();
 sg13g2_decap_8 FILLER_70_346 ();
 sg13g2_decap_8 FILLER_70_353 ();
 sg13g2_decap_8 FILLER_70_360 ();
 sg13g2_decap_8 FILLER_70_367 ();
 sg13g2_decap_8 FILLER_70_374 ();
 sg13g2_decap_8 FILLER_70_381 ();
 sg13g2_decap_8 FILLER_70_388 ();
 sg13g2_decap_8 FILLER_70_395 ();
 sg13g2_decap_8 FILLER_70_402 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_4 FILLER_71_140 ();
 sg13g2_fill_2 FILLER_71_144 ();
 sg13g2_fill_2 FILLER_71_262 ();
 sg13g2_decap_8 FILLER_71_317 ();
 sg13g2_decap_8 FILLER_71_324 ();
 sg13g2_decap_8 FILLER_71_331 ();
 sg13g2_decap_8 FILLER_71_338 ();
 sg13g2_decap_8 FILLER_71_345 ();
 sg13g2_decap_8 FILLER_71_352 ();
 sg13g2_decap_8 FILLER_71_359 ();
 sg13g2_decap_8 FILLER_71_366 ();
 sg13g2_decap_8 FILLER_71_373 ();
 sg13g2_decap_8 FILLER_71_380 ();
 sg13g2_decap_8 FILLER_71_387 ();
 sg13g2_decap_8 FILLER_71_394 ();
 sg13g2_decap_8 FILLER_71_401 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_4 FILLER_72_133 ();
 sg13g2_fill_2 FILLER_72_181 ();
 sg13g2_fill_2 FILLER_72_262 ();
 sg13g2_fill_1 FILLER_72_264 ();
 sg13g2_fill_2 FILLER_72_284 ();
 sg13g2_fill_1 FILLER_72_286 ();
 sg13g2_decap_8 FILLER_72_304 ();
 sg13g2_decap_8 FILLER_72_311 ();
 sg13g2_decap_8 FILLER_72_318 ();
 sg13g2_decap_8 FILLER_72_325 ();
 sg13g2_decap_8 FILLER_72_332 ();
 sg13g2_decap_8 FILLER_72_339 ();
 sg13g2_decap_8 FILLER_72_346 ();
 sg13g2_decap_8 FILLER_72_353 ();
 sg13g2_decap_8 FILLER_72_360 ();
 sg13g2_decap_8 FILLER_72_367 ();
 sg13g2_decap_8 FILLER_72_374 ();
 sg13g2_decap_8 FILLER_72_381 ();
 sg13g2_decap_8 FILLER_72_388 ();
 sg13g2_decap_8 FILLER_72_395 ();
 sg13g2_decap_8 FILLER_72_402 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_4 FILLER_73_140 ();
 sg13g2_fill_2 FILLER_73_199 ();
 sg13g2_fill_1 FILLER_73_219 ();
 sg13g2_fill_2 FILLER_73_246 ();
 sg13g2_decap_8 FILLER_73_296 ();
 sg13g2_decap_8 FILLER_73_303 ();
 sg13g2_decap_8 FILLER_73_310 ();
 sg13g2_decap_8 FILLER_73_317 ();
 sg13g2_decap_8 FILLER_73_324 ();
 sg13g2_decap_8 FILLER_73_331 ();
 sg13g2_decap_8 FILLER_73_338 ();
 sg13g2_decap_8 FILLER_73_345 ();
 sg13g2_decap_8 FILLER_73_352 ();
 sg13g2_decap_8 FILLER_73_359 ();
 sg13g2_decap_8 FILLER_73_366 ();
 sg13g2_decap_8 FILLER_73_373 ();
 sg13g2_decap_8 FILLER_73_380 ();
 sg13g2_decap_8 FILLER_73_387 ();
 sg13g2_decap_8 FILLER_73_394 ();
 sg13g2_decap_8 FILLER_73_401 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_4 FILLER_74_140 ();
 sg13g2_fill_1 FILLER_74_192 ();
 sg13g2_fill_1 FILLER_74_207 ();
 sg13g2_fill_2 FILLER_74_221 ();
 sg13g2_fill_2 FILLER_74_241 ();
 sg13g2_fill_1 FILLER_74_256 ();
 sg13g2_decap_8 FILLER_74_296 ();
 sg13g2_decap_8 FILLER_74_303 ();
 sg13g2_decap_8 FILLER_74_310 ();
 sg13g2_decap_8 FILLER_74_317 ();
 sg13g2_decap_8 FILLER_74_324 ();
 sg13g2_decap_8 FILLER_74_331 ();
 sg13g2_decap_8 FILLER_74_338 ();
 sg13g2_decap_8 FILLER_74_345 ();
 sg13g2_decap_8 FILLER_74_352 ();
 sg13g2_decap_8 FILLER_74_359 ();
 sg13g2_decap_8 FILLER_74_366 ();
 sg13g2_decap_8 FILLER_74_373 ();
 sg13g2_decap_8 FILLER_74_380 ();
 sg13g2_decap_8 FILLER_74_387 ();
 sg13g2_decap_8 FILLER_74_394 ();
 sg13g2_decap_8 FILLER_74_401 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_4 FILLER_75_140 ();
 sg13g2_fill_2 FILLER_75_144 ();
 sg13g2_fill_1 FILLER_75_168 ();
 sg13g2_fill_1 FILLER_75_178 ();
 sg13g2_fill_1 FILLER_75_187 ();
 sg13g2_fill_1 FILLER_75_205 ();
 sg13g2_fill_1 FILLER_75_232 ();
 sg13g2_decap_8 FILLER_75_309 ();
 sg13g2_decap_8 FILLER_75_316 ();
 sg13g2_decap_8 FILLER_75_323 ();
 sg13g2_decap_8 FILLER_75_330 ();
 sg13g2_decap_8 FILLER_75_337 ();
 sg13g2_decap_8 FILLER_75_344 ();
 sg13g2_decap_8 FILLER_75_351 ();
 sg13g2_decap_8 FILLER_75_358 ();
 sg13g2_decap_8 FILLER_75_365 ();
 sg13g2_decap_8 FILLER_75_372 ();
 sg13g2_decap_8 FILLER_75_379 ();
 sg13g2_decap_8 FILLER_75_386 ();
 sg13g2_decap_8 FILLER_75_393 ();
 sg13g2_decap_8 FILLER_75_400 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_4 FILLER_76_140 ();
 sg13g2_fill_2 FILLER_76_144 ();
 sg13g2_fill_2 FILLER_76_213 ();
 sg13g2_fill_1 FILLER_76_215 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_392 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_fill_2 FILLER_76_406 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_4 FILLER_77_140 ();
 sg13g2_fill_1 FILLER_77_144 ();
 sg13g2_fill_1 FILLER_77_176 ();
 sg13g2_fill_1 FILLER_77_217 ();
 sg13g2_fill_1 FILLER_77_281 ();
 sg13g2_decap_8 FILLER_77_297 ();
 sg13g2_decap_8 FILLER_77_304 ();
 sg13g2_decap_8 FILLER_77_311 ();
 sg13g2_decap_8 FILLER_77_318 ();
 sg13g2_decap_8 FILLER_77_325 ();
 sg13g2_decap_8 FILLER_77_332 ();
 sg13g2_decap_8 FILLER_77_339 ();
 sg13g2_decap_8 FILLER_77_346 ();
 sg13g2_decap_8 FILLER_77_353 ();
 sg13g2_decap_8 FILLER_77_360 ();
 sg13g2_decap_8 FILLER_77_367 ();
 sg13g2_decap_8 FILLER_77_374 ();
 sg13g2_decap_8 FILLER_77_381 ();
 sg13g2_decap_8 FILLER_77_388 ();
 sg13g2_decap_8 FILLER_77_395 ();
 sg13g2_decap_8 FILLER_77_402 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_fill_2 FILLER_78_147 ();
 sg13g2_fill_1 FILLER_78_149 ();
 sg13g2_fill_2 FILLER_78_267 ();
 sg13g2_fill_1 FILLER_78_269 ();
 sg13g2_decap_8 FILLER_78_305 ();
 sg13g2_decap_8 FILLER_78_312 ();
 sg13g2_decap_8 FILLER_78_319 ();
 sg13g2_decap_8 FILLER_78_326 ();
 sg13g2_decap_8 FILLER_78_333 ();
 sg13g2_decap_8 FILLER_78_340 ();
 sg13g2_decap_8 FILLER_78_347 ();
 sg13g2_decap_8 FILLER_78_354 ();
 sg13g2_decap_8 FILLER_78_361 ();
 sg13g2_decap_8 FILLER_78_368 ();
 sg13g2_decap_8 FILLER_78_375 ();
 sg13g2_decap_8 FILLER_78_382 ();
 sg13g2_decap_8 FILLER_78_389 ();
 sg13g2_decap_8 FILLER_78_396 ();
 sg13g2_decap_4 FILLER_78_403 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_4 FILLER_79_154 ();
 sg13g2_fill_1 FILLER_79_158 ();
 sg13g2_fill_2 FILLER_79_188 ();
 sg13g2_fill_2 FILLER_79_208 ();
 sg13g2_fill_1 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_296 ();
 sg13g2_decap_8 FILLER_79_303 ();
 sg13g2_decap_8 FILLER_79_310 ();
 sg13g2_decap_8 FILLER_79_317 ();
 sg13g2_decap_8 FILLER_79_324 ();
 sg13g2_decap_8 FILLER_79_331 ();
 sg13g2_decap_8 FILLER_79_338 ();
 sg13g2_decap_8 FILLER_79_345 ();
 sg13g2_decap_8 FILLER_79_352 ();
 sg13g2_decap_8 FILLER_79_359 ();
 sg13g2_decap_8 FILLER_79_366 ();
 sg13g2_decap_8 FILLER_79_373 ();
 sg13g2_decap_8 FILLER_79_380 ();
 sg13g2_decap_8 FILLER_79_387 ();
 sg13g2_decap_8 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_401 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_8 FILLER_80_124 ();
 sg13g2_decap_8 FILLER_80_131 ();
 sg13g2_decap_8 FILLER_80_138 ();
 sg13g2_decap_8 FILLER_80_145 ();
 sg13g2_decap_8 FILLER_80_152 ();
 sg13g2_decap_8 FILLER_80_159 ();
 sg13g2_fill_1 FILLER_80_166 ();
 sg13g2_fill_1 FILLER_80_214 ();
 sg13g2_fill_2 FILLER_80_235 ();
 sg13g2_fill_1 FILLER_80_237 ();
 sg13g2_fill_2 FILLER_80_247 ();
 sg13g2_fill_1 FILLER_80_267 ();
 sg13g2_decap_8 FILLER_80_294 ();
 sg13g2_decap_8 FILLER_80_301 ();
 sg13g2_decap_8 FILLER_80_308 ();
 sg13g2_decap_8 FILLER_80_315 ();
 sg13g2_decap_8 FILLER_80_322 ();
 sg13g2_decap_8 FILLER_80_329 ();
 sg13g2_decap_8 FILLER_80_336 ();
 sg13g2_fill_1 FILLER_80_343 ();
 sg13g2_decap_8 FILLER_80_348 ();
 sg13g2_decap_4 FILLER_80_355 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_decap_4 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_373 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net227;
 assign uio_oe[1] = net228;
 assign uio_oe[2] = net229;
 assign uio_oe[3] = net230;
 assign uio_oe[4] = net231;
 assign uio_oe[5] = net232;
 assign uio_oe[6] = net233;
 assign uio_oe[7] = net5;
 assign uio_out[7] = net6;
 assign uo_out[0] = net7;
 assign uo_out[1] = net8;
 assign uo_out[2] = net9;
 assign uo_out[3] = net10;
 assign uo_out[4] = net11;
 assign uo_out[5] = net12;
 assign uo_out[6] = net13;
 assign uo_out[7] = net14;
endmodule

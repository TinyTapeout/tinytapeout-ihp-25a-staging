module tt_um_tiny_ternary_tapeout (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire clknet_0_clk;
 wire \count[0] ;
 wire \count[1] ;
 wire \count[2] ;
 wire \count[3] ;
 wire \load_weights[0] ;
 wire \load_weights[10] ;
 wire \load_weights[11] ;
 wire \load_weights[12] ;
 wire \load_weights[13] ;
 wire \load_weights[14] ;
 wire \load_weights[15] ;
 wire \load_weights[16] ;
 wire \load_weights[17] ;
 wire \load_weights[18] ;
 wire \load_weights[19] ;
 wire \load_weights[1] ;
 wire \load_weights[2] ;
 wire \load_weights[3] ;
 wire \load_weights[4] ;
 wire \load_weights[5] ;
 wire \load_weights[6] ;
 wire \load_weights[7] ;
 wire \load_weights[8] ;
 wire \load_weights[9] ;
 wire state;
 wire \tt_um_load_inst.input_to_sr[0] ;
 wire \tt_um_load_inst.input_to_sr[10] ;
 wire \tt_um_load_inst.input_to_sr[11] ;
 wire \tt_um_load_inst.input_to_sr[12] ;
 wire \tt_um_load_inst.input_to_sr[13] ;
 wire \tt_um_load_inst.input_to_sr[14] ;
 wire \tt_um_load_inst.input_to_sr[15] ;
 wire \tt_um_load_inst.input_to_sr[16] ;
 wire \tt_um_load_inst.input_to_sr[17] ;
 wire \tt_um_load_inst.input_to_sr[18] ;
 wire \tt_um_load_inst.input_to_sr[19] ;
 wire \tt_um_load_inst.input_to_sr[1] ;
 wire \tt_um_load_inst.input_to_sr[2] ;
 wire \tt_um_load_inst.input_to_sr[3] ;
 wire \tt_um_load_inst.input_to_sr[4] ;
 wire \tt_um_load_inst.input_to_sr[5] ;
 wire \tt_um_load_inst.input_to_sr[6] ;
 wire \tt_um_load_inst.input_to_sr[7] ;
 wire \tt_um_load_inst.input_to_sr[8] ;
 wire \tt_um_load_inst.input_to_sr[9] ;
 wire \tt_um_load_inst.weights[20] ;
 wire \tt_um_load_inst.weights[21] ;
 wire \tt_um_load_inst.weights[22] ;
 wire \tt_um_load_inst.weights[23] ;
 wire \tt_um_load_inst.weights[24] ;
 wire \tt_um_load_inst.weights[25] ;
 wire \tt_um_load_inst.weights[26] ;
 wire \tt_um_load_inst.weights[27] ;
 wire \tt_um_load_inst.weights[28] ;
 wire \tt_um_load_inst.weights[29] ;
 wire \tt_um_load_inst.weights[30] ;
 wire \tt_um_load_inst.weights[31] ;
 wire \tt_um_load_inst.weights[32] ;
 wire \tt_um_load_inst.weights[33] ;
 wire \tt_um_load_inst.weights[34] ;
 wire \tt_um_load_inst.weights[35] ;
 wire \tt_um_load_inst.weights[36] ;
 wire \tt_um_load_inst.weights[37] ;
 wire \tt_um_load_inst.weights[38] ;
 wire \tt_um_load_inst.weights[39] ;
 wire \tt_um_load_inst.weights[40] ;
 wire \tt_um_load_inst.weights[41] ;
 wire \tt_um_load_inst.weights[42] ;
 wire \tt_um_load_inst.weights[43] ;
 wire \tt_um_load_inst.weights[44] ;
 wire \tt_um_load_inst.weights[45] ;
 wire \tt_um_load_inst.weights[46] ;
 wire \tt_um_load_inst.weights[47] ;
 wire \tt_um_load_inst.weights[48] ;
 wire \tt_um_load_inst.weights[49] ;
 wire \tt_um_load_inst.weights[50] ;
 wire \tt_um_load_inst.weights[51] ;
 wire \tt_um_load_inst.weights[52] ;
 wire \tt_um_load_inst.weights[53] ;
 wire \tt_um_load_inst.weights[54] ;
 wire \tt_um_load_inst.weights[55] ;
 wire \tt_um_load_inst.weights[56] ;
 wire \tt_um_load_inst.weights[57] ;
 wire \tt_um_load_inst.weights[58] ;
 wire \tt_um_load_inst.weights[59] ;
 wire \tt_um_load_inst.weights[60] ;
 wire \tt_um_load_inst.weights[61] ;
 wire \tt_um_load_inst.weights[62] ;
 wire \tt_um_load_inst.weights[63] ;
 wire \tt_um_load_inst.weights[64] ;
 wire \tt_um_load_inst.weights[65] ;
 wire \tt_um_load_inst.weights[66] ;
 wire \tt_um_load_inst.weights[67] ;
 wire \tt_um_load_inst.weights[68] ;
 wire \tt_um_load_inst.weights[69] ;
 wire \tt_um_load_inst.weights[70] ;
 wire \tt_um_load_inst.weights[71] ;
 wire \tt_um_load_inst.weights[72] ;
 wire \tt_um_load_inst.weights[73] ;
 wire \tt_um_load_inst.weights[74] ;
 wire \tt_um_load_inst.weights[75] ;
 wire \tt_um_load_inst.weights[76] ;
 wire \tt_um_load_inst.weights[77] ;
 wire \tt_um_load_inst.weights[78] ;
 wire \tt_um_load_inst.weights[79] ;
 wire \tt_um_load_inst.weights[80] ;
 wire \tt_um_load_inst.weights[81] ;
 wire \tt_um_load_inst.weights[82] ;
 wire \tt_um_load_inst.weights[83] ;
 wire \tt_um_load_inst.weights[84] ;
 wire \tt_um_load_inst.weights[85] ;
 wire \tt_um_load_inst.weights[86] ;
 wire \tt_um_load_inst.weights[87] ;
 wire \tt_um_load_inst.weights[88] ;
 wire \tt_um_load_inst.weights[89] ;
 wire \tt_um_load_inst.weights[90] ;
 wire \tt_um_load_inst.weights[91] ;
 wire \tt_um_load_inst.weights[92] ;
 wire \tt_um_load_inst.weights[93] ;
 wire \tt_um_load_inst.weights[94] ;
 wire \tt_um_load_inst.weights[95] ;
 wire \tt_um_load_inst.weights[96] ;
 wire \tt_um_load_inst.weights[97] ;
 wire \tt_um_load_inst.weights[98] ;
 wire \tt_um_load_inst.weights[99] ;
 wire \tt_um_mult_inst.pipe_out[0] ;
 wire \tt_um_mult_inst.pipe_out[10] ;
 wire \tt_um_mult_inst.pipe_out[11] ;
 wire \tt_um_mult_inst.pipe_out[12] ;
 wire \tt_um_mult_inst.pipe_out[13] ;
 wire \tt_um_mult_inst.pipe_out[14] ;
 wire \tt_um_mult_inst.pipe_out[15] ;
 wire \tt_um_mult_inst.pipe_out[16] ;
 wire \tt_um_mult_inst.pipe_out[17] ;
 wire \tt_um_mult_inst.pipe_out[18] ;
 wire \tt_um_mult_inst.pipe_out[19] ;
 wire \tt_um_mult_inst.pipe_out[1] ;
 wire \tt_um_mult_inst.pipe_out[20] ;
 wire \tt_um_mult_inst.pipe_out[21] ;
 wire \tt_um_mult_inst.pipe_out[22] ;
 wire \tt_um_mult_inst.pipe_out[23] ;
 wire \tt_um_mult_inst.pipe_out[24] ;
 wire \tt_um_mult_inst.pipe_out[25] ;
 wire \tt_um_mult_inst.pipe_out[26] ;
 wire \tt_um_mult_inst.pipe_out[27] ;
 wire \tt_um_mult_inst.pipe_out[28] ;
 wire \tt_um_mult_inst.pipe_out[29] ;
 wire \tt_um_mult_inst.pipe_out[2] ;
 wire \tt_um_mult_inst.pipe_out[30] ;
 wire \tt_um_mult_inst.pipe_out[31] ;
 wire \tt_um_mult_inst.pipe_out[32] ;
 wire \tt_um_mult_inst.pipe_out[33] ;
 wire \tt_um_mult_inst.pipe_out[34] ;
 wire \tt_um_mult_inst.pipe_out[35] ;
 wire \tt_um_mult_inst.pipe_out[36] ;
 wire \tt_um_mult_inst.pipe_out[37] ;
 wire \tt_um_mult_inst.pipe_out[38] ;
 wire \tt_um_mult_inst.pipe_out[39] ;
 wire \tt_um_mult_inst.pipe_out[3] ;
 wire \tt_um_mult_inst.pipe_out[4] ;
 wire \tt_um_mult_inst.pipe_out[5] ;
 wire \tt_um_mult_inst.pipe_out[6] ;
 wire \tt_um_mult_inst.pipe_out[7] ;
 wire \tt_um_mult_inst.pipe_out[8] ;
 wire \tt_um_mult_inst.pipe_out[9] ;
 wire \tt_um_mult_inst.temp_out[0] ;
 wire \tt_um_mult_inst.temp_out[10] ;
 wire \tt_um_mult_inst.temp_out[11] ;
 wire \tt_um_mult_inst.temp_out[12] ;
 wire \tt_um_mult_inst.temp_out[13] ;
 wire \tt_um_mult_inst.temp_out[14] ;
 wire \tt_um_mult_inst.temp_out[15] ;
 wire \tt_um_mult_inst.temp_out[16] ;
 wire \tt_um_mult_inst.temp_out[17] ;
 wire \tt_um_mult_inst.temp_out[18] ;
 wire \tt_um_mult_inst.temp_out[19] ;
 wire \tt_um_mult_inst.temp_out[1] ;
 wire \tt_um_mult_inst.temp_out[20] ;
 wire \tt_um_mult_inst.temp_out[21] ;
 wire \tt_um_mult_inst.temp_out[22] ;
 wire \tt_um_mult_inst.temp_out[23] ;
 wire \tt_um_mult_inst.temp_out[24] ;
 wire \tt_um_mult_inst.temp_out[25] ;
 wire \tt_um_mult_inst.temp_out[26] ;
 wire \tt_um_mult_inst.temp_out[27] ;
 wire \tt_um_mult_inst.temp_out[28] ;
 wire \tt_um_mult_inst.temp_out[29] ;
 wire \tt_um_mult_inst.temp_out[2] ;
 wire \tt_um_mult_inst.temp_out[30] ;
 wire \tt_um_mult_inst.temp_out[31] ;
 wire \tt_um_mult_inst.temp_out[32] ;
 wire \tt_um_mult_inst.temp_out[33] ;
 wire \tt_um_mult_inst.temp_out[34] ;
 wire \tt_um_mult_inst.temp_out[35] ;
 wire \tt_um_mult_inst.temp_out[36] ;
 wire \tt_um_mult_inst.temp_out[37] ;
 wire \tt_um_mult_inst.temp_out[38] ;
 wire \tt_um_mult_inst.temp_out[39] ;
 wire \tt_um_mult_inst.temp_out[3] ;
 wire \tt_um_mult_inst.temp_out[4] ;
 wire \tt_um_mult_inst.temp_out[5] ;
 wire \tt_um_mult_inst.temp_out[6] ;
 wire \tt_um_mult_inst.temp_out[7] ;
 wire \tt_um_mult_inst.temp_out[8] ;
 wire \tt_um_mult_inst.temp_out[9] ;
 wire \tt_um_mult_inst.temp_out_comb[0] ;
 wire \tt_um_mult_inst.temp_out_comb[10] ;
 wire \tt_um_mult_inst.temp_out_comb[11] ;
 wire \tt_um_mult_inst.temp_out_comb[12] ;
 wire \tt_um_mult_inst.temp_out_comb[13] ;
 wire \tt_um_mult_inst.temp_out_comb[14] ;
 wire \tt_um_mult_inst.temp_out_comb[15] ;
 wire \tt_um_mult_inst.temp_out_comb[16] ;
 wire \tt_um_mult_inst.temp_out_comb[17] ;
 wire \tt_um_mult_inst.temp_out_comb[18] ;
 wire \tt_um_mult_inst.temp_out_comb[19] ;
 wire \tt_um_mult_inst.temp_out_comb[1] ;
 wire \tt_um_mult_inst.temp_out_comb[20] ;
 wire \tt_um_mult_inst.temp_out_comb[21] ;
 wire \tt_um_mult_inst.temp_out_comb[22] ;
 wire \tt_um_mult_inst.temp_out_comb[23] ;
 wire \tt_um_mult_inst.temp_out_comb[24] ;
 wire \tt_um_mult_inst.temp_out_comb[25] ;
 wire \tt_um_mult_inst.temp_out_comb[26] ;
 wire \tt_um_mult_inst.temp_out_comb[27] ;
 wire \tt_um_mult_inst.temp_out_comb[28] ;
 wire \tt_um_mult_inst.temp_out_comb[29] ;
 wire \tt_um_mult_inst.temp_out_comb[2] ;
 wire \tt_um_mult_inst.temp_out_comb[30] ;
 wire \tt_um_mult_inst.temp_out_comb[31] ;
 wire \tt_um_mult_inst.temp_out_comb[32] ;
 wire \tt_um_mult_inst.temp_out_comb[33] ;
 wire \tt_um_mult_inst.temp_out_comb[34] ;
 wire \tt_um_mult_inst.temp_out_comb[35] ;
 wire \tt_um_mult_inst.temp_out_comb[36] ;
 wire \tt_um_mult_inst.temp_out_comb[37] ;
 wire \tt_um_mult_inst.temp_out_comb[38] ;
 wire \tt_um_mult_inst.temp_out_comb[39] ;
 wire \tt_um_mult_inst.temp_out_comb[3] ;
 wire \tt_um_mult_inst.temp_out_comb[4] ;
 wire \tt_um_mult_inst.temp_out_comb[5] ;
 wire \tt_um_mult_inst.temp_out_comb[6] ;
 wire \tt_um_mult_inst.temp_out_comb[7] ;
 wire \tt_um_mult_inst.temp_out_comb[8] ;
 wire \tt_um_mult_inst.temp_out_comb[9] ;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;

 sg13g2_inv_1 _0963_ (.Y(_0046_),
    .A(net1));
 sg13g2_inv_1 _0964_ (.Y(_0047_),
    .A(\tt_um_mult_inst.temp_out[0] ));
 sg13g2_inv_1 _0965_ (.Y(_0048_),
    .A(net389));
 sg13g2_inv_1 _0966_ (.Y(_0049_),
    .A(net442));
 sg13g2_inv_1 _0967_ (.Y(_0050_),
    .A(net438));
 sg13g2_inv_1 _0968_ (.Y(_0051_),
    .A(net4));
 sg13g2_inv_1 _0969_ (.Y(_0052_),
    .A(net5));
 sg13g2_inv_1 _0970_ (.Y(_0053_),
    .A(net336));
 sg13g2_nor2_1 _0971_ (.A(\count[3] ),
    .B(net110),
    .Y(_0054_));
 sg13g2_mux2_1 _0972_ (.A0(net431),
    .A1(net119),
    .S(net107),
    .X(\tt_um_load_inst.input_to_sr[0] ));
 sg13g2_mux2_1 _0973_ (.A0(net439),
    .A1(net117),
    .S(net108),
    .X(\tt_um_load_inst.input_to_sr[1] ));
 sg13g2_mux2_1 _0974_ (.A0(net430),
    .A1(net115),
    .S(net108),
    .X(\tt_um_load_inst.input_to_sr[2] ));
 sg13g2_mux2_1 _0975_ (.A0(net426),
    .A1(net114),
    .S(net107),
    .X(\tt_um_load_inst.input_to_sr[3] ));
 sg13g2_mux2_1 _0976_ (.A0(net435),
    .A1(net113),
    .S(net107),
    .X(\tt_um_load_inst.input_to_sr[4] ));
 sg13g2_mux2_1 _0977_ (.A0(net429),
    .A1(net112),
    .S(net107),
    .X(\tt_um_load_inst.input_to_sr[5] ));
 sg13g2_mux2_1 _0978_ (.A0(net433),
    .A1(net111),
    .S(net107),
    .X(\tt_um_load_inst.input_to_sr[6] ));
 sg13g2_mux2_1 _0979_ (.A0(net423),
    .A1(net14),
    .S(net107),
    .X(\tt_um_load_inst.input_to_sr[7] ));
 sg13g2_mux2_1 _0980_ (.A0(net414),
    .A1(net122),
    .S(net107),
    .X(\tt_um_load_inst.input_to_sr[8] ));
 sg13g2_mux2_1 _0981_ (.A0(net415),
    .A1(net120),
    .S(net107),
    .X(\tt_um_load_inst.input_to_sr[9] ));
 sg13g2_mux2_1 _0982_ (.A0(net8),
    .A1(net421),
    .S(net110),
    .X(\tt_um_load_inst.input_to_sr[10] ));
 sg13g2_mux2_1 _0983_ (.A0(net118),
    .A1(net419),
    .S(net110),
    .X(\tt_um_load_inst.input_to_sr[11] ));
 sg13g2_mux2_1 _0984_ (.A0(net9),
    .A1(net424),
    .S(net109),
    .X(\tt_um_load_inst.input_to_sr[12] ));
 sg13g2_mux2_1 _0985_ (.A0(net10),
    .A1(net408),
    .S(net109),
    .X(\tt_um_load_inst.input_to_sr[13] ));
 sg13g2_mux2_1 _0986_ (.A0(net113),
    .A1(net440),
    .S(net109),
    .X(\tt_um_load_inst.input_to_sr[14] ));
 sg13g2_mux2_1 _0987_ (.A0(net12),
    .A1(net412),
    .S(net109),
    .X(\tt_um_load_inst.input_to_sr[15] ));
 sg13g2_mux2_1 _0988_ (.A0(net111),
    .A1(net436),
    .S(net109),
    .X(\tt_um_load_inst.input_to_sr[16] ));
 sg13g2_mux2_1 _0989_ (.A0(net14),
    .A1(net416),
    .S(net109),
    .X(\tt_um_load_inst.input_to_sr[17] ));
 sg13g2_mux2_1 _0990_ (.A0(net122),
    .A1(net427),
    .S(net109),
    .X(\tt_um_load_inst.input_to_sr[18] ));
 sg13g2_mux2_1 _0991_ (.A0(net121),
    .A1(net410),
    .S(net109),
    .X(\tt_um_load_inst.input_to_sr[19] ));
 sg13g2_nor2_1 _0992_ (.A(net404),
    .B(net418),
    .Y(_0055_));
 sg13g2_nor3_1 _0993_ (.A(\count[1] ),
    .B(\count[0] ),
    .C(\count[2] ),
    .Y(_0056_));
 sg13g2_or3_2 _0994_ (.A(\count[1] ),
    .B(\count[0] ),
    .C(\count[2] ),
    .X(_0057_));
 sg13g2_nor2_1 _0995_ (.A(net379),
    .B(net105),
    .Y(_0058_));
 sg13g2_a21oi_1 _0996_ (.A1(_0047_),
    .A2(net104),
    .Y(_0000_),
    .B1(_0058_));
 sg13g2_mux2_1 _0997_ (.A0(net375),
    .A1(\tt_um_mult_inst.temp_out[1] ),
    .S(net104),
    .X(_0011_));
 sg13g2_mux2_1 _0998_ (.A0(net385),
    .A1(\tt_um_mult_inst.temp_out[2] ),
    .S(net105),
    .X(_0022_));
 sg13g2_mux2_1 _0999_ (.A0(net357),
    .A1(\tt_um_mult_inst.temp_out[3] ),
    .S(net105),
    .X(_0025_));
 sg13g2_mux2_1 _1000_ (.A0(net349),
    .A1(\tt_um_mult_inst.temp_out[4] ),
    .S(net105),
    .X(_0026_));
 sg13g2_mux2_1 _1001_ (.A0(net339),
    .A1(\tt_um_mult_inst.temp_out[5] ),
    .S(net100),
    .X(_0027_));
 sg13g2_mux2_1 _1002_ (.A0(net355),
    .A1(\tt_um_mult_inst.temp_out[6] ),
    .S(net100),
    .X(_0028_));
 sg13g2_mux2_1 _1003_ (.A0(net347),
    .A1(\tt_um_mult_inst.temp_out[7] ),
    .S(net100),
    .X(_0029_));
 sg13g2_nor2_1 _1004_ (.A(\tt_um_mult_inst.pipe_out[16] ),
    .B(net106),
    .Y(_0059_));
 sg13g2_a21oi_1 _1005_ (.A1(_0048_),
    .A2(net104),
    .Y(_0030_),
    .B1(_0059_));
 sg13g2_mux2_1 _1006_ (.A0(net367),
    .A1(\tt_um_mult_inst.temp_out[9] ),
    .S(net104),
    .X(_0031_));
 sg13g2_mux2_1 _1007_ (.A0(net395),
    .A1(\tt_um_mult_inst.temp_out[10] ),
    .S(net104),
    .X(_0001_));
 sg13g2_mux2_1 _1008_ (.A0(net397),
    .A1(\tt_um_mult_inst.temp_out[11] ),
    .S(net104),
    .X(_0002_));
 sg13g2_mux2_1 _1009_ (.A0(net334),
    .A1(\tt_um_mult_inst.temp_out[12] ),
    .S(net100),
    .X(_0003_));
 sg13g2_mux2_1 _1010_ (.A0(net373),
    .A1(\tt_um_mult_inst.temp_out[13] ),
    .S(net100),
    .X(_0004_));
 sg13g2_mux2_1 _1011_ (.A0(net351),
    .A1(\tt_um_mult_inst.temp_out[14] ),
    .S(net99),
    .X(_0005_));
 sg13g2_mux2_1 _1012_ (.A0(net381),
    .A1(\tt_um_mult_inst.temp_out[15] ),
    .S(net99),
    .X(_0006_));
 sg13g2_nor2_1 _1013_ (.A(net369),
    .B(net102),
    .Y(_0060_));
 sg13g2_a21oi_1 _1014_ (.A1(_0049_),
    .A2(net102),
    .Y(_0007_),
    .B1(_0060_));
 sg13g2_mux2_1 _1015_ (.A0(net383),
    .A1(\tt_um_mult_inst.temp_out[17] ),
    .S(net102),
    .X(_0008_));
 sg13g2_mux2_1 _1016_ (.A0(net363),
    .A1(\tt_um_mult_inst.temp_out[18] ),
    .S(net102),
    .X(_0009_));
 sg13g2_mux2_1 _1017_ (.A0(net377),
    .A1(\tt_um_mult_inst.temp_out[19] ),
    .S(net104),
    .X(_0010_));
 sg13g2_mux2_1 _1018_ (.A0(\tt_um_mult_inst.pipe_out[28] ),
    .A1(net399),
    .S(net100),
    .X(_0012_));
 sg13g2_mux2_1 _1019_ (.A0(net371),
    .A1(\tt_um_mult_inst.temp_out[21] ),
    .S(net99),
    .X(_0013_));
 sg13g2_mux2_1 _1020_ (.A0(net391),
    .A1(\tt_um_mult_inst.temp_out[22] ),
    .S(net99),
    .X(_0014_));
 sg13g2_mux2_1 _1021_ (.A0(net359),
    .A1(\tt_um_mult_inst.temp_out[23] ),
    .S(net99),
    .X(_0015_));
 sg13g2_nor2_1 _1022_ (.A(net345),
    .B(net102),
    .Y(_0061_));
 sg13g2_a21oi_1 _1023_ (.A1(_0050_),
    .A2(net102),
    .Y(_0016_),
    .B1(_0061_));
 sg13g2_mux2_1 _1024_ (.A0(net343),
    .A1(\tt_um_mult_inst.temp_out[25] ),
    .S(net102),
    .X(_0017_));
 sg13g2_mux2_1 _1025_ (.A0(net365),
    .A1(\tt_um_mult_inst.temp_out[26] ),
    .S(net103),
    .X(_0018_));
 sg13g2_mux2_1 _1026_ (.A0(net387),
    .A1(\tt_um_mult_inst.temp_out[27] ),
    .S(net103),
    .X(_0019_));
 sg13g2_mux2_1 _1027_ (.A0(net341),
    .A1(\tt_um_mult_inst.temp_out[28] ),
    .S(net101),
    .X(_0020_));
 sg13g2_mux2_1 _1028_ (.A0(net393),
    .A1(\tt_um_mult_inst.temp_out[29] ),
    .S(net101),
    .X(_0021_));
 sg13g2_mux2_1 _1029_ (.A0(net361),
    .A1(\tt_um_mult_inst.temp_out[30] ),
    .S(net99),
    .X(_0023_));
 sg13g2_mux2_1 _1030_ (.A0(net353),
    .A1(\tt_um_mult_inst.temp_out[31] ),
    .S(net99),
    .X(_0024_));
 sg13g2_nand2_1 _1031_ (.Y(_0062_),
    .A(net8),
    .B(net430));
 sg13g2_nand2_1 _1032_ (.Y(_0063_),
    .A(net123),
    .B(net434));
 sg13g2_nand4_1 _1033_ (.B(\load_weights[12] ),
    .C(net389),
    .A(net123),
    .Y(_0064_),
    .D(net97));
 sg13g2_o21ai_1 _1034_ (.B1(_0063_),
    .Y(_0065_),
    .A1(_0048_),
    .A2(net104));
 sg13g2_nand2_1 _1035_ (.Y(_0066_),
    .A(_0064_),
    .B(_0065_));
 sg13g2_xor2_1 _1036_ (.B(_0066_),
    .A(_0062_),
    .X(\tt_um_mult_inst.temp_out_comb[8] ));
 sg13g2_o21ai_1 _1037_ (.B1(_0064_),
    .Y(_0067_),
    .A1(_0062_),
    .A2(_0066_));
 sg13g2_and2_1 _1038_ (.A(\load_weights[2] ),
    .B(\load_weights[3] ),
    .X(_0068_));
 sg13g2_nand2_2 _1039_ (.Y(_0069_),
    .A(\load_weights[2] ),
    .B(\load_weights[3] ));
 sg13g2_nor2_1 _1040_ (.A(net119),
    .B(net117),
    .Y(_0070_));
 sg13g2_xor2_1 _1041_ (.B(net118),
    .A(net119),
    .X(_0071_));
 sg13g2_nor2b_2 _1042_ (.A(\load_weights[3] ),
    .B_N(\load_weights[2] ),
    .Y(_0072_));
 sg13g2_a22oi_1 _1043_ (.Y(_0073_),
    .B1(_0072_),
    .B2(net117),
    .A2(_0071_),
    .A1(_0068_));
 sg13g2_nand2_1 _1044_ (.Y(_0074_),
    .A(\tt_um_mult_inst.temp_out[9] ),
    .B(net97));
 sg13g2_and2_2 _1045_ (.A(\load_weights[12] ),
    .B(\load_weights[13] ),
    .X(_0075_));
 sg13g2_nand2_1 _1046_ (.Y(_0076_),
    .A(\load_weights[12] ),
    .B(\load_weights[13] ));
 sg13g2_xor2_1 _1047_ (.B(net120),
    .A(net123),
    .X(_0077_));
 sg13g2_nor2b_2 _1048_ (.A(\load_weights[13] ),
    .B_N(\load_weights[12] ),
    .Y(_0078_));
 sg13g2_a22oi_1 _1049_ (.Y(_0079_),
    .B1(_0078_),
    .B2(net121),
    .A2(_0077_),
    .A1(_0075_));
 sg13g2_or2_1 _1050_ (.X(_0080_),
    .B(_0079_),
    .A(_0074_));
 sg13g2_xnor2_1 _1051_ (.Y(_0081_),
    .A(_0074_),
    .B(_0079_));
 sg13g2_xor2_1 _1052_ (.B(_0081_),
    .A(_0073_),
    .X(_0082_));
 sg13g2_nand2_1 _1053_ (.Y(_0083_),
    .A(_0067_),
    .B(_0082_));
 sg13g2_o21ai_1 _1054_ (.B1(_0080_),
    .Y(_0084_),
    .A1(_0073_),
    .A2(_0081_));
 sg13g2_nor3_1 _1055_ (.A(net119),
    .B(net117),
    .C(net115),
    .Y(_0085_));
 sg13g2_xnor2_1 _1056_ (.Y(_0086_),
    .A(net115),
    .B(_0070_));
 sg13g2_xor2_1 _1057_ (.B(_0070_),
    .A(net116),
    .X(_0087_));
 sg13g2_nand2_1 _1058_ (.Y(_0088_),
    .A(net116),
    .B(_0072_));
 sg13g2_a22oi_1 _1059_ (.Y(_0089_),
    .B1(_0086_),
    .B2(_0068_),
    .A2(_0072_),
    .A1(net116));
 sg13g2_o21ai_1 _1060_ (.B1(_0088_),
    .Y(_0090_),
    .A1(_0069_),
    .A2(_0087_));
 sg13g2_nand2_1 _1061_ (.Y(_0091_),
    .A(\tt_um_mult_inst.temp_out[10] ),
    .B(net97));
 sg13g2_or3_2 _1062_ (.A(net123),
    .B(net121),
    .C(net2),
    .X(_0092_));
 sg13g2_o21ai_1 _1063_ (.B1(net2),
    .Y(_0093_),
    .A1(net123),
    .A2(net120));
 sg13g2_nand3_1 _1064_ (.B(_0092_),
    .C(_0093_),
    .A(_0075_),
    .Y(_0094_));
 sg13g2_nand2_1 _1065_ (.Y(_0095_),
    .A(net2),
    .B(_0078_));
 sg13g2_a21oi_1 _1066_ (.A1(_0094_),
    .A2(_0095_),
    .Y(_0096_),
    .B1(_0091_));
 sg13g2_a21o_1 _1067_ (.A2(_0095_),
    .A1(_0094_),
    .B1(_0091_),
    .X(_0097_));
 sg13g2_and3_1 _1068_ (.X(_0098_),
    .A(_0091_),
    .B(_0094_),
    .C(_0095_));
 sg13g2_nand3_1 _1069_ (.B(_0094_),
    .C(_0095_),
    .A(_0091_),
    .Y(_0099_));
 sg13g2_nor3_1 _1070_ (.A(_0089_),
    .B(_0096_),
    .C(_0098_),
    .Y(_0100_));
 sg13g2_nand3_1 _1071_ (.B(_0097_),
    .C(_0099_),
    .A(_0090_),
    .Y(_0101_));
 sg13g2_a21oi_1 _1072_ (.A1(_0097_),
    .A2(_0099_),
    .Y(_0102_),
    .B1(_0090_));
 sg13g2_o21ai_1 _1073_ (.B1(_0089_),
    .Y(_0103_),
    .A1(_0096_),
    .A2(_0098_));
 sg13g2_nand3_1 _1074_ (.B(_0101_),
    .C(_0103_),
    .A(_0084_),
    .Y(_0104_));
 sg13g2_a21oi_1 _1075_ (.A1(_0101_),
    .A2(_0103_),
    .Y(_0105_),
    .B1(_0084_));
 sg13g2_nor3_1 _1076_ (.A(_0084_),
    .B(_0100_),
    .C(_0102_),
    .Y(_0106_));
 sg13g2_o21ai_1 _1077_ (.B1(_0084_),
    .Y(_0107_),
    .A1(_0100_),
    .A2(_0102_));
 sg13g2_nand2b_1 _1078_ (.Y(_0108_),
    .B(_0107_),
    .A_N(_0106_));
 sg13g2_xnor2_1 _1079_ (.Y(\tt_um_mult_inst.temp_out_comb[10] ),
    .A(_0083_),
    .B(_0108_));
 sg13g2_o21ai_1 _1080_ (.B1(_0104_),
    .Y(_0109_),
    .A1(_0083_),
    .A2(_0105_));
 sg13g2_nor2_1 _1081_ (.A(_0096_),
    .B(_0100_),
    .Y(_0110_));
 sg13g2_or4_1 _1082_ (.A(net119),
    .B(net117),
    .C(net115),
    .D(net114),
    .X(_0111_));
 sg13g2_xor2_1 _1083_ (.B(_0085_),
    .A(net114),
    .X(_0112_));
 sg13g2_nand2_1 _1084_ (.Y(_0113_),
    .A(net114),
    .B(_0072_));
 sg13g2_o21ai_1 _1085_ (.B1(_0113_),
    .Y(_0114_),
    .A1(_0069_),
    .A2(_0112_));
 sg13g2_nand2_1 _1086_ (.Y(_0115_),
    .A(\tt_um_mult_inst.temp_out[11] ),
    .B(net97));
 sg13g2_nor4_2 _1087_ (.A(net123),
    .B(net120),
    .C(net2),
    .Y(_0116_),
    .D(net3));
 sg13g2_xnor2_1 _1088_ (.Y(_0117_),
    .A(net3),
    .B(_0092_));
 sg13g2_nand2_1 _1089_ (.Y(_0118_),
    .A(net3),
    .B(_0078_));
 sg13g2_o21ai_1 _1090_ (.B1(_0118_),
    .Y(_0119_),
    .A1(_0076_),
    .A2(_0117_));
 sg13g2_nor2b_1 _1091_ (.A(_0115_),
    .B_N(_0119_),
    .Y(_0120_));
 sg13g2_xnor2_1 _1092_ (.Y(_0121_),
    .A(_0115_),
    .B(_0119_));
 sg13g2_xnor2_1 _1093_ (.Y(_0122_),
    .A(_0114_),
    .B(_0121_));
 sg13g2_nor2_1 _1094_ (.A(_0110_),
    .B(_0122_),
    .Y(_0123_));
 sg13g2_xor2_1 _1095_ (.B(_0122_),
    .A(_0110_),
    .X(_0124_));
 sg13g2_xor2_1 _1096_ (.B(_0124_),
    .A(_0109_),
    .X(\tt_um_mult_inst.temp_out_comb[11] ));
 sg13g2_a21oi_2 _1097_ (.B1(_0123_),
    .Y(_0125_),
    .A2(_0124_),
    .A1(_0109_));
 sg13g2_xnor2_1 _1098_ (.Y(_0126_),
    .A(net11),
    .B(_0111_));
 sg13g2_nand2_1 _1099_ (.Y(_0127_),
    .A(net11),
    .B(_0072_));
 sg13g2_o21ai_1 _1100_ (.B1(_0127_),
    .Y(_0128_),
    .A1(_0069_),
    .A2(_0126_));
 sg13g2_nand2_1 _1101_ (.Y(_0129_),
    .A(\tt_um_mult_inst.temp_out[12] ),
    .B(net94));
 sg13g2_xnor2_1 _1102_ (.Y(_0130_),
    .A(net4),
    .B(_0116_));
 sg13g2_a22oi_1 _1103_ (.Y(_0131_),
    .B1(_0130_),
    .B2(_0075_),
    .A2(_0078_),
    .A1(net4));
 sg13g2_nor2_1 _1104_ (.A(_0129_),
    .B(_0131_),
    .Y(_0132_));
 sg13g2_nand2_1 _1105_ (.Y(_0133_),
    .A(_0129_),
    .B(_0131_));
 sg13g2_xor2_1 _1106_ (.B(_0131_),
    .A(_0129_),
    .X(_0134_));
 sg13g2_xnor2_1 _1107_ (.Y(_0135_),
    .A(_0128_),
    .B(_0134_));
 sg13g2_a21oi_2 _1108_ (.B1(_0120_),
    .Y(_0136_),
    .A2(_0121_),
    .A1(_0114_));
 sg13g2_nor2_1 _1109_ (.A(_0135_),
    .B(_0136_),
    .Y(_0137_));
 sg13g2_xnor2_1 _1110_ (.Y(_0138_),
    .A(_0135_),
    .B(_0136_));
 sg13g2_nor2_1 _1111_ (.A(_0125_),
    .B(_0138_),
    .Y(_0139_));
 sg13g2_xor2_1 _1112_ (.B(_0138_),
    .A(_0125_),
    .X(\tt_um_mult_inst.temp_out_comb[12] ));
 sg13g2_nor3_1 _1113_ (.A(net113),
    .B(net112),
    .C(_0111_),
    .Y(_0140_));
 sg13g2_o21ai_1 _1114_ (.B1(net112),
    .Y(_0141_),
    .A1(net113),
    .A2(_0111_));
 sg13g2_nand2b_2 _1115_ (.Y(_0142_),
    .B(_0141_),
    .A_N(_0140_));
 sg13g2_nand2_1 _1116_ (.Y(_0143_),
    .A(net112),
    .B(_0072_));
 sg13g2_o21ai_1 _1117_ (.B1(_0143_),
    .Y(_0144_),
    .A1(_0069_),
    .A2(_0142_));
 sg13g2_nand2_1 _1118_ (.Y(_0145_),
    .A(\tt_um_mult_inst.temp_out[13] ),
    .B(net94));
 sg13g2_nand3_1 _1119_ (.B(_0052_),
    .C(_0116_),
    .A(_0051_),
    .Y(_0146_));
 sg13g2_a21o_2 _1120_ (.A2(_0116_),
    .A1(_0051_),
    .B1(_0052_),
    .X(_0147_));
 sg13g2_nand3_1 _1121_ (.B(_0146_),
    .C(_0147_),
    .A(_0075_),
    .Y(_0148_));
 sg13g2_nand2_1 _1122_ (.Y(_0149_),
    .A(net5),
    .B(_0078_));
 sg13g2_a21oi_1 _1123_ (.A1(_0148_),
    .A2(_0149_),
    .Y(_0150_),
    .B1(_0145_));
 sg13g2_a21o_1 _1124_ (.A2(_0149_),
    .A1(_0148_),
    .B1(_0145_),
    .X(_0151_));
 sg13g2_nand3_1 _1125_ (.B(_0148_),
    .C(_0149_),
    .A(_0145_),
    .Y(_0152_));
 sg13g2_a21oi_1 _1126_ (.A1(_0151_),
    .A2(_0152_),
    .Y(_0153_),
    .B1(_0144_));
 sg13g2_and3_1 _1127_ (.X(_0154_),
    .A(_0144_),
    .B(_0151_),
    .C(_0152_));
 sg13g2_a21oi_1 _1128_ (.A1(_0128_),
    .A2(_0133_),
    .Y(_0155_),
    .B1(_0132_));
 sg13g2_nor3_1 _1129_ (.A(_0153_),
    .B(_0154_),
    .C(_0155_),
    .Y(_0156_));
 sg13g2_or3_1 _1130_ (.A(_0153_),
    .B(_0154_),
    .C(_0155_),
    .X(_0157_));
 sg13g2_o21ai_1 _1131_ (.B1(_0155_),
    .Y(_0158_),
    .A1(_0153_),
    .A2(_0154_));
 sg13g2_nand2_1 _1132_ (.Y(_0159_),
    .A(_0157_),
    .B(_0158_));
 sg13g2_nor2_1 _1133_ (.A(_0137_),
    .B(_0139_),
    .Y(_0160_));
 sg13g2_xor2_1 _1134_ (.B(_0160_),
    .A(_0159_),
    .X(\tt_um_mult_inst.temp_out_comb[13] ));
 sg13g2_nand3b_1 _1135_ (.B(_0157_),
    .C(_0158_),
    .Y(_0161_),
    .A_N(_0138_));
 sg13g2_o21ai_1 _1136_ (.B1(_0158_),
    .Y(_0162_),
    .A1(_0137_),
    .A2(_0156_));
 sg13g2_o21ai_1 _1137_ (.B1(_0162_),
    .Y(_0163_),
    .A1(_0125_),
    .A2(_0161_));
 sg13g2_nor2_1 _1138_ (.A(_0150_),
    .B(_0154_),
    .Y(_0164_));
 sg13g2_nor2b_1 _1139_ (.A(net13),
    .B_N(_0140_),
    .Y(_0165_));
 sg13g2_xnor2_1 _1140_ (.Y(_0166_),
    .A(net111),
    .B(_0140_));
 sg13g2_a22oi_1 _1141_ (.Y(_0167_),
    .B1(_0166_),
    .B2(_0068_),
    .A2(_0072_),
    .A1(net111));
 sg13g2_nand2_1 _1142_ (.Y(_0168_),
    .A(\tt_um_mult_inst.temp_out[14] ),
    .B(net93));
 sg13g2_nor2_1 _1143_ (.A(net6),
    .B(_0146_),
    .Y(_0169_));
 sg13g2_xor2_1 _1144_ (.B(_0146_),
    .A(net6),
    .X(_0170_));
 sg13g2_a22oi_1 _1145_ (.Y(_0171_),
    .B1(_0170_),
    .B2(_0075_),
    .A2(_0078_),
    .A1(net6));
 sg13g2_or2_1 _1146_ (.X(_0172_),
    .B(_0171_),
    .A(_0168_));
 sg13g2_xnor2_1 _1147_ (.Y(_0173_),
    .A(_0168_),
    .B(_0171_));
 sg13g2_xnor2_1 _1148_ (.Y(_0174_),
    .A(_0167_),
    .B(_0173_));
 sg13g2_nor2_1 _1149_ (.A(_0164_),
    .B(_0174_),
    .Y(_0175_));
 sg13g2_xor2_1 _1150_ (.B(_0174_),
    .A(_0164_),
    .X(_0176_));
 sg13g2_xor2_1 _1151_ (.B(_0176_),
    .A(_0163_),
    .X(\tt_um_mult_inst.temp_out_comb[14] ));
 sg13g2_a21oi_1 _1152_ (.A1(_0163_),
    .A2(_0176_),
    .Y(_0177_),
    .B1(_0175_));
 sg13g2_o21ai_1 _1153_ (.B1(_0172_),
    .Y(_0178_),
    .A1(_0167_),
    .A2(_0173_));
 sg13g2_nand2_1 _1154_ (.Y(_0179_),
    .A(net443),
    .B(net93));
 sg13g2_xnor2_1 _1155_ (.Y(_0180_),
    .A(net7),
    .B(_0169_));
 sg13g2_a22oi_1 _1156_ (.Y(_0181_),
    .B1(_0180_),
    .B2(_0075_),
    .A2(_0078_),
    .A1(net7));
 sg13g2_xnor2_1 _1157_ (.Y(_0182_),
    .A(net14),
    .B(_0165_));
 sg13g2_a22oi_1 _1158_ (.Y(_0183_),
    .B1(_0182_),
    .B2(_0068_),
    .A2(_0072_),
    .A1(net14));
 sg13g2_xnor2_1 _1159_ (.Y(_0184_),
    .A(_0181_),
    .B(_0183_));
 sg13g2_xnor2_1 _1160_ (.Y(_0185_),
    .A(_0179_),
    .B(_0184_));
 sg13g2_xnor2_1 _1161_ (.Y(_0186_),
    .A(_0178_),
    .B(_0185_));
 sg13g2_xnor2_1 _1162_ (.Y(\tt_um_mult_inst.temp_out_comb[15] ),
    .A(_0177_),
    .B(_0186_));
 sg13g2_xor2_1 _1163_ (.B(_0082_),
    .A(_0067_),
    .X(\tt_um_mult_inst.temp_out_comb[9] ));
 sg13g2_nand2_1 _1164_ (.Y(_0187_),
    .A(net8),
    .B(net431));
 sg13g2_nand2_1 _1165_ (.Y(_0188_),
    .A(net123),
    .B(\load_weights[10] ));
 sg13g2_nand4_1 _1166_ (.B(\load_weights[10] ),
    .C(net444),
    .A(net123),
    .Y(_0189_),
    .D(net98));
 sg13g2_o21ai_1 _1167_ (.B1(_0188_),
    .Y(_0190_),
    .A1(_0047_),
    .A2(net105));
 sg13g2_nand2_1 _1168_ (.Y(_0191_),
    .A(_0189_),
    .B(_0190_));
 sg13g2_xor2_1 _1169_ (.B(_0191_),
    .A(_0187_),
    .X(\tt_um_mult_inst.temp_out_comb[0] ));
 sg13g2_o21ai_1 _1170_ (.B1(_0189_),
    .Y(_0192_),
    .A1(_0187_),
    .A2(_0191_));
 sg13g2_and2_1 _1171_ (.A(\load_weights[0] ),
    .B(\load_weights[1] ),
    .X(_0193_));
 sg13g2_nand2_2 _1172_ (.Y(_0194_),
    .A(\load_weights[0] ),
    .B(\load_weights[1] ));
 sg13g2_nor2b_2 _1173_ (.A(\load_weights[1] ),
    .B_N(\load_weights[0] ),
    .Y(_0195_));
 sg13g2_a22oi_1 _1174_ (.Y(_0196_),
    .B1(_0195_),
    .B2(net118),
    .A2(_0193_),
    .A1(_0071_));
 sg13g2_nand2_1 _1175_ (.Y(_0197_),
    .A(\tt_um_mult_inst.temp_out[1] ),
    .B(net97));
 sg13g2_and2_2 _1176_ (.A(\load_weights[10] ),
    .B(\load_weights[11] ),
    .X(_0198_));
 sg13g2_nand2_1 _1177_ (.Y(_0199_),
    .A(\load_weights[10] ),
    .B(\load_weights[11] ));
 sg13g2_nor2b_2 _1178_ (.A(\load_weights[11] ),
    .B_N(\load_weights[10] ),
    .Y(_0200_));
 sg13g2_a22oi_1 _1179_ (.Y(_0201_),
    .B1(_0200_),
    .B2(net120),
    .A2(_0198_),
    .A1(_0077_));
 sg13g2_or2_1 _1180_ (.X(_0202_),
    .B(_0201_),
    .A(_0197_));
 sg13g2_xnor2_1 _1181_ (.Y(_0203_),
    .A(_0197_),
    .B(_0201_));
 sg13g2_xor2_1 _1182_ (.B(_0203_),
    .A(_0196_),
    .X(_0204_));
 sg13g2_nand2_1 _1183_ (.Y(_0205_),
    .A(_0192_),
    .B(_0204_));
 sg13g2_o21ai_1 _1184_ (.B1(_0202_),
    .Y(_0206_),
    .A1(_0196_),
    .A2(_0203_));
 sg13g2_nand2_1 _1185_ (.Y(_0207_),
    .A(net116),
    .B(_0195_));
 sg13g2_a22oi_1 _1186_ (.Y(_0208_),
    .B1(_0195_),
    .B2(net116),
    .A2(_0193_),
    .A1(_0086_));
 sg13g2_o21ai_1 _1187_ (.B1(_0207_),
    .Y(_0209_),
    .A1(_0087_),
    .A2(_0194_));
 sg13g2_nand2_1 _1188_ (.Y(_0210_),
    .A(\tt_um_mult_inst.temp_out[2] ),
    .B(net97));
 sg13g2_nand3_1 _1189_ (.B(_0093_),
    .C(_0198_),
    .A(_0092_),
    .Y(_0211_));
 sg13g2_nand2_1 _1190_ (.Y(_0212_),
    .A(net2),
    .B(_0200_));
 sg13g2_a21oi_1 _1191_ (.A1(_0211_),
    .A2(_0212_),
    .Y(_0213_),
    .B1(_0210_));
 sg13g2_a21o_1 _1192_ (.A2(_0212_),
    .A1(_0211_),
    .B1(_0210_),
    .X(_0214_));
 sg13g2_and3_1 _1193_ (.X(_0215_),
    .A(_0210_),
    .B(_0211_),
    .C(_0212_));
 sg13g2_nand3_1 _1194_ (.B(_0211_),
    .C(_0212_),
    .A(_0210_),
    .Y(_0216_));
 sg13g2_nor3_1 _1195_ (.A(_0208_),
    .B(_0213_),
    .C(_0215_),
    .Y(_0217_));
 sg13g2_nand3_1 _1196_ (.B(_0214_),
    .C(_0216_),
    .A(_0209_),
    .Y(_0218_));
 sg13g2_a21oi_1 _1197_ (.A1(_0214_),
    .A2(_0216_),
    .Y(_0219_),
    .B1(_0209_));
 sg13g2_o21ai_1 _1198_ (.B1(_0208_),
    .Y(_0220_),
    .A1(_0213_),
    .A2(_0215_));
 sg13g2_nand3_1 _1199_ (.B(_0218_),
    .C(_0220_),
    .A(_0206_),
    .Y(_0221_));
 sg13g2_a21oi_1 _1200_ (.A1(_0218_),
    .A2(_0220_),
    .Y(_0222_),
    .B1(_0206_));
 sg13g2_nor3_1 _1201_ (.A(_0206_),
    .B(_0217_),
    .C(_0219_),
    .Y(_0223_));
 sg13g2_o21ai_1 _1202_ (.B1(_0206_),
    .Y(_0224_),
    .A1(_0217_),
    .A2(_0219_));
 sg13g2_nand2b_1 _1203_ (.Y(_0225_),
    .B(_0224_),
    .A_N(_0223_));
 sg13g2_xnor2_1 _1204_ (.Y(\tt_um_mult_inst.temp_out_comb[2] ),
    .A(_0205_),
    .B(_0225_));
 sg13g2_o21ai_1 _1205_ (.B1(_0221_),
    .Y(_0226_),
    .A1(_0205_),
    .A2(_0222_));
 sg13g2_nor2_1 _1206_ (.A(_0213_),
    .B(_0217_),
    .Y(_0227_));
 sg13g2_nand2_1 _1207_ (.Y(_0228_),
    .A(net114),
    .B(_0195_));
 sg13g2_o21ai_1 _1208_ (.B1(_0228_),
    .Y(_0229_),
    .A1(_0112_),
    .A2(_0194_));
 sg13g2_nand2_1 _1209_ (.Y(_0230_),
    .A(\tt_um_mult_inst.temp_out[3] ),
    .B(net97));
 sg13g2_nand2_1 _1210_ (.Y(_0231_),
    .A(net3),
    .B(_0200_));
 sg13g2_o21ai_1 _1211_ (.B1(_0231_),
    .Y(_0232_),
    .A1(_0117_),
    .A2(_0199_));
 sg13g2_nor2b_1 _1212_ (.A(_0230_),
    .B_N(_0232_),
    .Y(_0233_));
 sg13g2_xnor2_1 _1213_ (.Y(_0234_),
    .A(_0230_),
    .B(_0232_));
 sg13g2_xnor2_1 _1214_ (.Y(_0235_),
    .A(_0229_),
    .B(_0234_));
 sg13g2_nor2_1 _1215_ (.A(_0227_),
    .B(_0235_),
    .Y(_0236_));
 sg13g2_xor2_1 _1216_ (.B(_0235_),
    .A(_0227_),
    .X(_0237_));
 sg13g2_xor2_1 _1217_ (.B(_0237_),
    .A(_0226_),
    .X(\tt_um_mult_inst.temp_out_comb[3] ));
 sg13g2_a21oi_2 _1218_ (.B1(_0236_),
    .Y(_0238_),
    .A2(_0237_),
    .A1(_0226_));
 sg13g2_nand2_1 _1219_ (.Y(_0239_),
    .A(net113),
    .B(_0195_));
 sg13g2_o21ai_1 _1220_ (.B1(_0239_),
    .Y(_0240_),
    .A1(_0126_),
    .A2(_0194_));
 sg13g2_nand2_1 _1221_ (.Y(_0241_),
    .A(\tt_um_mult_inst.temp_out[4] ),
    .B(net94));
 sg13g2_a22oi_1 _1222_ (.Y(_0242_),
    .B1(_0200_),
    .B2(net4),
    .A2(_0198_),
    .A1(_0130_));
 sg13g2_nor2_1 _1223_ (.A(_0241_),
    .B(_0242_),
    .Y(_0243_));
 sg13g2_nand2_1 _1224_ (.Y(_0244_),
    .A(_0241_),
    .B(_0242_));
 sg13g2_xor2_1 _1225_ (.B(_0242_),
    .A(_0241_),
    .X(_0245_));
 sg13g2_xnor2_1 _1226_ (.Y(_0246_),
    .A(_0240_),
    .B(_0245_));
 sg13g2_a21oi_1 _1227_ (.A1(_0229_),
    .A2(_0234_),
    .Y(_0247_),
    .B1(_0233_));
 sg13g2_nor2_1 _1228_ (.A(_0246_),
    .B(_0247_),
    .Y(_0248_));
 sg13g2_xnor2_1 _1229_ (.Y(_0249_),
    .A(_0246_),
    .B(_0247_));
 sg13g2_nor2_1 _1230_ (.A(_0238_),
    .B(_0249_),
    .Y(_0250_));
 sg13g2_xor2_1 _1231_ (.B(_0249_),
    .A(_0238_),
    .X(\tt_um_mult_inst.temp_out_comb[4] ));
 sg13g2_nand2_1 _1232_ (.Y(_0251_),
    .A(net112),
    .B(_0195_));
 sg13g2_o21ai_1 _1233_ (.B1(_0251_),
    .Y(_0252_),
    .A1(_0142_),
    .A2(_0194_));
 sg13g2_nand2_1 _1234_ (.Y(_0253_),
    .A(\tt_um_mult_inst.temp_out[5] ),
    .B(net94));
 sg13g2_nand3_1 _1235_ (.B(_0147_),
    .C(_0198_),
    .A(_0146_),
    .Y(_0254_));
 sg13g2_nand2_1 _1236_ (.Y(_0255_),
    .A(net5),
    .B(_0200_));
 sg13g2_a21oi_1 _1237_ (.A1(_0254_),
    .A2(_0255_),
    .Y(_0256_),
    .B1(_0253_));
 sg13g2_a21o_1 _1238_ (.A2(_0255_),
    .A1(_0254_),
    .B1(_0253_),
    .X(_0257_));
 sg13g2_nand3_1 _1239_ (.B(_0254_),
    .C(_0255_),
    .A(_0253_),
    .Y(_0258_));
 sg13g2_a21oi_1 _1240_ (.A1(_0257_),
    .A2(_0258_),
    .Y(_0259_),
    .B1(_0252_));
 sg13g2_and3_1 _1241_ (.X(_0260_),
    .A(_0252_),
    .B(_0257_),
    .C(_0258_));
 sg13g2_a21oi_1 _1242_ (.A1(_0240_),
    .A2(_0244_),
    .Y(_0261_),
    .B1(_0243_));
 sg13g2_nor3_1 _1243_ (.A(_0259_),
    .B(_0260_),
    .C(_0261_),
    .Y(_0262_));
 sg13g2_or3_1 _1244_ (.A(_0259_),
    .B(_0260_),
    .C(_0261_),
    .X(_0263_));
 sg13g2_o21ai_1 _1245_ (.B1(_0261_),
    .Y(_0264_),
    .A1(_0259_),
    .A2(_0260_));
 sg13g2_nand2_1 _1246_ (.Y(_0265_),
    .A(_0263_),
    .B(_0264_));
 sg13g2_nor2_1 _1247_ (.A(_0248_),
    .B(_0250_),
    .Y(_0266_));
 sg13g2_xor2_1 _1248_ (.B(_0266_),
    .A(_0265_),
    .X(\tt_um_mult_inst.temp_out_comb[5] ));
 sg13g2_nand3b_1 _1249_ (.B(_0263_),
    .C(_0264_),
    .Y(_0267_),
    .A_N(_0249_));
 sg13g2_o21ai_1 _1250_ (.B1(_0264_),
    .Y(_0268_),
    .A1(_0248_),
    .A2(_0262_));
 sg13g2_o21ai_1 _1251_ (.B1(_0268_),
    .Y(_0269_),
    .A1(_0238_),
    .A2(_0267_));
 sg13g2_nor2_1 _1252_ (.A(_0256_),
    .B(_0260_),
    .Y(_0270_));
 sg13g2_a22oi_1 _1253_ (.Y(_0271_),
    .B1(_0195_),
    .B2(net111),
    .A2(_0193_),
    .A1(_0166_));
 sg13g2_nand2_1 _1254_ (.Y(_0272_),
    .A(\tt_um_mult_inst.temp_out[6] ),
    .B(net94));
 sg13g2_a22oi_1 _1255_ (.Y(_0273_),
    .B1(_0200_),
    .B2(net6),
    .A2(_0198_),
    .A1(_0170_));
 sg13g2_or2_1 _1256_ (.X(_0274_),
    .B(_0273_),
    .A(_0272_));
 sg13g2_xnor2_1 _1257_ (.Y(_0275_),
    .A(_0272_),
    .B(_0273_));
 sg13g2_xnor2_1 _1258_ (.Y(_0276_),
    .A(_0271_),
    .B(_0275_));
 sg13g2_nor2_1 _1259_ (.A(_0270_),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_xor2_1 _1260_ (.B(_0276_),
    .A(_0270_),
    .X(_0278_));
 sg13g2_xor2_1 _1261_ (.B(_0278_),
    .A(_0269_),
    .X(\tt_um_mult_inst.temp_out_comb[6] ));
 sg13g2_a21oi_1 _1262_ (.A1(_0269_),
    .A2(_0278_),
    .Y(_0279_),
    .B1(_0277_));
 sg13g2_o21ai_1 _1263_ (.B1(_0274_),
    .Y(_0280_),
    .A1(_0271_),
    .A2(_0275_));
 sg13g2_nand2_1 _1264_ (.Y(_0281_),
    .A(\tt_um_mult_inst.temp_out[7] ),
    .B(net94));
 sg13g2_a22oi_1 _1265_ (.Y(_0282_),
    .B1(_0200_),
    .B2(net7),
    .A2(_0198_),
    .A1(_0180_));
 sg13g2_a22oi_1 _1266_ (.Y(_0283_),
    .B1(_0195_),
    .B2(net14),
    .A2(_0193_),
    .A1(_0182_));
 sg13g2_xnor2_1 _1267_ (.Y(_0284_),
    .A(_0282_),
    .B(_0283_));
 sg13g2_xnor2_1 _1268_ (.Y(_0285_),
    .A(_0281_),
    .B(_0284_));
 sg13g2_xnor2_1 _1269_ (.Y(_0286_),
    .A(_0280_),
    .B(_0285_));
 sg13g2_xnor2_1 _1270_ (.Y(\tt_um_mult_inst.temp_out_comb[7] ),
    .A(_0279_),
    .B(_0286_));
 sg13g2_xor2_1 _1271_ (.B(_0204_),
    .A(_0192_),
    .X(\tt_um_mult_inst.temp_out_comb[1] ));
 sg13g2_nand2_1 _1272_ (.Y(_0287_),
    .A(net119),
    .B(net433));
 sg13g2_nand2_1 _1273_ (.Y(_0288_),
    .A(net122),
    .B(\load_weights[16] ));
 sg13g2_nand4_1 _1274_ (.B(\load_weights[16] ),
    .C(net438),
    .A(net122),
    .Y(_0289_),
    .D(net96));
 sg13g2_o21ai_1 _1275_ (.B1(_0288_),
    .Y(_0290_),
    .A1(_0050_),
    .A2(net103));
 sg13g2_nand2_1 _1276_ (.Y(_0291_),
    .A(_0289_),
    .B(_0290_));
 sg13g2_xor2_1 _1277_ (.B(_0291_),
    .A(_0287_),
    .X(\tt_um_mult_inst.temp_out_comb[24] ));
 sg13g2_o21ai_1 _1278_ (.B1(_0289_),
    .Y(_0292_),
    .A1(_0287_),
    .A2(_0291_));
 sg13g2_and2_1 _1279_ (.A(\load_weights[6] ),
    .B(\load_weights[7] ),
    .X(_0293_));
 sg13g2_nand2_2 _1280_ (.Y(_0294_),
    .A(\load_weights[6] ),
    .B(\load_weights[7] ));
 sg13g2_nor2b_2 _1281_ (.A(\load_weights[7] ),
    .B_N(\load_weights[6] ),
    .Y(_0295_));
 sg13g2_a22oi_1 _1282_ (.Y(_0296_),
    .B1(_0295_),
    .B2(net117),
    .A2(_0293_),
    .A1(_0071_));
 sg13g2_nand2_1 _1283_ (.Y(_0297_),
    .A(\tt_um_mult_inst.temp_out[25] ),
    .B(net98));
 sg13g2_and2_2 _1284_ (.A(\load_weights[16] ),
    .B(\load_weights[17] ),
    .X(_0298_));
 sg13g2_nand2_1 _1285_ (.Y(_0299_),
    .A(\load_weights[16] ),
    .B(\load_weights[17] ));
 sg13g2_nor2b_2 _1286_ (.A(\load_weights[17] ),
    .B_N(\load_weights[16] ),
    .Y(_0300_));
 sg13g2_a22oi_1 _1287_ (.Y(_0301_),
    .B1(_0300_),
    .B2(net120),
    .A2(_0298_),
    .A1(_0077_));
 sg13g2_or2_1 _1288_ (.X(_0302_),
    .B(_0301_),
    .A(_0297_));
 sg13g2_xnor2_1 _1289_ (.Y(_0303_),
    .A(_0297_),
    .B(_0301_));
 sg13g2_xor2_1 _1290_ (.B(_0303_),
    .A(_0296_),
    .X(_0304_));
 sg13g2_nand2_1 _1291_ (.Y(_0305_),
    .A(_0292_),
    .B(_0304_));
 sg13g2_xor2_1 _1292_ (.B(_0304_),
    .A(_0292_),
    .X(\tt_um_mult_inst.temp_out_comb[25] ));
 sg13g2_o21ai_1 _1293_ (.B1(_0302_),
    .Y(_0306_),
    .A1(_0296_),
    .A2(_0303_));
 sg13g2_nand2_1 _1294_ (.Y(_0307_),
    .A(net115),
    .B(_0295_));
 sg13g2_a22oi_1 _1295_ (.Y(_0308_),
    .B1(_0295_),
    .B2(net115),
    .A2(_0293_),
    .A1(_0086_));
 sg13g2_o21ai_1 _1296_ (.B1(_0307_),
    .Y(_0309_),
    .A1(_0087_),
    .A2(_0294_));
 sg13g2_nand2_2 _1297_ (.Y(_0310_),
    .A(\tt_um_mult_inst.temp_out[26] ),
    .B(net96));
 sg13g2_nand3_1 _1298_ (.B(_0093_),
    .C(_0298_),
    .A(_0092_),
    .Y(_0311_));
 sg13g2_nand2_2 _1299_ (.Y(_0312_),
    .A(net2),
    .B(_0300_));
 sg13g2_a21oi_2 _1300_ (.B1(_0310_),
    .Y(_0313_),
    .A2(_0312_),
    .A1(_0311_));
 sg13g2_a21o_1 _1301_ (.A2(_0312_),
    .A1(_0311_),
    .B1(_0310_),
    .X(_0314_));
 sg13g2_and3_1 _1302_ (.X(_0315_),
    .A(_0310_),
    .B(_0311_),
    .C(_0312_));
 sg13g2_nand3_1 _1303_ (.B(_0311_),
    .C(_0312_),
    .A(_0310_),
    .Y(_0316_));
 sg13g2_nor3_2 _1304_ (.A(_0308_),
    .B(_0313_),
    .C(_0315_),
    .Y(_0317_));
 sg13g2_nand3_1 _1305_ (.B(_0314_),
    .C(_0316_),
    .A(_0309_),
    .Y(_0318_));
 sg13g2_a21oi_1 _1306_ (.A1(_0314_),
    .A2(_0316_),
    .Y(_0319_),
    .B1(_0309_));
 sg13g2_o21ai_1 _1307_ (.B1(_0308_),
    .Y(_0320_),
    .A1(_0313_),
    .A2(_0315_));
 sg13g2_nand3_1 _1308_ (.B(_0318_),
    .C(_0320_),
    .A(_0306_),
    .Y(_0321_));
 sg13g2_a21oi_1 _1309_ (.A1(_0318_),
    .A2(_0320_),
    .Y(_0322_),
    .B1(_0306_));
 sg13g2_nor3_1 _1310_ (.A(_0306_),
    .B(_0317_),
    .C(_0319_),
    .Y(_0323_));
 sg13g2_o21ai_1 _1311_ (.B1(_0306_),
    .Y(_0324_),
    .A1(_0317_),
    .A2(_0319_));
 sg13g2_nand2b_1 _1312_ (.Y(_0325_),
    .B(_0324_),
    .A_N(_0323_));
 sg13g2_xnor2_1 _1313_ (.Y(\tt_um_mult_inst.temp_out_comb[26] ),
    .A(_0305_),
    .B(_0325_));
 sg13g2_o21ai_1 _1314_ (.B1(_0321_),
    .Y(_0326_),
    .A1(_0305_),
    .A2(_0322_));
 sg13g2_nor2_1 _1315_ (.A(_0313_),
    .B(_0317_),
    .Y(_0327_));
 sg13g2_nand2_1 _1316_ (.Y(_0328_),
    .A(net114),
    .B(_0295_));
 sg13g2_o21ai_1 _1317_ (.B1(_0328_),
    .Y(_0329_),
    .A1(_0112_),
    .A2(_0294_));
 sg13g2_nand2_1 _1318_ (.Y(_0330_),
    .A(\tt_um_mult_inst.temp_out[27] ),
    .B(net96));
 sg13g2_nand2_1 _1319_ (.Y(_0331_),
    .A(net3),
    .B(_0300_));
 sg13g2_o21ai_1 _1320_ (.B1(_0331_),
    .Y(_0332_),
    .A1(_0117_),
    .A2(_0299_));
 sg13g2_nor2b_1 _1321_ (.A(_0330_),
    .B_N(_0332_),
    .Y(_0333_));
 sg13g2_xnor2_1 _1322_ (.Y(_0334_),
    .A(_0330_),
    .B(_0332_));
 sg13g2_xnor2_1 _1323_ (.Y(_0335_),
    .A(_0329_),
    .B(_0334_));
 sg13g2_nor2_1 _1324_ (.A(_0327_),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_xor2_1 _1325_ (.B(_0335_),
    .A(_0327_),
    .X(_0337_));
 sg13g2_xor2_1 _1326_ (.B(_0337_),
    .A(_0326_),
    .X(\tt_um_mult_inst.temp_out_comb[27] ));
 sg13g2_a21oi_2 _1327_ (.B1(_0336_),
    .Y(_0338_),
    .A2(_0337_),
    .A1(_0326_));
 sg13g2_nand2_1 _1328_ (.Y(_0339_),
    .A(net113),
    .B(_0295_));
 sg13g2_o21ai_1 _1329_ (.B1(_0339_),
    .Y(_0340_),
    .A1(_0126_),
    .A2(_0294_));
 sg13g2_nand2_1 _1330_ (.Y(_0341_),
    .A(\tt_um_mult_inst.temp_out[28] ),
    .B(net95));
 sg13g2_a22oi_1 _1331_ (.Y(_0342_),
    .B1(_0300_),
    .B2(net4),
    .A2(_0298_),
    .A1(_0130_));
 sg13g2_nor2_1 _1332_ (.A(_0341_),
    .B(_0342_),
    .Y(_0343_));
 sg13g2_nand2_1 _1333_ (.Y(_0344_),
    .A(_0341_),
    .B(_0342_));
 sg13g2_xor2_1 _1334_ (.B(_0342_),
    .A(_0341_),
    .X(_0345_));
 sg13g2_xnor2_1 _1335_ (.Y(_0346_),
    .A(_0340_),
    .B(_0345_));
 sg13g2_a21oi_2 _1336_ (.B1(_0333_),
    .Y(_0347_),
    .A2(_0334_),
    .A1(_0329_));
 sg13g2_nor2_1 _1337_ (.A(_0346_),
    .B(_0347_),
    .Y(_0348_));
 sg13g2_xor2_1 _1338_ (.B(_0347_),
    .A(_0346_),
    .X(_0349_));
 sg13g2_nor2b_1 _1339_ (.A(_0338_),
    .B_N(_0349_),
    .Y(_0350_));
 sg13g2_xnor2_1 _1340_ (.Y(\tt_um_mult_inst.temp_out_comb[28] ),
    .A(_0338_),
    .B(_0349_));
 sg13g2_a21oi_1 _1341_ (.A1(_0340_),
    .A2(_0344_),
    .Y(_0351_),
    .B1(_0343_));
 sg13g2_nand2_1 _1342_ (.Y(_0352_),
    .A(net112),
    .B(_0295_));
 sg13g2_o21ai_1 _1343_ (.B1(_0352_),
    .Y(_0353_),
    .A1(_0142_),
    .A2(_0294_));
 sg13g2_nand2_1 _1344_ (.Y(_0354_),
    .A(\tt_um_mult_inst.temp_out[29] ),
    .B(net95));
 sg13g2_nand3_1 _1345_ (.B(_0147_),
    .C(_0298_),
    .A(_0146_),
    .Y(_0355_));
 sg13g2_nand2_1 _1346_ (.Y(_0356_),
    .A(net5),
    .B(_0300_));
 sg13g2_a21oi_1 _1347_ (.A1(_0355_),
    .A2(_0356_),
    .Y(_0357_),
    .B1(_0354_));
 sg13g2_a21o_1 _1348_ (.A2(_0356_),
    .A1(_0355_),
    .B1(_0354_),
    .X(_0358_));
 sg13g2_nand3_1 _1349_ (.B(_0355_),
    .C(_0356_),
    .A(_0354_),
    .Y(_0359_));
 sg13g2_and3_1 _1350_ (.X(_0360_),
    .A(_0353_),
    .B(_0358_),
    .C(_0359_));
 sg13g2_a21oi_1 _1351_ (.A1(_0358_),
    .A2(_0359_),
    .Y(_0361_),
    .B1(_0353_));
 sg13g2_o21ai_1 _1352_ (.B1(_0351_),
    .Y(_0362_),
    .A1(_0360_),
    .A2(_0361_));
 sg13g2_nor3_1 _1353_ (.A(_0351_),
    .B(_0360_),
    .C(_0361_),
    .Y(_0363_));
 sg13g2_or3_1 _1354_ (.A(_0351_),
    .B(_0360_),
    .C(_0361_),
    .X(_0364_));
 sg13g2_and2_1 _1355_ (.A(_0362_),
    .B(_0364_),
    .X(_0365_));
 sg13g2_nor2_1 _1356_ (.A(_0348_),
    .B(_0350_),
    .Y(_0366_));
 sg13g2_xnor2_1 _1357_ (.Y(\tt_um_mult_inst.temp_out_comb[29] ),
    .A(_0365_),
    .B(_0366_));
 sg13g2_nand3b_1 _1358_ (.B(_0349_),
    .C(_0362_),
    .Y(_0367_),
    .A_N(_0363_));
 sg13g2_a21oi_1 _1359_ (.A1(_0348_),
    .A2(_0362_),
    .Y(_0368_),
    .B1(_0363_));
 sg13g2_o21ai_1 _1360_ (.B1(_0368_),
    .Y(_0369_),
    .A1(_0338_),
    .A2(_0367_));
 sg13g2_nor2_1 _1361_ (.A(_0357_),
    .B(_0360_),
    .Y(_0370_));
 sg13g2_a22oi_1 _1362_ (.Y(_0371_),
    .B1(_0295_),
    .B2(net111),
    .A2(_0293_),
    .A1(_0166_));
 sg13g2_nand2_1 _1363_ (.Y(_0372_),
    .A(\tt_um_mult_inst.temp_out[30] ),
    .B(net93));
 sg13g2_a22oi_1 _1364_ (.Y(_0373_),
    .B1(_0300_),
    .B2(net6),
    .A2(_0298_),
    .A1(_0170_));
 sg13g2_or2_1 _1365_ (.X(_0374_),
    .B(_0373_),
    .A(_0372_));
 sg13g2_xnor2_1 _1366_ (.Y(_0375_),
    .A(_0372_),
    .B(_0373_));
 sg13g2_xnor2_1 _1367_ (.Y(_0376_),
    .A(_0371_),
    .B(_0375_));
 sg13g2_nor2_1 _1368_ (.A(_0370_),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_xor2_1 _1369_ (.B(_0376_),
    .A(_0370_),
    .X(_0378_));
 sg13g2_xor2_1 _1370_ (.B(_0378_),
    .A(_0369_),
    .X(\tt_um_mult_inst.temp_out_comb[30] ));
 sg13g2_a21oi_1 _1371_ (.A1(_0369_),
    .A2(_0378_),
    .Y(_0379_),
    .B1(_0377_));
 sg13g2_o21ai_1 _1372_ (.B1(_0374_),
    .Y(_0380_),
    .A1(_0371_),
    .A2(_0375_));
 sg13g2_nand2_1 _1373_ (.Y(_0381_),
    .A(\tt_um_mult_inst.temp_out[31] ),
    .B(net93));
 sg13g2_a22oi_1 _1374_ (.Y(_0382_),
    .B1(_0300_),
    .B2(net7),
    .A2(_0298_),
    .A1(_0180_));
 sg13g2_a22oi_1 _1375_ (.Y(_0383_),
    .B1(_0295_),
    .B2(net14),
    .A2(_0293_),
    .A1(_0182_));
 sg13g2_xnor2_1 _1376_ (.Y(_0384_),
    .A(_0382_),
    .B(_0383_));
 sg13g2_xnor2_1 _1377_ (.Y(_0385_),
    .A(_0381_),
    .B(_0384_));
 sg13g2_xnor2_1 _1378_ (.Y(_0386_),
    .A(_0380_),
    .B(_0385_));
 sg13g2_xnor2_1 _1379_ (.Y(\tt_um_mult_inst.temp_out_comb[31] ),
    .A(_0379_),
    .B(_0386_));
 sg13g2_nand2_1 _1380_ (.Y(_0387_),
    .A(net119),
    .B(net414));
 sg13g2_nand2_1 _1381_ (.Y(_0388_),
    .A(net122),
    .B(\load_weights[18] ));
 sg13g2_nand4_1 _1382_ (.B(\load_weights[18] ),
    .C(net336),
    .A(net122),
    .Y(_0389_),
    .D(net96));
 sg13g2_o21ai_1 _1383_ (.B1(_0388_),
    .Y(_0390_),
    .A1(_0053_),
    .A2(net103));
 sg13g2_nand2_1 _1384_ (.Y(_0391_),
    .A(_0389_),
    .B(_0390_));
 sg13g2_xor2_1 _1385_ (.B(_0391_),
    .A(_0387_),
    .X(\tt_um_mult_inst.temp_out_comb[32] ));
 sg13g2_o21ai_1 _1386_ (.B1(_0389_),
    .Y(_0392_),
    .A1(_0387_),
    .A2(_0391_));
 sg13g2_and2_1 _1387_ (.A(\load_weights[8] ),
    .B(\load_weights[9] ),
    .X(_0393_));
 sg13g2_nand2_2 _1388_ (.Y(_0394_),
    .A(\load_weights[8] ),
    .B(\load_weights[9] ));
 sg13g2_nor2b_2 _1389_ (.A(\load_weights[9] ),
    .B_N(\load_weights[8] ),
    .Y(_0395_));
 sg13g2_a22oi_1 _1390_ (.Y(_0396_),
    .B1(_0395_),
    .B2(net117),
    .A2(_0393_),
    .A1(_0071_));
 sg13g2_nand2_1 _1391_ (.Y(_0397_),
    .A(\tt_um_mult_inst.temp_out[33] ),
    .B(net96));
 sg13g2_and2_2 _1392_ (.A(\load_weights[18] ),
    .B(\load_weights[19] ),
    .X(_0398_));
 sg13g2_nand2_1 _1393_ (.Y(_0399_),
    .A(\load_weights[18] ),
    .B(\load_weights[19] ));
 sg13g2_nor2b_2 _1394_ (.A(\load_weights[19] ),
    .B_N(\load_weights[18] ),
    .Y(_0400_));
 sg13g2_a22oi_1 _1395_ (.Y(_0401_),
    .B1(_0400_),
    .B2(net120),
    .A2(_0398_),
    .A1(_0077_));
 sg13g2_or2_1 _1396_ (.X(_0402_),
    .B(_0401_),
    .A(_0397_));
 sg13g2_xnor2_1 _1397_ (.Y(_0403_),
    .A(_0397_),
    .B(_0401_));
 sg13g2_xor2_1 _1398_ (.B(_0403_),
    .A(_0396_),
    .X(_0404_));
 sg13g2_nand2_1 _1399_ (.Y(_0405_),
    .A(_0392_),
    .B(_0404_));
 sg13g2_xor2_1 _1400_ (.B(_0404_),
    .A(_0392_),
    .X(\tt_um_mult_inst.temp_out_comb[33] ));
 sg13g2_o21ai_1 _1401_ (.B1(_0402_),
    .Y(_0406_),
    .A1(_0396_),
    .A2(_0403_));
 sg13g2_nand2_1 _1402_ (.Y(_0407_),
    .A(net115),
    .B(_0395_));
 sg13g2_a22oi_1 _1403_ (.Y(_0408_),
    .B1(_0395_),
    .B2(net115),
    .A2(_0393_),
    .A1(_0086_));
 sg13g2_o21ai_1 _1404_ (.B1(_0407_),
    .Y(_0409_),
    .A1(_0087_),
    .A2(_0394_));
 sg13g2_nand2_2 _1405_ (.Y(_0410_),
    .A(\tt_um_mult_inst.temp_out[34] ),
    .B(net96));
 sg13g2_nand3_1 _1406_ (.B(_0093_),
    .C(_0398_),
    .A(_0092_),
    .Y(_0411_));
 sg13g2_nand2_2 _1407_ (.Y(_0412_),
    .A(net2),
    .B(_0400_));
 sg13g2_a21oi_2 _1408_ (.B1(_0410_),
    .Y(_0413_),
    .A2(_0412_),
    .A1(_0411_));
 sg13g2_a21o_1 _1409_ (.A2(_0412_),
    .A1(_0411_),
    .B1(_0410_),
    .X(_0414_));
 sg13g2_and3_1 _1410_ (.X(_0415_),
    .A(_0410_),
    .B(_0411_),
    .C(_0412_));
 sg13g2_nand3_1 _1411_ (.B(_0411_),
    .C(_0412_),
    .A(_0410_),
    .Y(_0416_));
 sg13g2_nor3_2 _1412_ (.A(_0408_),
    .B(_0413_),
    .C(_0415_),
    .Y(_0417_));
 sg13g2_nand3_1 _1413_ (.B(_0414_),
    .C(_0416_),
    .A(_0409_),
    .Y(_0418_));
 sg13g2_a21oi_1 _1414_ (.A1(_0414_),
    .A2(_0416_),
    .Y(_0419_),
    .B1(_0409_));
 sg13g2_o21ai_1 _1415_ (.B1(_0408_),
    .Y(_0420_),
    .A1(_0413_),
    .A2(_0415_));
 sg13g2_nand3_1 _1416_ (.B(_0418_),
    .C(_0420_),
    .A(_0406_),
    .Y(_0421_));
 sg13g2_a21oi_1 _1417_ (.A1(_0418_),
    .A2(_0420_),
    .Y(_0422_),
    .B1(_0406_));
 sg13g2_nor3_1 _1418_ (.A(_0406_),
    .B(_0417_),
    .C(_0419_),
    .Y(_0423_));
 sg13g2_o21ai_1 _1419_ (.B1(_0406_),
    .Y(_0424_),
    .A1(_0417_),
    .A2(_0419_));
 sg13g2_nand2b_1 _1420_ (.Y(_0425_),
    .B(_0424_),
    .A_N(_0423_));
 sg13g2_xnor2_1 _1421_ (.Y(\tt_um_mult_inst.temp_out_comb[34] ),
    .A(_0405_),
    .B(_0425_));
 sg13g2_o21ai_1 _1422_ (.B1(_0421_),
    .Y(_0426_),
    .A1(_0405_),
    .A2(_0422_));
 sg13g2_nor2_1 _1423_ (.A(_0413_),
    .B(_0417_),
    .Y(_0427_));
 sg13g2_nand2_1 _1424_ (.Y(_0428_),
    .A(net114),
    .B(_0395_));
 sg13g2_o21ai_1 _1425_ (.B1(_0428_),
    .Y(_0429_),
    .A1(_0112_),
    .A2(_0394_));
 sg13g2_nand2_1 _1426_ (.Y(_0430_),
    .A(\tt_um_mult_inst.temp_out[35] ),
    .B(net95));
 sg13g2_nand2_1 _1427_ (.Y(_0431_),
    .A(net3),
    .B(_0400_));
 sg13g2_o21ai_1 _1428_ (.B1(_0431_),
    .Y(_0432_),
    .A1(_0117_),
    .A2(_0399_));
 sg13g2_nor2b_1 _1429_ (.A(_0430_),
    .B_N(_0432_),
    .Y(_0433_));
 sg13g2_xnor2_1 _1430_ (.Y(_0434_),
    .A(_0430_),
    .B(_0432_));
 sg13g2_xnor2_1 _1431_ (.Y(_0435_),
    .A(_0429_),
    .B(_0434_));
 sg13g2_nor2_1 _1432_ (.A(_0427_),
    .B(_0435_),
    .Y(_0436_));
 sg13g2_xor2_1 _1433_ (.B(_0435_),
    .A(_0427_),
    .X(_0437_));
 sg13g2_xor2_1 _1434_ (.B(_0437_),
    .A(_0426_),
    .X(\tt_um_mult_inst.temp_out_comb[35] ));
 sg13g2_a21oi_2 _1435_ (.B1(_0436_),
    .Y(_0438_),
    .A2(_0437_),
    .A1(_0426_));
 sg13g2_nand2_1 _1436_ (.Y(_0439_),
    .A(net113),
    .B(_0395_));
 sg13g2_o21ai_1 _1437_ (.B1(_0439_),
    .Y(_0440_),
    .A1(_0126_),
    .A2(_0394_));
 sg13g2_nand2_1 _1438_ (.Y(_0441_),
    .A(\tt_um_mult_inst.temp_out[36] ),
    .B(net95));
 sg13g2_a22oi_1 _1439_ (.Y(_0442_),
    .B1(_0400_),
    .B2(net4),
    .A2(_0398_),
    .A1(_0130_));
 sg13g2_nor2_1 _1440_ (.A(_0441_),
    .B(_0442_),
    .Y(_0443_));
 sg13g2_nand2_1 _1441_ (.Y(_0444_),
    .A(_0441_),
    .B(_0442_));
 sg13g2_xor2_1 _1442_ (.B(_0442_),
    .A(_0441_),
    .X(_0445_));
 sg13g2_xnor2_1 _1443_ (.Y(_0446_),
    .A(_0440_),
    .B(_0445_));
 sg13g2_a21oi_2 _1444_ (.B1(_0433_),
    .Y(_0447_),
    .A2(_0434_),
    .A1(_0429_));
 sg13g2_nor2_1 _1445_ (.A(_0446_),
    .B(_0447_),
    .Y(_0448_));
 sg13g2_xnor2_1 _1446_ (.Y(_0449_),
    .A(_0446_),
    .B(_0447_));
 sg13g2_nor2_1 _1447_ (.A(_0438_),
    .B(_0449_),
    .Y(_0450_));
 sg13g2_xor2_1 _1448_ (.B(_0449_),
    .A(_0438_),
    .X(\tt_um_mult_inst.temp_out_comb[36] ));
 sg13g2_a21oi_1 _1449_ (.A1(_0440_),
    .A2(_0444_),
    .Y(_0451_),
    .B1(_0443_));
 sg13g2_nand2_1 _1450_ (.Y(_0452_),
    .A(net112),
    .B(_0395_));
 sg13g2_o21ai_1 _1451_ (.B1(_0452_),
    .Y(_0453_),
    .A1(_0142_),
    .A2(_0394_));
 sg13g2_nand2_1 _1452_ (.Y(_0454_),
    .A(\tt_um_mult_inst.temp_out[37] ),
    .B(net95));
 sg13g2_nand3_1 _1453_ (.B(_0147_),
    .C(_0398_),
    .A(_0146_),
    .Y(_0455_));
 sg13g2_nand2_1 _1454_ (.Y(_0456_),
    .A(net5),
    .B(_0400_));
 sg13g2_a21oi_1 _1455_ (.A1(_0455_),
    .A2(_0456_),
    .Y(_0457_),
    .B1(_0454_));
 sg13g2_a21o_1 _1456_ (.A2(_0456_),
    .A1(_0455_),
    .B1(_0454_),
    .X(_0458_));
 sg13g2_nand3_1 _1457_ (.B(_0455_),
    .C(_0456_),
    .A(_0454_),
    .Y(_0459_));
 sg13g2_and3_1 _1458_ (.X(_0460_),
    .A(_0453_),
    .B(_0458_),
    .C(_0459_));
 sg13g2_a21oi_1 _1459_ (.A1(_0458_),
    .A2(_0459_),
    .Y(_0461_),
    .B1(_0453_));
 sg13g2_o21ai_1 _1460_ (.B1(_0451_),
    .Y(_0462_),
    .A1(_0460_),
    .A2(_0461_));
 sg13g2_nor3_1 _1461_ (.A(_0451_),
    .B(_0460_),
    .C(_0461_),
    .Y(_0463_));
 sg13g2_or3_1 _1462_ (.A(_0451_),
    .B(_0460_),
    .C(_0461_),
    .X(_0464_));
 sg13g2_nand2_1 _1463_ (.Y(_0465_),
    .A(_0462_),
    .B(_0464_));
 sg13g2_nor2_1 _1464_ (.A(_0448_),
    .B(_0450_),
    .Y(_0466_));
 sg13g2_xor2_1 _1465_ (.B(_0466_),
    .A(_0465_),
    .X(\tt_um_mult_inst.temp_out_comb[37] ));
 sg13g2_nand3b_1 _1466_ (.B(_0462_),
    .C(_0464_),
    .Y(_0467_),
    .A_N(_0449_));
 sg13g2_a21oi_1 _1467_ (.A1(_0448_),
    .A2(_0462_),
    .Y(_0468_),
    .B1(_0463_));
 sg13g2_o21ai_1 _1468_ (.B1(_0468_),
    .Y(_0469_),
    .A1(_0438_),
    .A2(_0467_));
 sg13g2_nor2_1 _1469_ (.A(_0457_),
    .B(_0460_),
    .Y(_0470_));
 sg13g2_a22oi_1 _1470_ (.Y(_0471_),
    .B1(_0395_),
    .B2(net111),
    .A2(_0393_),
    .A1(_0166_));
 sg13g2_nand2_1 _1471_ (.Y(_0472_),
    .A(\tt_um_mult_inst.temp_out[38] ),
    .B(net95));
 sg13g2_a22oi_1 _1472_ (.Y(_0473_),
    .B1(_0400_),
    .B2(net6),
    .A2(_0398_),
    .A1(_0170_));
 sg13g2_or2_1 _1473_ (.X(_0474_),
    .B(_0473_),
    .A(_0472_));
 sg13g2_xnor2_1 _1474_ (.Y(_0475_),
    .A(_0472_),
    .B(_0473_));
 sg13g2_xnor2_1 _1475_ (.Y(_0476_),
    .A(_0471_),
    .B(_0475_));
 sg13g2_nor2_1 _1476_ (.A(_0470_),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_xor2_1 _1477_ (.B(_0476_),
    .A(_0470_),
    .X(_0478_));
 sg13g2_xor2_1 _1478_ (.B(_0478_),
    .A(_0469_),
    .X(\tt_um_mult_inst.temp_out_comb[38] ));
 sg13g2_a21oi_1 _1479_ (.A1(_0469_),
    .A2(_0478_),
    .Y(_0479_),
    .B1(_0477_));
 sg13g2_o21ai_1 _1480_ (.B1(_0474_),
    .Y(_0480_),
    .A1(_0471_),
    .A2(_0475_));
 sg13g2_nand2_1 _1481_ (.Y(_0481_),
    .A(net333),
    .B(net95));
 sg13g2_a22oi_1 _1482_ (.Y(_0482_),
    .B1(_0400_),
    .B2(net7),
    .A2(_0398_),
    .A1(_0180_));
 sg13g2_a22oi_1 _1483_ (.Y(_0483_),
    .B1(_0395_),
    .B2(net14),
    .A2(_0393_),
    .A1(_0182_));
 sg13g2_xnor2_1 _1484_ (.Y(_0484_),
    .A(_0482_),
    .B(_0483_));
 sg13g2_xnor2_1 _1485_ (.Y(_0485_),
    .A(_0481_),
    .B(_0484_));
 sg13g2_xnor2_1 _1486_ (.Y(_0486_),
    .A(_0480_),
    .B(_0485_));
 sg13g2_xnor2_1 _1487_ (.Y(\tt_um_mult_inst.temp_out_comb[39] ),
    .A(_0479_),
    .B(_0486_));
 sg13g2_nand2_1 _1488_ (.Y(_0487_),
    .A(net119),
    .B(net435));
 sg13g2_nand2_1 _1489_ (.Y(_0488_),
    .A(net122),
    .B(\load_weights[14] ));
 sg13g2_nand4_1 _1490_ (.B(\load_weights[14] ),
    .C(net442),
    .A(net122),
    .Y(_0489_),
    .D(net96));
 sg13g2_o21ai_1 _1491_ (.B1(_0488_),
    .Y(_0490_),
    .A1(_0049_),
    .A2(net102));
 sg13g2_nand2_1 _1492_ (.Y(_0491_),
    .A(_0489_),
    .B(_0490_));
 sg13g2_xor2_1 _1493_ (.B(_0491_),
    .A(_0487_),
    .X(\tt_um_mult_inst.temp_out_comb[16] ));
 sg13g2_o21ai_1 _1494_ (.B1(_0489_),
    .Y(_0492_),
    .A1(_0487_),
    .A2(_0491_));
 sg13g2_and2_1 _1495_ (.A(\load_weights[4] ),
    .B(\load_weights[5] ),
    .X(_0493_));
 sg13g2_nand2_2 _1496_ (.Y(_0494_),
    .A(\load_weights[4] ),
    .B(\load_weights[5] ));
 sg13g2_nor2b_2 _1497_ (.A(\load_weights[5] ),
    .B_N(\load_weights[4] ),
    .Y(_0495_));
 sg13g2_a22oi_1 _1498_ (.Y(_0496_),
    .B1(_0495_),
    .B2(net117),
    .A2(_0493_),
    .A1(_0071_));
 sg13g2_nand2_1 _1499_ (.Y(_0497_),
    .A(\tt_um_mult_inst.temp_out[17] ),
    .B(net98));
 sg13g2_and2_2 _1500_ (.A(\load_weights[14] ),
    .B(\load_weights[15] ),
    .X(_0498_));
 sg13g2_nand2_1 _1501_ (.Y(_0499_),
    .A(\load_weights[14] ),
    .B(\load_weights[15] ));
 sg13g2_nor2b_2 _1502_ (.A(\load_weights[15] ),
    .B_N(\load_weights[14] ),
    .Y(_0500_));
 sg13g2_a22oi_1 _1503_ (.Y(_0501_),
    .B1(_0500_),
    .B2(net120),
    .A2(_0498_),
    .A1(_0077_));
 sg13g2_or2_1 _1504_ (.X(_0502_),
    .B(_0501_),
    .A(_0497_));
 sg13g2_xnor2_1 _1505_ (.Y(_0503_),
    .A(_0497_),
    .B(_0501_));
 sg13g2_xor2_1 _1506_ (.B(_0503_),
    .A(_0496_),
    .X(_0504_));
 sg13g2_nand2_1 _1507_ (.Y(_0505_),
    .A(_0492_),
    .B(_0504_));
 sg13g2_xor2_1 _1508_ (.B(_0504_),
    .A(_0492_),
    .X(\tt_um_mult_inst.temp_out_comb[17] ));
 sg13g2_o21ai_1 _1509_ (.B1(_0502_),
    .Y(_0506_),
    .A1(_0496_),
    .A2(_0503_));
 sg13g2_nand2_1 _1510_ (.Y(_0507_),
    .A(net116),
    .B(_0495_));
 sg13g2_a22oi_1 _1511_ (.Y(_0508_),
    .B1(_0495_),
    .B2(net116),
    .A2(_0493_),
    .A1(_0086_));
 sg13g2_o21ai_1 _1512_ (.B1(_0507_),
    .Y(_0509_),
    .A1(_0087_),
    .A2(_0494_));
 sg13g2_nand2_2 _1513_ (.Y(_0510_),
    .A(\tt_um_mult_inst.temp_out[18] ),
    .B(net98));
 sg13g2_nand3_1 _1514_ (.B(_0093_),
    .C(_0498_),
    .A(_0092_),
    .Y(_0511_));
 sg13g2_nand2_2 _1515_ (.Y(_0512_),
    .A(net2),
    .B(_0500_));
 sg13g2_a21oi_2 _1516_ (.B1(_0510_),
    .Y(_0513_),
    .A2(_0512_),
    .A1(_0511_));
 sg13g2_a21o_1 _1517_ (.A2(_0512_),
    .A1(_0511_),
    .B1(_0510_),
    .X(_0514_));
 sg13g2_and3_1 _1518_ (.X(_0515_),
    .A(_0510_),
    .B(_0511_),
    .C(_0512_));
 sg13g2_nand3_1 _1519_ (.B(_0511_),
    .C(_0512_),
    .A(_0510_),
    .Y(_0516_));
 sg13g2_nor3_2 _1520_ (.A(_0508_),
    .B(_0513_),
    .C(_0515_),
    .Y(_0517_));
 sg13g2_nand3_1 _1521_ (.B(_0514_),
    .C(_0516_),
    .A(_0509_),
    .Y(_0518_));
 sg13g2_a21oi_1 _1522_ (.A1(_0514_),
    .A2(_0516_),
    .Y(_0519_),
    .B1(_0509_));
 sg13g2_o21ai_1 _1523_ (.B1(_0508_),
    .Y(_0520_),
    .A1(_0513_),
    .A2(_0515_));
 sg13g2_nand3_1 _1524_ (.B(_0518_),
    .C(_0520_),
    .A(_0506_),
    .Y(_0521_));
 sg13g2_a21oi_1 _1525_ (.A1(_0518_),
    .A2(_0520_),
    .Y(_0522_),
    .B1(_0506_));
 sg13g2_nor3_1 _1526_ (.A(_0506_),
    .B(_0517_),
    .C(_0519_),
    .Y(_0523_));
 sg13g2_o21ai_1 _1527_ (.B1(_0506_),
    .Y(_0524_),
    .A1(_0517_),
    .A2(_0519_));
 sg13g2_nand2b_1 _1528_ (.Y(_0525_),
    .B(_0524_),
    .A_N(_0523_));
 sg13g2_xnor2_1 _1529_ (.Y(\tt_um_mult_inst.temp_out_comb[18] ),
    .A(_0505_),
    .B(_0525_));
 sg13g2_o21ai_1 _1530_ (.B1(_0521_),
    .Y(_0526_),
    .A1(_0505_),
    .A2(_0522_));
 sg13g2_nor2_1 _1531_ (.A(_0513_),
    .B(_0517_),
    .Y(_0527_));
 sg13g2_nand2_1 _1532_ (.Y(_0528_),
    .A(net114),
    .B(_0495_));
 sg13g2_o21ai_1 _1533_ (.B1(_0528_),
    .Y(_0529_),
    .A1(_0112_),
    .A2(_0494_));
 sg13g2_nand2_1 _1534_ (.Y(_0530_),
    .A(\tt_um_mult_inst.temp_out[19] ),
    .B(net97));
 sg13g2_nand2_1 _1535_ (.Y(_0531_),
    .A(net3),
    .B(_0500_));
 sg13g2_o21ai_1 _1536_ (.B1(_0531_),
    .Y(_0532_),
    .A1(_0117_),
    .A2(_0499_));
 sg13g2_nor2b_1 _1537_ (.A(_0530_),
    .B_N(_0532_),
    .Y(_0533_));
 sg13g2_xnor2_1 _1538_ (.Y(_0534_),
    .A(_0530_),
    .B(_0532_));
 sg13g2_xnor2_1 _1539_ (.Y(_0535_),
    .A(_0529_),
    .B(_0534_));
 sg13g2_nor2_1 _1540_ (.A(_0527_),
    .B(_0535_),
    .Y(_0536_));
 sg13g2_xor2_1 _1541_ (.B(_0535_),
    .A(_0527_),
    .X(_0537_));
 sg13g2_xor2_1 _1542_ (.B(_0537_),
    .A(_0526_),
    .X(\tt_um_mult_inst.temp_out_comb[19] ));
 sg13g2_a21oi_2 _1543_ (.B1(_0536_),
    .Y(_0538_),
    .A2(_0537_),
    .A1(_0526_));
 sg13g2_nand2_1 _1544_ (.Y(_0539_),
    .A(net113),
    .B(_0495_));
 sg13g2_o21ai_1 _1545_ (.B1(_0539_),
    .Y(_0540_),
    .A1(_0126_),
    .A2(_0494_));
 sg13g2_nand2_1 _1546_ (.Y(_0541_),
    .A(\tt_um_mult_inst.temp_out[20] ),
    .B(net93));
 sg13g2_a22oi_1 _1547_ (.Y(_0542_),
    .B1(_0500_),
    .B2(net4),
    .A2(_0498_),
    .A1(_0130_));
 sg13g2_nor2_1 _1548_ (.A(_0541_),
    .B(_0542_),
    .Y(_0543_));
 sg13g2_nand2_1 _1549_ (.Y(_0544_),
    .A(_0541_),
    .B(_0542_));
 sg13g2_xor2_1 _1550_ (.B(_0542_),
    .A(_0541_),
    .X(_0545_));
 sg13g2_xnor2_1 _1551_ (.Y(_0546_),
    .A(_0540_),
    .B(_0545_));
 sg13g2_a21oi_2 _1552_ (.B1(_0533_),
    .Y(_0547_),
    .A2(_0534_),
    .A1(_0529_));
 sg13g2_nor2_1 _1553_ (.A(_0546_),
    .B(_0547_),
    .Y(_0548_));
 sg13g2_xor2_1 _1554_ (.B(_0547_),
    .A(_0546_),
    .X(_0549_));
 sg13g2_nor2b_1 _1555_ (.A(_0538_),
    .B_N(_0549_),
    .Y(_0550_));
 sg13g2_xnor2_1 _1556_ (.Y(\tt_um_mult_inst.temp_out_comb[20] ),
    .A(_0538_),
    .B(_0549_));
 sg13g2_a21oi_1 _1557_ (.A1(_0540_),
    .A2(_0544_),
    .Y(_0551_),
    .B1(_0543_));
 sg13g2_nand2_1 _1558_ (.Y(_0552_),
    .A(net112),
    .B(_0495_));
 sg13g2_o21ai_1 _1559_ (.B1(_0552_),
    .Y(_0553_),
    .A1(_0142_),
    .A2(_0494_));
 sg13g2_nand2_1 _1560_ (.Y(_0554_),
    .A(\tt_um_mult_inst.temp_out[21] ),
    .B(net93));
 sg13g2_nand3_1 _1561_ (.B(_0147_),
    .C(_0498_),
    .A(_0146_),
    .Y(_0555_));
 sg13g2_nand2_1 _1562_ (.Y(_0556_),
    .A(net5),
    .B(_0500_));
 sg13g2_a21oi_1 _1563_ (.A1(_0555_),
    .A2(_0556_),
    .Y(_0557_),
    .B1(_0554_));
 sg13g2_a21o_1 _1564_ (.A2(_0556_),
    .A1(_0555_),
    .B1(_0554_),
    .X(_0558_));
 sg13g2_nand3_1 _1565_ (.B(_0555_),
    .C(_0556_),
    .A(_0554_),
    .Y(_0559_));
 sg13g2_and3_1 _1566_ (.X(_0560_),
    .A(_0553_),
    .B(_0558_),
    .C(_0559_));
 sg13g2_a21oi_1 _1567_ (.A1(_0558_),
    .A2(_0559_),
    .Y(_0561_),
    .B1(_0553_));
 sg13g2_o21ai_1 _1568_ (.B1(_0551_),
    .Y(_0562_),
    .A1(_0560_),
    .A2(_0561_));
 sg13g2_nor3_1 _1569_ (.A(_0551_),
    .B(_0560_),
    .C(_0561_),
    .Y(_0563_));
 sg13g2_or3_1 _1570_ (.A(_0551_),
    .B(_0560_),
    .C(_0561_),
    .X(_0564_));
 sg13g2_and2_1 _1571_ (.A(_0562_),
    .B(_0564_),
    .X(_0565_));
 sg13g2_nor2_1 _1572_ (.A(_0548_),
    .B(_0550_),
    .Y(_0566_));
 sg13g2_xnor2_1 _1573_ (.Y(\tt_um_mult_inst.temp_out_comb[21] ),
    .A(_0565_),
    .B(_0566_));
 sg13g2_nand3b_1 _1574_ (.B(_0549_),
    .C(_0562_),
    .Y(_0567_),
    .A_N(_0563_));
 sg13g2_a21oi_1 _1575_ (.A1(_0548_),
    .A2(_0562_),
    .Y(_0568_),
    .B1(_0563_));
 sg13g2_o21ai_1 _1576_ (.B1(_0568_),
    .Y(_0569_),
    .A1(_0538_),
    .A2(_0567_));
 sg13g2_nor2_1 _1577_ (.A(_0557_),
    .B(_0560_),
    .Y(_0570_));
 sg13g2_a22oi_1 _1578_ (.Y(_0571_),
    .B1(_0495_),
    .B2(net111),
    .A2(_0493_),
    .A1(_0166_));
 sg13g2_nand2_1 _1579_ (.Y(_0572_),
    .A(\tt_um_mult_inst.temp_out[22] ),
    .B(net93));
 sg13g2_a22oi_1 _1580_ (.Y(_0573_),
    .B1(_0500_),
    .B2(net6),
    .A2(_0498_),
    .A1(_0170_));
 sg13g2_or2_1 _1581_ (.X(_0574_),
    .B(_0573_),
    .A(_0572_));
 sg13g2_xnor2_1 _1582_ (.Y(_0575_),
    .A(_0572_),
    .B(_0573_));
 sg13g2_xnor2_1 _1583_ (.Y(_0576_),
    .A(_0571_),
    .B(_0575_));
 sg13g2_nor2_1 _1584_ (.A(_0570_),
    .B(_0576_),
    .Y(_0577_));
 sg13g2_xor2_1 _1585_ (.B(_0576_),
    .A(_0570_),
    .X(_0578_));
 sg13g2_xor2_1 _1586_ (.B(_0578_),
    .A(_0569_),
    .X(\tt_um_mult_inst.temp_out_comb[22] ));
 sg13g2_a21oi_1 _1587_ (.A1(_0569_),
    .A2(_0578_),
    .Y(_0579_),
    .B1(_0577_));
 sg13g2_o21ai_1 _1588_ (.B1(_0574_),
    .Y(_0580_),
    .A1(_0571_),
    .A2(_0575_));
 sg13g2_nand2_1 _1589_ (.Y(_0581_),
    .A(net445),
    .B(net93));
 sg13g2_a22oi_1 _1590_ (.Y(_0582_),
    .B1(_0500_),
    .B2(net7),
    .A2(_0498_),
    .A1(_0180_));
 sg13g2_a22oi_1 _1591_ (.Y(_0583_),
    .B1(_0495_),
    .B2(net14),
    .A2(_0493_),
    .A1(_0182_));
 sg13g2_xnor2_1 _1592_ (.Y(_0584_),
    .A(_0582_),
    .B(_0583_));
 sg13g2_xnor2_1 _1593_ (.Y(_0585_),
    .A(_0581_),
    .B(_0584_));
 sg13g2_xnor2_1 _1594_ (.Y(_0586_),
    .A(_0580_),
    .B(_0585_));
 sg13g2_xnor2_1 _1595_ (.Y(\tt_um_mult_inst.temp_out_comb[23] ),
    .A(_0579_),
    .B(_0586_));
 sg13g2_nor2_1 _1596_ (.A(_0053_),
    .B(net96),
    .Y(_0033_));
 sg13g2_and2_1 _1597_ (.A(net331),
    .B(net103),
    .X(_0034_));
 sg13g2_and2_1 _1598_ (.A(net337),
    .B(net103),
    .X(_0035_));
 sg13g2_and2_1 _1599_ (.A(net338),
    .B(net103),
    .X(_0036_));
 sg13g2_and2_1 _1600_ (.A(net329),
    .B(net101),
    .X(_0037_));
 sg13g2_and2_1 _1601_ (.A(net330),
    .B(net101),
    .X(_0038_));
 sg13g2_and2_1 _1602_ (.A(net332),
    .B(net101),
    .X(_0039_));
 sg13g2_and2_1 _1603_ (.A(net333),
    .B(net99),
    .X(_0040_));
 sg13g2_and2_1 _1604_ (.A(net404),
    .B(\count[0] ),
    .X(_0587_));
 sg13g2_nor3_1 _1605_ (.A(_0046_),
    .B(_0055_),
    .C(net405),
    .Y(_0041_));
 sg13g2_nand2_1 _1606_ (.Y(_0588_),
    .A(net401),
    .B(_0055_));
 sg13g2_nor2_1 _1607_ (.A(net401),
    .B(net405),
    .Y(_0589_));
 sg13g2_nand2_1 _1608_ (.Y(_0590_),
    .A(net401),
    .B(_0587_));
 sg13g2_nand3_1 _1609_ (.B(_0588_),
    .C(_0590_),
    .A(net1),
    .Y(_0591_));
 sg13g2_nor2_1 _1610_ (.A(_0589_),
    .B(_0591_),
    .Y(_0042_));
 sg13g2_xor2_1 _1611_ (.B(_0590_),
    .A(net406),
    .X(_0592_));
 sg13g2_a21oi_1 _1612_ (.A1(_0588_),
    .A2(_0592_),
    .Y(_0043_),
    .B1(_0046_));
 sg13g2_and3_1 _1613_ (.X(_0044_),
    .A(net1),
    .B(net327),
    .C(_0588_));
 sg13g2_a21oi_1 _1614_ (.A1(net401),
    .A2(_0055_),
    .Y(_0593_),
    .B1(net110));
 sg13g2_nor3_1 _1615_ (.A(_0046_),
    .B(net108),
    .C(net402),
    .Y(_0045_));
 sg13g2_dfrbp_1 _1616_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net42),
    .D(_0033_),
    .Q_N(_0606_),
    .Q(\tt_um_mult_inst.pipe_out[32] ));
 sg13g2_dfrbp_1 _1617_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net34),
    .D(_0034_),
    .Q_N(_0605_),
    .Q(\tt_um_mult_inst.pipe_out[33] ));
 sg13g2_dfrbp_1 _1618_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net33),
    .D(_0035_),
    .Q_N(_0604_),
    .Q(\tt_um_mult_inst.pipe_out[34] ));
 sg13g2_dfrbp_1 _1619_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net32),
    .D(_0036_),
    .Q_N(_0603_),
    .Q(\tt_um_mult_inst.pipe_out[35] ));
 sg13g2_dfrbp_1 _1620_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net31),
    .D(_0037_),
    .Q_N(_0602_),
    .Q(\tt_um_mult_inst.pipe_out[36] ));
 sg13g2_dfrbp_1 _1621_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net206),
    .D(_0038_),
    .Q_N(_0601_),
    .Q(\tt_um_mult_inst.pipe_out[37] ));
 sg13g2_dfrbp_1 _1622_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net173),
    .D(_0039_),
    .Q_N(_0600_),
    .Q(\tt_um_mult_inst.pipe_out[38] ));
 sg13g2_dfrbp_1 _1623_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net41),
    .D(_0040_),
    .Q_N(_0599_),
    .Q(\tt_um_mult_inst.pipe_out[39] ));
 sg13g2_dfrbp_1 _1624_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net40),
    .D(_0041_),
    .Q_N(_0598_),
    .Q(\count[1] ));
 sg13g2_dfrbp_1 _1625_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net39),
    .D(_0042_),
    .Q_N(_0597_),
    .Q(\count[2] ));
 sg13g2_dfrbp_1 _1626_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net43),
    .D(net407),
    .Q_N(_0607_),
    .Q(\count[3] ));
 sg13g2_dfrbp_1 _1627_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net44),
    .D(net256),
    .Q_N(_0608_),
    .Q(\load_weights[0] ));
 sg13g2_dfrbp_1 _1628_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net45),
    .D(net291),
    .Q_N(_0609_),
    .Q(\load_weights[1] ));
 sg13g2_dfrbp_1 _1629_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net46),
    .D(net263),
    .Q_N(_0610_),
    .Q(\load_weights[2] ));
 sg13g2_dfrbp_1 _1630_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net47),
    .D(net255),
    .Q_N(_0611_),
    .Q(\load_weights[3] ));
 sg13g2_dfrbp_1 _1631_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net48),
    .D(net277),
    .Q_N(_0612_),
    .Q(\load_weights[4] ));
 sg13g2_dfrbp_1 _1632_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net49),
    .D(net253),
    .Q_N(_0613_),
    .Q(\load_weights[5] ));
 sg13g2_dfrbp_1 _1633_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net50),
    .D(net286),
    .Q_N(_0614_),
    .Q(\load_weights[6] ));
 sg13g2_dfrbp_1 _1634_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net51),
    .D(net287),
    .Q_N(_0615_),
    .Q(\load_weights[7] ));
 sg13g2_dfrbp_1 _1635_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net52),
    .D(net254),
    .Q_N(_0616_),
    .Q(\load_weights[8] ));
 sg13g2_dfrbp_1 _1636_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net53),
    .D(net257),
    .Q_N(_0617_),
    .Q(\load_weights[9] ));
 sg13g2_dfrbp_1 _1637_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net54),
    .D(net311),
    .Q_N(_0618_),
    .Q(\load_weights[10] ));
 sg13g2_dfrbp_1 _1638_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net55),
    .D(net313),
    .Q_N(_0619_),
    .Q(\load_weights[11] ));
 sg13g2_dfrbp_1 _1639_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net56),
    .D(net301),
    .Q_N(_0620_),
    .Q(\load_weights[12] ));
 sg13g2_dfrbp_1 _1640_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net57),
    .D(net288),
    .Q_N(_0621_),
    .Q(\load_weights[13] ));
 sg13g2_dfrbp_1 _1641_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net58),
    .D(net251),
    .Q_N(_0622_),
    .Q(\load_weights[14] ));
 sg13g2_dfrbp_1 _1642_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net59),
    .D(net293),
    .Q_N(_0623_),
    .Q(\load_weights[15] ));
 sg13g2_dfrbp_1 _1643_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net60),
    .D(net285),
    .Q_N(_0624_),
    .Q(\load_weights[16] ));
 sg13g2_dfrbp_1 _1644_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net61),
    .D(net312),
    .Q_N(_0625_),
    .Q(\load_weights[17] ));
 sg13g2_dfrbp_1 _1645_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net62),
    .D(net305),
    .Q_N(_0626_),
    .Q(\load_weights[18] ));
 sg13g2_dfrbp_1 _1646_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net63),
    .D(net297),
    .Q_N(_0627_),
    .Q(\load_weights[19] ));
 sg13g2_dfrbp_1 _1647_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net64),
    .D(net248),
    .Q_N(_0628_),
    .Q(\tt_um_load_inst.weights[20] ));
 sg13g2_dfrbp_1 _1648_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net65),
    .D(net274),
    .Q_N(_0629_),
    .Q(\tt_um_load_inst.weights[21] ));
 sg13g2_dfrbp_1 _1649_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net66),
    .D(net317),
    .Q_N(_0630_),
    .Q(\tt_um_load_inst.weights[22] ));
 sg13g2_dfrbp_1 _1650_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net67),
    .D(net272),
    .Q_N(_0631_),
    .Q(\tt_um_load_inst.weights[23] ));
 sg13g2_dfrbp_1 _1651_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net68),
    .D(net278),
    .Q_N(_0632_),
    .Q(\tt_um_load_inst.weights[24] ));
 sg13g2_dfrbp_1 _1652_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net69),
    .D(net261),
    .Q_N(_0633_),
    .Q(\tt_um_load_inst.weights[25] ));
 sg13g2_dfrbp_1 _1653_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net70),
    .D(net276),
    .Q_N(_0634_),
    .Q(\tt_um_load_inst.weights[26] ));
 sg13g2_dfrbp_1 _1654_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net71),
    .D(net252),
    .Q_N(_0635_),
    .Q(\tt_um_load_inst.weights[27] ));
 sg13g2_dfrbp_1 _1655_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net72),
    .D(net318),
    .Q_N(_0636_),
    .Q(\tt_um_load_inst.weights[28] ));
 sg13g2_dfrbp_1 _1656_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net73),
    .D(net247),
    .Q_N(_0637_),
    .Q(\tt_um_load_inst.weights[29] ));
 sg13g2_dfrbp_1 _1657_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net74),
    .D(net307),
    .Q_N(_0638_),
    .Q(\tt_um_load_inst.weights[30] ));
 sg13g2_dfrbp_1 _1658_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net75),
    .D(net310),
    .Q_N(_0639_),
    .Q(\tt_um_load_inst.weights[31] ));
 sg13g2_dfrbp_1 _1659_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net76),
    .D(net290),
    .Q_N(_0640_),
    .Q(\tt_um_load_inst.weights[32] ));
 sg13g2_dfrbp_1 _1660_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net77),
    .D(net309),
    .Q_N(_0641_),
    .Q(\tt_um_load_inst.weights[33] ));
 sg13g2_dfrbp_1 _1661_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net78),
    .D(net281),
    .Q_N(_0642_),
    .Q(\tt_um_load_inst.weights[34] ));
 sg13g2_dfrbp_1 _1662_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net79),
    .D(net323),
    .Q_N(_0643_),
    .Q(\tt_um_load_inst.weights[35] ));
 sg13g2_dfrbp_1 _1663_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net80),
    .D(net275),
    .Q_N(_0644_),
    .Q(\tt_um_load_inst.weights[36] ));
 sg13g2_dfrbp_1 _1664_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net81),
    .D(net250),
    .Q_N(_0645_),
    .Q(\tt_um_load_inst.weights[37] ));
 sg13g2_dfrbp_1 _1665_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net82),
    .D(net322),
    .Q_N(_0646_),
    .Q(\tt_um_load_inst.weights[38] ));
 sg13g2_dfrbp_1 _1666_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net83),
    .D(net326),
    .Q_N(_0647_),
    .Q(\tt_um_load_inst.weights[39] ));
 sg13g2_dfrbp_1 _1667_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net84),
    .D(net260),
    .Q_N(_0648_),
    .Q(\tt_um_load_inst.weights[40] ));
 sg13g2_dfrbp_1 _1668_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net85),
    .D(net296),
    .Q_N(_0649_),
    .Q(\tt_um_load_inst.weights[41] ));
 sg13g2_dfrbp_1 _1669_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net86),
    .D(net271),
    .Q_N(_0650_),
    .Q(\tt_um_load_inst.weights[42] ));
 sg13g2_dfrbp_1 _1670_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net87),
    .D(net282),
    .Q_N(_0651_),
    .Q(\tt_um_load_inst.weights[43] ));
 sg13g2_dfrbp_1 _1671_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net88),
    .D(net284),
    .Q_N(_0652_),
    .Q(\tt_um_load_inst.weights[44] ));
 sg13g2_dfrbp_1 _1672_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net89),
    .D(net249),
    .Q_N(_0653_),
    .Q(\tt_um_load_inst.weights[45] ));
 sg13g2_dfrbp_1 _1673_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net90),
    .D(net280),
    .Q_N(_0654_),
    .Q(\tt_um_load_inst.weights[46] ));
 sg13g2_dfrbp_1 _1674_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net91),
    .D(net294),
    .Q_N(_0655_),
    .Q(\tt_um_load_inst.weights[47] ));
 sg13g2_dfrbp_1 _1675_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net92),
    .D(net299),
    .Q_N(_0656_),
    .Q(\tt_um_load_inst.weights[48] ));
 sg13g2_dfrbp_1 _1676_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net124),
    .D(net324),
    .Q_N(_0657_),
    .Q(\tt_um_load_inst.weights[49] ));
 sg13g2_dfrbp_1 _1677_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net125),
    .D(net295),
    .Q_N(_0658_),
    .Q(\tt_um_load_inst.weights[50] ));
 sg13g2_dfrbp_1 _1678_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net126),
    .D(net262),
    .Q_N(_0659_),
    .Q(\tt_um_load_inst.weights[51] ));
 sg13g2_dfrbp_1 _1679_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net127),
    .D(net300),
    .Q_N(_0660_),
    .Q(\tt_um_load_inst.weights[52] ));
 sg13g2_dfrbp_1 _1680_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net128),
    .D(net316),
    .Q_N(_0661_),
    .Q(\tt_um_load_inst.weights[53] ));
 sg13g2_dfrbp_1 _1681_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net129),
    .D(net267),
    .Q_N(_0662_),
    .Q(\tt_um_load_inst.weights[54] ));
 sg13g2_dfrbp_1 _1682_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net130),
    .D(net302),
    .Q_N(_0663_),
    .Q(\tt_um_load_inst.weights[55] ));
 sg13g2_dfrbp_1 _1683_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net131),
    .D(net270),
    .Q_N(_0664_),
    .Q(\tt_um_load_inst.weights[56] ));
 sg13g2_dfrbp_1 _1684_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net132),
    .D(net315),
    .Q_N(_0665_),
    .Q(\tt_um_load_inst.weights[57] ));
 sg13g2_dfrbp_1 _1685_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net133),
    .D(net308),
    .Q_N(_0666_),
    .Q(\tt_um_load_inst.weights[58] ));
 sg13g2_dfrbp_1 _1686_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net134),
    .D(net303),
    .Q_N(_0667_),
    .Q(\tt_um_load_inst.weights[59] ));
 sg13g2_dfrbp_1 _1687_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net135),
    .D(net292),
    .Q_N(_0668_),
    .Q(\tt_um_load_inst.weights[60] ));
 sg13g2_dfrbp_1 _1688_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net136),
    .D(net320),
    .Q_N(_0669_),
    .Q(\tt_um_load_inst.weights[61] ));
 sg13g2_dfrbp_1 _1689_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net137),
    .D(net258),
    .Q_N(_0670_),
    .Q(\tt_um_load_inst.weights[62] ));
 sg13g2_dfrbp_1 _1690_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net138),
    .D(net314),
    .Q_N(_0671_),
    .Q(\tt_um_load_inst.weights[63] ));
 sg13g2_dfrbp_1 _1691_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net139),
    .D(net268),
    .Q_N(_0672_),
    .Q(\tt_um_load_inst.weights[64] ));
 sg13g2_dfrbp_1 _1692_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net140),
    .D(net289),
    .Q_N(_0673_),
    .Q(\tt_um_load_inst.weights[65] ));
 sg13g2_dfrbp_1 _1693_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net141),
    .D(net273),
    .Q_N(_0674_),
    .Q(\tt_um_load_inst.weights[66] ));
 sg13g2_dfrbp_1 _1694_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net142),
    .D(net306),
    .Q_N(_0675_),
    .Q(\tt_um_load_inst.weights[67] ));
 sg13g2_dfrbp_1 _1695_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net143),
    .D(net259),
    .Q_N(_0676_),
    .Q(\tt_um_load_inst.weights[68] ));
 sg13g2_dfrbp_1 _1696_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net144),
    .D(net304),
    .Q_N(_0677_),
    .Q(\tt_um_load_inst.weights[69] ));
 sg13g2_dfrbp_1 _1697_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net145),
    .D(net319),
    .Q_N(_0678_),
    .Q(\tt_um_load_inst.weights[70] ));
 sg13g2_dfrbp_1 _1698_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net146),
    .D(net325),
    .Q_N(_0679_),
    .Q(\tt_um_load_inst.weights[71] ));
 sg13g2_dfrbp_1 _1699_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net147),
    .D(net265),
    .Q_N(_0680_),
    .Q(\tt_um_load_inst.weights[72] ));
 sg13g2_dfrbp_1 _1700_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net148),
    .D(net298),
    .Q_N(_0681_),
    .Q(\tt_um_load_inst.weights[73] ));
 sg13g2_dfrbp_1 _1701_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net149),
    .D(net321),
    .Q_N(_0682_),
    .Q(\tt_um_load_inst.weights[74] ));
 sg13g2_dfrbp_1 _1702_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net150),
    .D(net266),
    .Q_N(_0683_),
    .Q(\tt_um_load_inst.weights[75] ));
 sg13g2_dfrbp_1 _1703_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net151),
    .D(net279),
    .Q_N(_0684_),
    .Q(\tt_um_load_inst.weights[76] ));
 sg13g2_dfrbp_1 _1704_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net152),
    .D(net283),
    .Q_N(_0685_),
    .Q(\tt_um_load_inst.weights[77] ));
 sg13g2_dfrbp_1 _1705_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net153),
    .D(net269),
    .Q_N(_0686_),
    .Q(\tt_um_load_inst.weights[78] ));
 sg13g2_dfrbp_1 _1706_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net154),
    .D(net264),
    .Q_N(_0687_),
    .Q(\tt_um_load_inst.weights[79] ));
 sg13g2_dfrbp_1 _1707_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net155),
    .D(\tt_um_load_inst.input_to_sr[0] ),
    .Q_N(_0688_),
    .Q(\tt_um_load_inst.weights[80] ));
 sg13g2_dfrbp_1 _1708_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net156),
    .D(\tt_um_load_inst.input_to_sr[1] ),
    .Q_N(_0689_),
    .Q(\tt_um_load_inst.weights[81] ));
 sg13g2_dfrbp_1 _1709_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net157),
    .D(\tt_um_load_inst.input_to_sr[2] ),
    .Q_N(_0690_),
    .Q(\tt_um_load_inst.weights[82] ));
 sg13g2_dfrbp_1 _1710_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net158),
    .D(\tt_um_load_inst.input_to_sr[3] ),
    .Q_N(_0691_),
    .Q(\tt_um_load_inst.weights[83] ));
 sg13g2_dfrbp_1 _1711_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net159),
    .D(\tt_um_load_inst.input_to_sr[4] ),
    .Q_N(_0692_),
    .Q(\tt_um_load_inst.weights[84] ));
 sg13g2_dfrbp_1 _1712_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net160),
    .D(\tt_um_load_inst.input_to_sr[5] ),
    .Q_N(_0693_),
    .Q(\tt_um_load_inst.weights[85] ));
 sg13g2_dfrbp_1 _1713_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net161),
    .D(\tt_um_load_inst.input_to_sr[6] ),
    .Q_N(_0694_),
    .Q(\tt_um_load_inst.weights[86] ));
 sg13g2_dfrbp_1 _1714_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net162),
    .D(\tt_um_load_inst.input_to_sr[7] ),
    .Q_N(_0695_),
    .Q(\tt_um_load_inst.weights[87] ));
 sg13g2_dfrbp_1 _1715_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net163),
    .D(\tt_um_load_inst.input_to_sr[8] ),
    .Q_N(_0696_),
    .Q(\tt_um_load_inst.weights[88] ));
 sg13g2_dfrbp_1 _1716_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net164),
    .D(\tt_um_load_inst.input_to_sr[9] ),
    .Q_N(_0697_),
    .Q(\tt_um_load_inst.weights[89] ));
 sg13g2_dfrbp_1 _1717_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net165),
    .D(net422),
    .Q_N(_0698_),
    .Q(\tt_um_load_inst.weights[90] ));
 sg13g2_dfrbp_1 _1718_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net166),
    .D(net420),
    .Q_N(_0699_),
    .Q(\tt_um_load_inst.weights[91] ));
 sg13g2_dfrbp_1 _1719_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net167),
    .D(net425),
    .Q_N(_0700_),
    .Q(\tt_um_load_inst.weights[92] ));
 sg13g2_dfrbp_1 _1720_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net168),
    .D(net409),
    .Q_N(_0701_),
    .Q(\tt_um_load_inst.weights[93] ));
 sg13g2_dfrbp_1 _1721_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net169),
    .D(net441),
    .Q_N(_0702_),
    .Q(\tt_um_load_inst.weights[94] ));
 sg13g2_dfrbp_1 _1722_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net170),
    .D(net413),
    .Q_N(_0703_),
    .Q(\tt_um_load_inst.weights[95] ));
 sg13g2_dfrbp_1 _1723_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net171),
    .D(net437),
    .Q_N(_0704_),
    .Q(\tt_um_load_inst.weights[96] ));
 sg13g2_dfrbp_1 _1724_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net172),
    .D(net417),
    .Q_N(_0705_),
    .Q(\tt_um_load_inst.weights[97] ));
 sg13g2_dfrbp_1 _1725_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net174),
    .D(net428),
    .Q_N(_0706_),
    .Q(\tt_um_load_inst.weights[98] ));
 sg13g2_dfrbp_1 _1726_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net38),
    .D(net411),
    .Q_N(_0596_),
    .Q(\tt_um_load_inst.weights[99] ));
 sg13g2_dfrbp_1 _1727_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net175),
    .D(net328),
    .Q_N(_0032_),
    .Q(\count[0] ));
 sg13g2_dfrbp_1 _1728_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net176),
    .D(net380),
    .Q_N(_0707_),
    .Q(\tt_um_mult_inst.pipe_out[0] ));
 sg13g2_dfrbp_1 _1729_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net177),
    .D(net376),
    .Q_N(_0708_),
    .Q(\tt_um_mult_inst.pipe_out[1] ));
 sg13g2_dfrbp_1 _1730_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net178),
    .D(net386),
    .Q_N(_0709_),
    .Q(\tt_um_mult_inst.pipe_out[2] ));
 sg13g2_dfrbp_1 _1731_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net179),
    .D(net358),
    .Q_N(_0710_),
    .Q(\tt_um_mult_inst.pipe_out[3] ));
 sg13g2_dfrbp_1 _1732_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net180),
    .D(net350),
    .Q_N(_0711_),
    .Q(\tt_um_mult_inst.pipe_out[4] ));
 sg13g2_dfrbp_1 _1733_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net181),
    .D(net340),
    .Q_N(_0712_),
    .Q(\tt_um_mult_inst.pipe_out[5] ));
 sg13g2_dfrbp_1 _1734_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net182),
    .D(net356),
    .Q_N(_0713_),
    .Q(\tt_um_mult_inst.pipe_out[6] ));
 sg13g2_dfrbp_1 _1735_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net183),
    .D(net348),
    .Q_N(_0714_),
    .Q(\tt_um_mult_inst.pipe_out[7] ));
 sg13g2_dfrbp_1 _1736_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net184),
    .D(net390),
    .Q_N(_0715_),
    .Q(\tt_um_mult_inst.pipe_out[8] ));
 sg13g2_dfrbp_1 _1737_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net185),
    .D(net368),
    .Q_N(_0716_),
    .Q(\tt_um_mult_inst.pipe_out[9] ));
 sg13g2_dfrbp_1 _1738_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net186),
    .D(net396),
    .Q_N(_0717_),
    .Q(\tt_um_mult_inst.pipe_out[10] ));
 sg13g2_dfrbp_1 _1739_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net187),
    .D(net398),
    .Q_N(_0718_),
    .Q(\tt_um_mult_inst.pipe_out[11] ));
 sg13g2_dfrbp_1 _1740_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net188),
    .D(net335),
    .Q_N(_0719_),
    .Q(\tt_um_mult_inst.pipe_out[12] ));
 sg13g2_dfrbp_1 _1741_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net189),
    .D(net374),
    .Q_N(_0720_),
    .Q(\tt_um_mult_inst.pipe_out[13] ));
 sg13g2_dfrbp_1 _1742_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net190),
    .D(net352),
    .Q_N(_0721_),
    .Q(\tt_um_mult_inst.pipe_out[14] ));
 sg13g2_dfrbp_1 _1743_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net191),
    .D(net382),
    .Q_N(_0722_),
    .Q(\tt_um_mult_inst.pipe_out[15] ));
 sg13g2_dfrbp_1 _1744_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net192),
    .D(net370),
    .Q_N(_0723_),
    .Q(\tt_um_mult_inst.pipe_out[16] ));
 sg13g2_dfrbp_1 _1745_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net193),
    .D(net384),
    .Q_N(_0724_),
    .Q(\tt_um_mult_inst.pipe_out[17] ));
 sg13g2_dfrbp_1 _1746_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net194),
    .D(net364),
    .Q_N(_0725_),
    .Q(\tt_um_mult_inst.pipe_out[18] ));
 sg13g2_dfrbp_1 _1747_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net195),
    .D(net378),
    .Q_N(_0726_),
    .Q(\tt_um_mult_inst.pipe_out[19] ));
 sg13g2_dfrbp_1 _1748_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net196),
    .D(net400),
    .Q_N(_0727_),
    .Q(\tt_um_mult_inst.pipe_out[20] ));
 sg13g2_dfrbp_1 _1749_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net197),
    .D(net372),
    .Q_N(_0728_),
    .Q(\tt_um_mult_inst.pipe_out[21] ));
 sg13g2_dfrbp_1 _1750_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net198),
    .D(net392),
    .Q_N(_0729_),
    .Q(\tt_um_mult_inst.pipe_out[22] ));
 sg13g2_dfrbp_1 _1751_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net199),
    .D(net360),
    .Q_N(_0730_),
    .Q(\tt_um_mult_inst.pipe_out[23] ));
 sg13g2_dfrbp_1 _1752_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net200),
    .D(net346),
    .Q_N(_0731_),
    .Q(\tt_um_mult_inst.pipe_out[24] ));
 sg13g2_dfrbp_1 _1753_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net201),
    .D(net344),
    .Q_N(_0732_),
    .Q(\tt_um_mult_inst.pipe_out[25] ));
 sg13g2_dfrbp_1 _1754_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net202),
    .D(net366),
    .Q_N(_0733_),
    .Q(\tt_um_mult_inst.pipe_out[26] ));
 sg13g2_dfrbp_1 _1755_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net203),
    .D(net388),
    .Q_N(_0734_),
    .Q(\tt_um_mult_inst.pipe_out[27] ));
 sg13g2_dfrbp_1 _1756_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net204),
    .D(net342),
    .Q_N(_0735_),
    .Q(\tt_um_mult_inst.pipe_out[28] ));
 sg13g2_dfrbp_1 _1757_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net205),
    .D(net394),
    .Q_N(_0736_),
    .Q(\tt_um_mult_inst.pipe_out[29] ));
 sg13g2_dfrbp_1 _1758_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net207),
    .D(net362),
    .Q_N(_0737_),
    .Q(\tt_um_mult_inst.pipe_out[30] ));
 sg13g2_dfrbp_1 _1759_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net37),
    .D(net354),
    .Q_N(_0595_),
    .Q(\tt_um_mult_inst.pipe_out[31] ));
 sg13g2_dfrbp_1 _1760_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net208),
    .D(net403),
    .Q_N(_0738_),
    .Q(state));
 sg13g2_dfrbp_1 _1761_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net209),
    .D(net432),
    .Q_N(_0739_),
    .Q(\tt_um_mult_inst.temp_out[0] ));
 sg13g2_dfrbp_1 _1762_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net210),
    .D(\tt_um_mult_inst.temp_out_comb[1] ),
    .Q_N(_0740_),
    .Q(\tt_um_mult_inst.temp_out[1] ));
 sg13g2_dfrbp_1 _1763_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net211),
    .D(\tt_um_mult_inst.temp_out_comb[2] ),
    .Q_N(_0741_),
    .Q(\tt_um_mult_inst.temp_out[2] ));
 sg13g2_dfrbp_1 _1764_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net212),
    .D(\tt_um_mult_inst.temp_out_comb[3] ),
    .Q_N(_0742_),
    .Q(\tt_um_mult_inst.temp_out[3] ));
 sg13g2_dfrbp_1 _1765_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net213),
    .D(\tt_um_mult_inst.temp_out_comb[4] ),
    .Q_N(_0743_),
    .Q(\tt_um_mult_inst.temp_out[4] ));
 sg13g2_dfrbp_1 _1766_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net214),
    .D(\tt_um_mult_inst.temp_out_comb[5] ),
    .Q_N(_0744_),
    .Q(\tt_um_mult_inst.temp_out[5] ));
 sg13g2_dfrbp_1 _1767_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net215),
    .D(\tt_um_mult_inst.temp_out_comb[6] ),
    .Q_N(_0745_),
    .Q(\tt_um_mult_inst.temp_out[6] ));
 sg13g2_dfrbp_1 _1768_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net216),
    .D(\tt_um_mult_inst.temp_out_comb[7] ),
    .Q_N(_0746_),
    .Q(\tt_um_mult_inst.temp_out[7] ));
 sg13g2_dfrbp_1 _1769_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net217),
    .D(\tt_um_mult_inst.temp_out_comb[8] ),
    .Q_N(_0747_),
    .Q(\tt_um_mult_inst.temp_out[8] ));
 sg13g2_dfrbp_1 _1770_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net218),
    .D(\tt_um_mult_inst.temp_out_comb[9] ),
    .Q_N(_0748_),
    .Q(\tt_um_mult_inst.temp_out[9] ));
 sg13g2_dfrbp_1 _1771_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net219),
    .D(\tt_um_mult_inst.temp_out_comb[10] ),
    .Q_N(_0749_),
    .Q(\tt_um_mult_inst.temp_out[10] ));
 sg13g2_dfrbp_1 _1772_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net220),
    .D(\tt_um_mult_inst.temp_out_comb[11] ),
    .Q_N(_0750_),
    .Q(\tt_um_mult_inst.temp_out[11] ));
 sg13g2_dfrbp_1 _1773_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net221),
    .D(\tt_um_mult_inst.temp_out_comb[12] ),
    .Q_N(_0751_),
    .Q(\tt_um_mult_inst.temp_out[12] ));
 sg13g2_dfrbp_1 _1774_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net222),
    .D(\tt_um_mult_inst.temp_out_comb[13] ),
    .Q_N(_0752_),
    .Q(\tt_um_mult_inst.temp_out[13] ));
 sg13g2_dfrbp_1 _1775_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net223),
    .D(\tt_um_mult_inst.temp_out_comb[14] ),
    .Q_N(_0753_),
    .Q(\tt_um_mult_inst.temp_out[14] ));
 sg13g2_dfrbp_1 _1776_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net224),
    .D(\tt_um_mult_inst.temp_out_comb[15] ),
    .Q_N(_0754_),
    .Q(\tt_um_mult_inst.temp_out[15] ));
 sg13g2_dfrbp_1 _1777_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net225),
    .D(\tt_um_mult_inst.temp_out_comb[16] ),
    .Q_N(_0755_),
    .Q(\tt_um_mult_inst.temp_out[16] ));
 sg13g2_dfrbp_1 _1778_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net226),
    .D(\tt_um_mult_inst.temp_out_comb[17] ),
    .Q_N(_0756_),
    .Q(\tt_um_mult_inst.temp_out[17] ));
 sg13g2_dfrbp_1 _1779_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net227),
    .D(\tt_um_mult_inst.temp_out_comb[18] ),
    .Q_N(_0757_),
    .Q(\tt_um_mult_inst.temp_out[18] ));
 sg13g2_dfrbp_1 _1780_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net228),
    .D(\tt_um_mult_inst.temp_out_comb[19] ),
    .Q_N(_0758_),
    .Q(\tt_um_mult_inst.temp_out[19] ));
 sg13g2_dfrbp_1 _1781_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net229),
    .D(\tt_um_mult_inst.temp_out_comb[20] ),
    .Q_N(_0759_),
    .Q(\tt_um_mult_inst.temp_out[20] ));
 sg13g2_dfrbp_1 _1782_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net230),
    .D(\tt_um_mult_inst.temp_out_comb[21] ),
    .Q_N(_0760_),
    .Q(\tt_um_mult_inst.temp_out[21] ));
 sg13g2_dfrbp_1 _1783_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net231),
    .D(\tt_um_mult_inst.temp_out_comb[22] ),
    .Q_N(_0761_),
    .Q(\tt_um_mult_inst.temp_out[22] ));
 sg13g2_dfrbp_1 _1784_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net232),
    .D(\tt_um_mult_inst.temp_out_comb[23] ),
    .Q_N(_0762_),
    .Q(\tt_um_mult_inst.temp_out[23] ));
 sg13g2_dfrbp_1 _1785_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net233),
    .D(\tt_um_mult_inst.temp_out_comb[24] ),
    .Q_N(_0763_),
    .Q(\tt_um_mult_inst.temp_out[24] ));
 sg13g2_dfrbp_1 _1786_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net234),
    .D(\tt_um_mult_inst.temp_out_comb[25] ),
    .Q_N(_0764_),
    .Q(\tt_um_mult_inst.temp_out[25] ));
 sg13g2_dfrbp_1 _1787_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net235),
    .D(\tt_um_mult_inst.temp_out_comb[26] ),
    .Q_N(_0765_),
    .Q(\tt_um_mult_inst.temp_out[26] ));
 sg13g2_dfrbp_1 _1788_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net236),
    .D(\tt_um_mult_inst.temp_out_comb[27] ),
    .Q_N(_0766_),
    .Q(\tt_um_mult_inst.temp_out[27] ));
 sg13g2_dfrbp_1 _1789_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net237),
    .D(\tt_um_mult_inst.temp_out_comb[28] ),
    .Q_N(_0767_),
    .Q(\tt_um_mult_inst.temp_out[28] ));
 sg13g2_dfrbp_1 _1790_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net238),
    .D(\tt_um_mult_inst.temp_out_comb[29] ),
    .Q_N(_0768_),
    .Q(\tt_um_mult_inst.temp_out[29] ));
 sg13g2_dfrbp_1 _1791_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net239),
    .D(\tt_um_mult_inst.temp_out_comb[30] ),
    .Q_N(_0769_),
    .Q(\tt_um_mult_inst.temp_out[30] ));
 sg13g2_dfrbp_1 _1792_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net240),
    .D(\tt_um_mult_inst.temp_out_comb[31] ),
    .Q_N(_0770_),
    .Q(\tt_um_mult_inst.temp_out[31] ));
 sg13g2_dfrbp_1 _1793_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net241),
    .D(\tt_um_mult_inst.temp_out_comb[32] ),
    .Q_N(_0771_),
    .Q(\tt_um_mult_inst.temp_out[32] ));
 sg13g2_dfrbp_1 _1794_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net242),
    .D(\tt_um_mult_inst.temp_out_comb[33] ),
    .Q_N(_0772_),
    .Q(\tt_um_mult_inst.temp_out[33] ));
 sg13g2_dfrbp_1 _1795_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net243),
    .D(\tt_um_mult_inst.temp_out_comb[34] ),
    .Q_N(_0773_),
    .Q(\tt_um_mult_inst.temp_out[34] ));
 sg13g2_dfrbp_1 _1796_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net244),
    .D(\tt_um_mult_inst.temp_out_comb[35] ),
    .Q_N(_0774_),
    .Q(\tt_um_mult_inst.temp_out[35] ));
 sg13g2_dfrbp_1 _1797_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net245),
    .D(\tt_um_mult_inst.temp_out_comb[36] ),
    .Q_N(_0775_),
    .Q(\tt_um_mult_inst.temp_out[36] ));
 sg13g2_dfrbp_1 _1798_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net246),
    .D(\tt_um_mult_inst.temp_out_comb[37] ),
    .Q_N(_0776_),
    .Q(\tt_um_mult_inst.temp_out[37] ));
 sg13g2_dfrbp_1 _1799_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net35),
    .D(\tt_um_mult_inst.temp_out_comb[38] ),
    .Q_N(_0777_),
    .Q(\tt_um_mult_inst.temp_out[38] ));
 sg13g2_dfrbp_1 _1800_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net36),
    .D(\tt_um_mult_inst.temp_out_comb[39] ),
    .Q_N(_0594_),
    .Q(\tt_um_mult_inst.temp_out[39] ));
 sg13g2_tiehi _1619__32 (.L_HI(net32));
 sg13g2_tiehi _1618__33 (.L_HI(net33));
 sg13g2_tiehi _1617__34 (.L_HI(net34));
 sg13g2_tiehi _1799__35 (.L_HI(net35));
 sg13g2_tiehi _1800__36 (.L_HI(net36));
 sg13g2_tiehi _1759__37 (.L_HI(net37));
 sg13g2_tiehi _1726__38 (.L_HI(net38));
 sg13g2_tiehi _1625__39 (.L_HI(net39));
 sg13g2_tiehi _1624__40 (.L_HI(net40));
 sg13g2_tiehi _1623__41 (.L_HI(net41));
 sg13g2_tiehi _1616__42 (.L_HI(net42));
 sg13g2_tiehi _1626__43 (.L_HI(net43));
 sg13g2_tiehi _1627__44 (.L_HI(net44));
 sg13g2_tiehi _1628__45 (.L_HI(net45));
 sg13g2_tiehi _1629__46 (.L_HI(net46));
 sg13g2_tiehi _1630__47 (.L_HI(net47));
 sg13g2_tiehi _1631__48 (.L_HI(net48));
 sg13g2_tiehi _1632__49 (.L_HI(net49));
 sg13g2_tiehi _1633__50 (.L_HI(net50));
 sg13g2_tiehi _1634__51 (.L_HI(net51));
 sg13g2_tiehi _1635__52 (.L_HI(net52));
 sg13g2_tiehi _1636__53 (.L_HI(net53));
 sg13g2_tiehi _1637__54 (.L_HI(net54));
 sg13g2_tiehi _1638__55 (.L_HI(net55));
 sg13g2_tiehi _1639__56 (.L_HI(net56));
 sg13g2_tiehi _1640__57 (.L_HI(net57));
 sg13g2_tiehi _1641__58 (.L_HI(net58));
 sg13g2_tiehi _1642__59 (.L_HI(net59));
 sg13g2_tiehi _1643__60 (.L_HI(net60));
 sg13g2_tiehi _1644__61 (.L_HI(net61));
 sg13g2_tiehi _1645__62 (.L_HI(net62));
 sg13g2_tiehi _1646__63 (.L_HI(net63));
 sg13g2_tiehi _1647__64 (.L_HI(net64));
 sg13g2_tiehi _1648__65 (.L_HI(net65));
 sg13g2_tiehi _1649__66 (.L_HI(net66));
 sg13g2_tiehi _1650__67 (.L_HI(net67));
 sg13g2_tiehi _1651__68 (.L_HI(net68));
 sg13g2_tiehi _1652__69 (.L_HI(net69));
 sg13g2_tiehi _1653__70 (.L_HI(net70));
 sg13g2_tiehi _1654__71 (.L_HI(net71));
 sg13g2_tiehi _1655__72 (.L_HI(net72));
 sg13g2_tiehi _1656__73 (.L_HI(net73));
 sg13g2_tiehi _1657__74 (.L_HI(net74));
 sg13g2_tiehi _1658__75 (.L_HI(net75));
 sg13g2_tiehi _1659__76 (.L_HI(net76));
 sg13g2_tiehi _1660__77 (.L_HI(net77));
 sg13g2_tiehi _1661__78 (.L_HI(net78));
 sg13g2_tiehi _1662__79 (.L_HI(net79));
 sg13g2_tiehi _1663__80 (.L_HI(net80));
 sg13g2_tiehi _1664__81 (.L_HI(net81));
 sg13g2_tiehi _1665__82 (.L_HI(net82));
 sg13g2_tiehi _1666__83 (.L_HI(net83));
 sg13g2_tiehi _1667__84 (.L_HI(net84));
 sg13g2_tiehi _1668__85 (.L_HI(net85));
 sg13g2_tiehi _1669__86 (.L_HI(net86));
 sg13g2_tiehi _1670__87 (.L_HI(net87));
 sg13g2_tiehi _1671__88 (.L_HI(net88));
 sg13g2_tiehi _1672__89 (.L_HI(net89));
 sg13g2_tiehi _1673__90 (.L_HI(net90));
 sg13g2_tiehi _1674__91 (.L_HI(net91));
 sg13g2_tiehi _1675__92 (.L_HI(net92));
 sg13g2_tiehi _1676__93 (.L_HI(net124));
 sg13g2_tiehi _1677__94 (.L_HI(net125));
 sg13g2_tiehi _1678__95 (.L_HI(net126));
 sg13g2_tiehi _1679__96 (.L_HI(net127));
 sg13g2_tiehi _1680__97 (.L_HI(net128));
 sg13g2_tiehi _1681__98 (.L_HI(net129));
 sg13g2_tiehi _1682__99 (.L_HI(net130));
 sg13g2_tiehi _1683__100 (.L_HI(net131));
 sg13g2_tiehi _1684__101 (.L_HI(net132));
 sg13g2_tiehi _1685__102 (.L_HI(net133));
 sg13g2_tiehi _1686__103 (.L_HI(net134));
 sg13g2_tiehi _1687__104 (.L_HI(net135));
 sg13g2_tiehi _1688__105 (.L_HI(net136));
 sg13g2_tiehi _1689__106 (.L_HI(net137));
 sg13g2_tiehi _1690__107 (.L_HI(net138));
 sg13g2_tiehi _1691__108 (.L_HI(net139));
 sg13g2_tiehi _1692__109 (.L_HI(net140));
 sg13g2_tiehi _1693__110 (.L_HI(net141));
 sg13g2_tiehi _1694__111 (.L_HI(net142));
 sg13g2_tiehi _1695__112 (.L_HI(net143));
 sg13g2_tiehi _1696__113 (.L_HI(net144));
 sg13g2_tiehi _1697__114 (.L_HI(net145));
 sg13g2_tiehi _1698__115 (.L_HI(net146));
 sg13g2_tiehi _1699__116 (.L_HI(net147));
 sg13g2_tiehi _1700__117 (.L_HI(net148));
 sg13g2_tiehi _1701__118 (.L_HI(net149));
 sg13g2_tiehi _1702__119 (.L_HI(net150));
 sg13g2_tiehi _1703__120 (.L_HI(net151));
 sg13g2_tiehi _1704__121 (.L_HI(net152));
 sg13g2_tiehi _1705__122 (.L_HI(net153));
 sg13g2_tiehi _1706__123 (.L_HI(net154));
 sg13g2_tiehi _1707__124 (.L_HI(net155));
 sg13g2_tiehi _1708__125 (.L_HI(net156));
 sg13g2_tiehi _1709__126 (.L_HI(net157));
 sg13g2_tiehi _1710__127 (.L_HI(net158));
 sg13g2_tiehi _1711__128 (.L_HI(net159));
 sg13g2_tiehi _1712__129 (.L_HI(net160));
 sg13g2_tiehi _1713__130 (.L_HI(net161));
 sg13g2_tiehi _1714__131 (.L_HI(net162));
 sg13g2_tiehi _1715__132 (.L_HI(net163));
 sg13g2_tiehi _1716__133 (.L_HI(net164));
 sg13g2_tiehi _1717__134 (.L_HI(net165));
 sg13g2_tiehi _1718__135 (.L_HI(net166));
 sg13g2_tiehi _1719__136 (.L_HI(net167));
 sg13g2_tiehi _1720__137 (.L_HI(net168));
 sg13g2_tiehi _1721__138 (.L_HI(net169));
 sg13g2_tiehi _1722__139 (.L_HI(net170));
 sg13g2_tiehi _1723__140 (.L_HI(net171));
 sg13g2_tiehi _1724__141 (.L_HI(net172));
 sg13g2_tiehi _1622__142 (.L_HI(net173));
 sg13g2_tiehi _1725__143 (.L_HI(net174));
 sg13g2_tiehi _1727__144 (.L_HI(net175));
 sg13g2_tiehi _1728__145 (.L_HI(net176));
 sg13g2_tiehi _1729__146 (.L_HI(net177));
 sg13g2_tiehi _1730__147 (.L_HI(net178));
 sg13g2_tiehi _1731__148 (.L_HI(net179));
 sg13g2_tiehi _1732__149 (.L_HI(net180));
 sg13g2_tiehi _1733__150 (.L_HI(net181));
 sg13g2_tiehi _1734__151 (.L_HI(net182));
 sg13g2_tiehi _1735__152 (.L_HI(net183));
 sg13g2_tiehi _1736__153 (.L_HI(net184));
 sg13g2_tiehi _1737__154 (.L_HI(net185));
 sg13g2_tiehi _1738__155 (.L_HI(net186));
 sg13g2_tiehi _1739__156 (.L_HI(net187));
 sg13g2_tiehi _1740__157 (.L_HI(net188));
 sg13g2_tiehi _1741__158 (.L_HI(net189));
 sg13g2_tiehi _1742__159 (.L_HI(net190));
 sg13g2_tiehi _1743__160 (.L_HI(net191));
 sg13g2_tiehi _1744__161 (.L_HI(net192));
 sg13g2_tiehi _1745__162 (.L_HI(net193));
 sg13g2_tiehi _1746__163 (.L_HI(net194));
 sg13g2_tiehi _1747__164 (.L_HI(net195));
 sg13g2_tiehi _1748__165 (.L_HI(net196));
 sg13g2_tiehi _1749__166 (.L_HI(net197));
 sg13g2_tiehi _1750__167 (.L_HI(net198));
 sg13g2_tiehi _1751__168 (.L_HI(net199));
 sg13g2_tiehi _1752__169 (.L_HI(net200));
 sg13g2_tiehi _1753__170 (.L_HI(net201));
 sg13g2_tiehi _1754__171 (.L_HI(net202));
 sg13g2_tiehi _1755__172 (.L_HI(net203));
 sg13g2_tiehi _1756__173 (.L_HI(net204));
 sg13g2_tiehi _1757__174 (.L_HI(net205));
 sg13g2_tiehi _1621__175 (.L_HI(net206));
 sg13g2_tiehi _1758__176 (.L_HI(net207));
 sg13g2_tiehi _1760__177 (.L_HI(net208));
 sg13g2_tiehi _1761__178 (.L_HI(net209));
 sg13g2_tiehi _1762__179 (.L_HI(net210));
 sg13g2_tiehi _1763__180 (.L_HI(net211));
 sg13g2_tiehi _1764__181 (.L_HI(net212));
 sg13g2_tiehi _1765__182 (.L_HI(net213));
 sg13g2_tiehi _1766__183 (.L_HI(net214));
 sg13g2_tiehi _1767__184 (.L_HI(net215));
 sg13g2_tiehi _1768__185 (.L_HI(net216));
 sg13g2_tiehi _1769__186 (.L_HI(net217));
 sg13g2_tiehi _1770__187 (.L_HI(net218));
 sg13g2_tiehi _1771__188 (.L_HI(net219));
 sg13g2_tiehi _1772__189 (.L_HI(net220));
 sg13g2_tiehi _1773__190 (.L_HI(net221));
 sg13g2_tiehi _1774__191 (.L_HI(net222));
 sg13g2_tiehi _1775__192 (.L_HI(net223));
 sg13g2_tiehi _1776__193 (.L_HI(net224));
 sg13g2_tiehi _1777__194 (.L_HI(net225));
 sg13g2_tiehi _1778__195 (.L_HI(net226));
 sg13g2_tiehi _1779__196 (.L_HI(net227));
 sg13g2_tiehi _1780__197 (.L_HI(net228));
 sg13g2_tiehi _1781__198 (.L_HI(net229));
 sg13g2_tiehi _1782__199 (.L_HI(net230));
 sg13g2_tiehi _1783__200 (.L_HI(net231));
 sg13g2_tiehi _1784__201 (.L_HI(net232));
 sg13g2_tiehi _1785__202 (.L_HI(net233));
 sg13g2_tiehi _1786__203 (.L_HI(net234));
 sg13g2_tiehi _1787__204 (.L_HI(net235));
 sg13g2_tiehi _1788__205 (.L_HI(net236));
 sg13g2_tiehi _1789__206 (.L_HI(net237));
 sg13g2_tiehi _1790__207 (.L_HI(net238));
 sg13g2_tiehi _1791__208 (.L_HI(net239));
 sg13g2_tiehi _1792__209 (.L_HI(net240));
 sg13g2_tiehi _1793__210 (.L_HI(net241));
 sg13g2_tiehi _1794__211 (.L_HI(net242));
 sg13g2_tiehi _1795__212 (.L_HI(net243));
 sg13g2_tiehi _1796__213 (.L_HI(net244));
 sg13g2_tiehi _1797__214 (.L_HI(net245));
 sg13g2_tiehi _1798__215 (.L_HI(net246));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_16 (.L_LO(net16));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_17 (.L_LO(net17));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_18 (.L_LO(net18));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_19 (.L_LO(net19));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_20 (.L_LO(net20));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_21 (.L_LO(net21));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_22 (.L_LO(net22));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_23 (.L_LO(net23));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_24 (.L_LO(net24));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_25 (.L_LO(net25));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_26 (.L_LO(net26));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_27 (.L_LO(net27));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_28 (.L_LO(net28));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_29 (.L_LO(net29));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_30 (.L_LO(net30));
 sg13g2_tiehi _1620__31 (.L_HI(net31));
 sg13g2_buf_1 _2002_ (.A(\tt_um_mult_inst.pipe_out[0] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _2003_ (.A(\tt_um_mult_inst.pipe_out[1] ),
    .X(uo_out[1]));
 sg13g2_buf_1 _2004_ (.A(\tt_um_mult_inst.pipe_out[2] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _2005_ (.A(\tt_um_mult_inst.pipe_out[3] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _2006_ (.A(\tt_um_mult_inst.pipe_out[4] ),
    .X(uo_out[4]));
 sg13g2_buf_1 _2007_ (.A(\tt_um_mult_inst.pipe_out[5] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _2008_ (.A(\tt_um_mult_inst.pipe_out[6] ),
    .X(uo_out[6]));
 sg13g2_buf_1 _2009_ (.A(\tt_um_mult_inst.pipe_out[7] ),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout93 (.X(net93),
    .A(_0057_));
 sg13g2_buf_2 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_4 fanout95 (.X(net95),
    .A(_0057_));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(net98));
 sg13g2_buf_2 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_0057_),
    .X(net98));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(net101));
 sg13g2_buf_4 fanout100 (.X(net100),
    .A(net101));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(net106));
 sg13g2_buf_2 fanout102 (.A(net103),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(net106),
    .X(net103));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(net105));
 sg13g2_buf_2 fanout105 (.A(net106),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_0056_),
    .X(net106));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(net108));
 sg13g2_buf_2 fanout108 (.A(_0054_),
    .X(net108));
 sg13g2_buf_4 fanout109 (.X(net109),
    .A(state));
 sg13g2_buf_1 fanout110 (.A(state),
    .X(net110));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(net13));
 sg13g2_buf_2 fanout112 (.A(net12),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(net11),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(net10),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(net9),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(net9),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(net118),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(uio_in[1]),
    .X(net118));
 sg13g2_buf_4 fanout119 (.X(net119),
    .A(net8));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(net121));
 sg13g2_buf_2 fanout121 (.A(ui_in[1]),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(ui_in[0]),
    .X(net122));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(ui_in[0]));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[2]));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[3]));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[4]));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[5]));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[6]));
 sg13g2_buf_4 input7 (.X(net7),
    .A(ui_in[7]));
 sg13g2_buf_2 input8 (.A(uio_in[0]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[6]),
    .X(net13));
 sg13g2_buf_4 input14 (.X(net14),
    .A(uio_in[7]));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_15 (.L_LO(net15));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\tt_um_load_inst.weights[49] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold2 (.A(\tt_um_load_inst.weights[40] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold3 (.A(\tt_um_load_inst.weights[65] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold4 (.A(\tt_um_load_inst.weights[57] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold5 (.A(\tt_um_load_inst.weights[34] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold6 (.A(\tt_um_load_inst.weights[47] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold7 (.A(\tt_um_load_inst.weights[25] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold8 (.A(\tt_um_load_inst.weights[28] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold9 (.A(\tt_um_load_inst.weights[23] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold10 (.A(\tt_um_load_inst.weights[20] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold11 (.A(\tt_um_load_inst.weights[29] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold12 (.A(\tt_um_load_inst.weights[82] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold13 (.A(\tt_um_load_inst.weights[88] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold14 (.A(\tt_um_load_inst.weights[60] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold15 (.A(\tt_um_load_inst.weights[45] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold16 (.A(\tt_um_load_inst.weights[71] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold17 (.A(\tt_um_load_inst.weights[22] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold18 (.A(\tt_um_load_inst.weights[99] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold19 (.A(\tt_um_load_inst.weights[92] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold20 (.A(\tt_um_load_inst.weights[95] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold21 (.A(\tt_um_load_inst.weights[74] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold22 (.A(\tt_um_load_inst.weights[84] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold23 (.A(\tt_um_load_inst.weights[98] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold24 (.A(\tt_um_load_inst.weights[76] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold25 (.A(\tt_um_load_inst.weights[62] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold26 (.A(\tt_um_load_inst.weights[43] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold27 (.A(\tt_um_load_inst.weights[86] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold28 (.A(\tt_um_load_inst.weights[41] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold29 (.A(\tt_um_load_inst.weights[56] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold30 (.A(\tt_um_load_inst.weights[46] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold31 (.A(\tt_um_load_inst.weights[24] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold32 (.A(\tt_um_load_inst.weights[44] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold33 (.A(\tt_um_load_inst.weights[96] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold34 (.A(\tt_um_load_inst.weights[66] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold35 (.A(\tt_um_load_inst.weights[54] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold36 (.A(\tt_um_load_inst.weights[63] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold37 (.A(\tt_um_load_inst.weights[97] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold38 (.A(\tt_um_load_inst.weights[64] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold39 (.A(\tt_um_load_inst.weights[36] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold40 (.A(\tt_um_load_inst.weights[26] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold41 (.A(\tt_um_load_inst.weights[27] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold42 (.A(\tt_um_load_inst.weights[33] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold43 (.A(\tt_um_load_inst.weights[85] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold44 (.A(\tt_um_load_inst.weights[52] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold45 (.A(\tt_um_load_inst.weights[21] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold46 (.A(\tt_um_load_inst.weights[80] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold47 (.A(\tt_um_load_inst.weights[35] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold48 (.A(\tt_um_load_inst.weights[67] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold49 (.A(\tt_um_load_inst.weights[70] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold50 (.A(\tt_um_load_inst.weights[61] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold51 (.A(\tt_um_load_inst.weights[39] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold52 (.A(\tt_um_load_inst.weights[93] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold53 (.A(\tt_um_load_inst.weights[68] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold54 (.A(\tt_um_load_inst.weights[72] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold55 (.A(\tt_um_load_inst.weights[32] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold56 (.A(\tt_um_load_inst.weights[75] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold57 (.A(\tt_um_load_inst.weights[79] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold58 (.A(\tt_um_load_inst.weights[89] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold59 (.A(\tt_um_load_inst.weights[38] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold60 (.A(\tt_um_load_inst.weights[87] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold61 (.A(\tt_um_load_inst.weights[50] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold62 (.A(\tt_um_load_inst.weights[78] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold63 (.A(\tt_um_load_inst.weights[53] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold64 (.A(\tt_um_load_inst.weights[51] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold65 (.A(\tt_um_load_inst.weights[30] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold66 (.A(\tt_um_load_inst.weights[37] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold67 (.A(\tt_um_load_inst.weights[31] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold68 (.A(\tt_um_load_inst.weights[83] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold69 (.A(\tt_um_load_inst.weights[77] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold70 (.A(\tt_um_load_inst.weights[73] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold71 (.A(\tt_um_load_inst.weights[42] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold72 (.A(\tt_um_load_inst.weights[48] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold73 (.A(\tt_um_load_inst.weights[90] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold74 (.A(\tt_um_load_inst.weights[81] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold75 (.A(\tt_um_load_inst.weights[94] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold76 (.A(\tt_um_load_inst.weights[58] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold77 (.A(\tt_um_load_inst.weights[55] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold78 (.A(\tt_um_load_inst.weights[69] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold79 (.A(\tt_um_load_inst.weights[91] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold80 (.A(\tt_um_load_inst.weights[59] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0032_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0044_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold83 (.A(\tt_um_mult_inst.temp_out[36] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold84 (.A(\tt_um_mult_inst.temp_out[37] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold85 (.A(\tt_um_mult_inst.temp_out[33] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold86 (.A(\tt_um_mult_inst.temp_out[38] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold87 (.A(\tt_um_mult_inst.temp_out[39] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold88 (.A(\tt_um_mult_inst.pipe_out[20] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0003_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold90 (.A(\tt_um_mult_inst.temp_out[32] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold91 (.A(\tt_um_mult_inst.temp_out[34] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold92 (.A(\tt_um_mult_inst.temp_out[35] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold93 (.A(\tt_um_mult_inst.pipe_out[13] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0027_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold95 (.A(\tt_um_mult_inst.pipe_out[36] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0020_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold97 (.A(\tt_um_mult_inst.pipe_out[33] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0017_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold99 (.A(\tt_um_mult_inst.pipe_out[32] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0016_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold101 (.A(\tt_um_mult_inst.pipe_out[15] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0029_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold103 (.A(\tt_um_mult_inst.pipe_out[12] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0026_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold105 (.A(\tt_um_mult_inst.pipe_out[22] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0005_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold107 (.A(\tt_um_mult_inst.pipe_out[39] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0024_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold109 (.A(\tt_um_mult_inst.pipe_out[14] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0028_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold111 (.A(\tt_um_mult_inst.pipe_out[11] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0025_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold113 (.A(\tt_um_mult_inst.pipe_out[31] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0015_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold115 (.A(\tt_um_mult_inst.pipe_out[38] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0023_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold117 (.A(\tt_um_mult_inst.pipe_out[26] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0009_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold119 (.A(\tt_um_mult_inst.pipe_out[34] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0018_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold121 (.A(\tt_um_mult_inst.pipe_out[17] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0031_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold123 (.A(\tt_um_mult_inst.pipe_out[24] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0007_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold125 (.A(\tt_um_mult_inst.pipe_out[29] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0013_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold127 (.A(\tt_um_mult_inst.pipe_out[21] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0004_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold129 (.A(\tt_um_mult_inst.pipe_out[9] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0011_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold131 (.A(\tt_um_mult_inst.pipe_out[27] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0010_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold133 (.A(\tt_um_mult_inst.pipe_out[8] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0000_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold135 (.A(\tt_um_mult_inst.pipe_out[23] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0006_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold137 (.A(\tt_um_mult_inst.pipe_out[25] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0008_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold139 (.A(\tt_um_mult_inst.pipe_out[10] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0022_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold141 (.A(\tt_um_mult_inst.pipe_out[35] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0019_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold143 (.A(\tt_um_mult_inst.temp_out[8] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0030_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold145 (.A(\tt_um_mult_inst.pipe_out[30] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0014_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold147 (.A(\tt_um_mult_inst.pipe_out[37] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0021_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold149 (.A(\tt_um_mult_inst.pipe_out[18] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0001_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold151 (.A(\tt_um_mult_inst.pipe_out[19] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0002_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold153 (.A(\tt_um_mult_inst.temp_out[20] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0012_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold155 (.A(\count[2] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0593_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0045_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold158 (.A(\count[1] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0587_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold160 (.A(\count[3] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0043_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold162 (.A(\load_weights[13] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold163 (.A(\tt_um_load_inst.input_to_sr[13] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold164 (.A(\load_weights[19] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold165 (.A(\tt_um_load_inst.input_to_sr[19] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold166 (.A(\load_weights[15] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold167 (.A(\tt_um_load_inst.input_to_sr[15] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold168 (.A(\load_weights[8] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold169 (.A(\load_weights[9] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold170 (.A(\load_weights[17] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold171 (.A(\tt_um_load_inst.input_to_sr[17] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold172 (.A(\count[0] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold173 (.A(\load_weights[11] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold174 (.A(\tt_um_load_inst.input_to_sr[11] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold175 (.A(\load_weights[10] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold176 (.A(\tt_um_load_inst.input_to_sr[10] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold177 (.A(\load_weights[7] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold178 (.A(\load_weights[12] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold179 (.A(\tt_um_load_inst.input_to_sr[12] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold180 (.A(\load_weights[3] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold181 (.A(\load_weights[18] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold182 (.A(\tt_um_load_inst.input_to_sr[18] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold183 (.A(\load_weights[5] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold184 (.A(\load_weights[2] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold185 (.A(\load_weights[0] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold186 (.A(\tt_um_mult_inst.temp_out_comb[0] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold187 (.A(\load_weights[6] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold188 (.A(\load_weights[12] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold189 (.A(\load_weights[4] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold190 (.A(\load_weights[16] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold191 (.A(\tt_um_load_inst.input_to_sr[16] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold192 (.A(\tt_um_mult_inst.temp_out[24] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold193 (.A(\load_weights[1] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold194 (.A(\load_weights[14] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold195 (.A(\tt_um_load_inst.input_to_sr[14] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold196 (.A(\tt_um_mult_inst.temp_out[16] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold197 (.A(\tt_um_mult_inst.temp_out[15] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold198 (.A(\tt_um_mult_inst.temp_out[0] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold199 (.A(\tt_um_mult_inst.temp_out[23] ),
    .X(net445));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_fill_1 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_255 ();
 sg13g2_decap_8 FILLER_1_262 ();
 sg13g2_fill_2 FILLER_1_269 ();
 sg13g2_fill_1 FILLER_1_271 ();
 sg13g2_decap_8 FILLER_1_281 ();
 sg13g2_decap_8 FILLER_1_288 ();
 sg13g2_decap_8 FILLER_1_295 ();
 sg13g2_decap_8 FILLER_1_302 ();
 sg13g2_decap_8 FILLER_1_309 ();
 sg13g2_decap_8 FILLER_1_316 ();
 sg13g2_decap_8 FILLER_1_323 ();
 sg13g2_decap_8 FILLER_1_330 ();
 sg13g2_decap_8 FILLER_1_337 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_fill_2 FILLER_2_217 ();
 sg13g2_fill_1 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_307 ();
 sg13g2_decap_8 FILLER_2_314 ();
 sg13g2_decap_8 FILLER_2_321 ();
 sg13g2_decap_8 FILLER_2_328 ();
 sg13g2_decap_8 FILLER_2_335 ();
 sg13g2_decap_8 FILLER_2_342 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_4 FILLER_3_105 ();
 sg13g2_fill_2 FILLER_3_109 ();
 sg13g2_fill_2 FILLER_3_155 ();
 sg13g2_decap_8 FILLER_3_166 ();
 sg13g2_decap_8 FILLER_3_173 ();
 sg13g2_decap_8 FILLER_3_180 ();
 sg13g2_decap_4 FILLER_3_187 ();
 sg13g2_fill_1 FILLER_3_191 ();
 sg13g2_fill_1 FILLER_3_218 ();
 sg13g2_decap_4 FILLER_3_245 ();
 sg13g2_fill_1 FILLER_3_257 ();
 sg13g2_fill_1 FILLER_3_272 ();
 sg13g2_fill_2 FILLER_3_281 ();
 sg13g2_fill_1 FILLER_3_283 ();
 sg13g2_decap_8 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_330 ();
 sg13g2_decap_8 FILLER_3_337 ();
 sg13g2_decap_8 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_351 ();
 sg13g2_decap_8 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_fill_1 FILLER_4_98 ();
 sg13g2_decap_4 FILLER_4_125 ();
 sg13g2_fill_2 FILLER_4_129 ();
 sg13g2_decap_4 FILLER_4_196 ();
 sg13g2_fill_2 FILLER_4_200 ();
 sg13g2_decap_8 FILLER_4_323 ();
 sg13g2_decap_8 FILLER_4_330 ();
 sg13g2_decap_8 FILLER_4_337 ();
 sg13g2_decap_8 FILLER_4_344 ();
 sg13g2_decap_8 FILLER_4_351 ();
 sg13g2_decap_8 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_365 ();
 sg13g2_decap_8 FILLER_4_372 ();
 sg13g2_decap_8 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_386 ();
 sg13g2_decap_8 FILLER_4_393 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_4 FILLER_5_49 ();
 sg13g2_fill_2 FILLER_5_53 ();
 sg13g2_decap_4 FILLER_5_81 ();
 sg13g2_decap_4 FILLER_5_89 ();
 sg13g2_fill_1 FILLER_5_93 ();
 sg13g2_fill_1 FILLER_5_108 ();
 sg13g2_fill_2 FILLER_5_117 ();
 sg13g2_fill_1 FILLER_5_119 ();
 sg13g2_fill_2 FILLER_5_129 ();
 sg13g2_decap_8 FILLER_5_135 ();
 sg13g2_decap_4 FILLER_5_142 ();
 sg13g2_decap_8 FILLER_5_159 ();
 sg13g2_fill_2 FILLER_5_166 ();
 sg13g2_fill_2 FILLER_5_172 ();
 sg13g2_fill_1 FILLER_5_174 ();
 sg13g2_decap_4 FILLER_5_201 ();
 sg13g2_fill_1 FILLER_5_205 ();
 sg13g2_fill_2 FILLER_5_232 ();
 sg13g2_fill_1 FILLER_5_234 ();
 sg13g2_fill_1 FILLER_5_261 ();
 sg13g2_fill_1 FILLER_5_288 ();
 sg13g2_fill_2 FILLER_5_307 ();
 sg13g2_decap_8 FILLER_5_335 ();
 sg13g2_decap_8 FILLER_5_342 ();
 sg13g2_decap_8 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_356 ();
 sg13g2_decap_8 FILLER_5_363 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_4 FILLER_6_49 ();
 sg13g2_fill_2 FILLER_6_53 ();
 sg13g2_decap_8 FILLER_6_172 ();
 sg13g2_fill_1 FILLER_6_179 ();
 sg13g2_fill_2 FILLER_6_232 ();
 sg13g2_fill_2 FILLER_6_243 ();
 sg13g2_fill_1 FILLER_6_245 ();
 sg13g2_fill_2 FILLER_6_286 ();
 sg13g2_fill_1 FILLER_6_288 ();
 sg13g2_fill_1 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_324 ();
 sg13g2_decap_8 FILLER_6_331 ();
 sg13g2_decap_8 FILLER_6_338 ();
 sg13g2_decap_8 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_352 ();
 sg13g2_decap_8 FILLER_6_359 ();
 sg13g2_decap_8 FILLER_6_366 ();
 sg13g2_decap_8 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_fill_1 FILLER_7_58 ();
 sg13g2_decap_4 FILLER_7_68 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_fill_1 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_89 ();
 sg13g2_fill_1 FILLER_7_96 ();
 sg13g2_fill_2 FILLER_7_106 ();
 sg13g2_fill_1 FILLER_7_108 ();
 sg13g2_decap_8 FILLER_7_113 ();
 sg13g2_fill_2 FILLER_7_120 ();
 sg13g2_fill_1 FILLER_7_122 ();
 sg13g2_fill_1 FILLER_7_132 ();
 sg13g2_decap_4 FILLER_7_146 ();
 sg13g2_fill_1 FILLER_7_150 ();
 sg13g2_fill_2 FILLER_7_179 ();
 sg13g2_fill_1 FILLER_7_191 ();
 sg13g2_fill_2 FILLER_7_196 ();
 sg13g2_decap_4 FILLER_7_208 ();
 sg13g2_fill_2 FILLER_7_212 ();
 sg13g2_fill_2 FILLER_7_240 ();
 sg13g2_fill_1 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_325 ();
 sg13g2_decap_8 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_346 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_fill_2 FILLER_8_42 ();
 sg13g2_fill_1 FILLER_8_44 ();
 sg13g2_fill_2 FILLER_8_158 ();
 sg13g2_fill_2 FILLER_8_184 ();
 sg13g2_fill_1 FILLER_8_186 ();
 sg13g2_decap_4 FILLER_8_196 ();
 sg13g2_fill_2 FILLER_8_200 ();
 sg13g2_fill_2 FILLER_8_212 ();
 sg13g2_fill_1 FILLER_8_214 ();
 sg13g2_fill_1 FILLER_8_291 ();
 sg13g2_fill_2 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_37 ();
 sg13g2_decap_8 FILLER_9_44 ();
 sg13g2_fill_1 FILLER_9_55 ();
 sg13g2_fill_1 FILLER_9_183 ();
 sg13g2_fill_1 FILLER_9_262 ();
 sg13g2_fill_1 FILLER_9_289 ();
 sg13g2_fill_2 FILLER_9_337 ();
 sg13g2_decap_8 FILLER_9_348 ();
 sg13g2_decap_8 FILLER_9_355 ();
 sg13g2_decap_8 FILLER_9_362 ();
 sg13g2_decap_8 FILLER_9_369 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_119 ();
 sg13g2_decap_4 FILLER_10_143 ();
 sg13g2_fill_1 FILLER_10_147 ();
 sg13g2_fill_2 FILLER_10_153 ();
 sg13g2_decap_4 FILLER_10_174 ();
 sg13g2_decap_4 FILLER_10_188 ();
 sg13g2_fill_1 FILLER_10_264 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_4 FILLER_11_26 ();
 sg13g2_fill_1 FILLER_11_30 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_fill_2 FILLER_11_49 ();
 sg13g2_fill_1 FILLER_11_51 ();
 sg13g2_fill_2 FILLER_11_83 ();
 sg13g2_fill_1 FILLER_11_85 ();
 sg13g2_fill_1 FILLER_11_90 ();
 sg13g2_decap_8 FILLER_11_169 ();
 sg13g2_fill_1 FILLER_11_289 ();
 sg13g2_fill_2 FILLER_11_316 ();
 sg13g2_fill_1 FILLER_11_318 ();
 sg13g2_fill_1 FILLER_11_328 ();
 sg13g2_decap_8 FILLER_11_334 ();
 sg13g2_fill_2 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_fill_2 FILLER_11_396 ();
 sg13g2_fill_1 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_48 ();
 sg13g2_decap_4 FILLER_12_89 ();
 sg13g2_fill_1 FILLER_12_111 ();
 sg13g2_fill_2 FILLER_12_156 ();
 sg13g2_fill_2 FILLER_12_168 ();
 sg13g2_fill_1 FILLER_12_170 ();
 sg13g2_fill_2 FILLER_12_197 ();
 sg13g2_fill_2 FILLER_12_211 ();
 sg13g2_fill_1 FILLER_12_221 ();
 sg13g2_fill_1 FILLER_12_248 ();
 sg13g2_fill_1 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_307 ();
 sg13g2_decap_4 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_4 FILLER_12_391 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_10 ();
 sg13g2_decap_4 FILLER_13_15 ();
 sg13g2_fill_2 FILLER_13_19 ();
 sg13g2_fill_2 FILLER_13_30 ();
 sg13g2_fill_1 FILLER_13_32 ();
 sg13g2_fill_2 FILLER_13_68 ();
 sg13g2_fill_1 FILLER_13_70 ();
 sg13g2_fill_2 FILLER_13_133 ();
 sg13g2_decap_4 FILLER_13_165 ();
 sg13g2_fill_2 FILLER_13_186 ();
 sg13g2_fill_1 FILLER_13_188 ();
 sg13g2_decap_4 FILLER_13_233 ();
 sg13g2_fill_2 FILLER_13_241 ();
 sg13g2_fill_2 FILLER_13_269 ();
 sg13g2_fill_2 FILLER_13_290 ();
 sg13g2_fill_1 FILLER_13_296 ();
 sg13g2_fill_2 FILLER_13_327 ();
 sg13g2_fill_1 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_334 ();
 sg13g2_decap_4 FILLER_13_341 ();
 sg13g2_fill_2 FILLER_13_358 ();
 sg13g2_fill_1 FILLER_13_377 ();
 sg13g2_fill_1 FILLER_14_26 ();
 sg13g2_fill_2 FILLER_14_31 ();
 sg13g2_fill_1 FILLER_14_33 ();
 sg13g2_decap_8 FILLER_14_47 ();
 sg13g2_fill_2 FILLER_14_54 ();
 sg13g2_fill_2 FILLER_14_76 ();
 sg13g2_fill_1 FILLER_14_78 ();
 sg13g2_fill_2 FILLER_14_93 ();
 sg13g2_fill_1 FILLER_14_95 ();
 sg13g2_fill_2 FILLER_14_104 ();
 sg13g2_fill_1 FILLER_14_106 ();
 sg13g2_decap_4 FILLER_14_111 ();
 sg13g2_fill_2 FILLER_14_115 ();
 sg13g2_fill_1 FILLER_14_138 ();
 sg13g2_decap_4 FILLER_14_156 ();
 sg13g2_fill_1 FILLER_14_176 ();
 sg13g2_decap_4 FILLER_14_193 ();
 sg13g2_fill_2 FILLER_14_213 ();
 sg13g2_fill_1 FILLER_14_230 ();
 sg13g2_decap_4 FILLER_14_239 ();
 sg13g2_fill_2 FILLER_14_243 ();
 sg13g2_fill_1 FILLER_14_258 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_1 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_15 ();
 sg13g2_decap_4 FILLER_15_22 ();
 sg13g2_fill_2 FILLER_15_52 ();
 sg13g2_fill_2 FILLER_15_74 ();
 sg13g2_fill_2 FILLER_15_88 ();
 sg13g2_fill_1 FILLER_15_90 ();
 sg13g2_fill_1 FILLER_15_111 ();
 sg13g2_fill_1 FILLER_15_132 ();
 sg13g2_decap_8 FILLER_15_141 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_decap_8 FILLER_15_176 ();
 sg13g2_decap_8 FILLER_15_183 ();
 sg13g2_fill_2 FILLER_15_190 ();
 sg13g2_fill_1 FILLER_15_192 ();
 sg13g2_fill_1 FILLER_15_227 ();
 sg13g2_fill_2 FILLER_15_236 ();
 sg13g2_fill_1 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_247 ();
 sg13g2_fill_1 FILLER_15_294 ();
 sg13g2_fill_2 FILLER_15_309 ();
 sg13g2_fill_1 FILLER_15_346 ();
 sg13g2_fill_2 FILLER_15_369 ();
 sg13g2_fill_2 FILLER_15_380 ();
 sg13g2_fill_1 FILLER_15_382 ();
 sg13g2_decap_4 FILLER_16_26 ();
 sg13g2_fill_1 FILLER_16_30 ();
 sg13g2_fill_2 FILLER_16_54 ();
 sg13g2_fill_1 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_87 ();
 sg13g2_fill_1 FILLER_16_94 ();
 sg13g2_decap_8 FILLER_16_100 ();
 sg13g2_decap_8 FILLER_16_107 ();
 sg13g2_fill_2 FILLER_16_114 ();
 sg13g2_fill_2 FILLER_16_139 ();
 sg13g2_decap_8 FILLER_16_158 ();
 sg13g2_fill_2 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_191 ();
 sg13g2_decap_8 FILLER_16_216 ();
 sg13g2_decap_4 FILLER_16_236 ();
 sg13g2_fill_2 FILLER_16_240 ();
 sg13g2_decap_8 FILLER_16_255 ();
 sg13g2_fill_1 FILLER_16_274 ();
 sg13g2_fill_1 FILLER_16_315 ();
 sg13g2_fill_2 FILLER_16_397 ();
 sg13g2_fill_1 FILLER_16_399 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_4 ();
 sg13g2_decap_8 FILLER_17_58 ();
 sg13g2_fill_2 FILLER_17_65 ();
 sg13g2_decap_8 FILLER_17_94 ();
 sg13g2_fill_2 FILLER_17_101 ();
 sg13g2_fill_1 FILLER_17_123 ();
 sg13g2_fill_1 FILLER_17_164 ();
 sg13g2_decap_4 FILLER_17_170 ();
 sg13g2_fill_1 FILLER_17_196 ();
 sg13g2_decap_4 FILLER_17_218 ();
 sg13g2_fill_1 FILLER_17_231 ();
 sg13g2_fill_2 FILLER_17_248 ();
 sg13g2_fill_1 FILLER_17_250 ();
 sg13g2_fill_2 FILLER_17_286 ();
 sg13g2_fill_1 FILLER_17_298 ();
 sg13g2_fill_1 FILLER_17_345 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_4 ();
 sg13g2_decap_4 FILLER_18_36 ();
 sg13g2_fill_2 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_71 ();
 sg13g2_decap_8 FILLER_18_83 ();
 sg13g2_fill_1 FILLER_18_90 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_fill_1 FILLER_18_112 ();
 sg13g2_decap_4 FILLER_18_127 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_decap_8 FILLER_18_136 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_fill_1 FILLER_18_150 ();
 sg13g2_decap_8 FILLER_18_160 ();
 sg13g2_decap_8 FILLER_18_167 ();
 sg13g2_fill_2 FILLER_18_174 ();
 sg13g2_fill_1 FILLER_18_176 ();
 sg13g2_decap_8 FILLER_18_191 ();
 sg13g2_fill_2 FILLER_18_198 ();
 sg13g2_fill_1 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_240 ();
 sg13g2_decap_4 FILLER_18_269 ();
 sg13g2_fill_2 FILLER_18_299 ();
 sg13g2_fill_2 FILLER_18_332 ();
 sg13g2_fill_1 FILLER_18_334 ();
 sg13g2_fill_1 FILLER_18_342 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_36 ();
 sg13g2_fill_2 FILLER_19_54 ();
 sg13g2_fill_1 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_78 ();
 sg13g2_decap_4 FILLER_19_85 ();
 sg13g2_fill_2 FILLER_19_89 ();
 sg13g2_decap_8 FILLER_19_95 ();
 sg13g2_fill_1 FILLER_19_122 ();
 sg13g2_decap_4 FILLER_19_132 ();
 sg13g2_fill_2 FILLER_19_136 ();
 sg13g2_fill_2 FILLER_19_144 ();
 sg13g2_fill_2 FILLER_19_164 ();
 sg13g2_decap_4 FILLER_19_176 ();
 sg13g2_fill_2 FILLER_19_192 ();
 sg13g2_fill_1 FILLER_19_194 ();
 sg13g2_decap_4 FILLER_19_212 ();
 sg13g2_fill_1 FILLER_19_216 ();
 sg13g2_fill_1 FILLER_19_250 ();
 sg13g2_decap_8 FILLER_19_270 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_fill_2 FILLER_19_291 ();
 sg13g2_decap_8 FILLER_19_299 ();
 sg13g2_decap_4 FILLER_19_306 ();
 sg13g2_fill_1 FILLER_19_310 ();
 sg13g2_fill_2 FILLER_19_324 ();
 sg13g2_fill_1 FILLER_19_326 ();
 sg13g2_fill_2 FILLER_19_351 ();
 sg13g2_fill_2 FILLER_19_362 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_58 ();
 sg13g2_decap_4 FILLER_20_73 ();
 sg13g2_fill_1 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_82 ();
 sg13g2_decap_4 FILLER_20_89 ();
 sg13g2_fill_2 FILLER_20_99 ();
 sg13g2_fill_1 FILLER_20_101 ();
 sg13g2_fill_2 FILLER_20_132 ();
 sg13g2_fill_2 FILLER_20_148 ();
 sg13g2_fill_1 FILLER_20_150 ();
 sg13g2_decap_8 FILLER_20_165 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_fill_2 FILLER_20_179 ();
 sg13g2_decap_4 FILLER_20_224 ();
 sg13g2_fill_2 FILLER_20_240 ();
 sg13g2_fill_1 FILLER_20_242 ();
 sg13g2_fill_2 FILLER_20_316 ();
 sg13g2_fill_1 FILLER_20_335 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_43 ();
 sg13g2_fill_2 FILLER_21_50 ();
 sg13g2_fill_1 FILLER_21_52 ();
 sg13g2_fill_1 FILLER_21_66 ();
 sg13g2_fill_2 FILLER_21_117 ();
 sg13g2_fill_1 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_136 ();
 sg13g2_fill_2 FILLER_21_143 ();
 sg13g2_decap_4 FILLER_21_149 ();
 sg13g2_fill_2 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_167 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_4 FILLER_21_196 ();
 sg13g2_fill_2 FILLER_21_210 ();
 sg13g2_decap_4 FILLER_21_248 ();
 sg13g2_fill_2 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_270 ();
 sg13g2_decap_4 FILLER_21_277 ();
 sg13g2_fill_2 FILLER_21_281 ();
 sg13g2_fill_2 FILLER_21_287 ();
 sg13g2_fill_1 FILLER_21_289 ();
 sg13g2_fill_2 FILLER_21_298 ();
 sg13g2_fill_1 FILLER_21_300 ();
 sg13g2_fill_2 FILLER_21_318 ();
 sg13g2_fill_1 FILLER_21_320 ();
 sg13g2_fill_1 FILLER_21_380 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_fill_2 FILLER_22_54 ();
 sg13g2_decap_4 FILLER_22_77 ();
 sg13g2_decap_4 FILLER_22_86 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_fill_2 FILLER_22_101 ();
 sg13g2_fill_1 FILLER_22_103 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_116 ();
 sg13g2_fill_1 FILLER_22_118 ();
 sg13g2_decap_8 FILLER_22_122 ();
 sg13g2_decap_4 FILLER_22_129 ();
 sg13g2_fill_1 FILLER_22_133 ();
 sg13g2_decap_4 FILLER_22_160 ();
 sg13g2_fill_2 FILLER_22_164 ();
 sg13g2_fill_2 FILLER_22_179 ();
 sg13g2_decap_4 FILLER_22_191 ();
 sg13g2_fill_2 FILLER_22_195 ();
 sg13g2_decap_4 FILLER_22_205 ();
 sg13g2_fill_1 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_233 ();
 sg13g2_decap_4 FILLER_22_240 ();
 sg13g2_fill_1 FILLER_22_244 ();
 sg13g2_fill_1 FILLER_22_266 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_fill_2 FILLER_22_326 ();
 sg13g2_fill_2 FILLER_22_367 ();
 sg13g2_fill_1 FILLER_22_369 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_50 ();
 sg13g2_fill_1 FILLER_23_72 ();
 sg13g2_fill_2 FILLER_23_96 ();
 sg13g2_fill_1 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_4 FILLER_23_140 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_decap_8 FILLER_23_166 ();
 sg13g2_fill_2 FILLER_23_178 ();
 sg13g2_fill_2 FILLER_23_191 ();
 sg13g2_fill_2 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_244 ();
 sg13g2_decap_4 FILLER_23_261 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_4 FILLER_23_280 ();
 sg13g2_fill_2 FILLER_23_284 ();
 sg13g2_fill_2 FILLER_23_290 ();
 sg13g2_fill_2 FILLER_23_298 ();
 sg13g2_fill_1 FILLER_23_343 ();
 sg13g2_fill_2 FILLER_24_47 ();
 sg13g2_fill_1 FILLER_24_49 ();
 sg13g2_fill_2 FILLER_24_71 ();
 sg13g2_fill_1 FILLER_24_81 ();
 sg13g2_fill_1 FILLER_24_92 ();
 sg13g2_decap_4 FILLER_24_97 ();
 sg13g2_fill_2 FILLER_24_101 ();
 sg13g2_fill_1 FILLER_24_113 ();
 sg13g2_decap_8 FILLER_24_121 ();
 sg13g2_fill_2 FILLER_24_128 ();
 sg13g2_fill_1 FILLER_24_144 ();
 sg13g2_decap_8 FILLER_24_167 ();
 sg13g2_fill_2 FILLER_24_174 ();
 sg13g2_fill_1 FILLER_24_176 ();
 sg13g2_fill_1 FILLER_24_186 ();
 sg13g2_decap_4 FILLER_24_197 ();
 sg13g2_fill_2 FILLER_24_201 ();
 sg13g2_decap_8 FILLER_24_211 ();
 sg13g2_fill_2 FILLER_24_218 ();
 sg13g2_decap_4 FILLER_24_271 ();
 sg13g2_fill_2 FILLER_24_275 ();
 sg13g2_fill_2 FILLER_24_311 ();
 sg13g2_fill_1 FILLER_24_313 ();
 sg13g2_fill_1 FILLER_24_357 ();
 sg13g2_fill_2 FILLER_24_362 ();
 sg13g2_fill_1 FILLER_24_364 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_decap_4 FILLER_25_19 ();
 sg13g2_fill_2 FILLER_25_49 ();
 sg13g2_decap_4 FILLER_25_63 ();
 sg13g2_fill_1 FILLER_25_67 ();
 sg13g2_fill_2 FILLER_25_97 ();
 sg13g2_fill_1 FILLER_25_123 ();
 sg13g2_decap_8 FILLER_25_132 ();
 sg13g2_fill_2 FILLER_25_139 ();
 sg13g2_decap_4 FILLER_25_165 ();
 sg13g2_decap_4 FILLER_25_193 ();
 sg13g2_decap_8 FILLER_25_218 ();
 sg13g2_fill_2 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_227 ();
 sg13g2_fill_1 FILLER_25_259 ();
 sg13g2_fill_2 FILLER_25_286 ();
 sg13g2_fill_1 FILLER_25_382 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_4 ();
 sg13g2_fill_2 FILLER_26_36 ();
 sg13g2_decap_8 FILLER_26_59 ();
 sg13g2_fill_2 FILLER_26_114 ();
 sg13g2_decap_8 FILLER_26_125 ();
 sg13g2_decap_8 FILLER_26_132 ();
 sg13g2_decap_8 FILLER_26_139 ();
 sg13g2_fill_2 FILLER_26_146 ();
 sg13g2_fill_1 FILLER_26_148 ();
 sg13g2_decap_8 FILLER_26_159 ();
 sg13g2_decap_8 FILLER_26_166 ();
 sg13g2_decap_4 FILLER_26_173 ();
 sg13g2_fill_1 FILLER_26_177 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_192 ();
 sg13g2_decap_8 FILLER_26_199 ();
 sg13g2_decap_8 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_fill_1 FILLER_26_222 ();
 sg13g2_decap_4 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_246 ();
 sg13g2_fill_2 FILLER_26_257 ();
 sg13g2_fill_2 FILLER_26_275 ();
 sg13g2_fill_2 FILLER_26_282 ();
 sg13g2_fill_2 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_296 ();
 sg13g2_fill_2 FILLER_26_323 ();
 sg13g2_fill_2 FILLER_26_370 ();
 sg13g2_fill_1 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_27_70 ();
 sg13g2_fill_1 FILLER_27_72 ();
 sg13g2_fill_2 FILLER_27_99 ();
 sg13g2_fill_2 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_107 ();
 sg13g2_fill_2 FILLER_27_114 ();
 sg13g2_fill_1 FILLER_27_116 ();
 sg13g2_decap_4 FILLER_27_123 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_fill_1 FILLER_27_140 ();
 sg13g2_fill_2 FILLER_27_161 ();
 sg13g2_fill_1 FILLER_27_163 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_fill_2 FILLER_27_194 ();
 sg13g2_fill_1 FILLER_27_196 ();
 sg13g2_decap_4 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_206 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_270 ();
 sg13g2_fill_2 FILLER_27_305 ();
 sg13g2_fill_2 FILLER_27_380 ();
 sg13g2_fill_1 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_40 ();
 sg13g2_fill_1 FILLER_28_44 ();
 sg13g2_fill_1 FILLER_28_61 ();
 sg13g2_fill_1 FILLER_28_70 ();
 sg13g2_fill_2 FILLER_28_81 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_decap_4 FILLER_28_88 ();
 sg13g2_fill_2 FILLER_28_117 ();
 sg13g2_fill_1 FILLER_28_125 ();
 sg13g2_fill_1 FILLER_28_142 ();
 sg13g2_fill_2 FILLER_28_164 ();
 sg13g2_fill_2 FILLER_28_171 ();
 sg13g2_fill_1 FILLER_28_173 ();
 sg13g2_fill_2 FILLER_28_196 ();
 sg13g2_decap_4 FILLER_28_215 ();
 sg13g2_fill_2 FILLER_28_242 ();
 sg13g2_fill_1 FILLER_28_259 ();
 sg13g2_fill_1 FILLER_28_285 ();
 sg13g2_fill_1 FILLER_28_294 ();
 sg13g2_fill_2 FILLER_28_323 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_fill_2 FILLER_28_354 ();
 sg13g2_fill_1 FILLER_28_356 ();
 sg13g2_fill_2 FILLER_29_26 ();
 sg13g2_fill_1 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_42 ();
 sg13g2_fill_2 FILLER_29_55 ();
 sg13g2_fill_1 FILLER_29_57 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_4 FILLER_29_84 ();
 sg13g2_fill_1 FILLER_29_88 ();
 sg13g2_decap_8 FILLER_29_106 ();
 sg13g2_fill_1 FILLER_29_113 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_121 ();
 sg13g2_decap_8 FILLER_29_130 ();
 sg13g2_fill_2 FILLER_29_137 ();
 sg13g2_fill_1 FILLER_29_139 ();
 sg13g2_fill_2 FILLER_29_158 ();
 sg13g2_fill_1 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_172 ();
 sg13g2_fill_2 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_191 ();
 sg13g2_fill_2 FILLER_29_201 ();
 sg13g2_fill_1 FILLER_29_203 ();
 sg13g2_decap_4 FILLER_29_209 ();
 sg13g2_fill_2 FILLER_29_223 ();
 sg13g2_fill_2 FILLER_29_255 ();
 sg13g2_fill_1 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_fill_2 FILLER_29_366 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_72 ();
 sg13g2_fill_1 FILLER_30_79 ();
 sg13g2_fill_1 FILLER_30_108 ();
 sg13g2_decap_8 FILLER_30_134 ();
 sg13g2_decap_4 FILLER_30_141 ();
 sg13g2_fill_2 FILLER_30_178 ();
 sg13g2_fill_2 FILLER_30_184 ();
 sg13g2_fill_1 FILLER_30_186 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_4 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_fill_2 FILLER_30_244 ();
 sg13g2_fill_1 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_257 ();
 sg13g2_fill_2 FILLER_30_267 ();
 sg13g2_fill_2 FILLER_30_281 ();
 sg13g2_fill_1 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_299 ();
 sg13g2_fill_1 FILLER_30_346 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_15 ();
 sg13g2_fill_1 FILLER_31_22 ();
 sg13g2_fill_1 FILLER_31_32 ();
 sg13g2_decap_4 FILLER_31_67 ();
 sg13g2_fill_2 FILLER_31_71 ();
 sg13g2_decap_8 FILLER_31_99 ();
 sg13g2_fill_2 FILLER_31_106 ();
 sg13g2_fill_1 FILLER_31_120 ();
 sg13g2_decap_8 FILLER_31_129 ();
 sg13g2_decap_4 FILLER_31_136 ();
 sg13g2_fill_2 FILLER_31_140 ();
 sg13g2_decap_4 FILLER_31_158 ();
 sg13g2_fill_1 FILLER_31_162 ();
 sg13g2_decap_4 FILLER_31_171 ();
 sg13g2_fill_1 FILLER_31_175 ();
 sg13g2_fill_2 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_223 ();
 sg13g2_fill_2 FILLER_31_245 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_fill_1 FILLER_31_348 ();
 sg13g2_fill_1 FILLER_31_376 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_fill_1 FILLER_32_55 ();
 sg13g2_fill_2 FILLER_32_61 ();
 sg13g2_fill_1 FILLER_32_63 ();
 sg13g2_decap_4 FILLER_32_68 ();
 sg13g2_fill_2 FILLER_32_96 ();
 sg13g2_fill_1 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_104 ();
 sg13g2_fill_1 FILLER_32_111 ();
 sg13g2_fill_2 FILLER_32_128 ();
 sg13g2_fill_2 FILLER_32_142 ();
 sg13g2_fill_1 FILLER_32_144 ();
 sg13g2_decap_8 FILLER_32_162 ();
 sg13g2_decap_8 FILLER_32_169 ();
 sg13g2_decap_8 FILLER_32_195 ();
 sg13g2_decap_4 FILLER_32_202 ();
 sg13g2_fill_1 FILLER_32_206 ();
 sg13g2_fill_2 FILLER_32_233 ();
 sg13g2_fill_1 FILLER_32_235 ();
 sg13g2_fill_1 FILLER_32_248 ();
 sg13g2_fill_2 FILLER_32_261 ();
 sg13g2_fill_1 FILLER_32_267 ();
 sg13g2_fill_2 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_285 ();
 sg13g2_fill_2 FILLER_32_291 ();
 sg13g2_fill_2 FILLER_32_316 ();
 sg13g2_fill_1 FILLER_32_318 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_50 ();
 sg13g2_fill_1 FILLER_33_52 ();
 sg13g2_decap_8 FILLER_33_79 ();
 sg13g2_fill_2 FILLER_33_86 ();
 sg13g2_fill_1 FILLER_33_127 ();
 sg13g2_fill_2 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_157 ();
 sg13g2_decap_4 FILLER_33_164 ();
 sg13g2_fill_2 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_fill_1 FILLER_33_202 ();
 sg13g2_fill_2 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_230 ();
 sg13g2_fill_2 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_306 ();
 sg13g2_fill_1 FILLER_33_316 ();
 sg13g2_fill_2 FILLER_33_336 ();
 sg13g2_fill_1 FILLER_33_338 ();
 sg13g2_fill_2 FILLER_33_357 ();
 sg13g2_fill_1 FILLER_33_390 ();
 sg13g2_fill_2 FILLER_34_66 ();
 sg13g2_decap_4 FILLER_34_72 ();
 sg13g2_fill_2 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_104 ();
 sg13g2_fill_2 FILLER_34_122 ();
 sg13g2_fill_1 FILLER_34_152 ();
 sg13g2_fill_1 FILLER_34_165 ();
 sg13g2_fill_1 FILLER_34_191 ();
 sg13g2_fill_2 FILLER_34_200 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_2 FILLER_34_255 ();
 sg13g2_fill_2 FILLER_34_271 ();
 sg13g2_fill_2 FILLER_34_312 ();
 sg13g2_fill_1 FILLER_34_314 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_11 ();
 sg13g2_fill_1 FILLER_35_56 ();
 sg13g2_fill_1 FILLER_35_91 ();
 sg13g2_fill_2 FILLER_35_101 ();
 sg13g2_fill_1 FILLER_35_131 ();
 sg13g2_fill_1 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_165 ();
 sg13g2_fill_2 FILLER_35_188 ();
 sg13g2_fill_1 FILLER_35_190 ();
 sg13g2_fill_2 FILLER_35_225 ();
 sg13g2_fill_1 FILLER_35_227 ();
 sg13g2_fill_1 FILLER_35_371 ();
 sg13g2_fill_1 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_11 ();
 sg13g2_fill_1 FILLER_36_47 ();
 sg13g2_fill_2 FILLER_36_61 ();
 sg13g2_fill_1 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_76 ();
 sg13g2_fill_1 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_114 ();
 sg13g2_fill_2 FILLER_36_141 ();
 sg13g2_fill_1 FILLER_36_181 ();
 sg13g2_fill_1 FILLER_36_212 ();
 sg13g2_fill_2 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_225 ();
 sg13g2_fill_1 FILLER_36_239 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_18 ();
 sg13g2_fill_2 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_44 ();
 sg13g2_fill_2 FILLER_37_94 ();
 sg13g2_fill_2 FILLER_37_130 ();
 sg13g2_fill_1 FILLER_37_132 ();
 sg13g2_fill_2 FILLER_37_151 ();
 sg13g2_fill_1 FILLER_37_188 ();
 sg13g2_fill_1 FILLER_37_232 ();
 sg13g2_fill_1 FILLER_37_261 ();
 sg13g2_fill_1 FILLER_37_278 ();
 sg13g2_fill_2 FILLER_37_324 ();
 sg13g2_fill_1 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_99 ();
 sg13g2_fill_1 FILLER_38_101 ();
 sg13g2_fill_2 FILLER_38_128 ();
 sg13g2_fill_1 FILLER_38_130 ();
 sg13g2_fill_2 FILLER_38_217 ();
 sg13g2_fill_1 FILLER_38_219 ();
 sg13g2_fill_1 FILLER_38_246 ();
 assign uio_oe[0] = net15;
 assign uio_oe[1] = net16;
 assign uio_oe[2] = net17;
 assign uio_oe[3] = net18;
 assign uio_oe[4] = net19;
 assign uio_oe[5] = net20;
 assign uio_oe[6] = net21;
 assign uio_oe[7] = net22;
 assign uio_out[0] = net23;
 assign uio_out[1] = net24;
 assign uio_out[2] = net25;
 assign uio_out[3] = net26;
 assign uio_out[4] = net27;
 assign uio_out[5] = net28;
 assign uio_out[6] = net29;
 assign uio_out[7] = net30;
endmodule

module tt_um_benpayne_ps2_decoder (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire clknet_0_clk;
 wire cs_prev;
 wire cs_trigger;
 wire \memory.count[0] ;
 wire \memory.count[1] ;
 wire \memory.count[2] ;
 wire \memory.mem[0][0] ;
 wire \memory.mem[0][1] ;
 wire \memory.mem[0][2] ;
 wire \memory.mem[0][3] ;
 wire \memory.mem[0][4] ;
 wire \memory.mem[0][5] ;
 wire \memory.mem[0][6] ;
 wire \memory.mem[0][7] ;
 wire \memory.mem[1][0] ;
 wire \memory.mem[1][1] ;
 wire \memory.mem[1][2] ;
 wire \memory.mem[1][3] ;
 wire \memory.mem[1][4] ;
 wire \memory.mem[1][5] ;
 wire \memory.mem[1][6] ;
 wire \memory.mem[1][7] ;
 wire \memory.mem[2][0] ;
 wire \memory.mem[2][1] ;
 wire \memory.mem[2][2] ;
 wire \memory.mem[2][3] ;
 wire \memory.mem[2][4] ;
 wire \memory.mem[2][5] ;
 wire \memory.mem[2][6] ;
 wire \memory.mem[2][7] ;
 wire \memory.mem[3][0] ;
 wire \memory.mem[3][1] ;
 wire \memory.mem[3][2] ;
 wire \memory.mem[3][3] ;
 wire \memory.mem[3][4] ;
 wire \memory.mem[3][5] ;
 wire \memory.mem[3][6] ;
 wire \memory.mem[3][7] ;
 wire \memory.rd_ptr[0] ;
 wire \memory.rd_ptr[1] ;
 wire \memory.wr_ptr[0] ;
 wire \memory.wr_ptr[1] ;
 wire \ps2_clk_debounce.counter[0] ;
 wire \ps2_clk_debounce.counter[1] ;
 wire \ps2_clk_debounce.counter[2] ;
 wire \ps2_clk_debounce.counter[3] ;
 wire \ps2_clk_debounce.counter[4] ;
 wire \ps2_clk_debounce.counter[5] ;
 wire \ps2_clk_debounce.counter[6] ;
 wire \ps2_clk_debounce.counter[7] ;
 wire \ps2_clk_debounce.debounced_button ;
 wire \ps2_clk_debounce.last_button ;
 wire \ps2_data_debounce.counter[0] ;
 wire \ps2_data_debounce.counter[1] ;
 wire \ps2_data_debounce.counter[2] ;
 wire \ps2_data_debounce.counter[3] ;
 wire \ps2_data_debounce.counter[4] ;
 wire \ps2_data_debounce.counter[5] ;
 wire \ps2_data_debounce.counter[6] ;
 wire \ps2_data_debounce.counter[7] ;
 wire \ps2_data_debounce.debounced_button ;
 wire \ps2_data_debounce.last_button ;
 wire \ps2_decoder_inst.clk_timeout[0] ;
 wire \ps2_decoder_inst.clk_timeout[10] ;
 wire \ps2_decoder_inst.clk_timeout[11] ;
 wire \ps2_decoder_inst.clk_timeout[12] ;
 wire \ps2_decoder_inst.clk_timeout[1] ;
 wire \ps2_decoder_inst.clk_timeout[2] ;
 wire \ps2_decoder_inst.clk_timeout[3] ;
 wire \ps2_decoder_inst.clk_timeout[4] ;
 wire \ps2_decoder_inst.clk_timeout[5] ;
 wire \ps2_decoder_inst.clk_timeout[6] ;
 wire \ps2_decoder_inst.clk_timeout[7] ;
 wire \ps2_decoder_inst.clk_timeout[8] ;
 wire \ps2_decoder_inst.clk_timeout[9] ;
 wire \ps2_decoder_inst.int_reg ;
 wire \ps2_decoder_inst.ps2_clk_prev ;
 wire \ps2_decoder_inst.ps2_value[0] ;
 wire \ps2_decoder_inst.ps2_value[1] ;
 wire \ps2_decoder_inst.ps2_value[2] ;
 wire \ps2_decoder_inst.ps2_value[3] ;
 wire \ps2_decoder_inst.ps2_value[4] ;
 wire \ps2_decoder_inst.ps2_value[5] ;
 wire \ps2_decoder_inst.ps2_value[6] ;
 wire \ps2_decoder_inst.ps2_value[7] ;
 wire \ps2_decoder_inst.shift_reg[0] ;
 wire \ps2_decoder_inst.shift_reg[10] ;
 wire \ps2_decoder_inst.shift_reg[1] ;
 wire \ps2_decoder_inst.shift_reg[2] ;
 wire \ps2_decoder_inst.shift_reg[3] ;
 wire \ps2_decoder_inst.shift_reg[4] ;
 wire \ps2_decoder_inst.shift_reg[5] ;
 wire \ps2_decoder_inst.shift_reg[6] ;
 wire \ps2_decoder_inst.shift_reg[7] ;
 wire \ps2_decoder_inst.shift_reg[8] ;
 wire \ps2_decoder_inst.shift_reg[9] ;
 wire \ps2_decoder_inst.shift_reset ;
 wire \ps2_decoder_inst.state_reg[0] ;
 wire \ps2_decoder_inst.state_reg[1] ;
 wire \ps2_decoder_inst.valid_reg ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;

 sg13g2_inv_1 _443_ (.Y(_110_),
    .A(\memory.count[2] ));
 sg13g2_inv_1 _444_ (.Y(_111_),
    .A(cs_trigger));
 sg13g2_inv_2 _445_ (.Y(_112_),
    .A(\ps2_clk_debounce.debounced_button ));
 sg13g2_inv_1 _446_ (.Y(_113_),
    .A(net78));
 sg13g2_inv_1 _447_ (.Y(_114_),
    .A(net164));
 sg13g2_inv_1 _448_ (.Y(_115_),
    .A(\ps2_decoder_inst.clk_timeout[12] ));
 sg13g2_inv_1 _449_ (.Y(_116_),
    .A(net108));
 sg13g2_inv_1 _450_ (.Y(_117_),
    .A(\memory.wr_ptr[1] ));
 sg13g2_inv_1 _451_ (.Y(_118_),
    .A(net3));
 sg13g2_inv_1 _452_ (.Y(_119_),
    .A(net197));
 sg13g2_inv_1 _453_ (.Y(_120_),
    .A(net148));
 sg13g2_inv_1 _454_ (.Y(_121_),
    .A(net206));
 sg13g2_inv_1 _455_ (.Y(_122_),
    .A(net84));
 sg13g2_nor3_1 _456_ (.A(\memory.count[2] ),
    .B(\memory.count[1] ),
    .C(\memory.count[0] ),
    .Y(_123_));
 sg13g2_inv_1 _457_ (.Y(uo_out[2]),
    .A(_123_));
 sg13g2_nor2b_1 _458_ (.A(net43),
    .B_N(net4),
    .Y(_000_));
 sg13g2_xor2_1 _459_ (.B(net1),
    .A(\ps2_clk_debounce.last_button ),
    .X(_124_));
 sg13g2_nor2_1 _460_ (.A(net52),
    .B(_124_),
    .Y(_125_));
 sg13g2_or2_2 _461_ (.X(_126_),
    .B(_124_),
    .A(net52));
 sg13g2_and2_1 _462_ (.A(net131),
    .B(net75),
    .X(_127_));
 sg13g2_and3_1 _463_ (.X(_128_),
    .A(net82),
    .B(\ps2_clk_debounce.counter[3] ),
    .C(_127_));
 sg13g2_and2_1 _464_ (.A(net113),
    .B(_128_),
    .X(_129_));
 sg13g2_nand2_1 _465_ (.Y(_130_),
    .A(net113),
    .B(_128_));
 sg13g2_nand3_1 _466_ (.B(net148),
    .C(_129_),
    .A(net121),
    .Y(_131_));
 sg13g2_a21oi_1 _467_ (.A1(net52),
    .A2(_131_),
    .Y(_001_),
    .B1(_124_));
 sg13g2_nand2_1 _468_ (.Y(_132_),
    .A(net80),
    .B(net2));
 sg13g2_xor2_1 _469_ (.B(net2),
    .A(\ps2_data_debounce.last_button ),
    .X(_133_));
 sg13g2_nor2_1 _470_ (.A(net71),
    .B(_133_),
    .Y(_134_));
 sg13g2_or2_1 _471_ (.X(_135_),
    .B(_133_),
    .A(net71));
 sg13g2_and2_1 _472_ (.A(net127),
    .B(net116),
    .X(_136_));
 sg13g2_and3_1 _473_ (.X(_137_),
    .A(net123),
    .B(\ps2_data_debounce.counter[3] ),
    .C(_136_));
 sg13g2_and2_1 _474_ (.A(\ps2_data_debounce.counter[4] ),
    .B(_137_),
    .X(_138_));
 sg13g2_nand2_1 _475_ (.Y(_139_),
    .A(net133),
    .B(_137_));
 sg13g2_nand3_1 _476_ (.B(net84),
    .C(_138_),
    .A(\ps2_data_debounce.counter[5] ),
    .Y(_140_));
 sg13g2_a21oi_1 _477_ (.A1(net71),
    .A2(_140_),
    .Y(_002_),
    .B1(_133_));
 sg13g2_nor2b_2 _478_ (.A(\memory.count[2] ),
    .B_N(\ps2_decoder_inst.valid_reg ),
    .Y(_141_));
 sg13g2_nand2_2 _479_ (.Y(_142_),
    .A(\memory.wr_ptr[0] ),
    .B(_141_));
 sg13g2_nor3_2 _480_ (.A(_116_),
    .B(_117_),
    .C(_142_),
    .Y(_143_));
 sg13g2_mux2_1 _481_ (.A0(net191),
    .A1(\ps2_decoder_inst.ps2_value[0] ),
    .S(_143_),
    .X(_009_));
 sg13g2_mux2_1 _482_ (.A0(net144),
    .A1(\ps2_decoder_inst.ps2_value[1] ),
    .S(_143_),
    .X(_010_));
 sg13g2_mux2_1 _483_ (.A0(net160),
    .A1(\ps2_decoder_inst.ps2_value[2] ),
    .S(_143_),
    .X(_011_));
 sg13g2_mux2_1 _484_ (.A0(net136),
    .A1(\ps2_decoder_inst.ps2_value[3] ),
    .S(_143_),
    .X(_012_));
 sg13g2_mux2_1 _485_ (.A0(net185),
    .A1(\ps2_decoder_inst.ps2_value[4] ),
    .S(_143_),
    .X(_013_));
 sg13g2_mux2_1 _486_ (.A0(net138),
    .A1(\ps2_decoder_inst.ps2_value[5] ),
    .S(_143_),
    .X(_014_));
 sg13g2_mux2_1 _487_ (.A0(net125),
    .A1(\ps2_decoder_inst.ps2_value[6] ),
    .S(_143_),
    .X(_015_));
 sg13g2_mux2_1 _488_ (.A0(net175),
    .A1(\ps2_decoder_inst.ps2_value[7] ),
    .S(_143_),
    .X(_016_));
 sg13g2_nor2_2 _489_ (.A(\ps2_clk_debounce.counter[7] ),
    .B(_124_),
    .Y(_144_));
 sg13g2_and2_1 _490_ (.A(_126_),
    .B(_144_),
    .X(_145_));
 sg13g2_nor2_1 _491_ (.A(net131),
    .B(_145_),
    .Y(_146_));
 sg13g2_a21oi_1 _492_ (.A1(net131),
    .A2(_126_),
    .Y(_017_),
    .B1(_146_));
 sg13g2_nor3_1 _493_ (.A(\ps2_clk_debounce.counter[7] ),
    .B(_124_),
    .C(_127_),
    .Y(_147_));
 sg13g2_nor2_1 _494_ (.A(_125_),
    .B(_147_),
    .Y(_148_));
 sg13g2_a21oi_1 _495_ (.A1(\ps2_clk_debounce.counter[0] ),
    .A2(_126_),
    .Y(_149_),
    .B1(net75));
 sg13g2_nor2_1 _496_ (.A(_148_),
    .B(net76),
    .Y(_018_));
 sg13g2_a21oi_1 _497_ (.A1(_127_),
    .A2(_145_),
    .Y(_150_),
    .B1(net82));
 sg13g2_a21oi_1 _498_ (.A1(net82),
    .A2(_148_),
    .Y(_019_),
    .B1(_150_));
 sg13g2_nand3_1 _499_ (.B(_126_),
    .C(_127_),
    .A(net82),
    .Y(_151_));
 sg13g2_nand2b_1 _500_ (.Y(_152_),
    .B(_144_),
    .A_N(_128_));
 sg13g2_a22oi_1 _501_ (.Y(_020_),
    .B1(_152_),
    .B2(_126_),
    .A2(_151_),
    .A1(_119_));
 sg13g2_a21oi_1 _502_ (.A1(_130_),
    .A2(_144_),
    .Y(_153_),
    .B1(_125_));
 sg13g2_a21oi_1 _503_ (.A1(_126_),
    .A2(_128_),
    .Y(_154_),
    .B1(net113));
 sg13g2_nor2_1 _504_ (.A(_153_),
    .B(net114),
    .Y(_021_));
 sg13g2_a21oi_1 _505_ (.A1(_129_),
    .A2(_145_),
    .Y(_155_),
    .B1(net121));
 sg13g2_a21oi_1 _506_ (.A1(net121),
    .A2(_153_),
    .Y(_022_),
    .B1(_155_));
 sg13g2_nand2_1 _507_ (.Y(_156_),
    .A(_131_),
    .B(_144_));
 sg13g2_nand3_1 _508_ (.B(_126_),
    .C(_129_),
    .A(net121),
    .Y(_157_));
 sg13g2_a22oi_1 _509_ (.Y(_023_),
    .B1(_157_),
    .B2(_120_),
    .A2(_156_),
    .A1(_126_));
 sg13g2_nand3b_1 _510_ (.B(net1),
    .C(net210),
    .Y(_158_),
    .A_N(net52));
 sg13g2_o21ai_1 _511_ (.B1(_158_),
    .Y(_024_),
    .A1(_112_),
    .A2(_125_));
 sg13g2_nor2_2 _512_ (.A(\ps2_data_debounce.counter[7] ),
    .B(_133_),
    .Y(_159_));
 sg13g2_and2_1 _513_ (.A(_135_),
    .B(_159_),
    .X(_160_));
 sg13g2_nor2_1 _514_ (.A(net127),
    .B(_160_),
    .Y(_161_));
 sg13g2_a21oi_1 _515_ (.A1(net127),
    .A2(net94),
    .Y(_025_),
    .B1(_161_));
 sg13g2_nor3_1 _516_ (.A(\ps2_data_debounce.counter[7] ),
    .B(_133_),
    .C(_136_),
    .Y(_162_));
 sg13g2_nor2_1 _517_ (.A(_134_),
    .B(_162_),
    .Y(_163_));
 sg13g2_a21oi_1 _518_ (.A1(\ps2_data_debounce.counter[0] ),
    .A2(net94),
    .Y(_164_),
    .B1(net116));
 sg13g2_nor2_1 _519_ (.A(_163_),
    .B(net117),
    .Y(_026_));
 sg13g2_a21oi_1 _520_ (.A1(_136_),
    .A2(_160_),
    .Y(_165_),
    .B1(net123));
 sg13g2_a21oi_1 _521_ (.A1(net123),
    .A2(_163_),
    .Y(_027_),
    .B1(_165_));
 sg13g2_nand3_1 _522_ (.B(net94),
    .C(_136_),
    .A(net123),
    .Y(_166_));
 sg13g2_nand2b_1 _523_ (.Y(_167_),
    .B(_159_),
    .A_N(_137_));
 sg13g2_a22oi_1 _524_ (.Y(_028_),
    .B1(_167_),
    .B2(net94),
    .A2(_166_),
    .A1(_121_));
 sg13g2_a21oi_1 _525_ (.A1(_139_),
    .A2(_159_),
    .Y(_168_),
    .B1(_134_));
 sg13g2_a21oi_1 _526_ (.A1(net94),
    .A2(_137_),
    .Y(_169_),
    .B1(net133));
 sg13g2_nor2_1 _527_ (.A(_168_),
    .B(net134),
    .Y(_029_));
 sg13g2_a21oi_1 _528_ (.A1(_138_),
    .A2(_160_),
    .Y(_170_),
    .B1(net119));
 sg13g2_a21oi_1 _529_ (.A1(net119),
    .A2(_168_),
    .Y(_030_),
    .B1(_170_));
 sg13g2_nand2_1 _530_ (.Y(_171_),
    .A(_140_),
    .B(_159_));
 sg13g2_nand3_1 _531_ (.B(net94),
    .C(_138_),
    .A(\ps2_data_debounce.counter[5] ),
    .Y(_172_));
 sg13g2_a22oi_1 _532_ (.Y(_031_),
    .B1(_172_),
    .B2(_122_),
    .A2(_171_),
    .A1(net94));
 sg13g2_nand2_1 _533_ (.Y(_173_),
    .A(net203),
    .B(\ps2_decoder_inst.shift_reset ));
 sg13g2_o21ai_1 _534_ (.B1(net204),
    .Y(_032_),
    .A1(_112_),
    .A2(\ps2_decoder_inst.shift_reset ));
 sg13g2_nor3_2 _535_ (.A(_116_),
    .B(\memory.wr_ptr[1] ),
    .C(_142_),
    .Y(_174_));
 sg13g2_mux2_1 _536_ (.A0(net208),
    .A1(\ps2_decoder_inst.ps2_value[0] ),
    .S(_174_),
    .X(_033_));
 sg13g2_mux2_1 _537_ (.A0(net142),
    .A1(\ps2_decoder_inst.ps2_value[1] ),
    .S(_174_),
    .X(_034_));
 sg13g2_mux2_1 _538_ (.A0(net152),
    .A1(\ps2_decoder_inst.ps2_value[2] ),
    .S(_174_),
    .X(_035_));
 sg13g2_mux2_1 _539_ (.A0(net193),
    .A1(\ps2_decoder_inst.ps2_value[3] ),
    .S(_174_),
    .X(_036_));
 sg13g2_mux2_1 _540_ (.A0(net146),
    .A1(\ps2_decoder_inst.ps2_value[4] ),
    .S(_174_),
    .X(_037_));
 sg13g2_mux2_1 _541_ (.A0(net162),
    .A1(\ps2_decoder_inst.ps2_value[5] ),
    .S(_174_),
    .X(_038_));
 sg13g2_mux2_1 _542_ (.A0(net150),
    .A1(\ps2_decoder_inst.ps2_value[6] ),
    .S(_174_),
    .X(_039_));
 sg13g2_mux2_1 _543_ (.A0(net181),
    .A1(\ps2_decoder_inst.ps2_value[7] ),
    .S(_174_),
    .X(_040_));
 sg13g2_mux2_1 _544_ (.A0(\memory.wr_ptr[0] ),
    .A1(net54),
    .S(_141_),
    .X(_041_));
 sg13g2_xnor2_1 _545_ (.Y(_042_),
    .A(net239),
    .B(_142_));
 sg13g2_nand2b_1 _546_ (.Y(_175_),
    .B(cs_trigger),
    .A_N(_123_));
 sg13g2_mux2_1 _547_ (.A0(net46),
    .A1(\memory.rd_ptr[0] ),
    .S(net93),
    .X(_043_));
 sg13g2_and2_1 _548_ (.A(\memory.rd_ptr[0] ),
    .B(\memory.rd_ptr[1] ),
    .X(_176_));
 sg13g2_nor2_1 _549_ (.A(\memory.rd_ptr[0] ),
    .B(\memory.rd_ptr[1] ),
    .Y(_177_));
 sg13g2_nor2b_2 _550_ (.A(\memory.rd_ptr[1] ),
    .B_N(\memory.rd_ptr[0] ),
    .Y(_178_));
 sg13g2_nor2b_2 _551_ (.A(\memory.rd_ptr[0] ),
    .B_N(\memory.rd_ptr[1] ),
    .Y(_179_));
 sg13g2_nor3_1 _552_ (.A(net92),
    .B(net96),
    .C(net95),
    .Y(_180_));
 sg13g2_a21o_1 _553_ (.A2(net92),
    .A1(net249),
    .B1(_180_),
    .X(_044_));
 sg13g2_nand2_1 _554_ (.Y(_181_),
    .A(net108),
    .B(_141_));
 sg13g2_nor3_2 _555_ (.A(\memory.wr_ptr[0] ),
    .B(_117_),
    .C(_181_),
    .Y(_182_));
 sg13g2_mux2_1 _556_ (.A0(net201),
    .A1(\ps2_decoder_inst.ps2_value[0] ),
    .S(_182_),
    .X(_045_));
 sg13g2_mux2_1 _557_ (.A0(net199),
    .A1(\ps2_decoder_inst.ps2_value[1] ),
    .S(_182_),
    .X(_046_));
 sg13g2_mux2_1 _558_ (.A0(net173),
    .A1(\ps2_decoder_inst.ps2_value[2] ),
    .S(_182_),
    .X(_047_));
 sg13g2_mux2_1 _559_ (.A0(net171),
    .A1(\ps2_decoder_inst.ps2_value[3] ),
    .S(_182_),
    .X(_048_));
 sg13g2_mux2_1 _560_ (.A0(net158),
    .A1(\ps2_decoder_inst.ps2_value[4] ),
    .S(_182_),
    .X(_049_));
 sg13g2_mux2_1 _561_ (.A0(net189),
    .A1(\ps2_decoder_inst.ps2_value[5] ),
    .S(_182_),
    .X(_050_));
 sg13g2_mux2_1 _562_ (.A0(net177),
    .A1(\ps2_decoder_inst.ps2_value[6] ),
    .S(_182_),
    .X(_051_));
 sg13g2_mux2_1 _563_ (.A0(net154),
    .A1(\ps2_decoder_inst.ps2_value[7] ),
    .S(_182_),
    .X(_052_));
 sg13g2_nor3_2 _564_ (.A(\memory.wr_ptr[0] ),
    .B(\memory.wr_ptr[1] ),
    .C(_181_),
    .Y(_183_));
 sg13g2_mux2_1 _565_ (.A0(net140),
    .A1(\ps2_decoder_inst.ps2_value[0] ),
    .S(_183_),
    .X(_053_));
 sg13g2_mux2_1 _566_ (.A0(net187),
    .A1(\ps2_decoder_inst.ps2_value[1] ),
    .S(_183_),
    .X(_054_));
 sg13g2_mux2_1 _567_ (.A0(net168),
    .A1(\ps2_decoder_inst.ps2_value[2] ),
    .S(_183_),
    .X(_055_));
 sg13g2_mux2_1 _568_ (.A0(net129),
    .A1(\ps2_decoder_inst.ps2_value[3] ),
    .S(_183_),
    .X(_056_));
 sg13g2_mux2_1 _569_ (.A0(net166),
    .A1(\ps2_decoder_inst.ps2_value[4] ),
    .S(_183_),
    .X(_057_));
 sg13g2_mux2_1 _570_ (.A0(net156),
    .A1(\ps2_decoder_inst.ps2_value[5] ),
    .S(_183_),
    .X(_058_));
 sg13g2_mux2_1 _571_ (.A0(net195),
    .A1(\ps2_decoder_inst.ps2_value[6] ),
    .S(_183_),
    .X(_059_));
 sg13g2_mux2_1 _572_ (.A0(net183),
    .A1(\ps2_decoder_inst.ps2_value[7] ),
    .S(_183_),
    .X(_060_));
 sg13g2_a22oi_1 _573_ (.Y(_184_),
    .B1(_179_),
    .B2(net201),
    .A2(net96),
    .A1(net191));
 sg13g2_a22oi_1 _574_ (.Y(_185_),
    .B1(_178_),
    .B2(net208),
    .A2(_177_),
    .A1(net140));
 sg13g2_nand2_1 _575_ (.Y(_186_),
    .A(_184_),
    .B(_185_));
 sg13g2_mux2_1 _576_ (.A0(_186_),
    .A1(net241),
    .S(net93),
    .X(_061_));
 sg13g2_a22oi_1 _577_ (.Y(_187_),
    .B1(net95),
    .B2(net187),
    .A2(net96),
    .A1(net144));
 sg13g2_a22oi_1 _578_ (.Y(_188_),
    .B1(_179_),
    .B2(net199),
    .A2(_178_),
    .A1(net142));
 sg13g2_nand2_1 _579_ (.Y(_189_),
    .A(_187_),
    .B(_188_));
 sg13g2_mux2_1 _580_ (.A0(_189_),
    .A1(net250),
    .S(net93),
    .X(_062_));
 sg13g2_a22oi_1 _581_ (.Y(_190_),
    .B1(net95),
    .B2(net168),
    .A2(net96),
    .A1(net160));
 sg13g2_a22oi_1 _582_ (.Y(_191_),
    .B1(_179_),
    .B2(net173),
    .A2(_178_),
    .A1(net152));
 sg13g2_nand2_1 _583_ (.Y(_192_),
    .A(_190_),
    .B(_191_));
 sg13g2_mux2_1 _584_ (.A0(_192_),
    .A1(net244),
    .S(net92),
    .X(_063_));
 sg13g2_a22oi_1 _585_ (.Y(_193_),
    .B1(_178_),
    .B2(net193),
    .A2(net95),
    .A1(net129));
 sg13g2_a22oi_1 _586_ (.Y(_194_),
    .B1(_179_),
    .B2(net171),
    .A2(_176_),
    .A1(net136));
 sg13g2_nand2_1 _587_ (.Y(_195_),
    .A(_193_),
    .B(_194_));
 sg13g2_mux2_1 _588_ (.A0(_195_),
    .A1(net227),
    .S(net92),
    .X(_064_));
 sg13g2_a22oi_1 _589_ (.Y(_196_),
    .B1(_179_),
    .B2(net158),
    .A2(_178_),
    .A1(net146));
 sg13g2_a22oi_1 _590_ (.Y(_197_),
    .B1(net95),
    .B2(net166),
    .A2(net96),
    .A1(net185));
 sg13g2_nand2_1 _591_ (.Y(_198_),
    .A(_196_),
    .B(_197_));
 sg13g2_mux2_1 _592_ (.A0(_198_),
    .A1(net234),
    .S(net92),
    .X(_065_));
 sg13g2_a22oi_1 _593_ (.Y(_199_),
    .B1(_179_),
    .B2(net189),
    .A2(_178_),
    .A1(net162));
 sg13g2_a22oi_1 _594_ (.Y(_200_),
    .B1(net95),
    .B2(net156),
    .A2(net96),
    .A1(net138));
 sg13g2_nand2_1 _595_ (.Y(_201_),
    .A(_199_),
    .B(_200_));
 sg13g2_mux2_1 _596_ (.A0(_201_),
    .A1(net224),
    .S(net92),
    .X(_066_));
 sg13g2_a22oi_1 _597_ (.Y(_202_),
    .B1(net95),
    .B2(net195),
    .A2(net96),
    .A1(net125));
 sg13g2_a22oi_1 _598_ (.Y(_203_),
    .B1(_179_),
    .B2(net177),
    .A2(_178_),
    .A1(net150));
 sg13g2_nand2_1 _599_ (.Y(_204_),
    .A(_202_),
    .B(_203_));
 sg13g2_mux2_1 _600_ (.A0(_204_),
    .A1(net225),
    .S(net92),
    .X(_067_));
 sg13g2_a22oi_1 _601_ (.Y(_205_),
    .B1(_179_),
    .B2(net154),
    .A2(net96),
    .A1(net175));
 sg13g2_a22oi_1 _602_ (.Y(_206_),
    .B1(_178_),
    .B2(net181),
    .A2(net95),
    .A1(net183));
 sg13g2_nand2_1 _603_ (.Y(_207_),
    .A(_205_),
    .B(_206_));
 sg13g2_mux2_1 _604_ (.A0(_207_),
    .A1(net226),
    .S(net92),
    .X(_068_));
 sg13g2_nand2_2 _605_ (.Y(_208_),
    .A(_141_),
    .B(net93));
 sg13g2_xnor2_1 _606_ (.Y(_209_),
    .A(_141_),
    .B(net93));
 sg13g2_mux2_1 _607_ (.A0(\memory.count[0] ),
    .A1(net179),
    .S(_209_),
    .X(_069_));
 sg13g2_xor2_1 _608_ (.B(_208_),
    .A(\memory.count[1] ),
    .X(_210_));
 sg13g2_xnor2_1 _609_ (.Y(_211_),
    .A(net179),
    .B(_210_));
 sg13g2_mux2_1 _610_ (.A0(net260),
    .A1(_211_),
    .S(_209_),
    .X(_070_));
 sg13g2_o21ai_1 _611_ (.B1(net212),
    .Y(_212_),
    .A1(\memory.count[1] ),
    .A2(_208_));
 sg13g2_a22oi_1 _612_ (.Y(_213_),
    .B1(_208_),
    .B2(\memory.count[1] ),
    .A2(_111_),
    .A1(\memory.count[2] ));
 sg13g2_a22oi_1 _613_ (.Y(_071_),
    .B1(net213),
    .B2(_213_),
    .A2(_208_),
    .A1(_110_));
 sg13g2_nor2_1 _614_ (.A(\ps2_decoder_inst.clk_timeout[1] ),
    .B(\ps2_decoder_inst.clk_timeout[0] ),
    .Y(_214_));
 sg13g2_and2_1 _615_ (.A(\ps2_decoder_inst.clk_timeout[7] ),
    .B(\ps2_decoder_inst.clk_timeout[6] ),
    .X(_215_));
 sg13g2_and4_1 _616_ (.A(_113_),
    .B(\ps2_decoder_inst.clk_timeout[2] ),
    .C(_214_),
    .D(_215_),
    .X(_216_));
 sg13g2_nand2b_1 _617_ (.Y(_217_),
    .B(\ps2_decoder_inst.clk_timeout[11] ),
    .A_N(\ps2_decoder_inst.clk_timeout[10] ));
 sg13g2_or2_1 _618_ (.X(_218_),
    .B(\ps2_decoder_inst.clk_timeout[4] ),
    .A(\ps2_decoder_inst.clk_timeout[5] ));
 sg13g2_nand2b_1 _619_ (.Y(_219_),
    .B(\ps2_decoder_inst.clk_timeout[8] ),
    .A_N(\ps2_decoder_inst.clk_timeout[9] ));
 sg13g2_nor4_2 _620_ (.A(\ps2_decoder_inst.clk_timeout[12] ),
    .B(_217_),
    .C(_218_),
    .Y(_220_),
    .D(_219_));
 sg13g2_nor3_1 _621_ (.A(\ps2_decoder_inst.clk_timeout[4] ),
    .B(\ps2_decoder_inst.clk_timeout[9] ),
    .C(\ps2_decoder_inst.clk_timeout[10] ),
    .Y(_221_));
 sg13g2_nand2_1 _622_ (.Y(_222_),
    .A(\ps2_decoder_inst.clk_timeout[2] ),
    .B(_215_));
 sg13g2_nand2b_1 _623_ (.Y(_223_),
    .B(\ps2_decoder_inst.clk_timeout[8] ),
    .A_N(\ps2_decoder_inst.clk_timeout[5] ));
 sg13g2_nor4_1 _624_ (.A(_114_),
    .B(\ps2_decoder_inst.clk_timeout[12] ),
    .C(_222_),
    .D(_223_),
    .Y(_224_));
 sg13g2_nand4_1 _625_ (.B(_214_),
    .C(_221_),
    .A(_113_),
    .Y(_225_),
    .D(_224_));
 sg13g2_a21o_2 _626_ (.A2(_220_),
    .A1(_216_),
    .B1(_112_),
    .X(_226_));
 sg13g2_nand2_1 _627_ (.Y(_227_),
    .A(\ps2_clk_debounce.debounced_button ),
    .B(net98));
 sg13g2_a21oi_1 _628_ (.A1(_226_),
    .A2(_227_),
    .Y(_228_),
    .B1(net217));
 sg13g2_nand2b_1 _629_ (.Y(_229_),
    .B(net217),
    .A_N(net98));
 sg13g2_nand2_1 _630_ (.Y(_230_),
    .A(\ps2_clk_debounce.debounced_button ),
    .B(_229_));
 sg13g2_a21oi_1 _631_ (.A1(_226_),
    .A2(_230_),
    .Y(_072_),
    .B1(net218));
 sg13g2_nor2_1 _632_ (.A(net253),
    .B(_229_),
    .Y(_231_));
 sg13g2_a22oi_1 _633_ (.Y(_232_),
    .B1(_226_),
    .B2(_231_),
    .A2(net98),
    .A1(net235));
 sg13g2_inv_1 _634_ (.Y(_073_),
    .A(net254));
 sg13g2_nand3b_1 _635_ (.B(_216_),
    .C(_220_),
    .Y(_233_),
    .A_N(_003_));
 sg13g2_o21ai_1 _636_ (.B1(_233_),
    .Y(_234_),
    .A1(_115_),
    .A2(_226_));
 sg13g2_or2_1 _637_ (.X(_235_),
    .B(net88),
    .A(_112_));
 sg13g2_nand2_1 _638_ (.Y(_236_),
    .A(net248),
    .B(net88));
 sg13g2_o21ai_1 _639_ (.B1(_236_),
    .Y(_074_),
    .A1(net248),
    .A2(net86));
 sg13g2_nand2_1 _640_ (.Y(_237_),
    .A(net232),
    .B(net88));
 sg13g2_xnor2_1 _641_ (.Y(_238_),
    .A(net232),
    .B(\ps2_decoder_inst.clk_timeout[0] ));
 sg13g2_o21ai_1 _642_ (.B1(_237_),
    .Y(_075_),
    .A1(net86),
    .A2(_238_));
 sg13g2_a21oi_1 _643_ (.A1(\ps2_decoder_inst.clk_timeout[1] ),
    .A2(\ps2_decoder_inst.clk_timeout[0] ),
    .Y(_239_),
    .B1(net220));
 sg13g2_nand2_1 _644_ (.Y(_240_),
    .A(net220),
    .B(net88));
 sg13g2_nand3_1 _645_ (.B(\ps2_decoder_inst.clk_timeout[0] ),
    .C(\ps2_decoder_inst.clk_timeout[2] ),
    .A(\ps2_decoder_inst.clk_timeout[1] ),
    .Y(_241_));
 sg13g2_nand2b_1 _646_ (.Y(_242_),
    .B(_241_),
    .A_N(_239_));
 sg13g2_o21ai_1 _647_ (.B1(_240_),
    .Y(_076_),
    .A1(net86),
    .A2(_242_));
 sg13g2_nand2_1 _648_ (.Y(_243_),
    .A(net78),
    .B(net88));
 sg13g2_nor2_2 _649_ (.A(_113_),
    .B(_241_),
    .Y(_244_));
 sg13g2_xnor2_1 _650_ (.Y(_245_),
    .A(_113_),
    .B(_241_));
 sg13g2_o21ai_1 _651_ (.B1(_243_),
    .Y(_077_),
    .A1(net86),
    .A2(_245_));
 sg13g2_nand2_1 _652_ (.Y(_246_),
    .A(net265),
    .B(net89));
 sg13g2_xnor2_1 _653_ (.Y(_247_),
    .A(net265),
    .B(_244_));
 sg13g2_o21ai_1 _654_ (.B1(_246_),
    .Y(_078_),
    .A1(net86),
    .A2(_247_));
 sg13g2_nand2_1 _655_ (.Y(_248_),
    .A(net237),
    .B(net89));
 sg13g2_a21oi_1 _656_ (.A1(\ps2_decoder_inst.clk_timeout[4] ),
    .A2(_244_),
    .Y(_249_),
    .B1(net237));
 sg13g2_nand3_1 _657_ (.B(\ps2_decoder_inst.clk_timeout[4] ),
    .C(_244_),
    .A(\ps2_decoder_inst.clk_timeout[5] ),
    .Y(_250_));
 sg13g2_nand2b_1 _658_ (.Y(_251_),
    .B(_250_),
    .A_N(_249_));
 sg13g2_o21ai_1 _659_ (.B1(_248_),
    .Y(_079_),
    .A1(net86),
    .A2(_251_));
 sg13g2_nand2_1 _660_ (.Y(_252_),
    .A(net222),
    .B(net89));
 sg13g2_nand4_1 _661_ (.B(\ps2_decoder_inst.clk_timeout[4] ),
    .C(\ps2_decoder_inst.clk_timeout[6] ),
    .A(\ps2_decoder_inst.clk_timeout[5] ),
    .Y(_253_),
    .D(_244_));
 sg13g2_xor2_1 _662_ (.B(_250_),
    .A(net222),
    .X(_254_));
 sg13g2_o21ai_1 _663_ (.B1(_252_),
    .Y(_080_),
    .A1(net86),
    .A2(_254_));
 sg13g2_nand2_1 _664_ (.Y(_255_),
    .A(net170),
    .B(net88));
 sg13g2_nor2b_1 _665_ (.A(net170),
    .B_N(_253_),
    .Y(_256_));
 sg13g2_and4_2 _666_ (.A(\ps2_decoder_inst.clk_timeout[5] ),
    .B(\ps2_decoder_inst.clk_timeout[4] ),
    .C(_215_),
    .D(_244_),
    .X(_257_));
 sg13g2_or2_1 _667_ (.X(_258_),
    .B(_257_),
    .A(_256_));
 sg13g2_o21ai_1 _668_ (.B1(_255_),
    .Y(_081_),
    .A1(net87),
    .A2(_258_));
 sg13g2_nand2_1 _669_ (.Y(_259_),
    .A(net252),
    .B(net88));
 sg13g2_xnor2_1 _670_ (.Y(_260_),
    .A(net252),
    .B(_257_));
 sg13g2_o21ai_1 _671_ (.B1(_259_),
    .Y(_082_),
    .A1(net87),
    .A2(_260_));
 sg13g2_nand2_1 _672_ (.Y(_261_),
    .A(net230),
    .B(net88));
 sg13g2_nand3_1 _673_ (.B(\ps2_decoder_inst.clk_timeout[8] ),
    .C(_257_),
    .A(net230),
    .Y(_262_));
 sg13g2_a21o_1 _674_ (.A2(_257_),
    .A1(\ps2_decoder_inst.clk_timeout[8] ),
    .B1(net230),
    .X(_263_));
 sg13g2_nand2_1 _675_ (.Y(_264_),
    .A(_262_),
    .B(_263_));
 sg13g2_o21ai_1 _676_ (.B1(_261_),
    .Y(_083_),
    .A1(net87),
    .A2(_264_));
 sg13g2_nand2_1 _677_ (.Y(_265_),
    .A(net228),
    .B(net89));
 sg13g2_nand4_1 _678_ (.B(\ps2_decoder_inst.clk_timeout[8] ),
    .C(net228),
    .A(net230),
    .Y(_266_),
    .D(_257_));
 sg13g2_xor2_1 _679_ (.B(_262_),
    .A(net228),
    .X(_267_));
 sg13g2_o21ai_1 _680_ (.B1(_265_),
    .Y(_084_),
    .A1(net87),
    .A2(_267_));
 sg13g2_nand2_1 _681_ (.Y(_268_),
    .A(net164),
    .B(net89));
 sg13g2_xnor2_1 _682_ (.Y(_269_),
    .A(_114_),
    .B(_266_));
 sg13g2_o21ai_1 _683_ (.B1(_268_),
    .Y(_085_),
    .A1(net86),
    .A2(_269_));
 sg13g2_xor2_1 _684_ (.B(\ps2_decoder_inst.shift_reg[5] ),
    .A(\ps2_decoder_inst.shift_reg[4] ),
    .X(_270_));
 sg13g2_xnor2_1 _685_ (.Y(_271_),
    .A(\ps2_decoder_inst.shift_reg[6] ),
    .B(_270_));
 sg13g2_xor2_1 _686_ (.B(\ps2_decoder_inst.shift_reg[7] ),
    .A(\ps2_decoder_inst.shift_reg[3] ),
    .X(_272_));
 sg13g2_xor2_1 _687_ (.B(\ps2_decoder_inst.shift_reg[2] ),
    .A(\ps2_decoder_inst.shift_reg[1] ),
    .X(_273_));
 sg13g2_xnor2_1 _688_ (.Y(_274_),
    .A(_272_),
    .B(_273_));
 sg13g2_xnor2_1 _689_ (.Y(_275_),
    .A(\ps2_decoder_inst.shift_reg[8] ),
    .B(\ps2_decoder_inst.shift_reg[9] ));
 sg13g2_xnor2_1 _690_ (.Y(_276_),
    .A(_274_),
    .B(_275_));
 sg13g2_xnor2_1 _691_ (.Y(_277_),
    .A(_271_),
    .B(_276_));
 sg13g2_nor2b_1 _692_ (.A(\ps2_decoder_inst.state_reg[0] ),
    .B_N(net97),
    .Y(_278_));
 sg13g2_o21ai_1 _693_ (.B1(_226_),
    .Y(_279_),
    .A1(_230_),
    .A2(_278_));
 sg13g2_nand3b_1 _694_ (.B(net44),
    .C(net235),
    .Y(_280_),
    .A_N(\ps2_decoder_inst.shift_reg[10] ));
 sg13g2_nor4_1 _695_ (.A(_277_),
    .B(_278_),
    .C(_279_),
    .D(_280_),
    .Y(_281_));
 sg13g2_a21o_1 _696_ (.A2(_279_),
    .A1(net242),
    .B1(_281_),
    .X(_086_));
 sg13g2_a21oi_1 _697_ (.A1(_216_),
    .A2(_220_),
    .Y(_282_),
    .B1(\ps2_decoder_inst.clk_timeout[12] ));
 sg13g2_o21ai_1 _698_ (.B1(_282_),
    .Y(_283_),
    .A1(_114_),
    .A2(_266_));
 sg13g2_or3_1 _699_ (.A(_003_),
    .B(_225_),
    .C(_278_),
    .X(_284_));
 sg13g2_and3_1 _700_ (.X(_087_),
    .A(net235),
    .B(_283_),
    .C(_284_));
 sg13g2_nor2b_1 _701_ (.A(net98),
    .B_N(net60),
    .Y(_285_));
 sg13g2_nor3_2 _702_ (.A(net217),
    .B(_003_),
    .C(_225_),
    .Y(_286_));
 sg13g2_mux2_1 _703_ (.A0(net261),
    .A1(_285_),
    .S(net85),
    .X(_088_));
 sg13g2_nor2b_1 _704_ (.A(net98),
    .B_N(\ps2_decoder_inst.shift_reg[8] ),
    .Y(_287_));
 sg13g2_mux2_1 _705_ (.A0(net255),
    .A1(_287_),
    .S(net85),
    .X(_089_));
 sg13g2_nor2b_1 _706_ (.A(net97),
    .B_N(net48),
    .Y(_288_));
 sg13g2_mux2_1 _707_ (.A0(net251),
    .A1(_288_),
    .S(net85),
    .X(_090_));
 sg13g2_nor2b_1 _708_ (.A(net97),
    .B_N(net58),
    .Y(_289_));
 sg13g2_mux2_1 _709_ (.A0(net266),
    .A1(_289_),
    .S(net85),
    .X(_091_));
 sg13g2_nor2b_1 _710_ (.A(net97),
    .B_N(net56),
    .Y(_290_));
 sg13g2_mux2_1 _711_ (.A0(net268),
    .A1(_290_),
    .S(net85),
    .X(_092_));
 sg13g2_nor2b_1 _712_ (.A(net97),
    .B_N(net62),
    .Y(_291_));
 sg13g2_mux2_1 _713_ (.A0(net259),
    .A1(_291_),
    .S(net85),
    .X(_093_));
 sg13g2_nor2b_1 _714_ (.A(net97),
    .B_N(\ps2_decoder_inst.shift_reg[3] ),
    .Y(_292_));
 sg13g2_mux2_1 _715_ (.A0(net257),
    .A1(_292_),
    .S(net85),
    .X(_094_));
 sg13g2_nor2b_1 _716_ (.A(net97),
    .B_N(\ps2_decoder_inst.shift_reg[2] ),
    .Y(_293_));
 sg13g2_mux2_1 _717_ (.A0(net263),
    .A1(_293_),
    .S(net85),
    .X(_095_));
 sg13g2_a21o_1 _718_ (.A2(net215),
    .A1(_118_),
    .B1(\ps2_decoder_inst.valid_reg ),
    .X(_096_));
 sg13g2_nor2_1 _719_ (.A(_229_),
    .B(_233_),
    .Y(_294_));
 sg13g2_nor2_1 _720_ (.A(net245),
    .B(_294_),
    .Y(_295_));
 sg13g2_a21oi_1 _721_ (.A1(net97),
    .A2(_286_),
    .Y(_097_),
    .B1(net246));
 sg13g2_nand2_1 _722_ (.Y(_296_),
    .A(\ps2_data_debounce.debounced_button ),
    .B(net94));
 sg13g2_o21ai_1 _723_ (.B1(_296_),
    .Y(_098_),
    .A1(net71),
    .A2(_132_));
 sg13g2_a21oi_2 _724_ (.B1(\ps2_decoder_inst.shift_reset ),
    .Y(_297_),
    .A2(_112_),
    .A1(\ps2_decoder_inst.ps2_clk_prev ));
 sg13g2_nand2_1 _725_ (.Y(_298_),
    .A(net69),
    .B(net91));
 sg13g2_nand3b_1 _726_ (.B(\ps2_decoder_inst.ps2_clk_prev ),
    .C(_112_),
    .Y(_299_),
    .A_N(\ps2_decoder_inst.shift_reset ));
 sg13g2_o21ai_1 _727_ (.B1(_298_),
    .Y(_099_),
    .A1(\ps2_data_debounce.debounced_button ),
    .A2(_299_));
 sg13g2_nand2_1 _728_ (.Y(_300_),
    .A(_401_),
    .B(_297_));
 sg13g2_o21ai_1 _729_ (.B1(_300_),
    .Y(_100_),
    .A1(net44),
    .A2(net90));
 sg13g2_nand2_1 _730_ (.Y(_301_),
    .A(_402_),
    .B(net91));
 sg13g2_o21ai_1 _731_ (.B1(_301_),
    .Y(_101_),
    .A1(net50),
    .A2(net90));
 sg13g2_nand2_1 _732_ (.Y(_302_),
    .A(net73),
    .B(net91));
 sg13g2_o21ai_1 _733_ (.B1(_302_),
    .Y(_102_),
    .A1(\ps2_decoder_inst.shift_reg[2] ),
    .A2(net90));
 sg13g2_nand2_1 _734_ (.Y(_303_),
    .A(net67),
    .B(net91));
 sg13g2_o21ai_1 _735_ (.B1(_303_),
    .Y(_103_),
    .A1(\ps2_decoder_inst.shift_reg[3] ),
    .A2(net90));
 sg13g2_nand2_1 _736_ (.Y(_304_),
    .A(_405_),
    .B(net91));
 sg13g2_o21ai_1 _737_ (.B1(_304_),
    .Y(_104_),
    .A1(net62),
    .A2(net90));
 sg13g2_nand2_1 _738_ (.Y(_305_),
    .A(_406_),
    .B(net91));
 sg13g2_o21ai_1 _739_ (.B1(_305_),
    .Y(_105_),
    .A1(net56),
    .A2(net90));
 sg13g2_nand2_1 _740_ (.Y(_306_),
    .A(_407_),
    .B(net91));
 sg13g2_o21ai_1 _741_ (.B1(_306_),
    .Y(_106_),
    .A1(net58),
    .A2(net90));
 sg13g2_nand2_1 _742_ (.Y(_307_),
    .A(_408_),
    .B(net91));
 sg13g2_o21ai_1 _743_ (.B1(_307_),
    .Y(_107_),
    .A1(net48),
    .A2(net90));
 sg13g2_nand2_1 _744_ (.Y(_308_),
    .A(net64),
    .B(_297_));
 sg13g2_o21ai_1 _745_ (.B1(net65),
    .Y(_108_),
    .A1(\ps2_decoder_inst.shift_reg[8] ),
    .A2(_299_));
 sg13g2_nand2_1 _746_ (.Y(_309_),
    .A(_410_),
    .B(_297_));
 sg13g2_o21ai_1 _747_ (.B1(_309_),
    .Y(_109_),
    .A1(net60),
    .A2(_299_));
 sg13g2_dfrbp_1 _748_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net21),
    .D(net192),
    .Q_N(_394_),
    .Q(\memory.mem[3][0] ));
 sg13g2_dfrbp_1 _749_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net28),
    .D(net145),
    .Q_N(_393_),
    .Q(\memory.mem[3][1] ));
 sg13g2_dfrbp_1 _750_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net27),
    .D(net161),
    .Q_N(_392_),
    .Q(\memory.mem[3][2] ));
 sg13g2_dfrbp_1 _751_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net26),
    .D(net137),
    .Q_N(_391_),
    .Q(\memory.mem[3][3] ));
 sg13g2_dfrbp_1 _752_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net25),
    .D(net186),
    .Q_N(_390_),
    .Q(\memory.mem[3][4] ));
 sg13g2_dfrbp_1 _753_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net24),
    .D(net139),
    .Q_N(_389_),
    .Q(\memory.mem[3][5] ));
 sg13g2_dfrbp_1 _754_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net23),
    .D(net126),
    .Q_N(_388_),
    .Q(\memory.mem[3][6] ));
 sg13g2_dfrbp_1 _755_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net22),
    .D(net176),
    .Q_N(_387_),
    .Q(\memory.mem[3][7] ));
 sg13g2_dfrbp_1 _756_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net106),
    .D(net132),
    .Q_N(_386_),
    .Q(\ps2_clk_debounce.counter[0] ));
 sg13g2_dfrbp_1 _757_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net106),
    .D(net77),
    .Q_N(_385_),
    .Q(\ps2_clk_debounce.counter[1] ));
 sg13g2_dfrbp_1 _758_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net106),
    .D(net83),
    .Q_N(_384_),
    .Q(\ps2_clk_debounce.counter[2] ));
 sg13g2_dfrbp_1 _759_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net106),
    .D(net198),
    .Q_N(_383_),
    .Q(\ps2_clk_debounce.counter[3] ));
 sg13g2_dfrbp_1 _760_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net109),
    .D(net115),
    .Q_N(_382_),
    .Q(\ps2_clk_debounce.counter[4] ));
 sg13g2_dfrbp_1 _761_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net109),
    .D(net122),
    .Q_N(_381_),
    .Q(\ps2_clk_debounce.counter[5] ));
 sg13g2_dfrbp_1 _762_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net109),
    .D(net149),
    .Q_N(_395_),
    .Q(\ps2_clk_debounce.counter[6] ));
 sg13g2_dfrbp_1 _763_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net109),
    .D(net1),
    .Q_N(_396_),
    .Q(\ps2_clk_debounce.last_button ));
 sg13g2_dfrbp_1 _764_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net101),
    .D(net5),
    .Q_N(_397_),
    .Q(cs_prev));
 sg13g2_dfrbp_1 _765_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net108),
    .D(_000_),
    .Q_N(_380_),
    .Q(cs_trigger));
 sg13g2_dfrbp_1 _766_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net104),
    .D(net211),
    .Q_N(_003_),
    .Q(\ps2_clk_debounce.debounced_button ));
 sg13g2_dfrbp_1 _767_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net109),
    .D(net128),
    .Q_N(_379_),
    .Q(\ps2_data_debounce.counter[0] ));
 sg13g2_dfrbp_1 _768_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net109),
    .D(net118),
    .Q_N(_378_),
    .Q(\ps2_data_debounce.counter[1] ));
 sg13g2_dfrbp_1 _769_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net109),
    .D(net124),
    .Q_N(_377_),
    .Q(\ps2_data_debounce.counter[2] ));
 sg13g2_dfrbp_1 _770_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net110),
    .D(net207),
    .Q_N(_376_),
    .Q(\ps2_data_debounce.counter[3] ));
 sg13g2_dfrbp_1 _771_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net110),
    .D(net135),
    .Q_N(_375_),
    .Q(\ps2_data_debounce.counter[4] ));
 sg13g2_dfrbp_1 _772_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net110),
    .D(net120),
    .Q_N(_374_),
    .Q(\ps2_data_debounce.counter[5] ));
 sg13g2_dfrbp_1 _773_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net110),
    .D(net112),
    .Q_N(_398_),
    .Q(\ps2_data_debounce.counter[6] ));
 sg13g2_dfrbp_1 _774_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net110),
    .D(net2),
    .Q_N(_373_),
    .Q(\ps2_data_debounce.last_button ));
 sg13g2_dfrbp_1 _775_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net103),
    .D(net205),
    .Q_N(_372_),
    .Q(\ps2_decoder_inst.ps2_clk_prev ));
 sg13g2_dfrbp_1 _776_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net20),
    .D(net209),
    .Q_N(_371_),
    .Q(\memory.mem[1][0] ));
 sg13g2_dfrbp_1 _777_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net19),
    .D(net143),
    .Q_N(_370_),
    .Q(\memory.mem[1][1] ));
 sg13g2_dfrbp_1 _778_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net18),
    .D(net153),
    .Q_N(_369_),
    .Q(\memory.mem[1][2] ));
 sg13g2_dfrbp_1 _779_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net17),
    .D(net194),
    .Q_N(_368_),
    .Q(\memory.mem[1][3] ));
 sg13g2_dfrbp_1 _780_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net16),
    .D(net147),
    .Q_N(_367_),
    .Q(\memory.mem[1][4] ));
 sg13g2_dfrbp_1 _781_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net15),
    .D(net163),
    .Q_N(_366_),
    .Q(\memory.mem[1][5] ));
 sg13g2_dfrbp_1 _782_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net14),
    .D(net151),
    .Q_N(_365_),
    .Q(\memory.mem[1][6] ));
 sg13g2_dfrbp_1 _783_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net13),
    .D(net182),
    .Q_N(_364_),
    .Q(\memory.mem[1][7] ));
 sg13g2_dfrbp_1 _784_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net108),
    .D(net55),
    .Q_N(_008_),
    .Q(\memory.wr_ptr[0] ));
 sg13g2_dfrbp_1 _785_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net108),
    .D(net240),
    .Q_N(_363_),
    .Q(\memory.wr_ptr[1] ));
 sg13g2_dfrbp_1 _786_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net101),
    .D(net47),
    .Q_N(_007_),
    .Q(\memory.rd_ptr[0] ));
 sg13g2_dfrbp_1 _787_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net101),
    .D(_044_),
    .Q_N(_362_),
    .Q(\memory.rd_ptr[1] ));
 sg13g2_dfrbp_1 _788_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net12),
    .D(net202),
    .Q_N(_361_),
    .Q(\memory.mem[2][0] ));
 sg13g2_dfrbp_1 _789_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net11),
    .D(net200),
    .Q_N(_360_),
    .Q(\memory.mem[2][1] ));
 sg13g2_dfrbp_1 _790_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net42),
    .D(net174),
    .Q_N(_359_),
    .Q(\memory.mem[2][2] ));
 sg13g2_dfrbp_1 _791_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net41),
    .D(net172),
    .Q_N(_358_),
    .Q(\memory.mem[2][3] ));
 sg13g2_dfrbp_1 _792_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net40),
    .D(net159),
    .Q_N(_357_),
    .Q(\memory.mem[2][4] ));
 sg13g2_dfrbp_1 _793_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net39),
    .D(net190),
    .Q_N(_356_),
    .Q(\memory.mem[2][5] ));
 sg13g2_dfrbp_1 _794_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net38),
    .D(net178),
    .Q_N(_355_),
    .Q(\memory.mem[2][6] ));
 sg13g2_dfrbp_1 _795_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net37),
    .D(net155),
    .Q_N(_354_),
    .Q(\memory.mem[2][7] ));
 sg13g2_dfrbp_1 _796_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net36),
    .D(net141),
    .Q_N(_353_),
    .Q(\memory.mem[0][0] ));
 sg13g2_dfrbp_1 _797_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net35),
    .D(net188),
    .Q_N(_352_),
    .Q(\memory.mem[0][1] ));
 sg13g2_dfrbp_1 _798_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net34),
    .D(net169),
    .Q_N(_351_),
    .Q(\memory.mem[0][2] ));
 sg13g2_dfrbp_1 _799_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net33),
    .D(net130),
    .Q_N(_350_),
    .Q(\memory.mem[0][3] ));
 sg13g2_dfrbp_1 _800_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net32),
    .D(net167),
    .Q_N(_349_),
    .Q(\memory.mem[0][4] ));
 sg13g2_dfrbp_1 _801_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net31),
    .D(net157),
    .Q_N(_348_),
    .Q(\memory.mem[0][5] ));
 sg13g2_dfrbp_1 _802_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net30),
    .D(net196),
    .Q_N(_347_),
    .Q(\memory.mem[0][6] ));
 sg13g2_dfrbp_1 _803_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net29),
    .D(net184),
    .Q_N(_346_),
    .Q(\memory.mem[0][7] ));
 sg13g2_dfrbp_1 _804_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net102),
    .D(_061_),
    .Q_N(_345_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _805_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net102),
    .D(_062_),
    .Q_N(_344_),
    .Q(uio_out[1]));
 sg13g2_dfrbp_1 _806_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net102),
    .D(_063_),
    .Q_N(_343_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _807_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net101),
    .D(_064_),
    .Q_N(_342_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _808_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net101),
    .D(_065_),
    .Q_N(_341_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _809_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net101),
    .D(_066_),
    .Q_N(_340_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _810_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net101),
    .D(_067_),
    .Q_N(_339_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _811_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net101),
    .D(_068_),
    .Q_N(_338_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _812_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net108),
    .D(net180),
    .Q_N(_006_),
    .Q(\memory.count[0] ));
 sg13g2_dfrbp_1 _813_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net111),
    .D(_070_),
    .Q_N(_337_),
    .Q(\memory.count[1] ));
 sg13g2_dfrbp_1 _814_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net108),
    .D(net214),
    .Q_N(_336_),
    .Q(\memory.count[2] ));
 sg13g2_dfrbp_1 _815_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net104),
    .D(net219),
    .Q_N(_335_),
    .Q(\ps2_decoder_inst.state_reg[0] ));
 sg13g2_dfrbp_1 _816_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net103),
    .D(_073_),
    .Q_N(_399_),
    .Q(\ps2_decoder_inst.state_reg[1] ));
 sg13g2_dfrbp_1 _817_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net106),
    .D(net53),
    .Q_N(_004_),
    .Q(\ps2_clk_debounce.counter[7] ));
 sg13g2_dfrbp_1 _818_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net110),
    .D(net72),
    .Q_N(_005_),
    .Q(\ps2_data_debounce.counter[7] ));
 sg13g2_dfrbp_1 _819_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net103),
    .D(_074_),
    .Q_N(_334_),
    .Q(\ps2_decoder_inst.clk_timeout[0] ));
 sg13g2_dfrbp_1 _820_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net103),
    .D(net233),
    .Q_N(_333_),
    .Q(\ps2_decoder_inst.clk_timeout[1] ));
 sg13g2_dfrbp_1 _821_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net105),
    .D(net221),
    .Q_N(_332_),
    .Q(\ps2_decoder_inst.clk_timeout[2] ));
 sg13g2_dfrbp_1 _822_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net103),
    .D(net79),
    .Q_N(_331_),
    .Q(\ps2_decoder_inst.clk_timeout[3] ));
 sg13g2_dfrbp_1 _823_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net105),
    .D(_078_),
    .Q_N(_330_),
    .Q(\ps2_decoder_inst.clk_timeout[4] ));
 sg13g2_dfrbp_1 _824_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net105),
    .D(net238),
    .Q_N(_329_),
    .Q(\ps2_decoder_inst.clk_timeout[5] ));
 sg13g2_dfrbp_1 _825_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net105),
    .D(net223),
    .Q_N(_328_),
    .Q(\ps2_decoder_inst.clk_timeout[6] ));
 sg13g2_dfrbp_1 _826_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net105),
    .D(_081_),
    .Q_N(_327_),
    .Q(\ps2_decoder_inst.clk_timeout[7] ));
 sg13g2_dfrbp_1 _827_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net105),
    .D(_082_),
    .Q_N(_326_),
    .Q(\ps2_decoder_inst.clk_timeout[8] ));
 sg13g2_dfrbp_1 _828_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net105),
    .D(net231),
    .Q_N(_325_),
    .Q(\ps2_decoder_inst.clk_timeout[9] ));
 sg13g2_dfrbp_1 _829_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net106),
    .D(net229),
    .Q_N(_324_),
    .Q(\ps2_decoder_inst.clk_timeout[10] ));
 sg13g2_dfrbp_1 _830_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net106),
    .D(net165),
    .Q_N(_323_),
    .Q(\ps2_decoder_inst.clk_timeout[11] ));
 sg13g2_dfrbp_1 _831_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net103),
    .D(net243),
    .Q_N(_322_),
    .Q(\ps2_decoder_inst.valid_reg ));
 sg13g2_dfrbp_1 _832_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net105),
    .D(net236),
    .Q_N(_321_),
    .Q(\ps2_decoder_inst.clk_timeout[12] ));
 sg13g2_dfrbp_1 _833_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net104),
    .D(net262),
    .Q_N(_320_),
    .Q(\ps2_decoder_inst.ps2_value[0] ));
 sg13g2_dfrbp_1 _834_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net100),
    .D(net256),
    .Q_N(_319_),
    .Q(\ps2_decoder_inst.ps2_value[1] ));
 sg13g2_dfrbp_1 _835_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net100),
    .D(_090_),
    .Q_N(_318_),
    .Q(\ps2_decoder_inst.ps2_value[2] ));
 sg13g2_dfrbp_1 _836_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net99),
    .D(net267),
    .Q_N(_317_),
    .Q(\ps2_decoder_inst.ps2_value[3] ));
 sg13g2_dfrbp_1 _837_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net100),
    .D(_092_),
    .Q_N(_316_),
    .Q(\ps2_decoder_inst.ps2_value[4] ));
 sg13g2_dfrbp_1 _838_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net99),
    .D(_093_),
    .Q_N(_315_),
    .Q(\ps2_decoder_inst.ps2_value[5] ));
 sg13g2_dfrbp_1 _839_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net99),
    .D(net258),
    .Q_N(_314_),
    .Q(\ps2_decoder_inst.ps2_value[6] ));
 sg13g2_dfrbp_1 _840_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net99),
    .D(net264),
    .Q_N(_313_),
    .Q(\ps2_decoder_inst.ps2_value[7] ));
 sg13g2_dfrbp_1 _841_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net108),
    .D(net216),
    .Q_N(_312_),
    .Q(\ps2_decoder_inst.int_reg ));
 sg13g2_dfrbp_1 _842_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net103),
    .D(net247),
    .Q_N(_311_),
    .Q(\ps2_decoder_inst.shift_reset ));
 sg13g2_dfrbp_1 _843_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net109),
    .D(net81),
    .Q_N(_310_),
    .Q(\ps2_data_debounce.debounced_button ));
 sg13g2_dfrbp_1 _844_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net103),
    .D(net70),
    .Q_N(\ps2_decoder_inst.shift_reg[0] ),
    .Q(_400_));
 sg13g2_dfrbp_1 _845_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net100),
    .D(net45),
    .Q_N(\ps2_decoder_inst.shift_reg[1] ),
    .Q(_401_));
 sg13g2_dfrbp_1 _846_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net100),
    .D(net51),
    .Q_N(\ps2_decoder_inst.shift_reg[2] ),
    .Q(_402_));
 sg13g2_dfrbp_1 _847_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net99),
    .D(net74),
    .Q_N(\ps2_decoder_inst.shift_reg[3] ),
    .Q(_403_));
 sg13g2_dfrbp_1 _848_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net99),
    .D(net68),
    .Q_N(\ps2_decoder_inst.shift_reg[4] ),
    .Q(_404_));
 sg13g2_dfrbp_1 _849_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net99),
    .D(net63),
    .Q_N(\ps2_decoder_inst.shift_reg[5] ),
    .Q(_405_));
 sg13g2_dfrbp_1 _850_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net100),
    .D(net57),
    .Q_N(\ps2_decoder_inst.shift_reg[6] ),
    .Q(_406_));
 sg13g2_dfrbp_1 _851_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net99),
    .D(net59),
    .Q_N(\ps2_decoder_inst.shift_reg[7] ),
    .Q(_407_));
 sg13g2_dfrbp_1 _852_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net102),
    .D(net49),
    .Q_N(\ps2_decoder_inst.shift_reg[8] ),
    .Q(_408_));
 sg13g2_dfrbp_1 _853_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net100),
    .D(net66),
    .Q_N(\ps2_decoder_inst.shift_reg[9] ),
    .Q(_409_));
 sg13g2_dfrbp_1 _854_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net104),
    .D(net61),
    .Q_N(\ps2_decoder_inst.shift_reg[10] ),
    .Q(_410_));
 sg13g2_tiehi _788__12 (.L_HI(net12));
 sg13g2_tiehi _783__13 (.L_HI(net13));
 sg13g2_tiehi _782__14 (.L_HI(net14));
 sg13g2_tiehi _781__15 (.L_HI(net15));
 sg13g2_tiehi _780__16 (.L_HI(net16));
 sg13g2_tiehi _779__17 (.L_HI(net17));
 sg13g2_tiehi _778__18 (.L_HI(net18));
 sg13g2_tiehi _777__19 (.L_HI(net19));
 sg13g2_tiehi _776__20 (.L_HI(net20));
 sg13g2_tiehi _748__21 (.L_HI(net21));
 sg13g2_tiehi _755__22 (.L_HI(net22));
 sg13g2_tiehi _754__23 (.L_HI(net23));
 sg13g2_tiehi _753__24 (.L_HI(net24));
 sg13g2_tiehi _752__25 (.L_HI(net25));
 sg13g2_tiehi _751__26 (.L_HI(net26));
 sg13g2_tiehi _750__27 (.L_HI(net27));
 sg13g2_tiehi _749__28 (.L_HI(net28));
 sg13g2_tiehi _803__29 (.L_HI(net29));
 sg13g2_tiehi _802__30 (.L_HI(net30));
 sg13g2_tiehi _801__31 (.L_HI(net31));
 sg13g2_tiehi _800__32 (.L_HI(net32));
 sg13g2_tiehi _799__33 (.L_HI(net33));
 sg13g2_tiehi _798__34 (.L_HI(net34));
 sg13g2_tiehi _797__35 (.L_HI(net35));
 sg13g2_tiehi _796__36 (.L_HI(net36));
 sg13g2_tiehi _795__37 (.L_HI(net37));
 sg13g2_tiehi _794__38 (.L_HI(net38));
 sg13g2_tiehi _793__39 (.L_HI(net39));
 sg13g2_tiehi _792__40 (.L_HI(net40));
 sg13g2_tiehi _791__41 (.L_HI(net41));
 sg13g2_tiehi _790__42 (.L_HI(net42));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_benpayne_ps2_decoder_7 (.L_LO(net7));
 sg13g2_tielo tt_um_benpayne_ps2_decoder_8 (.L_LO(net8));
 sg13g2_tielo tt_um_benpayne_ps2_decoder_9 (.L_LO(net9));
 sg13g2_tielo tt_um_benpayne_ps2_decoder_10 (.L_LO(net10));
 sg13g2_tiehi _789__11 (.L_HI(net11));
 sg13g2_buf_1 _892_ (.A(net5),
    .X(uio_oe[0]));
 sg13g2_buf_1 _893_ (.A(net5),
    .X(uio_oe[1]));
 sg13g2_buf_1 _894_ (.A(net5),
    .X(uio_oe[2]));
 sg13g2_buf_1 _895_ (.A(net5),
    .X(uio_oe[3]));
 sg13g2_buf_1 _896_ (.A(net5),
    .X(uio_oe[4]));
 sg13g2_buf_1 _897_ (.A(net5),
    .X(uio_oe[5]));
 sg13g2_buf_1 _898_ (.A(net5),
    .X(uio_oe[6]));
 sg13g2_buf_1 _899_ (.A(net4),
    .X(uio_oe[7]));
 sg13g2_buf_1 _900_ (.A(\ps2_decoder_inst.valid_reg ),
    .X(uo_out[0]));
 sg13g2_buf_1 _901_ (.A(\ps2_decoder_inst.int_reg ),
    .X(uo_out[1]));
 sg13g2_buf_4 fanout85 (.X(net85),
    .A(_286_));
 sg13g2_buf_2 fanout86 (.A(_235_),
    .X(net86));
 sg13g2_buf_1 fanout87 (.A(_235_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_234_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_234_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_299_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_297_),
    .X(net91));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(net93));
 sg13g2_buf_2 fanout93 (.A(_175_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_135_),
    .X(net94));
 sg13g2_buf_4 fanout95 (.X(net95),
    .A(_177_));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(_176_));
 sg13g2_buf_2 fanout97 (.A(\ps2_decoder_inst.state_reg[1] ),
    .X(net97));
 sg13g2_buf_1 fanout98 (.A(\ps2_decoder_inst.state_reg[1] ),
    .X(net98));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(net100));
 sg13g2_buf_4 fanout100 (.X(net100),
    .A(net102));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(net102));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(rst_n));
 sg13g2_buf_4 fanout103 (.X(net103),
    .A(net107));
 sg13g2_buf_2 fanout104 (.A(net107),
    .X(net104));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(net107));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(net107));
 sg13g2_buf_2 fanout107 (.A(rst_n),
    .X(net107));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(net111));
 sg13g2_buf_4 fanout109 (.X(net109),
    .A(net111));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(net111));
 sg13g2_buf_2 fanout111 (.A(rst_n),
    .X(net111));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 fanout5 (.A(net4),
    .X(net5));
 sg13g2_tielo tt_um_benpayne_ps2_decoder_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(cs_prev),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold2 (.A(\ps2_decoder_inst.shift_reg[0] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold3 (.A(_100_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold4 (.A(_007_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold5 (.A(_043_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold6 (.A(\ps2_decoder_inst.shift_reg[7] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold7 (.A(_107_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold8 (.A(\ps2_decoder_inst.shift_reg[1] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold9 (.A(_101_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold10 (.A(_004_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold11 (.A(_001_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold12 (.A(_008_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold13 (.A(_041_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold14 (.A(\ps2_decoder_inst.shift_reg[5] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold15 (.A(_105_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold16 (.A(\ps2_decoder_inst.shift_reg[6] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold17 (.A(_106_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold18 (.A(\ps2_decoder_inst.shift_reg[9] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold19 (.A(_109_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold20 (.A(\ps2_decoder_inst.shift_reg[4] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold21 (.A(_104_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold22 (.A(_409_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold23 (.A(_308_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold24 (.A(_108_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold25 (.A(_404_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold26 (.A(_103_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold27 (.A(_400_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold28 (.A(_099_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold29 (.A(_005_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold30 (.A(_002_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold31 (.A(_403_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold32 (.A(_102_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold33 (.A(\ps2_clk_debounce.counter[1] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold34 (.A(_149_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold35 (.A(_018_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold36 (.A(\ps2_decoder_inst.clk_timeout[3] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold37 (.A(_077_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold38 (.A(\ps2_data_debounce.last_button ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold39 (.A(_098_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold40 (.A(\ps2_clk_debounce.counter[2] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold41 (.A(_019_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold42 (.A(\ps2_data_debounce.counter[6] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold43 (.A(_031_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold44 (.A(\ps2_clk_debounce.counter[4] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold45 (.A(_154_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold46 (.A(_021_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold47 (.A(\ps2_data_debounce.counter[1] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold48 (.A(_164_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold49 (.A(_026_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold50 (.A(\ps2_data_debounce.counter[5] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold51 (.A(_030_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold52 (.A(\ps2_clk_debounce.counter[5] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold53 (.A(_022_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold54 (.A(\ps2_data_debounce.counter[2] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold55 (.A(_027_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold56 (.A(\memory.mem[3][6] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold57 (.A(_015_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold58 (.A(\ps2_data_debounce.counter[0] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold59 (.A(_025_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold60 (.A(\memory.mem[0][3] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold61 (.A(_056_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold62 (.A(\ps2_clk_debounce.counter[0] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold63 (.A(_017_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold64 (.A(\ps2_data_debounce.counter[4] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold65 (.A(_169_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold66 (.A(_029_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold67 (.A(\memory.mem[3][3] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold68 (.A(_012_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold69 (.A(\memory.mem[3][5] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold70 (.A(_014_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold71 (.A(\memory.mem[0][0] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold72 (.A(_053_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold73 (.A(\memory.mem[1][1] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold74 (.A(_034_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold75 (.A(\memory.mem[3][1] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold76 (.A(_010_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold77 (.A(\memory.mem[1][4] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold78 (.A(_037_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold79 (.A(\ps2_clk_debounce.counter[6] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold80 (.A(_023_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold81 (.A(\memory.mem[1][6] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold82 (.A(_039_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold83 (.A(\memory.mem[1][2] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold84 (.A(_035_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold85 (.A(\memory.mem[2][7] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold86 (.A(_052_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold87 (.A(\memory.mem[0][5] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold88 (.A(_058_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold89 (.A(\memory.mem[2][4] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold90 (.A(_049_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold91 (.A(\memory.mem[3][2] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold92 (.A(_011_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold93 (.A(\memory.mem[1][5] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold94 (.A(_038_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold95 (.A(\ps2_decoder_inst.clk_timeout[11] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold96 (.A(_085_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold97 (.A(\memory.mem[0][4] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold98 (.A(_057_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold99 (.A(\memory.mem[0][2] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold100 (.A(_055_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold101 (.A(\ps2_decoder_inst.clk_timeout[7] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold102 (.A(\memory.mem[2][3] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold103 (.A(_048_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold104 (.A(\memory.mem[2][2] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold105 (.A(_047_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold106 (.A(\memory.mem[3][7] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold107 (.A(_016_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold108 (.A(\memory.mem[2][6] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold109 (.A(_051_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold110 (.A(_006_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold111 (.A(_069_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold112 (.A(\memory.mem[1][7] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold113 (.A(_040_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold114 (.A(\memory.mem[0][7] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold115 (.A(_060_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold116 (.A(\memory.mem[3][4] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold117 (.A(_013_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold118 (.A(\memory.mem[0][1] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold119 (.A(_054_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold120 (.A(\memory.mem[2][5] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold121 (.A(_050_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold122 (.A(\memory.mem[3][0] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold123 (.A(_009_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold124 (.A(\memory.mem[1][3] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold125 (.A(_036_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold126 (.A(\memory.mem[0][6] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold127 (.A(_059_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold128 (.A(\ps2_clk_debounce.counter[3] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold129 (.A(_020_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold130 (.A(\memory.mem[2][1] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold131 (.A(_046_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold132 (.A(\memory.mem[2][0] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold133 (.A(_045_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold134 (.A(\ps2_decoder_inst.ps2_clk_prev ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold135 (.A(_173_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold136 (.A(_032_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold137 (.A(\ps2_data_debounce.counter[3] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold138 (.A(_028_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold139 (.A(\memory.mem[1][0] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold140 (.A(_033_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold141 (.A(\ps2_clk_debounce.last_button ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold142 (.A(_024_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold143 (.A(\memory.count[0] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold144 (.A(_212_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold145 (.A(_071_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold146 (.A(\ps2_decoder_inst.int_reg ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold147 (.A(_096_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold148 (.A(\ps2_decoder_inst.state_reg[0] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold149 (.A(_228_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold150 (.A(_072_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold151 (.A(\ps2_decoder_inst.clk_timeout[2] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold152 (.A(_076_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold153 (.A(\ps2_decoder_inst.clk_timeout[6] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold154 (.A(_080_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold155 (.A(uio_out[5]),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold156 (.A(uio_out[6]),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold157 (.A(uio_out[7]),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold158 (.A(uio_out[3]),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold159 (.A(\ps2_decoder_inst.clk_timeout[10] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold160 (.A(_084_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold161 (.A(\ps2_decoder_inst.clk_timeout[9] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold162 (.A(_083_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold163 (.A(\ps2_decoder_inst.clk_timeout[1] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold164 (.A(_075_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold165 (.A(uio_out[4]),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold166 (.A(\ps2_clk_debounce.debounced_button ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold167 (.A(_087_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold168 (.A(\ps2_decoder_inst.clk_timeout[5] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold169 (.A(_079_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold170 (.A(\memory.wr_ptr[1] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold171 (.A(_042_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold172 (.A(uio_out[0]),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold173 (.A(\ps2_decoder_inst.valid_reg ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold174 (.A(_086_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold175 (.A(uio_out[2]),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold176 (.A(\ps2_decoder_inst.shift_reset ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold177 (.A(_295_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold178 (.A(_097_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold179 (.A(\ps2_decoder_inst.clk_timeout[0] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold180 (.A(\memory.rd_ptr[1] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold181 (.A(uio_out[1]),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold182 (.A(\ps2_decoder_inst.ps2_value[2] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold183 (.A(\ps2_decoder_inst.clk_timeout[8] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold184 (.A(_003_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold185 (.A(_232_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold186 (.A(\ps2_decoder_inst.ps2_value[1] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold187 (.A(_089_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold188 (.A(\ps2_decoder_inst.ps2_value[6] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold189 (.A(_094_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold190 (.A(\ps2_decoder_inst.ps2_value[5] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold191 (.A(\memory.count[1] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold192 (.A(\ps2_decoder_inst.ps2_value[0] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold193 (.A(_088_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold194 (.A(\ps2_decoder_inst.ps2_value[7] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold195 (.A(_095_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold196 (.A(\ps2_decoder_inst.clk_timeout[4] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold197 (.A(\ps2_decoder_inst.ps2_value[3] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold198 (.A(_091_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold199 (.A(\ps2_decoder_inst.ps2_value[4] ),
    .X(net268));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_4 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_316 ();
 sg13g2_decap_8 FILLER_14_323 ();
 sg13g2_decap_8 FILLER_14_330 ();
 sg13g2_fill_2 FILLER_14_337 ();
 sg13g2_decap_4 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_365 ();
 sg13g2_decap_8 FILLER_14_372 ();
 sg13g2_decap_8 FILLER_14_379 ();
 sg13g2_decap_8 FILLER_14_386 ();
 sg13g2_decap_8 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_fill_2 FILLER_15_287 ();
 sg13g2_fill_1 FILLER_15_289 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_4 FILLER_16_245 ();
 sg13g2_fill_2 FILLER_16_249 ();
 sg13g2_fill_1 FILLER_16_277 ();
 sg13g2_fill_1 FILLER_16_292 ();
 sg13g2_fill_2 FILLER_16_316 ();
 sg13g2_fill_2 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_4 FILLER_17_231 ();
 sg13g2_fill_1 FILLER_17_244 ();
 sg13g2_fill_2 FILLER_17_313 ();
 sg13g2_fill_1 FILLER_17_315 ();
 sg13g2_fill_2 FILLER_17_336 ();
 sg13g2_fill_1 FILLER_17_338 ();
 sg13g2_fill_2 FILLER_17_354 ();
 sg13g2_fill_1 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_4 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_129 ();
 sg13g2_decap_8 FILLER_18_136 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_decap_8 FILLER_18_150 ();
 sg13g2_decap_8 FILLER_18_157 ();
 sg13g2_decap_8 FILLER_18_164 ();
 sg13g2_decap_8 FILLER_18_171 ();
 sg13g2_decap_8 FILLER_18_178 ();
 sg13g2_decap_8 FILLER_18_185 ();
 sg13g2_decap_8 FILLER_18_192 ();
 sg13g2_decap_8 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_206 ();
 sg13g2_decap_8 FILLER_18_213 ();
 sg13g2_decap_8 FILLER_18_220 ();
 sg13g2_fill_2 FILLER_18_227 ();
 sg13g2_fill_2 FILLER_18_236 ();
 sg13g2_fill_1 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_257 ();
 sg13g2_fill_2 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_291 ();
 sg13g2_fill_2 FILLER_18_305 ();
 sg13g2_fill_1 FILLER_18_335 ();
 sg13g2_fill_2 FILLER_18_359 ();
 sg13g2_fill_2 FILLER_18_375 ();
 sg13g2_fill_1 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_fill_2 FILLER_19_119 ();
 sg13g2_fill_1 FILLER_19_121 ();
 sg13g2_decap_4 FILLER_19_153 ();
 sg13g2_fill_2 FILLER_19_170 ();
 sg13g2_fill_1 FILLER_19_172 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_fill_2 FILLER_19_207 ();
 sg13g2_decap_4 FILLER_19_214 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_fill_2 FILLER_19_306 ();
 sg13g2_fill_1 FILLER_19_328 ();
 sg13g2_fill_2 FILLER_19_350 ();
 sg13g2_fill_1 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_fill_2 FILLER_20_91 ();
 sg13g2_fill_1 FILLER_20_124 ();
 sg13g2_fill_2 FILLER_20_190 ();
 sg13g2_fill_1 FILLER_20_192 ();
 sg13g2_fill_2 FILLER_20_224 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_fill_1 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_4 FILLER_21_77 ();
 sg13g2_fill_2 FILLER_21_81 ();
 sg13g2_decap_4 FILLER_21_139 ();
 sg13g2_decap_4 FILLER_21_170 ();
 sg13g2_fill_1 FILLER_21_174 ();
 sg13g2_fill_1 FILLER_21_188 ();
 sg13g2_fill_2 FILLER_21_197 ();
 sg13g2_fill_1 FILLER_21_199 ();
 sg13g2_fill_1 FILLER_21_218 ();
 sg13g2_fill_2 FILLER_21_250 ();
 sg13g2_fill_2 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_278 ();
 sg13g2_fill_2 FILLER_21_314 ();
 sg13g2_fill_2 FILLER_21_354 ();
 sg13g2_fill_1 FILLER_21_370 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_4 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_67 ();
 sg13g2_fill_1 FILLER_22_113 ();
 sg13g2_fill_2 FILLER_22_132 ();
 sg13g2_fill_1 FILLER_22_142 ();
 sg13g2_fill_2 FILLER_22_231 ();
 sg13g2_fill_2 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_290 ();
 sg13g2_fill_1 FILLER_22_325 ();
 sg13g2_fill_1 FILLER_22_352 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_4 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_67 ();
 sg13g2_fill_1 FILLER_23_97 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_fill_2 FILLER_23_125 ();
 sg13g2_fill_1 FILLER_23_127 ();
 sg13g2_decap_4 FILLER_23_154 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_fill_1 FILLER_23_258 ();
 sg13g2_fill_2 FILLER_23_312 ();
 sg13g2_fill_1 FILLER_23_314 ();
 sg13g2_fill_2 FILLER_23_346 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_fill_2 FILLER_24_63 ();
 sg13g2_fill_1 FILLER_24_65 ();
 sg13g2_fill_1 FILLER_24_92 ();
 sg13g2_fill_2 FILLER_24_124 ();
 sg13g2_fill_1 FILLER_24_126 ();
 sg13g2_decap_4 FILLER_24_178 ();
 sg13g2_decap_4 FILLER_24_191 ();
 sg13g2_fill_2 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_244 ();
 sg13g2_fill_2 FILLER_24_314 ();
 sg13g2_fill_1 FILLER_24_316 ();
 sg13g2_fill_1 FILLER_24_339 ();
 sg13g2_fill_1 FILLER_24_349 ();
 sg13g2_fill_2 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_110 ();
 sg13g2_fill_1 FILLER_25_112 ();
 sg13g2_decap_4 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_165 ();
 sg13g2_fill_1 FILLER_25_195 ();
 sg13g2_fill_1 FILLER_25_236 ();
 sg13g2_fill_2 FILLER_25_272 ();
 sg13g2_fill_1 FILLER_25_288 ();
 sg13g2_fill_2 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_322 ();
 sg13g2_fill_1 FILLER_25_324 ();
 sg13g2_fill_2 FILLER_25_356 ();
 sg13g2_fill_1 FILLER_25_367 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_4 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_148 ();
 sg13g2_fill_1 FILLER_26_175 ();
 sg13g2_fill_1 FILLER_26_208 ();
 sg13g2_decap_4 FILLER_26_219 ();
 sg13g2_fill_1 FILLER_26_233 ();
 sg13g2_fill_2 FILLER_26_270 ();
 sg13g2_fill_1 FILLER_26_272 ();
 sg13g2_fill_2 FILLER_26_299 ();
 sg13g2_fill_2 FILLER_26_325 ();
 sg13g2_fill_2 FILLER_26_349 ();
 sg13g2_fill_1 FILLER_26_351 ();
 sg13g2_fill_1 FILLER_26_368 ();
 sg13g2_fill_2 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_99 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_fill_2 FILLER_27_152 ();
 sg13g2_fill_2 FILLER_27_187 ();
 sg13g2_fill_1 FILLER_27_189 ();
 sg13g2_fill_1 FILLER_27_257 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_1 FILLER_27_286 ();
 sg13g2_fill_2 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_350 ();
 sg13g2_fill_1 FILLER_27_361 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_4 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_81 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_fill_2 FILLER_28_109 ();
 sg13g2_fill_1 FILLER_28_111 ();
 sg13g2_fill_2 FILLER_28_131 ();
 sg13g2_fill_1 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_216 ();
 sg13g2_fill_1 FILLER_28_284 ();
 sg13g2_fill_2 FILLER_28_327 ();
 sg13g2_fill_1 FILLER_28_338 ();
 sg13g2_fill_2 FILLER_28_359 ();
 sg13g2_fill_2 FILLER_28_381 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_72 ();
 sg13g2_fill_2 FILLER_29_95 ();
 sg13g2_fill_1 FILLER_29_175 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_fill_2 FILLER_29_310 ();
 sg13g2_fill_1 FILLER_29_312 ();
 sg13g2_fill_1 FILLER_29_339 ();
 sg13g2_fill_2 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_4 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_39 ();
 sg13g2_fill_1 FILLER_30_94 ();
 sg13g2_fill_1 FILLER_30_122 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_150 ();
 sg13g2_fill_1 FILLER_30_152 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_fill_2 FILLER_30_191 ();
 sg13g2_fill_2 FILLER_30_197 ();
 sg13g2_decap_4 FILLER_30_225 ();
 sg13g2_fill_1 FILLER_30_242 ();
 sg13g2_fill_2 FILLER_30_274 ();
 sg13g2_fill_1 FILLER_30_276 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_4 FILLER_31_35 ();
 sg13g2_fill_1 FILLER_31_39 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_fill_2 FILLER_31_203 ();
 sg13g2_fill_1 FILLER_31_205 ();
 sg13g2_fill_1 FILLER_31_219 ();
 sg13g2_fill_2 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_fill_2 FILLER_32_35 ();
 sg13g2_fill_1 FILLER_32_37 ();
 sg13g2_fill_1 FILLER_32_73 ();
 sg13g2_fill_1 FILLER_32_147 ();
 sg13g2_fill_1 FILLER_32_161 ();
 sg13g2_fill_2 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_fill_2 FILLER_32_350 ();
 sg13g2_fill_2 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_4 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_46 ();
 sg13g2_fill_2 FILLER_33_89 ();
 sg13g2_fill_1 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_171 ();
 sg13g2_fill_2 FILLER_33_233 ();
 sg13g2_fill_1 FILLER_33_235 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_decap_4 FILLER_33_319 ();
 sg13g2_fill_2 FILLER_33_323 ();
 sg13g2_fill_1 FILLER_33_348 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_4 FILLER_34_42 ();
 sg13g2_fill_2 FILLER_34_46 ();
 sg13g2_fill_2 FILLER_34_91 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_fill_1 FILLER_34_104 ();
 sg13g2_fill_1 FILLER_34_182 ();
 sg13g2_fill_2 FILLER_34_207 ();
 sg13g2_fill_1 FILLER_34_209 ();
 sg13g2_decap_4 FILLER_34_225 ();
 sg13g2_fill_2 FILLER_34_229 ();
 sg13g2_fill_2 FILLER_34_241 ();
 sg13g2_fill_1 FILLER_34_243 ();
 sg13g2_fill_1 FILLER_34_346 ();
 sg13g2_fill_2 FILLER_34_352 ();
 sg13g2_fill_1 FILLER_34_354 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_138 ();
 sg13g2_fill_2 FILLER_35_181 ();
 sg13g2_decap_8 FILLER_35_209 ();
 sg13g2_fill_2 FILLER_35_278 ();
 sg13g2_fill_1 FILLER_35_354 ();
 sg13g2_decap_8 FILLER_35_398 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_4 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_67 ();
 sg13g2_fill_1 FILLER_36_152 ();
 sg13g2_fill_1 FILLER_36_176 ();
 sg13g2_fill_1 FILLER_36_199 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_decap_8 FILLER_36_242 ();
 sg13g2_fill_2 FILLER_36_249 ();
 sg13g2_fill_2 FILLER_36_300 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_fill_1 FILLER_36_366 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_fill_1 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_93 ();
 sg13g2_fill_1 FILLER_37_201 ();
 sg13g2_fill_1 FILLER_37_232 ();
 sg13g2_fill_2 FILLER_37_369 ();
 sg13g2_fill_2 FILLER_37_380 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_fill_1 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_fill_1 FILLER_38_178 ();
 sg13g2_fill_2 FILLER_38_192 ();
 sg13g2_fill_1 FILLER_38_194 ();
 sg13g2_fill_1 FILLER_38_228 ();
 sg13g2_fill_1 FILLER_38_242 ();
 sg13g2_fill_2 FILLER_38_261 ();
 sg13g2_fill_2 FILLER_38_319 ();
 sg13g2_fill_1 FILLER_38_353 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uo_out[3] = net6;
 assign uo_out[4] = net7;
 assign uo_out[5] = net8;
 assign uo_out[6] = net9;
 assign uo_out[7] = net10;
endmodule

module tt_um_sushi_demo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire clknet_0_clk;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire h_sync;
 wire \pix_x[0] ;
 wire \pix_x[1] ;
 wire \pix_x[2] ;
 wire \pix_x[3] ;
 wire \pix_x[4] ;
 wire \pix_x[5] ;
 wire \pix_x[6] ;
 wire \pix_x[7] ;
 wire \pix_x[8] ;
 wire \pix_x[9] ;
 wire \pix_y[0] ;
 wire \pix_y[1] ;
 wire \pix_y[2] ;
 wire \pix_y[3] ;
 wire \pix_y[4] ;
 wire \pix_y[5] ;
 wire \pix_y[6] ;
 wire \pix_y[7] ;
 wire \pix_y[8] ;
 wire \pix_y[9] ;
 wire \sprite_x[0] ;
 wire \sprite_x[1] ;
 wire \sprite_x[2] ;
 wire \sprite_x[3] ;
 wire \sprite_x[4] ;
 wire \sprite_x[5] ;
 wire \sprite_x[6] ;
 wire \sprite_x[7] ;
 wire \sprite_x[8] ;
 wire \sprite_x[9] ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire v_sync;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net1;
 wire net2;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;

 sg13g2_inv_1 _0809_ (.Y(_0727_),
    .A(net93));
 sg13g2_inv_1 _0810_ (.Y(_0728_),
    .A(net63));
 sg13g2_inv_2 _0811_ (.Y(_0729_),
    .A(net255));
 sg13g2_inv_1 _0812_ (.Y(_0730_),
    .A(\pix_x[8] ));
 sg13g2_inv_1 _0813_ (.Y(_0731_),
    .A(\sprite_x[3] ));
 sg13g2_inv_1 _0814_ (.Y(_0732_),
    .A(\sprite_x[7] ));
 sg13g2_inv_1 _0815_ (.Y(_0733_),
    .A(\counter[4] ));
 sg13g2_inv_1 _0816_ (.Y(_0734_),
    .A(\counter[3] ));
 sg13g2_inv_1 _0817_ (.Y(_0055_),
    .A(net61));
 sg13g2_or4_1 _0818_ (.A(_0730_),
    .B(\pix_x[7] ),
    .C(net252),
    .D(net253),
    .X(_0056_));
 sg13g2_and3_1 _0819_ (.X(_0057_),
    .A(\pix_x[1] ),
    .B(net78),
    .C(net68));
 sg13g2_and2_1 _0820_ (.A(net87),
    .B(_0057_),
    .X(_0058_));
 sg13g2_and2_1 _0821_ (.A(net92),
    .B(_0058_),
    .X(_0059_));
 sg13g2_o21ai_1 _0822_ (.B1(\pix_x[9] ),
    .Y(_0060_),
    .A1(_0056_),
    .A2(_0059_));
 sg13g2_a21oi_2 _0823_ (.B1(_0060_),
    .Y(_0061_),
    .A2(_0056_),
    .A1(net103));
 sg13g2_nand2b_1 _0824_ (.Y(_0062_),
    .B(net255),
    .A_N(_0061_));
 sg13g2_nor2_1 _0825_ (.A(_0055_),
    .B(_0062_),
    .Y(_0012_));
 sg13g2_xnor2_1 _0826_ (.Y(_0063_),
    .A(\pix_x[1] ),
    .B(net78));
 sg13g2_nor2_1 _0827_ (.A(net246),
    .B(net79),
    .Y(_0013_));
 sg13g2_a21oi_1 _0828_ (.A1(\pix_x[1] ),
    .A2(\pix_x[0] ),
    .Y(_0064_),
    .B1(net68));
 sg13g2_nor3_1 _0829_ (.A(_0057_),
    .B(net246),
    .C(net69),
    .Y(_0014_));
 sg13g2_nor2_1 _0830_ (.A(net87),
    .B(_0057_),
    .Y(_0065_));
 sg13g2_nor3_1 _0831_ (.A(_0058_),
    .B(net246),
    .C(net88),
    .Y(_0015_));
 sg13g2_nor2_1 _0832_ (.A(net92),
    .B(_0058_),
    .Y(_0066_));
 sg13g2_nor3_1 _0833_ (.A(_0059_),
    .B(net246),
    .C(_0066_),
    .Y(_0016_));
 sg13g2_nor2b_1 _0834_ (.A(net76),
    .B_N(_0058_),
    .Y(_0067_));
 sg13g2_xnor2_1 _0835_ (.Y(_0068_),
    .A(\pix_x[5] ),
    .B(_0067_));
 sg13g2_nor2_1 _0836_ (.A(_0062_),
    .B(net77),
    .Y(_0017_));
 sg13g2_and3_1 _0837_ (.X(_0069_),
    .A(net252),
    .B(net80),
    .C(_0059_));
 sg13g2_a21oi_1 _0838_ (.A1(net80),
    .A2(_0059_),
    .Y(_0070_),
    .B1(net252));
 sg13g2_nor3_1 _0839_ (.A(net246),
    .B(_0069_),
    .C(net81),
    .Y(_0018_));
 sg13g2_nand2_1 _0840_ (.Y(_0071_),
    .A(net95),
    .B(_0069_));
 sg13g2_xnor2_1 _0841_ (.Y(_0072_),
    .A(net251),
    .B(_0069_));
 sg13g2_nor2_1 _0842_ (.A(net246),
    .B(_0072_),
    .Y(_0019_));
 sg13g2_xnor2_1 _0843_ (.Y(_0073_),
    .A(_0730_),
    .B(_0071_));
 sg13g2_nor2_1 _0844_ (.A(net246),
    .B(net96),
    .Y(_0020_));
 sg13g2_nor2_1 _0845_ (.A(net82),
    .B(_0071_),
    .Y(_0074_));
 sg13g2_nor2_1 _0846_ (.A(\pix_x[9] ),
    .B(net83),
    .Y(_0075_));
 sg13g2_nor2_1 _0847_ (.A(net246),
    .B(net84),
    .Y(_0021_));
 sg13g2_nor2_1 _0848_ (.A(net247),
    .B(\pix_y[2] ),
    .Y(_0076_));
 sg13g2_or2_1 _0849_ (.X(_0077_),
    .B(net248),
    .A(net247));
 sg13g2_nor3_1 _0850_ (.A(\pix_y[4] ),
    .B(net247),
    .C(net248),
    .Y(_0078_));
 sg13g2_nor2b_1 _0851_ (.A(_0078_),
    .B_N(\pix_y[5] ),
    .Y(_0079_));
 sg13g2_nand2_1 _0852_ (.Y(_0080_),
    .A(\pix_y[6] ),
    .B(_0079_));
 sg13g2_o21ai_1 _0853_ (.B1(_0007_),
    .Y(_0081_),
    .A1(\pix_y[7] ),
    .A2(_0080_));
 sg13g2_or2_1 _0854_ (.X(_0082_),
    .B(_0081_),
    .A(\pix_y[8] ));
 sg13g2_nand2_2 _0855_ (.Y(_0083_),
    .A(net247),
    .B(net248));
 sg13g2_a21oi_1 _0856_ (.A1(net247),
    .A2(net248),
    .Y(_0084_),
    .B1(_0006_));
 sg13g2_a21oi_2 _0857_ (.B1(_0084_),
    .Y(_0085_),
    .A2(_0077_),
    .A1(_0006_));
 sg13g2_xnor2_1 _0858_ (.Y(_0086_),
    .A(_0005_),
    .B(_0078_));
 sg13g2_nand2b_1 _0859_ (.Y(_0087_),
    .B(_0086_),
    .A_N(_0085_));
 sg13g2_xnor2_1 _0860_ (.Y(_0088_),
    .A(\pix_y[6] ),
    .B(_0079_));
 sg13g2_nand2b_1 _0861_ (.Y(_0089_),
    .B(_0088_),
    .A_N(_0087_));
 sg13g2_xor2_1 _0862_ (.B(_0080_),
    .A(\pix_y[7] ),
    .X(_0090_));
 sg13g2_nand2_1 _0863_ (.Y(_0091_),
    .A(_0089_),
    .B(_0090_));
 sg13g2_xor2_1 _0864_ (.B(_0081_),
    .A(\pix_y[8] ),
    .X(_0092_));
 sg13g2_nand2_1 _0865_ (.Y(_0093_),
    .A(_0091_),
    .B(_0092_));
 sg13g2_xnor2_1 _0866_ (.Y(_0094_),
    .A(_0727_),
    .B(_0082_));
 sg13g2_nand3_1 _0867_ (.B(_0092_),
    .C(_0094_),
    .A(_0091_),
    .Y(_0095_));
 sg13g2_o21ai_1 _0868_ (.B1(_0095_),
    .Y(_0096_),
    .A1(\pix_y[9] ),
    .A2(_0082_));
 sg13g2_nand2_2 _0869_ (.Y(_0097_),
    .A(_0077_),
    .B(_0083_));
 sg13g2_a21oi_2 _0870_ (.B1(_0085_),
    .Y(_0098_),
    .A2(_0083_),
    .A1(_0006_));
 sg13g2_a21o_1 _0871_ (.A2(_0083_),
    .A1(_0006_),
    .B1(_0085_),
    .X(_0099_));
 sg13g2_nand2b_2 _0872_ (.Y(_0100_),
    .B(\pix_x[9] ),
    .A_N(\sprite_x[9] ));
 sg13g2_nor2b_1 _0873_ (.A(\pix_x[9] ),
    .B_N(\sprite_x[9] ),
    .Y(_0101_));
 sg13g2_xor2_1 _0874_ (.B(\sprite_x[9] ),
    .A(\pix_x[9] ),
    .X(_0102_));
 sg13g2_nand2b_1 _0875_ (.Y(_0103_),
    .B(\pix_x[8] ),
    .A_N(\sprite_x[8] ));
 sg13g2_xnor2_1 _0876_ (.Y(_0104_),
    .A(\pix_x[8] ),
    .B(\sprite_x[8] ));
 sg13g2_nor2b_1 _0877_ (.A(\sprite_x[2] ),
    .B_N(\pix_x[2] ),
    .Y(_0105_));
 sg13g2_xnor2_1 _0878_ (.Y(_0106_),
    .A(\pix_x[2] ),
    .B(\sprite_x[2] ));
 sg13g2_nand2b_1 _0879_ (.Y(_0107_),
    .B(\pix_x[1] ),
    .A_N(\sprite_x[1] ));
 sg13g2_nor2b_1 _0880_ (.A(\pix_x[0] ),
    .B_N(\sprite_x[0] ),
    .Y(_0108_));
 sg13g2_nor2b_1 _0881_ (.A(\pix_x[1] ),
    .B_N(\sprite_x[1] ),
    .Y(_0109_));
 sg13g2_o21ai_1 _0882_ (.B1(_0107_),
    .Y(_0110_),
    .A1(_0108_),
    .A2(_0109_));
 sg13g2_a221oi_1 _0883_ (.B2(_0110_),
    .C1(_0105_),
    .B1(_0106_),
    .A1(\pix_x[3] ),
    .Y(_0111_),
    .A2(_0731_));
 sg13g2_nor2_2 _0884_ (.A(\pix_x[3] ),
    .B(_0731_),
    .Y(_0112_));
 sg13g2_nand2_1 _0885_ (.Y(_0113_),
    .A(net251),
    .B(_0732_));
 sg13g2_xor2_1 _0886_ (.B(\sprite_x[7] ),
    .A(net251),
    .X(_0114_));
 sg13g2_nor2b_1 _0887_ (.A(\sprite_x[6] ),
    .B_N(net252),
    .Y(_0115_));
 sg13g2_xor2_1 _0888_ (.B(\sprite_x[6] ),
    .A(net252),
    .X(_0116_));
 sg13g2_nor2_1 _0889_ (.A(_0114_),
    .B(_0116_),
    .Y(_0117_));
 sg13g2_nand2b_2 _0890_ (.Y(_0118_),
    .B(net253),
    .A_N(\sprite_x[5] ));
 sg13g2_nor2b_1 _0891_ (.A(net253),
    .B_N(\sprite_x[5] ),
    .Y(_0119_));
 sg13g2_inv_1 _0892_ (.Y(_0120_),
    .A(_0119_));
 sg13g2_xnor2_1 _0893_ (.Y(_0121_),
    .A(net253),
    .B(\sprite_x[5] ));
 sg13g2_nor2b_1 _0894_ (.A(\sprite_x[4] ),
    .B_N(\pix_x[4] ),
    .Y(_0122_));
 sg13g2_nand2b_1 _0895_ (.Y(_0123_),
    .B(\pix_x[4] ),
    .A_N(\sprite_x[4] ));
 sg13g2_xnor2_1 _0896_ (.Y(_0124_),
    .A(\pix_x[4] ),
    .B(\sprite_x[4] ));
 sg13g2_inv_1 _0897_ (.Y(_0125_),
    .A(_0124_));
 sg13g2_nand3_1 _0898_ (.B(_0121_),
    .C(_0124_),
    .A(_0117_),
    .Y(_0126_));
 sg13g2_nor3_1 _0899_ (.A(_0111_),
    .B(_0112_),
    .C(_0126_),
    .Y(_0127_));
 sg13g2_o21ai_1 _0900_ (.B1(_0118_),
    .Y(_0128_),
    .A1(_0119_),
    .A2(_0123_));
 sg13g2_nand2_1 _0901_ (.Y(_0129_),
    .A(_0117_),
    .B(_0128_));
 sg13g2_o21ai_1 _0902_ (.B1(_0115_),
    .Y(_0130_),
    .A1(net251),
    .A2(_0732_));
 sg13g2_nand3_1 _0903_ (.B(_0129_),
    .C(_0130_),
    .A(_0113_),
    .Y(_0131_));
 sg13g2_nor2_1 _0904_ (.A(_0127_),
    .B(_0131_),
    .Y(_0132_));
 sg13g2_o21ai_1 _0905_ (.B1(_0104_),
    .Y(_0133_),
    .A1(_0127_),
    .A2(_0131_));
 sg13g2_a21o_1 _0906_ (.A2(_0133_),
    .A1(_0103_),
    .B1(_0102_),
    .X(_0134_));
 sg13g2_nand3_1 _0907_ (.B(_0103_),
    .C(_0133_),
    .A(_0102_),
    .Y(_0135_));
 sg13g2_a21oi_2 _0908_ (.B1(_0098_),
    .Y(_0136_),
    .A2(_0135_),
    .A1(_0134_));
 sg13g2_nand2_2 _0909_ (.Y(_0137_),
    .A(_0100_),
    .B(_0134_));
 sg13g2_xor2_1 _0910_ (.B(_0086_),
    .A(_0085_),
    .X(_0138_));
 sg13g2_a21oi_1 _0911_ (.A1(_0100_),
    .A2(_0134_),
    .Y(_0139_),
    .B1(_0138_));
 sg13g2_xnor2_1 _0912_ (.Y(_0140_),
    .A(_0137_),
    .B(_0138_));
 sg13g2_and2_1 _0913_ (.A(_0136_),
    .B(_0140_),
    .X(_0141_));
 sg13g2_xnor2_1 _0914_ (.Y(_0142_),
    .A(_0136_),
    .B(_0140_));
 sg13g2_nor2_1 _0915_ (.A(_0096_),
    .B(_0142_),
    .Y(_0143_));
 sg13g2_xor2_1 _0916_ (.B(_0142_),
    .A(_0096_),
    .X(_0144_));
 sg13g2_and3_1 _0917_ (.X(_0145_),
    .A(_0098_),
    .B(_0134_),
    .C(_0135_));
 sg13g2_xnor2_1 _0918_ (.Y(_0146_),
    .A(_0104_),
    .B(_0132_));
 sg13g2_nor3_1 _0919_ (.A(_0136_),
    .B(_0145_),
    .C(_0146_),
    .Y(_0147_));
 sg13g2_or3_1 _0920_ (.A(_0136_),
    .B(_0145_),
    .C(_0146_),
    .X(_0148_));
 sg13g2_xnor2_1 _0921_ (.Y(_0149_),
    .A(_0093_),
    .B(_0094_));
 sg13g2_o21ai_1 _0922_ (.B1(_0146_),
    .Y(_0150_),
    .A1(_0136_),
    .A2(_0145_));
 sg13g2_nand3_1 _0923_ (.B(_0149_),
    .C(_0150_),
    .A(_0148_),
    .Y(_0151_));
 sg13g2_a21oi_1 _0924_ (.A1(_0149_),
    .A2(_0150_),
    .Y(_0152_),
    .B1(_0147_));
 sg13g2_nand2b_1 _0925_ (.Y(_0153_),
    .B(_0144_),
    .A_N(_0152_));
 sg13g2_xor2_1 _0926_ (.B(_0152_),
    .A(_0144_),
    .X(_0154_));
 sg13g2_xnor2_1 _0927_ (.Y(_0155_),
    .A(_0089_),
    .B(_0090_));
 sg13g2_nor3_2 _0928_ (.A(_0111_),
    .B(_0112_),
    .C(_0125_),
    .Y(_0156_));
 sg13g2_nor2_1 _0929_ (.A(_0122_),
    .B(_0156_),
    .Y(_0157_));
 sg13g2_o21ai_1 _0930_ (.B1(_0120_),
    .Y(_0158_),
    .A1(_0122_),
    .A2(_0156_));
 sg13g2_a21oi_1 _0931_ (.A1(_0118_),
    .A2(_0158_),
    .Y(_0159_),
    .B1(_0116_));
 sg13g2_a21o_1 _0932_ (.A2(_0158_),
    .A1(_0118_),
    .B1(_0116_),
    .X(_0160_));
 sg13g2_or3_1 _0933_ (.A(_0114_),
    .B(_0115_),
    .C(_0159_),
    .X(_0161_));
 sg13g2_o21ai_1 _0934_ (.B1(_0114_),
    .Y(_0162_),
    .A1(_0115_),
    .A2(_0159_));
 sg13g2_nand3_1 _0935_ (.B(_0161_),
    .C(_0162_),
    .A(_0155_),
    .Y(_0163_));
 sg13g2_xnor2_1 _0936_ (.Y(_0164_),
    .A(_0091_),
    .B(_0092_));
 sg13g2_nor2b_1 _0937_ (.A(_0164_),
    .B_N(_0097_),
    .Y(_0165_));
 sg13g2_xnor2_1 _0938_ (.Y(_0166_),
    .A(_0097_),
    .B(_0164_));
 sg13g2_xnor2_1 _0939_ (.Y(_0167_),
    .A(_0146_),
    .B(_0166_));
 sg13g2_or2_1 _0940_ (.X(_0168_),
    .B(_0167_),
    .A(_0163_));
 sg13g2_a21o_1 _0941_ (.A2(_0150_),
    .A1(_0148_),
    .B1(_0149_),
    .X(_0169_));
 sg13g2_a21o_1 _0942_ (.A2(_0166_),
    .A1(_0146_),
    .B1(_0165_),
    .X(_0170_));
 sg13g2_and3_1 _0943_ (.X(_0171_),
    .A(_0151_),
    .B(_0169_),
    .C(_0170_));
 sg13g2_a21oi_1 _0944_ (.A1(_0151_),
    .A2(_0169_),
    .Y(_0172_),
    .B1(_0170_));
 sg13g2_or3_2 _0945_ (.A(_0168_),
    .B(_0171_),
    .C(_0172_),
    .X(_0173_));
 sg13g2_or2_1 _0946_ (.X(_0174_),
    .B(_0173_),
    .A(_0154_));
 sg13g2_xor2_1 _0947_ (.B(_0088_),
    .A(_0087_),
    .X(_0175_));
 sg13g2_nand3_1 _0948_ (.B(_0118_),
    .C(_0158_),
    .A(_0116_),
    .Y(_0176_));
 sg13g2_a21oi_1 _0949_ (.A1(_0160_),
    .A2(_0176_),
    .Y(_0177_),
    .B1(_0175_));
 sg13g2_a21o_1 _0950_ (.A2(_0176_),
    .A1(_0160_),
    .B1(_0175_),
    .X(_0178_));
 sg13g2_a21o_1 _0951_ (.A2(_0162_),
    .A1(_0161_),
    .B1(_0155_),
    .X(_0179_));
 sg13g2_and3_2 _0952_ (.X(_0180_),
    .A(_0163_),
    .B(_0177_),
    .C(_0179_));
 sg13g2_xor2_1 _0953_ (.B(_0167_),
    .A(_0163_),
    .X(_0181_));
 sg13g2_nand2_1 _0954_ (.Y(_0182_),
    .A(_0180_),
    .B(_0181_));
 sg13g2_o21ai_1 _0955_ (.B1(_0168_),
    .Y(_0183_),
    .A1(_0171_),
    .A2(_0172_));
 sg13g2_and4_1 _0956_ (.A(_0173_),
    .B(_0180_),
    .C(_0181_),
    .D(_0183_),
    .X(_0184_));
 sg13g2_xor2_1 _0957_ (.B(_0157_),
    .A(_0121_),
    .X(_0185_));
 sg13g2_nor2b_1 _0958_ (.A(_0138_),
    .B_N(_0185_),
    .Y(_0186_));
 sg13g2_nand3_1 _0959_ (.B(_0175_),
    .C(_0176_),
    .A(_0160_),
    .Y(_0187_));
 sg13g2_and3_1 _0960_ (.X(_0188_),
    .A(_0178_),
    .B(_0186_),
    .C(_0187_));
 sg13g2_nand3_1 _0961_ (.B(_0186_),
    .C(_0187_),
    .A(_0178_),
    .Y(_0189_));
 sg13g2_a21oi_2 _0962_ (.B1(_0177_),
    .Y(_0190_),
    .A2(_0179_),
    .A1(_0163_));
 sg13g2_nor3_1 _0963_ (.A(_0180_),
    .B(_0189_),
    .C(_0190_),
    .Y(_0191_));
 sg13g2_xor2_1 _0964_ (.B(_0181_),
    .A(_0180_),
    .X(_0192_));
 sg13g2_nand2_1 _0965_ (.Y(_0193_),
    .A(_0191_),
    .B(_0192_));
 sg13g2_xnor2_1 _0966_ (.Y(_0194_),
    .A(_0138_),
    .B(_0185_));
 sg13g2_nand2b_1 _0967_ (.Y(_0195_),
    .B(_0111_),
    .A_N(_0112_));
 sg13g2_and2_1 _0968_ (.A(\pix_x[3] ),
    .B(\sprite_x[3] ),
    .X(_0196_));
 sg13g2_a21oi_1 _0969_ (.A1(_0106_),
    .A2(_0110_),
    .Y(_0197_),
    .B1(_0105_));
 sg13g2_nor2_1 _0970_ (.A(\pix_x[3] ),
    .B(\sprite_x[3] ),
    .Y(_0198_));
 sg13g2_or2_1 _0971_ (.X(_0199_),
    .B(_0198_),
    .A(_0197_));
 sg13g2_o21ai_1 _0972_ (.B1(_0195_),
    .Y(_0200_),
    .A1(_0196_),
    .A2(_0199_));
 sg13g2_o21ai_1 _0973_ (.B1(_0125_),
    .Y(_0201_),
    .A1(_0111_),
    .A2(_0112_));
 sg13g2_nor2b_1 _0974_ (.A(_0156_),
    .B_N(_0201_),
    .Y(_0202_));
 sg13g2_nor2_1 _0975_ (.A(_0200_),
    .B(_0202_),
    .Y(_0203_));
 sg13g2_xor2_1 _0976_ (.B(_0202_),
    .A(_0200_),
    .X(_0204_));
 sg13g2_a21oi_2 _0977_ (.B1(_0203_),
    .Y(_0205_),
    .A2(_0204_),
    .A1(_0099_));
 sg13g2_nand2b_1 _0978_ (.Y(_0206_),
    .B(_0194_),
    .A_N(_0205_));
 sg13g2_a21oi_1 _0979_ (.A1(_0178_),
    .A2(_0187_),
    .Y(_0207_),
    .B1(_0186_));
 sg13g2_or3_1 _0980_ (.A(_0188_),
    .B(_0206_),
    .C(_0207_),
    .X(_0208_));
 sg13g2_nor3_1 _0981_ (.A(_0180_),
    .B(_0190_),
    .C(_0208_),
    .Y(_0209_));
 sg13g2_and2_1 _0982_ (.A(_0097_),
    .B(_0200_),
    .X(_0210_));
 sg13g2_xnor2_1 _0983_ (.Y(_0211_),
    .A(_0098_),
    .B(_0204_));
 sg13g2_nand2_1 _0984_ (.Y(_0212_),
    .A(_0210_),
    .B(_0211_));
 sg13g2_xnor2_1 _0985_ (.Y(_0213_),
    .A(_0194_),
    .B(_0205_));
 sg13g2_nor2b_1 _0986_ (.A(_0212_),
    .B_N(_0213_),
    .Y(_0214_));
 sg13g2_o21ai_1 _0987_ (.B1(_0206_),
    .Y(_0215_),
    .A1(_0188_),
    .A2(_0207_));
 sg13g2_and2_2 _0988_ (.A(_0208_),
    .B(_0215_),
    .X(_0216_));
 sg13g2_nand3_1 _0989_ (.B(_0214_),
    .C(_0215_),
    .A(_0208_),
    .Y(_0217_));
 sg13g2_o21ai_1 _0990_ (.B1(_0189_),
    .Y(_0218_),
    .A1(_0206_),
    .A2(_0207_));
 sg13g2_o21ai_1 _0991_ (.B1(_0218_),
    .Y(_0219_),
    .A1(_0180_),
    .A2(_0190_));
 sg13g2_or3_1 _0992_ (.A(_0180_),
    .B(_0190_),
    .C(_0218_),
    .X(_0220_));
 sg13g2_and2_1 _0993_ (.A(_0219_),
    .B(_0220_),
    .X(_0221_));
 sg13g2_a21oi_1 _0994_ (.A1(_0219_),
    .A2(_0220_),
    .Y(_0222_),
    .B1(_0217_));
 sg13g2_nor2_1 _0995_ (.A(_0209_),
    .B(_0222_),
    .Y(_0223_));
 sg13g2_xor2_1 _0996_ (.B(_0192_),
    .A(_0191_),
    .X(_0224_));
 sg13g2_o21ai_1 _0997_ (.B1(_0224_),
    .Y(_0225_),
    .A1(_0209_),
    .A2(_0222_));
 sg13g2_and2_1 _0998_ (.A(_0193_),
    .B(_0225_),
    .X(_0226_));
 sg13g2_nand3_1 _0999_ (.B(_0182_),
    .C(_0183_),
    .A(_0173_),
    .Y(_0227_));
 sg13g2_a21o_1 _1000_ (.A2(_0183_),
    .A1(_0173_),
    .B1(_0182_),
    .X(_0228_));
 sg13g2_and2_1 _1001_ (.A(_0227_),
    .B(_0228_),
    .X(_0229_));
 sg13g2_a22oi_1 _1002_ (.Y(_0230_),
    .B1(_0227_),
    .B2(_0228_),
    .A2(_0225_),
    .A1(_0193_));
 sg13g2_nand2b_1 _1003_ (.Y(_0231_),
    .B(_0171_),
    .A_N(_0154_));
 sg13g2_nand2b_1 _1004_ (.Y(_0232_),
    .B(_0173_),
    .A_N(_0171_));
 sg13g2_xnor2_1 _1005_ (.Y(_0233_),
    .A(_0154_),
    .B(_0232_));
 sg13g2_xor2_1 _1006_ (.B(_0232_),
    .A(_0154_),
    .X(_0234_));
 sg13g2_o21ai_1 _1007_ (.B1(_0233_),
    .Y(_0235_),
    .A1(_0184_),
    .A2(_0230_));
 sg13g2_nand2_1 _1008_ (.Y(_0236_),
    .A(_0174_),
    .B(_0235_));
 sg13g2_nor2_1 _1009_ (.A(_0141_),
    .B(_0143_),
    .Y(_0237_));
 sg13g2_nand2_1 _1010_ (.Y(_0238_),
    .A(_0137_),
    .B(_0175_));
 sg13g2_xnor2_1 _1011_ (.Y(_0239_),
    .A(_0137_),
    .B(_0175_));
 sg13g2_nor2_1 _1012_ (.A(_0139_),
    .B(_0239_),
    .Y(_0240_));
 sg13g2_nand2_1 _1013_ (.Y(_0241_),
    .A(_0139_),
    .B(_0175_));
 sg13g2_o21ai_1 _1014_ (.B1(_0241_),
    .Y(_0242_),
    .A1(_0139_),
    .A2(_0239_));
 sg13g2_nor2_1 _1015_ (.A(_0096_),
    .B(_0240_),
    .Y(_0243_));
 sg13g2_xor2_1 _1016_ (.B(_0242_),
    .A(_0096_),
    .X(_0244_));
 sg13g2_nand2b_1 _1017_ (.Y(_0245_),
    .B(_0244_),
    .A_N(_0237_));
 sg13g2_nor3_1 _1018_ (.A(_0141_),
    .B(_0143_),
    .C(_0244_),
    .Y(_0246_));
 sg13g2_xnor2_1 _1019_ (.Y(_0247_),
    .A(_0237_),
    .B(_0244_));
 sg13g2_nand2_1 _1020_ (.Y(_0248_),
    .A(_0153_),
    .B(_0231_));
 sg13g2_nor2b_1 _1021_ (.A(_0231_),
    .B_N(_0247_),
    .Y(_0249_));
 sg13g2_xnor2_1 _1022_ (.Y(_0250_),
    .A(_0247_),
    .B(_0248_));
 sg13g2_a21oi_1 _1023_ (.A1(_0174_),
    .A2(_0235_),
    .Y(_0251_),
    .B1(_0250_));
 sg13g2_xnor2_1 _1024_ (.Y(_0252_),
    .A(_0236_),
    .B(_0250_));
 sg13g2_xor2_1 _1025_ (.B(_0250_),
    .A(_0236_),
    .X(_0253_));
 sg13g2_o21ai_1 _1026_ (.B1(_0245_),
    .Y(_0254_),
    .A1(_0153_),
    .A2(_0246_));
 sg13g2_a21oi_1 _1027_ (.A1(_0096_),
    .A2(_0241_),
    .Y(_0255_),
    .B1(_0243_));
 sg13g2_xor2_1 _1028_ (.B(_0238_),
    .A(_0155_),
    .X(_0256_));
 sg13g2_xnor2_1 _1029_ (.Y(_0257_),
    .A(_0255_),
    .B(_0256_));
 sg13g2_xnor2_1 _1030_ (.Y(_0258_),
    .A(_0254_),
    .B(_0257_));
 sg13g2_inv_1 _1031_ (.Y(_0259_),
    .A(_0258_));
 sg13g2_o21ai_1 _1032_ (.B1(_0259_),
    .Y(_0260_),
    .A1(_0249_),
    .A2(_0251_));
 sg13g2_or3_2 _1033_ (.A(_0249_),
    .B(_0251_),
    .C(_0259_),
    .X(_0261_));
 sg13g2_nand2_1 _1034_ (.Y(_0262_),
    .A(_0260_),
    .B(_0261_));
 sg13g2_a21oi_2 _1035_ (.B1(_0253_),
    .Y(_0263_),
    .A2(_0261_),
    .A1(_0260_));
 sg13g2_nand2_1 _1036_ (.Y(_0264_),
    .A(_0252_),
    .B(_0262_));
 sg13g2_xor2_1 _1037_ (.B(_0221_),
    .A(_0217_),
    .X(_0265_));
 sg13g2_inv_1 _1038_ (.Y(_0266_),
    .A(_0265_));
 sg13g2_xor2_1 _1039_ (.B(_0224_),
    .A(_0223_),
    .X(_0267_));
 sg13g2_and2_1 _1040_ (.A(_0266_),
    .B(_0267_),
    .X(_0268_));
 sg13g2_or3_2 _1041_ (.A(_0184_),
    .B(_0230_),
    .C(_0233_),
    .X(_0269_));
 sg13g2_or3_1 _1042_ (.A(_0184_),
    .B(_0230_),
    .C(_0234_),
    .X(_0270_));
 sg13g2_o21ai_1 _1043_ (.B1(_0234_),
    .Y(_0271_),
    .A1(_0184_),
    .A2(_0230_));
 sg13g2_xor2_1 _1044_ (.B(_0229_),
    .A(_0226_),
    .X(_0272_));
 sg13g2_xnor2_1 _1045_ (.Y(_0273_),
    .A(_0226_),
    .B(_0229_));
 sg13g2_and4_1 _1046_ (.A(_0268_),
    .B(net226),
    .C(net225),
    .D(_0272_),
    .X(_0274_));
 sg13g2_xor2_1 _1047_ (.B(_0200_),
    .A(_0097_),
    .X(_0275_));
 sg13g2_xnor2_1 _1048_ (.Y(_0276_),
    .A(_0097_),
    .B(_0200_));
 sg13g2_xnor2_1 _1049_ (.Y(_0277_),
    .A(_0210_),
    .B(_0211_));
 sg13g2_nor2_2 _1050_ (.A(_0211_),
    .B(_0276_),
    .Y(_0278_));
 sg13g2_inv_1 _1051_ (.Y(_0279_),
    .A(_0278_));
 sg13g2_and2_1 _1052_ (.A(_0276_),
    .B(net245),
    .X(_0280_));
 sg13g2_nand2_2 _1053_ (.Y(_0281_),
    .A(_0276_),
    .B(net245));
 sg13g2_xnor2_1 _1054_ (.Y(_0282_),
    .A(_0212_),
    .B(_0213_));
 sg13g2_nand2_2 _1055_ (.Y(_0283_),
    .A(_0216_),
    .B(net243));
 sg13g2_nor2_1 _1056_ (.A(_0281_),
    .B(_0283_),
    .Y(_0284_));
 sg13g2_nor2_1 _1057_ (.A(net244),
    .B(_0283_),
    .Y(_0285_));
 sg13g2_a21oi_2 _1058_ (.B1(_0283_),
    .Y(_0286_),
    .A2(_0281_),
    .A1(_0279_));
 sg13g2_nor2b_2 _1059_ (.A(_0216_),
    .B_N(net243),
    .Y(_0287_));
 sg13g2_nand2b_2 _1060_ (.Y(_0288_),
    .B(net243),
    .A_N(_0216_));
 sg13g2_and2_1 _1061_ (.A(_0211_),
    .B(_0275_),
    .X(_0289_));
 sg13g2_nand2_2 _1062_ (.Y(_0290_),
    .A(_0211_),
    .B(_0275_));
 sg13g2_nor2_2 _1063_ (.A(_0280_),
    .B(_0288_),
    .Y(_0291_));
 sg13g2_nand2_1 _1064_ (.Y(_0292_),
    .A(_0281_),
    .B(_0287_));
 sg13g2_nor2_2 _1065_ (.A(_0289_),
    .B(_0292_),
    .Y(_0293_));
 sg13g2_or2_1 _1066_ (.X(_0294_),
    .B(_0293_),
    .A(_0286_));
 sg13g2_and2_1 _1067_ (.A(_0265_),
    .B(_0267_),
    .X(_0295_));
 sg13g2_and4_1 _1068_ (.A(net226),
    .B(net225),
    .C(net224),
    .D(_0295_),
    .X(_0296_));
 sg13g2_nor2_2 _1069_ (.A(net245),
    .B(_0283_),
    .Y(_0297_));
 sg13g2_nor2_1 _1070_ (.A(_0275_),
    .B(net245),
    .Y(_0298_));
 sg13g2_nor2b_2 _1071_ (.A(_0283_),
    .B_N(_0298_),
    .Y(_0299_));
 sg13g2_a22oi_1 _1072_ (.Y(_0300_),
    .B1(net220),
    .B2(_0299_),
    .A2(_0294_),
    .A1(net221));
 sg13g2_nor2_1 _1073_ (.A(_0266_),
    .B(_0267_),
    .Y(_0301_));
 sg13g2_and4_2 _1074_ (.A(net227),
    .B(_0269_),
    .C(_0272_),
    .D(_0301_),
    .X(_0302_));
 sg13g2_xor2_1 _1075_ (.B(_0216_),
    .A(_0214_),
    .X(_0303_));
 sg13g2_nand2b_1 _1076_ (.Y(_0304_),
    .B(_0303_),
    .A_N(net243));
 sg13g2_nor2_1 _1077_ (.A(net244),
    .B(net237),
    .Y(_0305_));
 sg13g2_nor2_2 _1078_ (.A(_0281_),
    .B(net237),
    .Y(_0306_));
 sg13g2_or2_2 _1079_ (.X(_0307_),
    .B(_0304_),
    .A(_0281_));
 sg13g2_a21oi_1 _1080_ (.A1(net244),
    .A2(_0281_),
    .Y(_0308_),
    .B1(net237));
 sg13g2_nand2b_1 _1081_ (.Y(_0309_),
    .B(_0288_),
    .A_N(_0308_));
 sg13g2_and4_2 _1082_ (.A(net227),
    .B(_0269_),
    .C(_0272_),
    .D(_0295_),
    .X(_0310_));
 sg13g2_nor2_2 _1083_ (.A(net243),
    .B(_0303_),
    .Y(_0311_));
 sg13g2_and2_1 _1084_ (.A(_0298_),
    .B(_0311_),
    .X(_0312_));
 sg13g2_nand2_2 _1085_ (.Y(_0313_),
    .A(_0292_),
    .B(_0307_));
 sg13g2_or3_1 _1086_ (.A(_0291_),
    .B(_0308_),
    .C(net231),
    .X(_0314_));
 sg13g2_a22oi_1 _1087_ (.Y(_0315_),
    .B1(_0310_),
    .B2(_0314_),
    .A2(_0309_),
    .A1(_0302_));
 sg13g2_nor3_2 _1088_ (.A(_0281_),
    .B(_0282_),
    .C(_0303_),
    .Y(_0316_));
 sg13g2_nand2_1 _1089_ (.Y(_0317_),
    .A(_0280_),
    .B(_0311_));
 sg13g2_and4_1 _1090_ (.A(net226),
    .B(net225),
    .C(_0272_),
    .D(_0301_),
    .X(_0318_));
 sg13g2_nor2_1 _1091_ (.A(_0265_),
    .B(_0267_),
    .Y(_0319_));
 sg13g2_and4_1 _1092_ (.A(net226),
    .B(net225),
    .C(_0272_),
    .D(_0319_),
    .X(_0320_));
 sg13g2_nand2b_1 _1093_ (.Y(_0321_),
    .B(_0307_),
    .A_N(_0286_));
 sg13g2_a22oi_1 _1094_ (.Y(_0322_),
    .B1(net215),
    .B2(_0321_),
    .A2(_0318_),
    .A1(_0316_));
 sg13g2_nor3_2 _1095_ (.A(_0216_),
    .B(net244),
    .C(net243),
    .Y(_0323_));
 sg13g2_or2_2 _1096_ (.X(_0324_),
    .B(_0323_),
    .A(net231));
 sg13g2_nor3_2 _1097_ (.A(_0282_),
    .B(_0290_),
    .C(_0303_),
    .Y(_0325_));
 sg13g2_and2_2 _1098_ (.A(_0277_),
    .B(_0287_),
    .X(_0326_));
 sg13g2_nor2_2 _1099_ (.A(_0281_),
    .B(_0288_),
    .Y(_0327_));
 sg13g2_or2_2 _1100_ (.X(_0328_),
    .B(_0327_),
    .A(net235));
 sg13g2_o21ai_1 _1101_ (.B1(net219),
    .Y(_0329_),
    .A1(_0324_),
    .A2(_0328_));
 sg13g2_and4_1 _1102_ (.A(net227),
    .B(_0268_),
    .C(_0269_),
    .D(net224),
    .X(_0330_));
 sg13g2_and4_1 _1103_ (.A(net226),
    .B(net225),
    .C(net224),
    .D(_0301_),
    .X(_0331_));
 sg13g2_nor2_1 _1104_ (.A(_0290_),
    .B(_0304_),
    .Y(_0332_));
 sg13g2_or2_1 _1105_ (.X(_0333_),
    .B(net229),
    .A(net241));
 sg13g2_a22oi_1 _1106_ (.Y(_0334_),
    .B1(net212),
    .B2(net223),
    .A2(net213),
    .A1(net232));
 sg13g2_nor2_2 _1107_ (.A(_0288_),
    .B(_0290_),
    .Y(_0335_));
 sg13g2_nand2_1 _1108_ (.Y(_0336_),
    .A(_0287_),
    .B(_0289_));
 sg13g2_nand2_2 _1109_ (.Y(_0337_),
    .A(_0307_),
    .B(_0336_));
 sg13g2_nand2_1 _1110_ (.Y(_0338_),
    .A(net220),
    .B(_0313_));
 sg13g2_nand2_2 _1111_ (.Y(_0339_),
    .A(_0302_),
    .B(net235));
 sg13g2_nor2_2 _1112_ (.A(net245),
    .B(net237),
    .Y(_0340_));
 sg13g2_nor3_2 _1113_ (.A(_0275_),
    .B(net245),
    .C(net237),
    .Y(_0341_));
 sg13g2_and2_1 _1114_ (.A(_0265_),
    .B(_0341_),
    .X(_0342_));
 sg13g2_and4_1 _1115_ (.A(net226),
    .B(net225),
    .C(net224),
    .D(_0342_),
    .X(_0343_));
 sg13g2_and4_1 _1116_ (.A(net226),
    .B(net225),
    .C(_0272_),
    .D(_0295_),
    .X(_0344_));
 sg13g2_and4_1 _1117_ (.A(net227),
    .B(_0269_),
    .C(net224),
    .D(_0301_),
    .X(_0345_));
 sg13g2_nand2_1 _1118_ (.Y(_0346_),
    .A(net235),
    .B(net207));
 sg13g2_and4_1 _1119_ (.A(net227),
    .B(_0269_),
    .C(net224),
    .D(_0295_),
    .X(_0347_));
 sg13g2_and4_1 _1120_ (.A(net226),
    .B(net225),
    .C(net224),
    .D(_0319_),
    .X(_0348_));
 sg13g2_nor2_1 _1121_ (.A(_0283_),
    .B(_0290_),
    .Y(_0349_));
 sg13g2_or2_2 _1122_ (.X(_0350_),
    .B(_0323_),
    .A(_0316_));
 sg13g2_nand2_1 _1123_ (.Y(_0351_),
    .A(net211),
    .B(_0350_));
 sg13g2_and4_1 _1124_ (.A(_0268_),
    .B(_0270_),
    .C(_0271_),
    .D(_0273_),
    .X(_0352_));
 sg13g2_nand3_1 _1125_ (.B(_0311_),
    .C(net201),
    .A(_0276_),
    .Y(_0353_));
 sg13g2_a22oi_1 _1126_ (.Y(_0354_),
    .B1(net211),
    .B2(net234),
    .A2(_0316_),
    .A1(net222));
 sg13g2_a22oi_1 _1127_ (.Y(_0355_),
    .B1(net231),
    .B2(net209),
    .A2(net239),
    .A1(net222));
 sg13g2_a22oi_1 _1128_ (.Y(_0356_),
    .B1(net234),
    .B2(net220),
    .A2(net202),
    .A1(_0323_));
 sg13g2_nand3_1 _1129_ (.B(_0353_),
    .C(_0356_),
    .A(_0351_),
    .Y(_0357_));
 sg13g2_nand3b_1 _1130_ (.B(_0311_),
    .C(net202),
    .Y(_0358_),
    .A_N(net245));
 sg13g2_nand3_1 _1131_ (.B(_0355_),
    .C(_0358_),
    .A(_0354_),
    .Y(_0359_));
 sg13g2_nor2_1 _1132_ (.A(_0357_),
    .B(_0359_),
    .Y(_0360_));
 sg13g2_o21ai_1 _1133_ (.B1(_0336_),
    .Y(_0361_),
    .A1(_0279_),
    .A2(net237));
 sg13g2_a22oi_1 _1134_ (.Y(_0362_),
    .B1(net211),
    .B2(_0361_),
    .A2(net232),
    .A1(net220));
 sg13g2_nor2_2 _1135_ (.A(net245),
    .B(_0288_),
    .Y(_0363_));
 sg13g2_and2_1 _1136_ (.A(net242),
    .B(_0298_),
    .X(_0364_));
 sg13g2_o21ai_1 _1137_ (.B1(net209),
    .Y(_0365_),
    .A1(_0350_),
    .A2(_0364_));
 sg13g2_or2_2 _1138_ (.X(_0366_),
    .B(net238),
    .A(net240));
 sg13g2_nand2_1 _1139_ (.Y(_0367_),
    .A(_0286_),
    .B(net203));
 sg13g2_a22oi_1 _1140_ (.Y(_0368_),
    .B1(_0366_),
    .B2(net211),
    .A2(net200),
    .A1(net234));
 sg13g2_nand3_1 _1141_ (.B(_0367_),
    .C(_0368_),
    .A(_0365_),
    .Y(_0369_));
 sg13g2_nand3_1 _1142_ (.B(_0290_),
    .C(net208),
    .A(net242),
    .Y(_0370_));
 sg13g2_a22oi_1 _1143_ (.Y(_0371_),
    .B1(net234),
    .B2(net214),
    .A2(net206),
    .A1(net236));
 sg13g2_nand2_2 _1144_ (.Y(_0372_),
    .A(_0370_),
    .B(_0371_));
 sg13g2_a22oi_1 _1145_ (.Y(_0373_),
    .B1(_0326_),
    .B2(net209),
    .A2(net216),
    .A1(_0297_));
 sg13g2_nand2_1 _1146_ (.Y(_0374_),
    .A(_0337_),
    .B(net206));
 sg13g2_nand2_1 _1147_ (.Y(_0375_),
    .A(_0337_),
    .B(net208));
 sg13g2_nand4_1 _1148_ (.B(_0315_),
    .C(_0322_),
    .A(_0300_),
    .Y(_0376_),
    .D(_0329_));
 sg13g2_a22oi_1 _1149_ (.Y(_0377_),
    .B1(net204),
    .B2(net239),
    .A2(net217),
    .A1(_0291_));
 sg13g2_a22oi_1 _1150_ (.Y(_0378_),
    .B1(_0323_),
    .B2(net221),
    .A2(net219),
    .A1(_0286_));
 sg13g2_a22oi_1 _1151_ (.Y(_0379_),
    .B1(net207),
    .B2(_0316_),
    .A2(_0324_),
    .A1(net217));
 sg13g2_nand4_1 _1152_ (.B(_0377_),
    .C(_0378_),
    .A(_0334_),
    .Y(_0380_),
    .D(_0379_));
 sg13g2_a221oi_1 _1153_ (.B2(net208),
    .C1(_0343_),
    .B1(net236),
    .A1(net219),
    .Y(_0381_),
    .A2(_0313_));
 sg13g2_a22oi_1 _1154_ (.Y(_0382_),
    .B1(net206),
    .B2(_0293_),
    .A2(net209),
    .A1(net228));
 sg13g2_a22oi_1 _1155_ (.Y(_0383_),
    .B1(net206),
    .B2(_0312_),
    .A2(net230),
    .A1(net220));
 sg13g2_nand4_1 _1156_ (.B(_0381_),
    .C(_0382_),
    .A(_0339_),
    .Y(_0384_),
    .D(_0383_));
 sg13g2_nor4_2 _1157_ (.A(_0369_),
    .B(_0376_),
    .C(_0380_),
    .Y(_0385_),
    .D(_0384_));
 sg13g2_nand4_1 _1158_ (.B(_0373_),
    .C(_0374_),
    .A(_0362_),
    .Y(_0386_),
    .D(_0375_));
 sg13g2_nor4_1 _1159_ (.A(_0357_),
    .B(_0359_),
    .C(_0372_),
    .D(_0386_),
    .Y(_0387_));
 sg13g2_a21oi_2 _1160_ (.B1(_0264_),
    .Y(_0388_),
    .A2(_0387_),
    .A1(_0385_));
 sg13g2_nor2_2 _1161_ (.A(_0252_),
    .B(_0262_),
    .Y(_0389_));
 sg13g2_nand2_1 _1162_ (.Y(_0390_),
    .A(_0306_),
    .B(net212));
 sg13g2_nand3_1 _1163_ (.B(_0362_),
    .C(_0390_),
    .A(_0338_),
    .Y(_0391_));
 sg13g2_nand4_1 _1164_ (.B(_0260_),
    .C(_0261_),
    .A(_0253_),
    .Y(_0392_),
    .D(_0391_));
 sg13g2_a21oi_1 _1165_ (.A1(_0260_),
    .A2(_0261_),
    .Y(_0393_),
    .B1(_0252_));
 sg13g2_inv_1 _1166_ (.Y(_0394_),
    .A(net197));
 sg13g2_o21ai_1 _1167_ (.B1(_0310_),
    .Y(_0395_),
    .A1(net240),
    .A2(net239));
 sg13g2_nand2_1 _1168_ (.Y(_0396_),
    .A(_0302_),
    .B(_0366_));
 sg13g2_and4_2 _1169_ (.A(net227),
    .B(_0269_),
    .C(_0272_),
    .D(_0319_),
    .X(_0397_));
 sg13g2_o21ai_1 _1170_ (.B1(_0397_),
    .Y(_0398_),
    .A1(_0316_),
    .A2(net233));
 sg13g2_nand3_1 _1171_ (.B(_0396_),
    .C(_0398_),
    .A(_0395_),
    .Y(_0399_));
 sg13g2_nand2_1 _1172_ (.Y(_0400_),
    .A(_0302_),
    .B(net228));
 sg13g2_nor3_1 _1173_ (.A(net241),
    .B(net233),
    .C(_0350_),
    .Y(_0401_));
 sg13g2_nand2b_1 _1174_ (.Y(_0402_),
    .B(_0302_),
    .A_N(_0401_));
 sg13g2_nand2_1 _1175_ (.Y(_0403_),
    .A(_0310_),
    .B(net228));
 sg13g2_nand3_1 _1176_ (.B(_0402_),
    .C(_0403_),
    .A(_0400_),
    .Y(_0404_));
 sg13g2_or2_1 _1177_ (.X(_0405_),
    .B(net229),
    .A(net231));
 sg13g2_or2_1 _1178_ (.X(_0406_),
    .B(net223),
    .A(_0328_));
 sg13g2_a22oi_1 _1179_ (.Y(_0407_),
    .B1(_0406_),
    .B2(_0310_),
    .A2(_0405_),
    .A1(_0302_));
 sg13g2_nand2_1 _1180_ (.Y(_0408_),
    .A(_0315_),
    .B(_0407_));
 sg13g2_nor3_2 _1181_ (.A(_0399_),
    .B(_0404_),
    .C(_0408_),
    .Y(_0409_));
 sg13g2_o21ai_1 _1182_ (.B1(_0392_),
    .Y(_0410_),
    .A1(_0394_),
    .A2(_0409_));
 sg13g2_o21ai_1 _1183_ (.B1(net205),
    .Y(_0411_),
    .A1(net228),
    .A2(_0350_));
 sg13g2_and4_2 _1184_ (.A(net227),
    .B(_0269_),
    .C(net224),
    .D(_0319_),
    .X(_0412_));
 sg13g2_a22oi_1 _1185_ (.Y(_0413_),
    .B1(net233),
    .B2(net198),
    .A2(net214),
    .A1(net240));
 sg13g2_nand2_2 _1186_ (.Y(_0414_),
    .A(_0411_),
    .B(_0413_));
 sg13g2_and2_1 _1187_ (.A(_0366_),
    .B(_0412_),
    .X(_0415_));
 sg13g2_o21ai_1 _1188_ (.B1(_0317_),
    .Y(_0416_),
    .A1(net244),
    .A2(net243));
 sg13g2_nor4_1 _1189_ (.A(_0333_),
    .B(_0337_),
    .C(_0341_),
    .D(_0416_),
    .Y(_0417_));
 sg13g2_nor2b_1 _1190_ (.A(_0417_),
    .B_N(net208),
    .Y(_0418_));
 sg13g2_nor4_2 _1191_ (.A(_0372_),
    .B(_0414_),
    .C(_0415_),
    .Y(_0419_),
    .D(_0418_));
 sg13g2_nor2_1 _1192_ (.A(_0394_),
    .B(_0419_),
    .Y(_0420_));
 sg13g2_a22oi_1 _1193_ (.Y(_0421_),
    .B1(_0350_),
    .B2(_0310_),
    .A2(net207),
    .A1(net231));
 sg13g2_and4_2 _1194_ (.A(net227),
    .B(_0268_),
    .C(_0269_),
    .D(_0272_),
    .X(_0422_));
 sg13g2_a22oi_1 _1195_ (.Y(_0423_),
    .B1(_0422_),
    .B2(net239),
    .A2(net207),
    .A1(net240));
 sg13g2_nand3_1 _1196_ (.B(_0421_),
    .C(_0423_),
    .A(_0346_),
    .Y(_0424_));
 sg13g2_nand2_1 _1197_ (.Y(_0425_),
    .A(net197),
    .B(_0424_));
 sg13g2_o21ai_1 _1198_ (.B1(net218),
    .Y(_0426_),
    .A1(_0306_),
    .A2(_0416_));
 sg13g2_a22oi_1 _1199_ (.Y(_0427_),
    .B1(_0335_),
    .B2(_0344_),
    .A2(_0286_),
    .A1(net222));
 sg13g2_nand2_1 _1200_ (.Y(_0428_),
    .A(_0426_),
    .B(_0427_));
 sg13g2_a22oi_1 _1201_ (.Y(_0429_),
    .B1(net214),
    .B2(_0299_),
    .A2(net216),
    .A1(_0286_));
 sg13g2_nand2_1 _1202_ (.Y(_0430_),
    .A(_0284_),
    .B(net203));
 sg13g2_nand2_1 _1203_ (.Y(_0431_),
    .A(_0429_),
    .B(_0430_));
 sg13g2_o21ai_1 _1204_ (.B1(net197),
    .Y(_0432_),
    .A1(_0428_),
    .A2(_0431_));
 sg13g2_a22oi_1 _1205_ (.Y(_0433_),
    .B1(net206),
    .B2(_0312_),
    .A2(net216),
    .A1(net239));
 sg13g2_nand2b_1 _1206_ (.Y(_0434_),
    .B(net197),
    .A_N(_0433_));
 sg13g2_nand4_1 _1207_ (.B(_0425_),
    .C(_0432_),
    .A(_0733_),
    .Y(_0435_),
    .D(_0434_));
 sg13g2_nor4_2 _1208_ (.A(_0388_),
    .B(_0410_),
    .C(_0420_),
    .Y(_0436_),
    .D(_0435_));
 sg13g2_nand2_1 _1209_ (.Y(_0437_),
    .A(net242),
    .B(net206));
 sg13g2_nand3_1 _1210_ (.B(net206),
    .C(net196),
    .A(net242),
    .Y(_0438_));
 sg13g2_or2_2 _1211_ (.X(_0439_),
    .B(net228),
    .A(net232));
 sg13g2_a21oi_2 _1212_ (.B1(net237),
    .Y(_0440_),
    .A2(net244),
    .A1(_0275_));
 sg13g2_o21ai_1 _1213_ (.B1(net221),
    .Y(_0441_),
    .A1(_0306_),
    .A2(_0363_));
 sg13g2_a22oi_1 _1214_ (.Y(_0442_),
    .B1(net205),
    .B2(_0299_),
    .A2(net210),
    .A1(net223));
 sg13g2_a22oi_1 _1215_ (.Y(_0443_),
    .B1(_0440_),
    .B2(net215),
    .A2(net233),
    .A1(net217));
 sg13g2_nand3_1 _1216_ (.B(_0442_),
    .C(_0443_),
    .A(_0441_),
    .Y(_0444_));
 sg13g2_nand2_1 _1217_ (.Y(_0445_),
    .A(net195),
    .B(_0444_));
 sg13g2_o21ai_1 _1218_ (.B1(net195),
    .Y(_0446_),
    .A1(_0424_),
    .A2(_0444_));
 sg13g2_nand4_1 _1219_ (.B(_0434_),
    .C(_0438_),
    .A(\counter[4] ),
    .Y(_0447_),
    .D(_0446_));
 sg13g2_a22oi_1 _1220_ (.Y(_0448_),
    .B1(net205),
    .B2(_0308_),
    .A2(net217),
    .A1(_0291_));
 sg13g2_a22oi_1 _1221_ (.Y(_0449_),
    .B1(net198),
    .B2(net241),
    .A2(net235),
    .A1(net218));
 sg13g2_nor2_1 _1222_ (.A(_0276_),
    .B(net237),
    .Y(_0450_));
 sg13g2_a22oi_1 _1223_ (.Y(_0451_),
    .B1(net208),
    .B2(net233),
    .A2(net229),
    .A1(net213));
 sg13g2_a22oi_1 _1224_ (.Y(_0452_),
    .B1(net229),
    .B2(net215),
    .A2(net213),
    .A1(net241));
 sg13g2_nand4_1 _1225_ (.B(_0449_),
    .C(_0451_),
    .A(_0448_),
    .Y(_0453_),
    .D(_0452_));
 sg13g2_nand2_1 _1226_ (.Y(_0454_),
    .A(net195),
    .B(_0453_));
 sg13g2_o21ai_1 _1227_ (.B1(_0454_),
    .Y(_0455_),
    .A1(_0394_),
    .A2(_0419_));
 sg13g2_nor4_2 _1228_ (.A(_0388_),
    .B(_0410_),
    .C(_0447_),
    .Y(_0456_),
    .D(_0455_));
 sg13g2_nand2_1 _1229_ (.Y(_0457_),
    .A(\sprite_x[3] ),
    .B(\sprite_x[4] ));
 sg13g2_nand4_1 _1230_ (.B(\sprite_x[4] ),
    .C(\sprite_x[5] ),
    .A(\sprite_x[3] ),
    .Y(_0458_),
    .D(\sprite_x[6] ));
 sg13g2_nor2_1 _1231_ (.A(_0002_),
    .B(_0458_),
    .Y(_0459_));
 sg13g2_xnor2_1 _1232_ (.Y(_0460_),
    .A(\sprite_x[8] ),
    .B(_0459_));
 sg13g2_nor2_1 _1233_ (.A(_0730_),
    .B(_0460_),
    .Y(_0461_));
 sg13g2_xnor2_1 _1234_ (.Y(_0462_),
    .A(_0002_),
    .B(_0458_));
 sg13g2_nand2_1 _1235_ (.Y(_0463_),
    .A(net251),
    .B(_0462_));
 sg13g2_nor2_1 _1236_ (.A(_0003_),
    .B(_0457_),
    .Y(_0464_));
 sg13g2_xnor2_1 _1237_ (.Y(_0465_),
    .A(\sprite_x[6] ),
    .B(_0464_));
 sg13g2_nor2_1 _1238_ (.A(net252),
    .B(_0465_),
    .Y(_0466_));
 sg13g2_xor2_1 _1239_ (.B(\sprite_x[4] ),
    .A(\sprite_x[3] ),
    .X(_0467_));
 sg13g2_nor2b_1 _1240_ (.A(_0196_),
    .B_N(_0199_),
    .Y(_0468_));
 sg13g2_o21ai_1 _1241_ (.B1(_0468_),
    .Y(_0469_),
    .A1(_0004_),
    .A2(_0467_));
 sg13g2_xnor2_1 _1242_ (.Y(_0470_),
    .A(_0003_),
    .B(_0457_));
 sg13g2_o21ai_1 _1243_ (.B1(_0469_),
    .Y(_0471_),
    .A1(net253),
    .A2(_0470_));
 sg13g2_a21oi_1 _1244_ (.A1(_0004_),
    .A2(_0467_),
    .Y(_0472_),
    .B1(_0471_));
 sg13g2_a221oi_1 _1245_ (.B2(net253),
    .C1(_0472_),
    .B1(_0470_),
    .A1(net252),
    .Y(_0473_),
    .A2(_0465_));
 sg13g2_o21ai_1 _1246_ (.B1(_0463_),
    .Y(_0474_),
    .A1(_0466_),
    .A2(_0473_));
 sg13g2_nor2_1 _1247_ (.A(net251),
    .B(_0462_),
    .Y(_0475_));
 sg13g2_xnor2_1 _1248_ (.Y(_0476_),
    .A(_0000_),
    .B(_0460_));
 sg13g2_nor2_1 _1249_ (.A(_0475_),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_a21oi_1 _1250_ (.A1(_0474_),
    .A2(_0477_),
    .Y(_0478_),
    .B1(_0461_));
 sg13g2_nand2b_1 _1251_ (.Y(_0479_),
    .B(\sprite_x[7] ),
    .A_N(\sprite_x[8] ));
 sg13g2_o21ai_1 _1252_ (.B1(_0001_),
    .Y(_0480_),
    .A1(_0458_),
    .A2(_0479_));
 sg13g2_o21ai_1 _1253_ (.B1(_0100_),
    .Y(_0481_),
    .A1(_0101_),
    .A2(_0480_));
 sg13g2_nand2b_1 _1254_ (.Y(_0482_),
    .B(_0481_),
    .A_N(_0478_));
 sg13g2_nor2b_1 _1255_ (.A(\pix_y[4] ),
    .B_N(net71),
    .Y(_0483_));
 sg13g2_nor3_1 _1256_ (.A(\pix_y[3] ),
    .B(\pix_y[1] ),
    .C(\pix_y[0] ),
    .Y(_0484_));
 sg13g2_nand2_1 _1257_ (.Y(_0485_),
    .A(_0483_),
    .B(_0484_));
 sg13g2_a22oi_1 _1258_ (.Y(_0486_),
    .B1(_0485_),
    .B2(_0005_),
    .A2(_0483_),
    .A1(_0076_));
 sg13g2_a21oi_1 _1259_ (.A1(\pix_y[6] ),
    .A2(_0486_),
    .Y(_0487_),
    .B1(\pix_y[7] ));
 sg13g2_o21ai_1 _1260_ (.B1(\pix_x[9] ),
    .Y(_0488_),
    .A1(\pix_x[8] ),
    .A2(net251));
 sg13g2_nor2_1 _1261_ (.A(net93),
    .B(_0729_),
    .Y(_0489_));
 sg13g2_nand3b_1 _1262_ (.B(_0488_),
    .C(_0489_),
    .Y(_0490_),
    .A_N(\pix_y[8] ));
 sg13g2_and2_1 _1263_ (.A(\pix_y[7] ),
    .B(\pix_y[6] ),
    .X(_0491_));
 sg13g2_and4_1 _1264_ (.A(net71),
    .B(net85),
    .C(net247),
    .D(net248),
    .X(_0492_));
 sg13g2_nand2_1 _1265_ (.Y(_0493_),
    .A(_0491_),
    .B(_0492_));
 sg13g2_o21ai_1 _1266_ (.B1(_0493_),
    .Y(_0494_),
    .A1(_0100_),
    .A2(_0480_));
 sg13g2_nor3_1 _1267_ (.A(_0487_),
    .B(_0490_),
    .C(_0494_),
    .Y(_0495_));
 sg13g2_nand3_1 _1268_ (.B(_0482_),
    .C(_0495_),
    .A(_0137_),
    .Y(_0496_));
 sg13g2_nor3_1 _1269_ (.A(_0436_),
    .B(_0456_),
    .C(_0496_),
    .Y(_0022_));
 sg13g2_nand3_1 _1270_ (.B(_0311_),
    .C(net201),
    .A(_0275_),
    .Y(_0497_));
 sg13g2_o21ai_1 _1271_ (.B1(_0317_),
    .Y(_0498_),
    .A1(net244),
    .A2(_0288_));
 sg13g2_nand2_1 _1272_ (.Y(_0499_),
    .A(net219),
    .B(_0316_));
 sg13g2_nand2_1 _1273_ (.Y(_0500_),
    .A(net202),
    .B(_0498_));
 sg13g2_nand3_1 _1274_ (.B(_0499_),
    .C(_0500_),
    .A(_0497_),
    .Y(_0501_));
 sg13g2_nand2_2 _1275_ (.Y(_0502_),
    .A(_0326_),
    .B(net199));
 sg13g2_nand2_2 _1276_ (.Y(_0503_),
    .A(net241),
    .B(net199));
 sg13g2_nand2_1 _1277_ (.Y(_0504_),
    .A(_0502_),
    .B(_0503_));
 sg13g2_o21ai_1 _1278_ (.B1(_0307_),
    .Y(_0505_),
    .A1(_0278_),
    .A2(_0288_));
 sg13g2_a22oi_1 _1279_ (.Y(_0506_),
    .B1(net202),
    .B2(_0505_),
    .A2(net209),
    .A1(_0326_));
 sg13g2_a22oi_1 _1280_ (.Y(_0507_),
    .B1(net211),
    .B2(net231),
    .A2(_0328_),
    .A1(net222));
 sg13g2_nand2_1 _1281_ (.Y(_0508_),
    .A(_0506_),
    .B(_0507_));
 sg13g2_a22oi_1 _1282_ (.Y(_0509_),
    .B1(net202),
    .B2(net239),
    .A2(net211),
    .A1(_0328_));
 sg13g2_a22oi_1 _1283_ (.Y(_0510_),
    .B1(net199),
    .B2(_0366_),
    .A2(net202),
    .A1(_0340_));
 sg13g2_o21ai_1 _1284_ (.B1(net219),
    .Y(_0511_),
    .A1(_0285_),
    .A2(_0324_));
 sg13g2_nand4_1 _1285_ (.B(_0509_),
    .C(_0510_),
    .A(_0300_),
    .Y(_0512_),
    .D(_0511_));
 sg13g2_nor4_1 _1286_ (.A(_0501_),
    .B(_0504_),
    .C(_0508_),
    .D(_0512_),
    .Y(_0513_));
 sg13g2_a22oi_1 _1287_ (.Y(_0514_),
    .B1(net200),
    .B2(_0364_),
    .A2(net203),
    .A1(_0305_));
 sg13g2_o21ai_1 _1288_ (.B1(net199),
    .Y(_0515_),
    .A1(net232),
    .A2(_0337_));
 sg13g2_and2_1 _1289_ (.A(_0514_),
    .B(_0515_),
    .X(_0516_));
 sg13g2_nor4_1 _1290_ (.A(_0324_),
    .B(net230),
    .C(_0337_),
    .D(_0439_),
    .Y(_0517_));
 sg13g2_nor2b_1 _1291_ (.A(_0517_),
    .B_N(net221),
    .Y(_0518_));
 sg13g2_a221oi_1 _1292_ (.B2(_0340_),
    .C1(_0518_),
    .B1(net199),
    .A1(net236),
    .Y(_0519_),
    .A2(net210));
 sg13g2_nor2b_1 _1293_ (.A(_0369_),
    .B_N(_0519_),
    .Y(_0520_));
 sg13g2_nand4_1 _1294_ (.B(_0513_),
    .C(_0516_),
    .A(_0360_),
    .Y(_0521_),
    .D(_0520_));
 sg13g2_nand2_2 _1295_ (.Y(_0522_),
    .A(net205),
    .B(net233));
 sg13g2_nand2_1 _1296_ (.Y(_0523_),
    .A(_0397_),
    .B(_0439_));
 sg13g2_nor3_1 _1297_ (.A(net242),
    .B(_0306_),
    .C(net223),
    .Y(_0524_));
 sg13g2_nor2b_1 _1298_ (.A(_0524_),
    .B_N(_0397_),
    .Y(_0525_));
 sg13g2_nand2_1 _1299_ (.Y(_0526_),
    .A(_0286_),
    .B(net205));
 sg13g2_o21ai_1 _1300_ (.B1(_0422_),
    .Y(_0527_),
    .A1(net242),
    .A2(_0440_));
 sg13g2_or2_1 _1301_ (.X(_0528_),
    .B(net235),
    .A(net231));
 sg13g2_nand2_1 _1302_ (.Y(_0529_),
    .A(_0422_),
    .B(_0528_));
 sg13g2_a22oi_1 _1303_ (.Y(_0530_),
    .B1(net205),
    .B2(net229),
    .A2(net207),
    .A1(net238));
 sg13g2_a22oi_1 _1304_ (.Y(_0531_),
    .B1(_0412_),
    .B2(_0328_),
    .A2(_0363_),
    .A1(net213));
 sg13g2_a22oi_1 _1305_ (.Y(_0532_),
    .B1(_0422_),
    .B2(_0323_),
    .A2(net198),
    .A1(net231));
 sg13g2_or2_1 _1306_ (.X(_0533_),
    .B(net235),
    .A(_0324_));
 sg13g2_a22oi_1 _1307_ (.Y(_0534_),
    .B1(_0533_),
    .B2(_0397_),
    .A2(_0422_),
    .A1(_0316_));
 sg13g2_nand4_1 _1308_ (.B(_0531_),
    .C(_0532_),
    .A(_0530_),
    .Y(_0535_),
    .D(_0534_));
 sg13g2_nand2_1 _1309_ (.Y(_0536_),
    .A(net241),
    .B(net207));
 sg13g2_o21ai_1 _1310_ (.B1(_0412_),
    .Y(_0537_),
    .A1(_0313_),
    .A2(_0350_));
 sg13g2_nand3_1 _1311_ (.B(_0529_),
    .C(_0537_),
    .A(_0523_),
    .Y(_0538_));
 sg13g2_nand3_1 _1312_ (.B(_0527_),
    .C(_0536_),
    .A(_0526_),
    .Y(_0539_));
 sg13g2_nor4_1 _1313_ (.A(_0399_),
    .B(_0525_),
    .C(_0538_),
    .D(_0539_),
    .Y(_0540_));
 sg13g2_a22oi_1 _1314_ (.Y(_0541_),
    .B1(_0366_),
    .B2(net198),
    .A2(net205),
    .A1(net238));
 sg13g2_nand4_1 _1315_ (.B(_0423_),
    .C(_0522_),
    .A(_0402_),
    .Y(_0542_),
    .D(_0541_));
 sg13g2_nor2_1 _1316_ (.A(_0535_),
    .B(_0542_),
    .Y(_0543_));
 sg13g2_nand3_1 _1317_ (.B(_0540_),
    .C(_0543_),
    .A(_0451_),
    .Y(_0544_));
 sg13g2_a22oi_1 _1318_ (.Y(_0545_),
    .B1(_0544_),
    .B2(_0263_),
    .A2(_0521_),
    .A1(_0389_));
 sg13g2_o21ai_1 _1319_ (.B1(net214),
    .Y(_0546_),
    .A1(net236),
    .A2(_0326_));
 sg13g2_nand2_1 _1320_ (.Y(_0547_),
    .A(_0316_),
    .B(net214));
 sg13g2_nand2_1 _1321_ (.Y(_0548_),
    .A(net222),
    .B(net232));
 sg13g2_o21ai_1 _1322_ (.B1(net216),
    .Y(_0549_),
    .A1(_0327_),
    .A2(_0341_));
 sg13g2_a22oi_1 _1323_ (.Y(_0550_),
    .B1(_0324_),
    .B2(net214),
    .A2(_0318_),
    .A1(_0285_));
 sg13g2_a22oi_1 _1324_ (.Y(_0551_),
    .B1(_0337_),
    .B2(net203),
    .A2(net218),
    .A1(_0297_));
 sg13g2_and4_1 _1325_ (.A(_0546_),
    .B(_0547_),
    .C(_0548_),
    .D(_0551_),
    .X(_0552_));
 sg13g2_nand4_1 _1326_ (.B(_0549_),
    .C(_0550_),
    .A(_0516_),
    .Y(_0553_),
    .D(_0552_));
 sg13g2_and2_1 _1327_ (.A(net195),
    .B(_0525_),
    .X(_0554_));
 sg13g2_o21ai_1 _1328_ (.B1(_0317_),
    .Y(_0555_),
    .A1(_0216_),
    .A2(net244));
 sg13g2_a22oi_1 _1329_ (.Y(_0556_),
    .B1(_0555_),
    .B2(net216),
    .A2(net233),
    .A1(net209));
 sg13g2_nand2_1 _1330_ (.Y(_0557_),
    .A(net215),
    .B(_0363_));
 sg13g2_nand2_1 _1331_ (.Y(_0558_),
    .A(net215),
    .B(_0528_));
 sg13g2_nand3_1 _1332_ (.B(_0557_),
    .C(_0558_),
    .A(_0556_),
    .Y(_0559_));
 sg13g2_or4_1 _1333_ (.A(net238),
    .B(_0327_),
    .C(net228),
    .D(_0450_),
    .X(_0560_));
 sg13g2_nand2_1 _1334_ (.Y(_0561_),
    .A(net210),
    .B(_0366_));
 sg13g2_a22oi_1 _1335_ (.Y(_0562_),
    .B1(_0560_),
    .B2(net215),
    .A2(_0324_),
    .A1(net217));
 sg13g2_nand3_1 _1336_ (.B(net239),
    .C(net215),
    .A(_0275_),
    .Y(_0563_));
 sg13g2_nand4_1 _1337_ (.B(_0561_),
    .C(_0562_),
    .A(_0322_),
    .Y(_0564_),
    .D(_0563_));
 sg13g2_or2_1 _1338_ (.X(_0565_),
    .B(_0564_),
    .A(_0559_));
 sg13g2_a221oi_1 _1339_ (.B2(_0389_),
    .C1(_0554_),
    .B1(_0565_),
    .A1(_0263_),
    .Y(_0566_),
    .A2(_0553_));
 sg13g2_o21ai_1 _1340_ (.B1(net212),
    .Y(_0567_),
    .A1(_0366_),
    .A2(_0439_));
 sg13g2_nand3_1 _1341_ (.B(net242),
    .C(net204),
    .A(_0278_),
    .Y(_0568_));
 sg13g2_o21ai_1 _1342_ (.B1(net221),
    .Y(_0569_),
    .A1(net232),
    .A2(_0326_));
 sg13g2_nand3_1 _1343_ (.B(_0568_),
    .C(_0569_),
    .A(_0567_),
    .Y(_0570_));
 sg13g2_a22oi_1 _1344_ (.Y(_0571_),
    .B1(net198),
    .B2(net229),
    .A2(net228),
    .A1(net213));
 sg13g2_a22oi_1 _1345_ (.Y(_0572_),
    .B1(net213),
    .B2(_0306_),
    .A2(net217),
    .A1(net241));
 sg13g2_nand2_1 _1346_ (.Y(_0573_),
    .A(_0571_),
    .B(_0572_));
 sg13g2_a22oi_1 _1347_ (.Y(_0574_),
    .B1(_0350_),
    .B2(net198),
    .A2(net210),
    .A1(net235));
 sg13g2_nand3_1 _1348_ (.B(_0561_),
    .C(_0574_),
    .A(_0557_),
    .Y(_0575_));
 sg13g2_nand3_1 _1349_ (.B(_0550_),
    .C(_0556_),
    .A(_0506_),
    .Y(_0576_));
 sg13g2_nand2_1 _1350_ (.Y(_0577_),
    .A(_0334_),
    .B(_0532_));
 sg13g2_or4_1 _1351_ (.A(_0570_),
    .B(_0573_),
    .C(_0575_),
    .D(_0577_),
    .X(_0578_));
 sg13g2_o21ai_1 _1352_ (.B1(net195),
    .Y(_0579_),
    .A1(_0576_),
    .A2(_0578_));
 sg13g2_o21ai_1 _1353_ (.B1(_0327_),
    .Y(_0580_),
    .A1(net216),
    .A2(net212));
 sg13g2_nand4_1 _1354_ (.B(_0514_),
    .C(_0531_),
    .A(_0354_),
    .Y(_0581_),
    .D(_0580_));
 sg13g2_nor3_1 _1355_ (.A(_0291_),
    .B(net239),
    .C(net223),
    .Y(_0582_));
 sg13g2_nand2b_1 _1356_ (.Y(_0583_),
    .B(net219),
    .A_N(_0582_));
 sg13g2_o21ai_1 _1357_ (.B1(net198),
    .Y(_0584_),
    .A1(_0291_),
    .A2(_0440_));
 sg13g2_a22oi_1 _1358_ (.Y(_0585_),
    .B1(_0533_),
    .B2(net221),
    .A2(net233),
    .A1(net204));
 sg13g2_nand3_1 _1359_ (.B(_0584_),
    .C(_0585_),
    .A(_0583_),
    .Y(_0586_));
 sg13g2_nand4_1 _1360_ (.B(_0529_),
    .C(_0546_),
    .A(_0502_),
    .Y(_0587_),
    .D(_0558_));
 sg13g2_a22oi_1 _1361_ (.Y(_0588_),
    .B1(_0311_),
    .B2(net202),
    .A2(net219),
    .A1(net240));
 sg13g2_nand3_1 _1362_ (.B(_0390_),
    .C(_0588_),
    .A(_0351_),
    .Y(_0589_));
 sg13g2_or3_1 _1363_ (.A(_0586_),
    .B(_0587_),
    .C(_0589_),
    .X(_0590_));
 sg13g2_o21ai_1 _1364_ (.B1(net196),
    .Y(_0591_),
    .A1(_0581_),
    .A2(_0590_));
 sg13g2_o21ai_1 _1365_ (.B1(net199),
    .Y(_0592_),
    .A1(_0311_),
    .A2(_0337_));
 sg13g2_nand2_1 _1366_ (.Y(_0593_),
    .A(net230),
    .B(_0422_));
 sg13g2_nand4_1 _1367_ (.B(_0527_),
    .C(_0592_),
    .A(_0329_),
    .Y(_0594_),
    .D(_0593_));
 sg13g2_nand2_1 _1368_ (.Y(_0595_),
    .A(net195),
    .B(_0594_));
 sg13g2_o21ai_1 _1369_ (.B1(net199),
    .Y(_0596_),
    .A1(_0297_),
    .A2(net232));
 sg13g2_a22oi_1 _1370_ (.Y(_0597_),
    .B1(_0528_),
    .B2(net212),
    .A2(_0440_),
    .A1(net219));
 sg13g2_nand3_1 _1371_ (.B(_0596_),
    .C(_0597_),
    .A(_0499_),
    .Y(_0598_));
 sg13g2_nand2_1 _1372_ (.Y(_0599_),
    .A(net238),
    .B(net218));
 sg13g2_nand3_1 _1373_ (.B(_0547_),
    .C(_0599_),
    .A(_0522_),
    .Y(_0600_));
 sg13g2_o21ai_1 _1374_ (.B1(net195),
    .Y(_0601_),
    .A1(_0598_),
    .A2(_0600_));
 sg13g2_and3_1 _1375_ (.X(_0602_),
    .A(_0445_),
    .B(_0595_),
    .C(_0601_));
 sg13g2_and4_1 _1376_ (.A(_0566_),
    .B(_0579_),
    .C(_0591_),
    .D(_0602_),
    .X(_0603_));
 sg13g2_a21oi_1 _1377_ (.A1(_0545_),
    .A2(_0603_),
    .Y(_0604_),
    .B1(\counter[4] ));
 sg13g2_and4_1 _1378_ (.A(_0253_),
    .B(_0260_),
    .C(_0261_),
    .D(_0343_),
    .X(_0605_));
 sg13g2_o21ai_1 _1379_ (.B1(net232),
    .Y(_0606_),
    .A1(net209),
    .A2(net206));
 sg13g2_nand3_1 _1380_ (.B(_0403_),
    .C(_0606_),
    .A(_0390_),
    .Y(_0607_));
 sg13g2_nand2_1 _1381_ (.Y(_0608_),
    .A(_0327_),
    .B(net204));
 sg13g2_a22oi_1 _1382_ (.Y(_0609_),
    .B1(net207),
    .B2(_0439_),
    .A2(net217),
    .A1(_0306_));
 sg13g2_nand3_1 _1383_ (.B(_0608_),
    .C(_0609_),
    .A(_0400_),
    .Y(_0610_));
 sg13g2_or3_1 _1384_ (.A(_0501_),
    .B(_0607_),
    .C(_0610_),
    .X(_0611_));
 sg13g2_nand3b_1 _1385_ (.B(_0298_),
    .C(net218),
    .Y(_0612_),
    .A_N(net243));
 sg13g2_nand2_1 _1386_ (.Y(_0613_),
    .A(net240),
    .B(net203));
 sg13g2_nand4_1 _1387_ (.B(_0437_),
    .C(_0612_),
    .A(_0339_),
    .Y(_0614_),
    .D(_0613_));
 sg13g2_a221oi_1 _1388_ (.B2(net196),
    .C1(_0605_),
    .B1(_0614_),
    .A1(_0263_),
    .Y(_0615_),
    .A2(_0611_));
 sg13g2_and2_1 _1389_ (.A(_0339_),
    .B(_0530_),
    .X(_0616_));
 sg13g2_nand4_1 _1390_ (.B(_0522_),
    .C(_0547_),
    .A(_0429_),
    .Y(_0617_),
    .D(_0616_));
 sg13g2_a221oi_1 _1391_ (.B2(net196),
    .C1(_0605_),
    .B1(_0617_),
    .A1(_0263_),
    .Y(_0618_),
    .A2(_0611_));
 sg13g2_a22oi_1 _1392_ (.Y(_0619_),
    .B1(_0618_),
    .B2(_0456_),
    .A2(_0615_),
    .A1(_0436_));
 sg13g2_a22oi_1 _1393_ (.Y(_0620_),
    .B1(_0340_),
    .B2(net200),
    .A2(_0335_),
    .A1(net211));
 sg13g2_o21ai_1 _1394_ (.B1(net203),
    .Y(_0621_),
    .A1(net238),
    .A2(_0340_));
 sg13g2_nand2_1 _1395_ (.Y(_0622_),
    .A(_0306_),
    .B(net209));
 sg13g2_a22oi_1 _1396_ (.Y(_0623_),
    .B1(net200),
    .B2(net240),
    .A2(net212),
    .A1(_0293_));
 sg13g2_nand4_1 _1397_ (.B(_0621_),
    .C(_0622_),
    .A(_0620_),
    .Y(_0624_),
    .D(_0623_));
 sg13g2_nand2_1 _1398_ (.Y(_0625_),
    .A(net196),
    .B(_0624_));
 sg13g2_nand2_1 _1399_ (.Y(_0626_),
    .A(_0367_),
    .B(_0503_));
 sg13g2_o21ai_1 _1400_ (.B1(net195),
    .Y(_0627_),
    .A1(_0598_),
    .A2(_0626_));
 sg13g2_and3_1 _1401_ (.X(_0628_),
    .A(_0595_),
    .B(_0625_),
    .C(_0627_));
 sg13g2_and3_1 _1402_ (.X(_0629_),
    .A(_0566_),
    .B(_0591_),
    .C(_0628_));
 sg13g2_a21oi_1 _1403_ (.A1(_0545_),
    .A2(_0629_),
    .Y(_0630_),
    .B1(_0733_));
 sg13g2_or4_1 _1404_ (.A(_0496_),
    .B(_0604_),
    .C(_0619_),
    .D(_0630_),
    .X(_0023_));
 sg13g2_nand3_1 _1405_ (.B(_0545_),
    .C(_0629_),
    .A(_0456_),
    .Y(_0631_));
 sg13g2_nand3_1 _1406_ (.B(_0545_),
    .C(_0603_),
    .A(_0436_),
    .Y(_0632_));
 sg13g2_a21o_1 _1407_ (.A2(_0632_),
    .A1(_0631_),
    .B1(_0496_),
    .X(_0024_));
 sg13g2_nor2b_1 _1408_ (.A(_0496_),
    .B_N(_0619_),
    .Y(_0025_));
 sg13g2_o21ai_1 _1409_ (.B1(net212),
    .Y(_0633_),
    .A1(_0293_),
    .A2(net223));
 sg13g2_o21ai_1 _1410_ (.B1(net220),
    .Y(_0634_),
    .A1(_0328_),
    .A2(net223));
 sg13g2_nand2_1 _1411_ (.Y(_0635_),
    .A(_0633_),
    .B(_0634_));
 sg13g2_a22oi_1 _1412_ (.Y(_0636_),
    .B1(_0397_),
    .B2(net240),
    .A2(_0327_),
    .A1(net218));
 sg13g2_a22oi_1 _1413_ (.Y(_0637_),
    .B1(_0422_),
    .B2(_0286_),
    .A2(_0340_),
    .A1(net221));
 sg13g2_nand2_1 _1414_ (.Y(_0638_),
    .A(_0636_),
    .B(_0637_));
 sg13g2_nor4_2 _1415_ (.A(_0414_),
    .B(_0559_),
    .C(_0573_),
    .Y(_0639_),
    .D(_0638_));
 sg13g2_o21ai_1 _1416_ (.B1(_0439_),
    .Y(_0640_),
    .A1(net218),
    .A2(net198));
 sg13g2_nand3_1 _1417_ (.B(net242),
    .C(net205),
    .A(_0280_),
    .Y(_0641_));
 sg13g2_nand3_1 _1418_ (.B(_0640_),
    .C(_0641_),
    .A(_0421_),
    .Y(_0642_));
 sg13g2_a22oi_1 _1419_ (.Y(_0643_),
    .B1(net210),
    .B2(net235),
    .A2(net213),
    .A1(net238));
 sg13g2_a22oi_1 _1420_ (.Y(_0644_),
    .B1(_0450_),
    .B2(net215),
    .A2(net213),
    .A1(net241));
 sg13g2_nand4_1 _1421_ (.B(_0449_),
    .C(_0643_),
    .A(_0407_),
    .Y(_0645_),
    .D(_0644_));
 sg13g2_o21ai_1 _1422_ (.B1(net207),
    .Y(_0646_),
    .A1(_0323_),
    .A2(net229));
 sg13g2_o21ai_1 _1423_ (.B1(net210),
    .Y(_0647_),
    .A1(net223),
    .A2(_0337_));
 sg13g2_nand2_1 _1424_ (.Y(_0648_),
    .A(net221),
    .B(_0306_));
 sg13g2_nand3_1 _1425_ (.B(_0647_),
    .C(_0648_),
    .A(_0646_),
    .Y(_0649_));
 sg13g2_nand2_1 _1426_ (.Y(_0650_),
    .A(net217),
    .B(net229));
 sg13g2_nand2_1 _1427_ (.Y(_0651_),
    .A(net238),
    .B(_0397_));
 sg13g2_nand4_1 _1428_ (.B(_0593_),
    .C(_0650_),
    .A(_0561_),
    .Y(_0652_),
    .D(_0651_));
 sg13g2_nor4_2 _1429_ (.A(_0642_),
    .B(_0645_),
    .C(_0649_),
    .Y(_0653_),
    .D(_0652_));
 sg13g2_a21oi_1 _1430_ (.A1(_0639_),
    .A2(_0653_),
    .Y(_0654_),
    .B1(_0264_));
 sg13g2_a21o_1 _1431_ (.A2(_0635_),
    .A1(_0389_),
    .B1(_0654_),
    .X(_0655_));
 sg13g2_nand4_1 _1432_ (.B(_0355_),
    .C(_0365_),
    .A(_0253_),
    .Y(_0656_),
    .D(_0534_));
 sg13g2_nand2_1 _1433_ (.Y(_0657_),
    .A(net210),
    .B(_0439_));
 sg13g2_nand4_1 _1434_ (.B(_0650_),
    .C(_0651_),
    .A(_0526_),
    .Y(_0658_),
    .D(_0657_));
 sg13g2_or3_1 _1435_ (.A(_0638_),
    .B(_0656_),
    .C(_0658_),
    .X(_0659_));
 sg13g2_or2_1 _1436_ (.X(_0660_),
    .B(_0364_),
    .A(net228));
 sg13g2_a22oi_1 _1437_ (.Y(_0661_),
    .B1(_0660_),
    .B2(net202),
    .A2(_0366_),
    .A1(net199));
 sg13g2_nand4_1 _1438_ (.B(_0502_),
    .C(_0503_),
    .A(_0252_),
    .Y(_0662_),
    .D(_0661_));
 sg13g2_and2_1 _1439_ (.A(_0262_),
    .B(_0662_),
    .X(_0663_));
 sg13g2_nand2_1 _1440_ (.Y(_0664_),
    .A(_0647_),
    .B(_0657_));
 sg13g2_o21ai_1 _1441_ (.B1(net211),
    .Y(_0665_),
    .A1(_0293_),
    .A2(_0328_));
 sg13g2_nand2_1 _1442_ (.Y(_0666_),
    .A(net230),
    .B(net203));
 sg13g2_o21ai_1 _1443_ (.B1(net222),
    .Y(_0667_),
    .A1(_0312_),
    .A2(_0335_));
 sg13g2_nand4_1 _1444_ (.B(_0665_),
    .C(_0666_),
    .A(_0507_),
    .Y(_0668_),
    .D(_0667_));
 sg13g2_and2_1 _1445_ (.A(_0263_),
    .B(_0668_),
    .X(_0669_));
 sg13g2_a221oi_1 _1446_ (.B2(_0389_),
    .C1(_0669_),
    .B1(_0664_),
    .A1(_0659_),
    .Y(_0670_),
    .A2(_0663_));
 sg13g2_and2_1 _1447_ (.A(_0599_),
    .B(_0612_),
    .X(_0671_));
 sg13g2_inv_1 _1448_ (.Y(_0672_),
    .A(_0671_));
 sg13g2_o21ai_1 _1449_ (.B1(net196),
    .Y(_0673_),
    .A1(_0428_),
    .A2(_0672_));
 sg13g2_nand4_1 _1450_ (.B(_0618_),
    .C(_0670_),
    .A(_0579_),
    .Y(_0674_),
    .D(_0673_));
 sg13g2_o21ai_1 _1451_ (.B1(_0456_),
    .Y(_0675_),
    .A1(_0655_),
    .A2(_0674_));
 sg13g2_nand2_1 _1452_ (.Y(_0676_),
    .A(_0503_),
    .B(_0530_));
 sg13g2_o21ai_1 _1453_ (.B1(net196),
    .Y(_0677_),
    .A1(_0624_),
    .A2(_0676_));
 sg13g2_nand4_1 _1454_ (.B(_0615_),
    .C(_0670_),
    .A(_0454_),
    .Y(_0678_),
    .D(_0677_));
 sg13g2_o21ai_1 _1455_ (.B1(_0436_),
    .Y(_0679_),
    .A1(_0655_),
    .A2(_0678_));
 sg13g2_a21o_1 _1456_ (.A2(_0679_),
    .A1(_0675_),
    .B1(_0496_),
    .X(_0026_));
 sg13g2_and2_1 _1457_ (.A(net254),
    .B(_0010_),
    .X(_0028_));
 sg13g2_o21ai_1 _1458_ (.B1(net254),
    .Y(_0680_),
    .A1(\sprite_x[0] ),
    .A2(\sprite_x[1] ));
 sg13g2_a21oi_1 _1459_ (.A1(\sprite_x[0] ),
    .A2(\sprite_x[1] ),
    .Y(_0029_),
    .B1(_0680_));
 sg13g2_nand3_1 _1460_ (.B(\sprite_x[1] ),
    .C(\sprite_x[2] ),
    .A(\sprite_x[0] ),
    .Y(_0681_));
 sg13g2_inv_1 _1461_ (.Y(_0682_),
    .A(_0681_));
 sg13g2_a21oi_1 _1462_ (.A1(\sprite_x[0] ),
    .A2(\sprite_x[1] ),
    .Y(_0683_),
    .B1(\sprite_x[2] ));
 sg13g2_o21ai_1 _1463_ (.B1(net254),
    .Y(_0030_),
    .A1(_0682_),
    .A2(_0683_));
 sg13g2_xnor2_1 _1464_ (.Y(_0684_),
    .A(_0731_),
    .B(_0681_));
 sg13g2_nor2_1 _1465_ (.A(_0729_),
    .B(_0684_),
    .Y(_0031_));
 sg13g2_a21oi_1 _1466_ (.A1(\sprite_x[3] ),
    .A2(_0682_),
    .Y(_0685_),
    .B1(\sprite_x[4] ));
 sg13g2_nor2_1 _1467_ (.A(_0457_),
    .B(_0681_),
    .Y(_0686_));
 sg13g2_nor3_1 _1468_ (.A(_0729_),
    .B(_0685_),
    .C(_0686_),
    .Y(_0032_));
 sg13g2_xnor2_1 _1469_ (.Y(_0687_),
    .A(\sprite_x[5] ),
    .B(_0686_));
 sg13g2_nand2_1 _1470_ (.Y(_0033_),
    .A(net254),
    .B(_0687_));
 sg13g2_nor2_1 _1471_ (.A(_0458_),
    .B(_0681_),
    .Y(_0688_));
 sg13g2_a21oi_1 _1472_ (.A1(\sprite_x[5] ),
    .A2(_0686_),
    .Y(_0689_),
    .B1(\sprite_x[6] ));
 sg13g2_o21ai_1 _1473_ (.B1(net254),
    .Y(_0034_),
    .A1(_0688_),
    .A2(_0689_));
 sg13g2_o21ai_1 _1474_ (.B1(_0732_),
    .Y(_0690_),
    .A1(_0458_),
    .A2(_0681_));
 sg13g2_nand2_1 _1475_ (.Y(_0691_),
    .A(\sprite_x[7] ),
    .B(_0688_));
 sg13g2_and3_1 _1476_ (.X(_0035_),
    .A(net255),
    .B(_0690_),
    .C(_0691_));
 sg13g2_xor2_1 _1477_ (.B(_0691_),
    .A(\sprite_x[8] ),
    .X(_0692_));
 sg13g2_nor2_1 _1478_ (.A(_0729_),
    .B(_0692_),
    .Y(_0036_));
 sg13g2_nor2_1 _1479_ (.A(_0001_),
    .B(_0691_),
    .Y(_0693_));
 sg13g2_o21ai_1 _1480_ (.B1(net255),
    .Y(_0694_),
    .A1(\sprite_x[9] ),
    .A2(_0693_));
 sg13g2_a21oi_1 _1481_ (.A1(\sprite_x[9] ),
    .A2(_0693_),
    .Y(_0037_),
    .B1(_0694_));
 sg13g2_and2_1 _1482_ (.A(net254),
    .B(_0009_),
    .X(_0038_));
 sg13g2_o21ai_1 _1483_ (.B1(net1),
    .Y(_0695_),
    .A1(\counter[0] ),
    .A2(\counter[1] ));
 sg13g2_a21oi_1 _1484_ (.A1(\counter[0] ),
    .A2(\counter[1] ),
    .Y(_0039_),
    .B1(_0695_));
 sg13g2_a21oi_1 _1485_ (.A1(\counter[0] ),
    .A2(\counter[1] ),
    .Y(_0696_),
    .B1(\counter[2] ));
 sg13g2_nand3_1 _1486_ (.B(\counter[1] ),
    .C(\counter[2] ),
    .A(\counter[0] ),
    .Y(_0697_));
 sg13g2_nand2_1 _1487_ (.Y(_0698_),
    .A(net254),
    .B(_0697_));
 sg13g2_nor2_1 _1488_ (.A(_0696_),
    .B(_0698_),
    .Y(_0040_));
 sg13g2_and2_1 _1489_ (.A(_0734_),
    .B(_0697_),
    .X(_0699_));
 sg13g2_nor2_1 _1490_ (.A(_0734_),
    .B(_0697_),
    .Y(_0700_));
 sg13g2_nor3_1 _1491_ (.A(_0729_),
    .B(_0699_),
    .C(_0700_),
    .Y(_0041_));
 sg13g2_o21ai_1 _1492_ (.B1(net254),
    .Y(_0701_),
    .A1(\counter[4] ),
    .A2(_0700_));
 sg13g2_a21oi_1 _1493_ (.A1(\counter[4] ),
    .A2(_0700_),
    .Y(_0042_),
    .B1(_0701_));
 sg13g2_nor3_1 _1494_ (.A(net252),
    .B(net253),
    .C(net92),
    .Y(_0702_));
 sg13g2_nand3_1 _1495_ (.B(net253),
    .C(\pix_x[4] ),
    .A(net100),
    .Y(_0703_));
 sg13g2_nand4_1 _1496_ (.B(net251),
    .C(\pix_x[9] ),
    .A(_0730_),
    .Y(_0704_),
    .D(_0703_));
 sg13g2_o21ai_1 _1497_ (.B1(net255),
    .Y(_0043_),
    .A1(_0702_),
    .A2(net101));
 sg13g2_nand3b_1 _1498_ (.B(net65),
    .C(net247),
    .Y(_0705_),
    .A_N(net248));
 sg13g2_nand4_1 _1499_ (.B(net73),
    .C(_0483_),
    .A(_0727_),
    .Y(_0706_),
    .D(_0491_));
 sg13g2_o21ai_1 _1500_ (.B1(net255),
    .Y(_0044_),
    .A1(_0705_),
    .A2(net74));
 sg13g2_nor3_1 _1501_ (.A(\pix_y[6] ),
    .B(\pix_y[5] ),
    .C(\pix_y[4] ),
    .Y(_0707_));
 sg13g2_nand2_1 _1502_ (.Y(_0708_),
    .A(net255),
    .B(_0707_));
 sg13g2_nor3_1 _1503_ (.A(\pix_y[8] ),
    .B(\pix_y[7] ),
    .C(_0708_),
    .Y(_0709_));
 sg13g2_a21oi_2 _1504_ (.B1(_0489_),
    .Y(_0710_),
    .A2(_0709_),
    .A1(_0083_));
 sg13g2_inv_1 _1505_ (.Y(_0711_),
    .A(_0710_));
 sg13g2_o21ai_1 _1506_ (.B1(_0711_),
    .Y(_0712_),
    .A1(\pix_y[0] ),
    .A2(_0061_));
 sg13g2_a21oi_1 _1507_ (.A1(_0728_),
    .A2(_0061_),
    .Y(_0045_),
    .B1(_0712_));
 sg13g2_a21oi_1 _1508_ (.A1(\pix_y[0] ),
    .A2(_0061_),
    .Y(_0713_),
    .B1(net65));
 sg13g2_and3_2 _1509_ (.X(_0714_),
    .A(net65),
    .B(\pix_y[0] ),
    .C(_0061_));
 sg13g2_nor3_1 _1510_ (.A(_0710_),
    .B(net66),
    .C(_0714_),
    .Y(_0046_));
 sg13g2_nor2_1 _1511_ (.A(net248),
    .B(_0714_),
    .Y(_0715_));
 sg13g2_and2_1 _1512_ (.A(net248),
    .B(_0714_),
    .X(_0716_));
 sg13g2_nor3_1 _1513_ (.A(_0710_),
    .B(net99),
    .C(_0716_),
    .Y(_0047_));
 sg13g2_nor2b_1 _1514_ (.A(_0083_),
    .B_N(_0714_),
    .Y(_0717_));
 sg13g2_o21ai_1 _1515_ (.B1(_0711_),
    .Y(_0718_),
    .A1(net247),
    .A2(_0716_));
 sg13g2_nor2_1 _1516_ (.A(_0717_),
    .B(_0718_),
    .Y(_0048_));
 sg13g2_xnor2_1 _1517_ (.Y(_0719_),
    .A(net85),
    .B(_0717_));
 sg13g2_nor2_1 _1518_ (.A(_0710_),
    .B(_0719_),
    .Y(_0049_));
 sg13g2_nor2b_1 _1519_ (.A(_0006_),
    .B_N(_0717_),
    .Y(_0720_));
 sg13g2_o21ai_1 _1520_ (.B1(_0711_),
    .Y(_0721_),
    .A1(net71),
    .A2(_0720_));
 sg13g2_a21oi_1 _1521_ (.A1(net71),
    .A2(_0720_),
    .Y(_0050_),
    .B1(_0721_));
 sg13g2_a21oi_1 _1522_ (.A1(_0492_),
    .A2(_0714_),
    .Y(_0722_),
    .B1(net89));
 sg13g2_and3_1 _1523_ (.X(_0723_),
    .A(\pix_y[6] ),
    .B(_0492_),
    .C(_0714_));
 sg13g2_nor3_1 _1524_ (.A(_0710_),
    .B(net90),
    .C(_0723_),
    .Y(_0051_));
 sg13g2_xnor2_1 _1525_ (.Y(_0724_),
    .A(net97),
    .B(_0723_));
 sg13g2_nor2_1 _1526_ (.A(_0710_),
    .B(_0724_),
    .Y(_0052_));
 sg13g2_a21o_1 _1527_ (.A2(_0723_),
    .A1(net97),
    .B1(net73),
    .X(_0725_));
 sg13g2_nand3_1 _1528_ (.B(\pix_y[7] ),
    .C(_0723_),
    .A(net73),
    .Y(_0726_));
 sg13g2_and3_1 _1529_ (.X(_0053_),
    .A(_0711_),
    .B(_0725_),
    .C(_0726_));
 sg13g2_a21oi_1 _1530_ (.A1(_0727_),
    .A2(_0726_),
    .Y(_0054_),
    .B1(_0710_));
 sg13g2_nor2b_1 _1531_ (.A(_0496_),
    .B_N(_0619_),
    .Y(_0027_));
 sg13g2_dfrbp_1 _1532_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net35),
    .D(net62),
    .Q_N(_0011_),
    .Q(\pix_x[0] ));
 sg13g2_dfrbp_1 _1533_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net29),
    .D(_0013_),
    .Q_N(_0765_),
    .Q(\pix_x[1] ));
 sg13g2_dfrbp_1 _1534_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net28),
    .D(net70),
    .Q_N(_0764_),
    .Q(\pix_x[2] ));
 sg13g2_dfrbp_1 _1535_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net27),
    .D(_0015_),
    .Q_N(_0763_),
    .Q(\pix_x[3] ));
 sg13g2_dfrbp_1 _1536_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net26),
    .D(_0016_),
    .Q_N(_0004_),
    .Q(\pix_x[4] ));
 sg13g2_dfrbp_1 _1537_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net25),
    .D(_0017_),
    .Q_N(_0762_),
    .Q(\pix_x[5] ));
 sg13g2_dfrbp_1 _1538_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net24),
    .D(_0018_),
    .Q_N(_0761_),
    .Q(\pix_x[6] ));
 sg13g2_dfrbp_1 _1539_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net23),
    .D(_0019_),
    .Q_N(_0760_),
    .Q(\pix_x[7] ));
 sg13g2_dfrbp_1 _1540_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net22),
    .D(_0020_),
    .Q_N(_0000_),
    .Q(\pix_x[8] ));
 sg13g2_dfrbp_1 _1541_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net21),
    .D(_0021_),
    .Q_N(_0759_),
    .Q(\pix_x[9] ));
 sg13g2_dfrbp_1 _1542_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net20),
    .D(_0022_),
    .Q_N(_0758_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1543_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net19),
    .D(_0023_),
    .Q_N(_0757_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1544_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net18),
    .D(_0024_),
    .Q_N(_0756_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1545_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net60),
    .D(_0025_),
    .Q_N(_0755_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1546_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net59),
    .D(_0026_),
    .Q_N(_0754_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1547_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net58),
    .D(_0027_),
    .Q_N(_0753_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1548_ (.CLK(net250),
    .RESET_B(net57),
    .D(_0028_),
    .Q_N(_0010_),
    .Q(\sprite_x[0] ));
 sg13g2_dfrbp_1 _1549_ (.CLK(net250),
    .RESET_B(net56),
    .D(_0029_),
    .Q_N(_0752_),
    .Q(\sprite_x[1] ));
 sg13g2_dfrbp_1 _1550_ (.CLK(net250),
    .RESET_B(net55),
    .D(_0030_),
    .Q_N(_0751_),
    .Q(\sprite_x[2] ));
 sg13g2_dfrbp_1 _1551_ (.CLK(net250),
    .RESET_B(net54),
    .D(_0031_),
    .Q_N(_0750_),
    .Q(\sprite_x[3] ));
 sg13g2_dfrbp_1 _1552_ (.CLK(net250),
    .RESET_B(net53),
    .D(_0032_),
    .Q_N(_0749_),
    .Q(\sprite_x[4] ));
 sg13g2_dfrbp_1 _1553_ (.CLK(net249),
    .RESET_B(net52),
    .D(_0033_),
    .Q_N(_0003_),
    .Q(\sprite_x[5] ));
 sg13g2_dfrbp_1 _1554_ (.CLK(net249),
    .RESET_B(net51),
    .D(_0034_),
    .Q_N(_0748_),
    .Q(\sprite_x[6] ));
 sg13g2_dfrbp_1 _1555_ (.CLK(net249),
    .RESET_B(net50),
    .D(_0035_),
    .Q_N(_0002_),
    .Q(\sprite_x[7] ));
 sg13g2_dfrbp_1 _1556_ (.CLK(net249),
    .RESET_B(net49),
    .D(_0036_),
    .Q_N(_0001_),
    .Q(\sprite_x[8] ));
 sg13g2_dfrbp_1 _1557_ (.CLK(net249),
    .RESET_B(net48),
    .D(_0037_),
    .Q_N(_0747_),
    .Q(\sprite_x[9] ));
 sg13g2_dfrbp_1 _1558_ (.CLK(net249),
    .RESET_B(net47),
    .D(_0038_),
    .Q_N(_0009_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _1559_ (.CLK(v_sync),
    .RESET_B(net46),
    .D(_0039_),
    .Q_N(_0746_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _1560_ (.CLK(net250),
    .RESET_B(net45),
    .D(_0040_),
    .Q_N(_0745_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _1561_ (.CLK(net249),
    .RESET_B(net44),
    .D(_0041_),
    .Q_N(_0744_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _1562_ (.CLK(net250),
    .RESET_B(net43),
    .D(_0042_),
    .Q_N(_0743_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _1563_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net42),
    .D(_0043_),
    .Q_N(_0742_),
    .Q(h_sync));
 sg13g2_dfrbp_1 _1564_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net41),
    .D(net75),
    .Q_N(_0741_),
    .Q(v_sync));
 sg13g2_dfrbp_1 _1565_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net40),
    .D(net64),
    .Q_N(_0008_),
    .Q(\pix_y[0] ));
 sg13g2_dfrbp_1 _1566_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net38),
    .D(net67),
    .Q_N(_0740_),
    .Q(\pix_y[1] ));
 sg13g2_dfrbp_1 _1567_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net36),
    .D(_0047_),
    .Q_N(_0739_),
    .Q(\pix_y[2] ));
 sg13g2_dfrbp_1 _1568_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net34),
    .D(_0048_),
    .Q_N(_0738_),
    .Q(\pix_y[3] ));
 sg13g2_dfrbp_1 _1569_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net32),
    .D(net86),
    .Q_N(_0006_),
    .Q(\pix_y[4] ));
 sg13g2_dfrbp_1 _1570_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net30),
    .D(net72),
    .Q_N(_0005_),
    .Q(\pix_y[5] ));
 sg13g2_dfrbp_1 _1571_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net37),
    .D(net91),
    .Q_N(_0737_),
    .Q(\pix_y[6] ));
 sg13g2_dfrbp_1 _1572_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net33),
    .D(_0052_),
    .Q_N(_0007_),
    .Q(\pix_y[7] ));
 sg13g2_dfrbp_1 _1573_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net39),
    .D(_0053_),
    .Q_N(_0736_),
    .Q(\pix_y[8] ));
 sg13g2_dfrbp_1 _1574_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net31),
    .D(net94),
    .Q_N(_0735_),
    .Q(\pix_y[9] ));
 sg13g2_tiehi _1543__19 (.L_HI(net19));
 sg13g2_tiehi _1542__20 (.L_HI(net20));
 sg13g2_tiehi _1541__21 (.L_HI(net21));
 sg13g2_tiehi _1540__22 (.L_HI(net22));
 sg13g2_tiehi _1539__23 (.L_HI(net23));
 sg13g2_tiehi _1538__24 (.L_HI(net24));
 sg13g2_tiehi _1537__25 (.L_HI(net25));
 sg13g2_tiehi _1536__26 (.L_HI(net26));
 sg13g2_tiehi _1535__27 (.L_HI(net27));
 sg13g2_tiehi _1534__28 (.L_HI(net28));
 sg13g2_tiehi _1533__29 (.L_HI(net29));
 sg13g2_tiehi _1570__30 (.L_HI(net30));
 sg13g2_tiehi _1574__31 (.L_HI(net31));
 sg13g2_tiehi _1569__32 (.L_HI(net32));
 sg13g2_tiehi _1572__33 (.L_HI(net33));
 sg13g2_tiehi _1568__34 (.L_HI(net34));
 sg13g2_tiehi _1532__35 (.L_HI(net35));
 sg13g2_tiehi _1567__36 (.L_HI(net36));
 sg13g2_tiehi _1571__37 (.L_HI(net37));
 sg13g2_tiehi _1566__38 (.L_HI(net38));
 sg13g2_tiehi _1573__39 (.L_HI(net39));
 sg13g2_tiehi _1565__40 (.L_HI(net40));
 sg13g2_tiehi _1564__41 (.L_HI(net41));
 sg13g2_tiehi _1563__42 (.L_HI(net42));
 sg13g2_tiehi _1562__43 (.L_HI(net43));
 sg13g2_tiehi _1561__44 (.L_HI(net44));
 sg13g2_tiehi _1560__45 (.L_HI(net45));
 sg13g2_tiehi _1559__46 (.L_HI(net46));
 sg13g2_tiehi _1558__47 (.L_HI(net47));
 sg13g2_tiehi _1557__48 (.L_HI(net48));
 sg13g2_tiehi _1556__49 (.L_HI(net49));
 sg13g2_tiehi _1555__50 (.L_HI(net50));
 sg13g2_tiehi _1554__51 (.L_HI(net51));
 sg13g2_tiehi _1553__52 (.L_HI(net52));
 sg13g2_tiehi _1552__53 (.L_HI(net53));
 sg13g2_tiehi _1551__54 (.L_HI(net54));
 sg13g2_tiehi _1550__55 (.L_HI(net55));
 sg13g2_tiehi _1549__56 (.L_HI(net56));
 sg13g2_tiehi _1548__57 (.L_HI(net57));
 sg13g2_tiehi _1547__58 (.L_HI(net58));
 sg13g2_tiehi _1546__59 (.L_HI(net59));
 sg13g2_tiehi _1545__60 (.L_HI(net60));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_sushi_demo_3 (.L_LO(net3));
 sg13g2_tielo tt_um_sushi_demo_4 (.L_LO(net4));
 sg13g2_tielo tt_um_sushi_demo_5 (.L_LO(net5));
 sg13g2_tielo tt_um_sushi_demo_6 (.L_LO(net6));
 sg13g2_tielo tt_um_sushi_demo_7 (.L_LO(net7));
 sg13g2_tielo tt_um_sushi_demo_8 (.L_LO(net8));
 sg13g2_tielo tt_um_sushi_demo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_sushi_demo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_sushi_demo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_sushi_demo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_sushi_demo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_sushi_demo_14 (.L_LO(net14));
 sg13g2_tielo tt_um_sushi_demo_15 (.L_LO(net15));
 sg13g2_tielo tt_um_sushi_demo_16 (.L_LO(net16));
 sg13g2_tielo tt_um_sushi_demo_17 (.L_LO(net17));
 sg13g2_tiehi _1544__18 (.L_HI(net18));
 sg13g2_buf_1 _1634_ (.A(net249),
    .X(uo_out[3]));
 sg13g2_buf_1 _1635_ (.A(h_sync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout195 (.A(net196),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_0393_),
    .X(net196));
 sg13g2_buf_1 fanout197 (.A(_0393_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_0412_),
    .X(net198));
 sg13g2_buf_4 fanout199 (.X(net199),
    .A(net201));
 sg13g2_buf_1 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_1 fanout201 (.A(_0352_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(net204),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(net204),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_0348_),
    .X(net204));
 sg13g2_buf_4 fanout205 (.X(net205),
    .A(_0347_));
 sg13g2_buf_4 fanout206 (.X(net206),
    .A(_0347_));
 sg13g2_buf_2 fanout207 (.A(net208),
    .X(net207));
 sg13g2_buf_4 fanout208 (.X(net208),
    .A(_0345_));
 sg13g2_buf_2 fanout209 (.A(net210),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_0344_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(net212),
    .X(net211));
 sg13g2_buf_4 fanout212 (.X(net212),
    .A(_0331_));
 sg13g2_buf_2 fanout213 (.A(net214),
    .X(net213));
 sg13g2_buf_4 fanout214 (.X(net214),
    .A(_0330_));
 sg13g2_buf_4 fanout215 (.X(net215),
    .A(_0320_));
 sg13g2_buf_2 fanout216 (.A(_0320_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(net218),
    .X(net217));
 sg13g2_buf_4 fanout218 (.X(net218),
    .A(_0318_));
 sg13g2_buf_2 fanout219 (.A(_0296_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_0296_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_0274_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_0274_),
    .X(net222));
 sg13g2_buf_4 fanout223 (.X(net223),
    .A(_0333_));
 sg13g2_buf_2 fanout224 (.A(_0273_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_0271_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_0270_),
    .X(net226));
 sg13g2_buf_1 fanout227 (.A(_0235_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_0341_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(net230),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_0332_),
    .X(net230));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(_0312_));
 sg13g2_buf_2 fanout232 (.A(_0305_),
    .X(net232));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(_0349_));
 sg13g2_buf_1 fanout234 (.A(_0349_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_0325_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_0325_),
    .X(net236));
 sg13g2_buf_4 fanout237 (.X(net237),
    .A(_0304_));
 sg13g2_buf_2 fanout238 (.A(_0299_),
    .X(net238));
 sg13g2_buf_4 fanout239 (.X(net239),
    .A(_0297_));
 sg13g2_buf_4 fanout240 (.X(net240),
    .A(_0285_));
 sg13g2_buf_2 fanout241 (.A(_0284_),
    .X(net241));
 sg13g2_buf_4 fanout242 (.X(net242),
    .A(_0287_));
 sg13g2_buf_4 fanout243 (.X(net243),
    .A(_0282_));
 sg13g2_buf_2 fanout244 (.A(_0279_),
    .X(net244));
 sg13g2_buf_4 fanout245 (.X(net245),
    .A(_0277_));
 sg13g2_buf_2 fanout246 (.A(_0062_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(net102),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(net98),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(net250),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(v_sync),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(net95),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(\pix_x[6] ),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(\pix_x[5] ),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(net255),
    .X(net254));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(net1));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_tielo tt_um_sushi_demo_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0011_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0012_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0008_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0045_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold5 (.A(\pix_y[1] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0713_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0046_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold8 (.A(\pix_x[2] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0064_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0014_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold11 (.A(\pix_y[5] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0050_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold13 (.A(\pix_y[8] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0706_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0044_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0004_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0068_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold18 (.A(\pix_x[0] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0063_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold20 (.A(\pix_x[5] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0070_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0000_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0074_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0075_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold25 (.A(\pix_y[4] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0049_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold27 (.A(\pix_x[3] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0065_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold29 (.A(\pix_y[6] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0722_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0051_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold32 (.A(\pix_x[4] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold33 (.A(\pix_y[9] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0054_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold35 (.A(\pix_x[7] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0073_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold37 (.A(\pix_y[7] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold38 (.A(\pix_y[2] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0715_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold40 (.A(\pix_x[6] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0704_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold42 (.A(\pix_y[3] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0000_),
    .X(net103));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_4 FILLER_12_273 ();
 sg13g2_fill_2 FILLER_12_277 ();
 sg13g2_decap_4 FILLER_12_287 ();
 sg13g2_fill_2 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_302 ();
 sg13g2_decap_8 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_316 ();
 sg13g2_fill_1 FILLER_12_323 ();
 sg13g2_fill_2 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_fill_1 FILLER_13_252 ();
 sg13g2_decap_4 FILLER_13_271 ();
 sg13g2_fill_1 FILLER_13_305 ();
 sg13g2_fill_2 FILLER_13_321 ();
 sg13g2_fill_2 FILLER_13_349 ();
 sg13g2_fill_1 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_4 FILLER_14_231 ();
 sg13g2_fill_1 FILLER_14_235 ();
 sg13g2_decap_8 FILLER_14_240 ();
 sg13g2_fill_2 FILLER_14_247 ();
 sg13g2_fill_2 FILLER_14_294 ();
 sg13g2_fill_1 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_fill_1 FILLER_15_224 ();
 sg13g2_fill_2 FILLER_15_337 ();
 sg13g2_fill_1 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_fill_1 FILLER_16_217 ();
 sg13g2_fill_1 FILLER_16_222 ();
 sg13g2_fill_2 FILLER_16_250 ();
 sg13g2_fill_2 FILLER_16_260 ();
 sg13g2_fill_1 FILLER_16_262 ();
 sg13g2_fill_2 FILLER_16_271 ();
 sg13g2_fill_2 FILLER_16_323 ();
 sg13g2_fill_1 FILLER_16_325 ();
 sg13g2_fill_2 FILLER_16_342 ();
 sg13g2_fill_1 FILLER_16_344 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_4 FILLER_17_203 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_217 ();
 sg13g2_fill_2 FILLER_17_240 ();
 sg13g2_fill_1 FILLER_17_242 ();
 sg13g2_fill_2 FILLER_17_256 ();
 sg13g2_fill_1 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_268 ();
 sg13g2_fill_2 FILLER_17_275 ();
 sg13g2_fill_1 FILLER_17_277 ();
 sg13g2_decap_4 FILLER_17_291 ();
 sg13g2_fill_2 FILLER_17_350 ();
 sg13g2_fill_1 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_fill_2 FILLER_18_182 ();
 sg13g2_decap_4 FILLER_18_194 ();
 sg13g2_fill_1 FILLER_18_198 ();
 sg13g2_decap_8 FILLER_18_212 ();
 sg13g2_decap_4 FILLER_18_219 ();
 sg13g2_decap_8 FILLER_18_269 ();
 sg13g2_fill_2 FILLER_18_276 ();
 sg13g2_fill_1 FILLER_18_278 ();
 sg13g2_fill_1 FILLER_18_315 ();
 sg13g2_fill_2 FILLER_18_321 ();
 sg13g2_fill_1 FILLER_18_323 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_4 FILLER_19_112 ();
 sg13g2_fill_2 FILLER_19_116 ();
 sg13g2_fill_2 FILLER_19_132 ();
 sg13g2_fill_1 FILLER_19_134 ();
 sg13g2_decap_8 FILLER_19_152 ();
 sg13g2_decap_8 FILLER_19_164 ();
 sg13g2_decap_4 FILLER_19_171 ();
 sg13g2_fill_2 FILLER_19_183 ();
 sg13g2_fill_1 FILLER_19_185 ();
 sg13g2_decap_4 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_218 ();
 sg13g2_decap_8 FILLER_19_239 ();
 sg13g2_fill_2 FILLER_19_246 ();
 sg13g2_decap_8 FILLER_19_253 ();
 sg13g2_decap_8 FILLER_19_260 ();
 sg13g2_fill_2 FILLER_19_267 ();
 sg13g2_fill_1 FILLER_19_269 ();
 sg13g2_fill_1 FILLER_19_291 ();
 sg13g2_fill_2 FILLER_19_307 ();
 sg13g2_decap_4 FILLER_19_339 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_fill_1 FILLER_19_354 ();
 sg13g2_fill_1 FILLER_19_372 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_fill_1 FILLER_20_134 ();
 sg13g2_fill_2 FILLER_20_147 ();
 sg13g2_decap_4 FILLER_20_171 ();
 sg13g2_fill_1 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_191 ();
 sg13g2_fill_2 FILLER_20_198 ();
 sg13g2_fill_1 FILLER_20_200 ();
 sg13g2_fill_2 FILLER_20_208 ();
 sg13g2_fill_1 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_225 ();
 sg13g2_decap_4 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_244 ();
 sg13g2_fill_1 FILLER_20_260 ();
 sg13g2_fill_2 FILLER_20_276 ();
 sg13g2_fill_1 FILLER_20_278 ();
 sg13g2_fill_2 FILLER_20_292 ();
 sg13g2_decap_4 FILLER_20_318 ();
 sg13g2_fill_1 FILLER_20_322 ();
 sg13g2_decap_4 FILLER_20_327 ();
 sg13g2_fill_2 FILLER_20_331 ();
 sg13g2_fill_2 FILLER_20_390 ();
 sg13g2_fill_1 FILLER_20_392 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_4 FILLER_21_77 ();
 sg13g2_fill_2 FILLER_21_93 ();
 sg13g2_decap_8 FILLER_21_130 ();
 sg13g2_fill_2 FILLER_21_137 ();
 sg13g2_fill_1 FILLER_21_147 ();
 sg13g2_decap_4 FILLER_21_161 ();
 sg13g2_fill_1 FILLER_21_170 ();
 sg13g2_decap_4 FILLER_21_183 ();
 sg13g2_fill_1 FILLER_21_195 ();
 sg13g2_decap_4 FILLER_21_223 ();
 sg13g2_fill_1 FILLER_21_227 ();
 sg13g2_decap_4 FILLER_21_256 ();
 sg13g2_fill_2 FILLER_21_271 ();
 sg13g2_fill_1 FILLER_21_273 ();
 sg13g2_decap_4 FILLER_21_291 ();
 sg13g2_fill_1 FILLER_21_295 ();
 sg13g2_decap_4 FILLER_21_313 ();
 sg13g2_fill_2 FILLER_21_317 ();
 sg13g2_fill_2 FILLER_21_327 ();
 sg13g2_fill_1 FILLER_21_329 ();
 sg13g2_fill_2 FILLER_21_335 ();
 sg13g2_fill_2 FILLER_21_351 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_fill_2 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_37 ();
 sg13g2_decap_8 FILLER_22_47 ();
 sg13g2_decap_8 FILLER_22_54 ();
 sg13g2_fill_1 FILLER_22_61 ();
 sg13g2_decap_4 FILLER_22_66 ();
 sg13g2_fill_1 FILLER_22_70 ();
 sg13g2_fill_1 FILLER_22_83 ();
 sg13g2_decap_4 FILLER_22_97 ();
 sg13g2_decap_4 FILLER_22_139 ();
 sg13g2_fill_2 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_2 FILLER_22_176 ();
 sg13g2_fill_1 FILLER_22_188 ();
 sg13g2_decap_4 FILLER_22_194 ();
 sg13g2_fill_2 FILLER_22_198 ();
 sg13g2_fill_1 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_216 ();
 sg13g2_decap_8 FILLER_22_223 ();
 sg13g2_decap_4 FILLER_22_230 ();
 sg13g2_fill_2 FILLER_22_234 ();
 sg13g2_decap_8 FILLER_22_241 ();
 sg13g2_decap_4 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_265 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_4 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_295 ();
 sg13g2_decap_8 FILLER_22_302 ();
 sg13g2_fill_2 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_fill_2 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_2 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_30 ();
 sg13g2_fill_2 FILLER_23_57 ();
 sg13g2_fill_2 FILLER_23_77 ();
 sg13g2_fill_1 FILLER_23_79 ();
 sg13g2_fill_1 FILLER_23_88 ();
 sg13g2_fill_2 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_107 ();
 sg13g2_decap_8 FILLER_23_127 ();
 sg13g2_decap_8 FILLER_23_134 ();
 sg13g2_decap_8 FILLER_23_141 ();
 sg13g2_decap_8 FILLER_23_148 ();
 sg13g2_fill_2 FILLER_23_155 ();
 sg13g2_decap_4 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_195 ();
 sg13g2_decap_4 FILLER_23_209 ();
 sg13g2_decap_4 FILLER_23_226 ();
 sg13g2_fill_2 FILLER_23_230 ();
 sg13g2_decap_4 FILLER_23_248 ();
 sg13g2_fill_1 FILLER_23_252 ();
 sg13g2_fill_2 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_330 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_fill_2 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_32 ();
 sg13g2_decap_4 FILLER_24_58 ();
 sg13g2_fill_2 FILLER_24_62 ();
 sg13g2_decap_8 FILLER_24_85 ();
 sg13g2_decap_8 FILLER_24_92 ();
 sg13g2_decap_4 FILLER_24_99 ();
 sg13g2_fill_1 FILLER_24_103 ();
 sg13g2_decap_8 FILLER_24_108 ();
 sg13g2_decap_4 FILLER_24_135 ();
 sg13g2_fill_2 FILLER_24_139 ();
 sg13g2_decap_4 FILLER_24_178 ();
 sg13g2_fill_1 FILLER_24_194 ();
 sg13g2_fill_2 FILLER_24_203 ();
 sg13g2_fill_1 FILLER_24_205 ();
 sg13g2_fill_2 FILLER_24_211 ();
 sg13g2_fill_1 FILLER_24_213 ();
 sg13g2_decap_4 FILLER_24_219 ();
 sg13g2_fill_1 FILLER_24_223 ();
 sg13g2_decap_8 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_256 ();
 sg13g2_fill_2 FILLER_24_263 ();
 sg13g2_decap_4 FILLER_24_280 ();
 sg13g2_fill_2 FILLER_24_292 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_4 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_317 ();
 sg13g2_fill_1 FILLER_24_336 ();
 sg13g2_fill_2 FILLER_24_345 ();
 sg13g2_fill_1 FILLER_24_347 ();
 sg13g2_fill_1 FILLER_24_353 ();
 sg13g2_fill_2 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_fill_2 FILLER_25_35 ();
 sg13g2_fill_1 FILLER_25_37 ();
 sg13g2_fill_2 FILLER_25_46 ();
 sg13g2_fill_1 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_68 ();
 sg13g2_fill_1 FILLER_25_70 ();
 sg13g2_fill_2 FILLER_25_92 ();
 sg13g2_fill_1 FILLER_25_104 ();
 sg13g2_fill_2 FILLER_25_115 ();
 sg13g2_fill_1 FILLER_25_117 ();
 sg13g2_fill_2 FILLER_25_122 ();
 sg13g2_fill_1 FILLER_25_124 ();
 sg13g2_decap_4 FILLER_25_138 ();
 sg13g2_decap_8 FILLER_25_153 ();
 sg13g2_decap_4 FILLER_25_160 ();
 sg13g2_fill_1 FILLER_25_164 ();
 sg13g2_fill_1 FILLER_25_178 ();
 sg13g2_fill_2 FILLER_25_191 ();
 sg13g2_fill_2 FILLER_25_201 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_218 ();
 sg13g2_decap_4 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_294 ();
 sg13g2_fill_1 FILLER_25_300 ();
 sg13g2_fill_2 FILLER_25_342 ();
 sg13g2_fill_1 FILLER_25_344 ();
 sg13g2_fill_1 FILLER_25_358 ();
 sg13g2_fill_1 FILLER_25_364 ();
 sg13g2_fill_2 FILLER_25_398 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_fill_2 FILLER_26_21 ();
 sg13g2_fill_2 FILLER_26_58 ();
 sg13g2_fill_2 FILLER_26_79 ();
 sg13g2_fill_1 FILLER_26_81 ();
 sg13g2_fill_1 FILLER_26_109 ();
 sg13g2_fill_1 FILLER_26_120 ();
 sg13g2_decap_4 FILLER_26_147 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_fill_1 FILLER_26_179 ();
 sg13g2_fill_2 FILLER_26_185 ();
 sg13g2_fill_1 FILLER_26_187 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_207 ();
 sg13g2_fill_2 FILLER_26_218 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_decap_8 FILLER_26_246 ();
 sg13g2_decap_4 FILLER_26_253 ();
 sg13g2_fill_1 FILLER_26_257 ();
 sg13g2_decap_8 FILLER_26_262 ();
 sg13g2_fill_2 FILLER_26_269 ();
 sg13g2_fill_1 FILLER_26_271 ();
 sg13g2_fill_2 FILLER_26_276 ();
 sg13g2_fill_1 FILLER_26_278 ();
 sg13g2_fill_1 FILLER_26_312 ();
 sg13g2_decap_4 FILLER_26_326 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_fill_1 FILLER_26_346 ();
 sg13g2_fill_1 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_43 ();
 sg13g2_fill_1 FILLER_27_45 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_decap_4 FILLER_27_57 ();
 sg13g2_fill_1 FILLER_27_61 ();
 sg13g2_fill_2 FILLER_27_73 ();
 sg13g2_fill_2 FILLER_27_80 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_101 ();
 sg13g2_fill_1 FILLER_27_103 ();
 sg13g2_decap_4 FILLER_27_113 ();
 sg13g2_fill_1 FILLER_27_117 ();
 sg13g2_fill_2 FILLER_27_131 ();
 sg13g2_fill_2 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_185 ();
 sg13g2_decap_8 FILLER_27_194 ();
 sg13g2_decap_8 FILLER_27_201 ();
 sg13g2_decap_8 FILLER_27_220 ();
 sg13g2_fill_1 FILLER_27_227 ();
 sg13g2_decap_4 FILLER_27_244 ();
 sg13g2_fill_2 FILLER_27_248 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_decap_8 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_fill_1 FILLER_27_327 ();
 sg13g2_fill_2 FILLER_27_336 ();
 sg13g2_fill_1 FILLER_27_338 ();
 sg13g2_fill_1 FILLER_27_368 ();
 sg13g2_fill_2 FILLER_27_378 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_23 ();
 sg13g2_fill_2 FILLER_28_27 ();
 sg13g2_fill_1 FILLER_28_67 ();
 sg13g2_decap_4 FILLER_28_76 ();
 sg13g2_fill_1 FILLER_28_80 ();
 sg13g2_fill_2 FILLER_28_100 ();
 sg13g2_fill_1 FILLER_28_102 ();
 sg13g2_decap_4 FILLER_28_120 ();
 sg13g2_fill_1 FILLER_28_124 ();
 sg13g2_fill_2 FILLER_28_130 ();
 sg13g2_fill_1 FILLER_28_132 ();
 sg13g2_fill_2 FILLER_28_142 ();
 sg13g2_fill_1 FILLER_28_154 ();
 sg13g2_decap_4 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_165 ();
 sg13g2_decap_8 FILLER_28_177 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_fill_2 FILLER_28_192 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_244 ();
 sg13g2_decap_4 FILLER_28_251 ();
 sg13g2_fill_2 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_265 ();
 sg13g2_decap_8 FILLER_28_272 ();
 sg13g2_fill_2 FILLER_28_279 ();
 sg13g2_decap_8 FILLER_28_323 ();
 sg13g2_decap_4 FILLER_28_330 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_9 ();
 sg13g2_fill_2 FILLER_29_31 ();
 sg13g2_fill_1 FILLER_29_33 ();
 sg13g2_decap_4 FILLER_29_55 ();
 sg13g2_fill_2 FILLER_29_59 ();
 sg13g2_decap_4 FILLER_29_71 ();
 sg13g2_decap_4 FILLER_29_85 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_112 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_150 ();
 sg13g2_fill_2 FILLER_29_157 ();
 sg13g2_decap_4 FILLER_29_164 ();
 sg13g2_fill_2 FILLER_29_173 ();
 sg13g2_fill_2 FILLER_29_180 ();
 sg13g2_fill_2 FILLER_29_197 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_fill_2 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_226 ();
 sg13g2_fill_1 FILLER_29_243 ();
 sg13g2_decap_4 FILLER_29_274 ();
 sg13g2_fill_2 FILLER_29_278 ();
 sg13g2_fill_2 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_fill_2 FILLER_29_322 ();
 sg13g2_fill_1 FILLER_29_324 ();
 sg13g2_fill_2 FILLER_29_336 ();
 sg13g2_fill_2 FILLER_29_359 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_22 ();
 sg13g2_fill_2 FILLER_30_27 ();
 sg13g2_fill_1 FILLER_30_29 ();
 sg13g2_fill_2 FILLER_30_47 ();
 sg13g2_fill_1 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_78 ();
 sg13g2_fill_1 FILLER_30_80 ();
 sg13g2_decap_4 FILLER_30_127 ();
 sg13g2_decap_8 FILLER_30_139 ();
 sg13g2_decap_4 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_150 ();
 sg13g2_fill_2 FILLER_30_167 ();
 sg13g2_decap_4 FILLER_30_187 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_fill_2 FILLER_30_208 ();
 sg13g2_decap_8 FILLER_30_214 ();
 sg13g2_fill_1 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_236 ();
 sg13g2_decap_8 FILLER_30_243 ();
 sg13g2_decap_8 FILLER_30_250 ();
 sg13g2_fill_2 FILLER_30_257 ();
 sg13g2_fill_2 FILLER_30_285 ();
 sg13g2_fill_1 FILLER_30_296 ();
 sg13g2_fill_2 FILLER_30_336 ();
 sg13g2_decap_4 FILLER_30_342 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_fill_1 FILLER_30_372 ();
 sg13g2_fill_2 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_33 ();
 sg13g2_fill_1 FILLER_31_37 ();
 sg13g2_decap_8 FILLER_31_55 ();
 sg13g2_decap_4 FILLER_31_62 ();
 sg13g2_decap_8 FILLER_31_72 ();
 sg13g2_decap_4 FILLER_31_85 ();
 sg13g2_fill_2 FILLER_31_89 ();
 sg13g2_decap_8 FILLER_31_110 ();
 sg13g2_decap_4 FILLER_31_117 ();
 sg13g2_fill_1 FILLER_31_121 ();
 sg13g2_decap_4 FILLER_31_127 ();
 sg13g2_fill_2 FILLER_31_131 ();
 sg13g2_fill_2 FILLER_31_147 ();
 sg13g2_fill_1 FILLER_31_149 ();
 sg13g2_decap_4 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_189 ();
 sg13g2_fill_1 FILLER_31_191 ();
 sg13g2_fill_2 FILLER_31_198 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_219 ();
 sg13g2_fill_1 FILLER_31_221 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_fill_2 FILLER_31_237 ();
 sg13g2_fill_1 FILLER_31_239 ();
 sg13g2_decap_4 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_278 ();
 sg13g2_decap_4 FILLER_31_285 ();
 sg13g2_fill_2 FILLER_31_289 ();
 sg13g2_decap_4 FILLER_31_321 ();
 sg13g2_fill_2 FILLER_31_325 ();
 sg13g2_decap_8 FILLER_31_358 ();
 sg13g2_fill_2 FILLER_31_370 ();
 sg13g2_fill_1 FILLER_31_372 ();
 sg13g2_fill_2 FILLER_31_391 ();
 sg13g2_fill_1 FILLER_31_393 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_4 ();
 sg13g2_fill_1 FILLER_32_22 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_fill_2 FILLER_32_46 ();
 sg13g2_fill_2 FILLER_32_64 ();
 sg13g2_fill_2 FILLER_32_77 ();
 sg13g2_fill_1 FILLER_32_79 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_136 ();
 sg13g2_fill_1 FILLER_32_138 ();
 sg13g2_fill_2 FILLER_32_149 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_175 ();
 sg13g2_fill_1 FILLER_32_177 ();
 sg13g2_decap_4 FILLER_32_197 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_4 FILLER_32_224 ();
 sg13g2_fill_2 FILLER_32_237 ();
 sg13g2_decap_4 FILLER_32_255 ();
 sg13g2_fill_2 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_265 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_fill_2 FILLER_32_299 ();
 sg13g2_decap_4 FILLER_32_315 ();
 sg13g2_decap_4 FILLER_32_324 ();
 sg13g2_fill_1 FILLER_32_328 ();
 sg13g2_decap_8 FILLER_32_333 ();
 sg13g2_decap_4 FILLER_32_340 ();
 sg13g2_fill_1 FILLER_32_344 ();
 sg13g2_fill_2 FILLER_32_389 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_4 ();
 sg13g2_decap_4 FILLER_33_27 ();
 sg13g2_fill_1 FILLER_33_31 ();
 sg13g2_fill_2 FILLER_33_53 ();
 sg13g2_fill_2 FILLER_33_71 ();
 sg13g2_fill_1 FILLER_33_102 ();
 sg13g2_decap_8 FILLER_33_113 ();
 sg13g2_decap_8 FILLER_33_124 ();
 sg13g2_decap_4 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_135 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_fill_1 FILLER_33_184 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_fill_1 FILLER_33_208 ();
 sg13g2_fill_2 FILLER_33_216 ();
 sg13g2_fill_1 FILLER_33_218 ();
 sg13g2_decap_8 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_decap_4 FILLER_33_288 ();
 sg13g2_fill_2 FILLER_33_292 ();
 sg13g2_fill_1 FILLER_33_306 ();
 sg13g2_fill_1 FILLER_33_317 ();
 sg13g2_decap_4 FILLER_33_344 ();
 sg13g2_fill_2 FILLER_33_348 ();
 sg13g2_fill_2 FILLER_33_355 ();
 sg13g2_fill_1 FILLER_33_374 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_9 ();
 sg13g2_fill_2 FILLER_34_26 ();
 sg13g2_decap_4 FILLER_34_34 ();
 sg13g2_fill_1 FILLER_34_38 ();
 sg13g2_fill_2 FILLER_34_43 ();
 sg13g2_fill_1 FILLER_34_45 ();
 sg13g2_fill_2 FILLER_34_51 ();
 sg13g2_fill_1 FILLER_34_58 ();
 sg13g2_decap_4 FILLER_34_70 ();
 sg13g2_fill_1 FILLER_34_83 ();
 sg13g2_fill_2 FILLER_34_88 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_fill_1 FILLER_34_95 ();
 sg13g2_fill_2 FILLER_34_101 ();
 sg13g2_fill_1 FILLER_34_103 ();
 sg13g2_decap_4 FILLER_34_116 ();
 sg13g2_fill_1 FILLER_34_120 ();
 sg13g2_fill_2 FILLER_34_131 ();
 sg13g2_fill_1 FILLER_34_133 ();
 sg13g2_fill_2 FILLER_34_157 ();
 sg13g2_fill_1 FILLER_34_159 ();
 sg13g2_fill_2 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_181 ();
 sg13g2_fill_1 FILLER_34_189 ();
 sg13g2_fill_1 FILLER_34_194 ();
 sg13g2_decap_4 FILLER_34_203 ();
 sg13g2_decap_4 FILLER_34_235 ();
 sg13g2_decap_4 FILLER_34_244 ();
 sg13g2_decap_8 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_283 ();
 sg13g2_decap_8 FILLER_34_288 ();
 sg13g2_fill_1 FILLER_34_295 ();
 sg13g2_decap_4 FILLER_34_306 ();
 sg13g2_decap_4 FILLER_34_314 ();
 sg13g2_fill_1 FILLER_34_318 ();
 sg13g2_fill_1 FILLER_34_345 ();
 sg13g2_fill_2 FILLER_34_354 ();
 sg13g2_fill_1 FILLER_34_356 ();
 sg13g2_fill_2 FILLER_34_361 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_decap_8 FILLER_34_379 ();
 sg13g2_decap_8 FILLER_34_386 ();
 sg13g2_decap_8 FILLER_34_393 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_43 ();
 sg13g2_fill_1 FILLER_35_45 ();
 sg13g2_fill_1 FILLER_35_58 ();
 sg13g2_fill_1 FILLER_35_69 ();
 sg13g2_fill_2 FILLER_35_82 ();
 sg13g2_fill_1 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_106 ();
 sg13g2_fill_2 FILLER_35_133 ();
 sg13g2_fill_1 FILLER_35_135 ();
 sg13g2_decap_8 FILLER_35_157 ();
 sg13g2_fill_2 FILLER_35_164 ();
 sg13g2_fill_1 FILLER_35_166 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_fill_2 FILLER_35_211 ();
 sg13g2_fill_1 FILLER_35_238 ();
 sg13g2_fill_1 FILLER_35_257 ();
 sg13g2_fill_2 FILLER_35_262 ();
 sg13g2_fill_1 FILLER_35_326 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_fill_2 FILLER_35_343 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_decap_8 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_14 ();
 sg13g2_fill_2 FILLER_36_22 ();
 sg13g2_fill_1 FILLER_36_24 ();
 sg13g2_decap_8 FILLER_36_37 ();
 sg13g2_fill_2 FILLER_36_53 ();
 sg13g2_decap_8 FILLER_36_64 ();
 sg13g2_fill_1 FILLER_36_71 ();
 sg13g2_decap_8 FILLER_36_81 ();
 sg13g2_fill_2 FILLER_36_98 ();
 sg13g2_decap_4 FILLER_36_131 ();
 sg13g2_fill_1 FILLER_36_145 ();
 sg13g2_decap_4 FILLER_36_160 ();
 sg13g2_decap_4 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_191 ();
 sg13g2_decap_8 FILLER_36_198 ();
 sg13g2_decap_8 FILLER_36_205 ();
 sg13g2_fill_2 FILLER_36_212 ();
 sg13g2_decap_4 FILLER_36_223 ();
 sg13g2_fill_2 FILLER_36_227 ();
 sg13g2_decap_4 FILLER_36_232 ();
 sg13g2_fill_2 FILLER_36_236 ();
 sg13g2_decap_4 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_decap_8 FILLER_36_302 ();
 sg13g2_decap_8 FILLER_36_309 ();
 sg13g2_decap_8 FILLER_36_316 ();
 sg13g2_decap_8 FILLER_36_323 ();
 sg13g2_decap_8 FILLER_36_330 ();
 sg13g2_decap_8 FILLER_36_337 ();
 sg13g2_decap_8 FILLER_36_344 ();
 sg13g2_decap_8 FILLER_36_351 ();
 sg13g2_decap_8 FILLER_36_358 ();
 sg13g2_decap_8 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_124 ();
 sg13g2_decap_8 FILLER_37_131 ();
 sg13g2_fill_1 FILLER_37_138 ();
 sg13g2_decap_8 FILLER_37_158 ();
 sg13g2_decap_4 FILLER_37_165 ();
 sg13g2_decap_8 FILLER_37_174 ();
 sg13g2_decap_8 FILLER_37_181 ();
 sg13g2_decap_8 FILLER_37_188 ();
 sg13g2_decap_8 FILLER_37_195 ();
 sg13g2_decap_8 FILLER_37_202 ();
 sg13g2_decap_8 FILLER_37_209 ();
 sg13g2_decap_8 FILLER_37_216 ();
 sg13g2_decap_8 FILLER_37_223 ();
 sg13g2_decap_8 FILLER_37_230 ();
 sg13g2_decap_8 FILLER_37_237 ();
 sg13g2_decap_8 FILLER_37_244 ();
 sg13g2_decap_4 FILLER_37_251 ();
 sg13g2_fill_1 FILLER_37_255 ();
 sg13g2_decap_8 FILLER_37_260 ();
 sg13g2_decap_8 FILLER_37_267 ();
 sg13g2_decap_8 FILLER_37_274 ();
 sg13g2_decap_4 FILLER_37_281 ();
 sg13g2_fill_2 FILLER_37_285 ();
 sg13g2_decap_8 FILLER_37_291 ();
 sg13g2_decap_8 FILLER_37_298 ();
 sg13g2_decap_8 FILLER_37_305 ();
 sg13g2_decap_8 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_decap_8 FILLER_37_333 ();
 sg13g2_decap_8 FILLER_37_340 ();
 sg13g2_decap_8 FILLER_37_347 ();
 sg13g2_decap_8 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_37_361 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_decap_8 FILLER_38_285 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_decap_8 FILLER_38_299 ();
 sg13g2_decap_8 FILLER_38_306 ();
 sg13g2_decap_8 FILLER_38_313 ();
 sg13g2_decap_8 FILLER_38_320 ();
 sg13g2_decap_8 FILLER_38_327 ();
 sg13g2_decap_8 FILLER_38_334 ();
 sg13g2_decap_8 FILLER_38_341 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_decap_8 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_362 ();
 sg13g2_decap_8 FILLER_38_369 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
endmodule

module tt_um_htfab_checkers (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire clknet_0_clk;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;

 sg13g2_inv_1 _0501_ (.Y(_0443_),
    .A(net87));
 sg13g2_inv_1 _0502_ (.Y(_0444_),
    .A(\counter[7] ));
 sg13g2_inv_2 _0503_ (.Y(_0445_),
    .A(net165));
 sg13g2_inv_1 _0504_ (.Y(_0446_),
    .A(net170));
 sg13g2_inv_1 _0505_ (.Y(_0447_),
    .A(net175));
 sg13g2_inv_1 _0506_ (.Y(_0448_),
    .A(net58));
 sg13g2_inv_1 _0507_ (.Y(_0449_),
    .A(net155));
 sg13g2_inv_1 _0508_ (.Y(_0450_),
    .A(net146));
 sg13g2_inv_1 _0509_ (.Y(_0046_),
    .A(net148));
 sg13g2_inv_1 _0510_ (.Y(_0047_),
    .A(net75));
 sg13g2_inv_1 _0511_ (.Y(_0048_),
    .A(net187));
 sg13g2_inv_1 _0512_ (.Y(_0049_),
    .A(net3));
 sg13g2_inv_1 _0513_ (.Y(_0050_),
    .A(_0005_));
 sg13g2_inv_1 _0514_ (.Y(_0051_),
    .A(_0007_));
 sg13g2_inv_1 _0515_ (.Y(_0052_),
    .A(net90));
 sg13g2_inv_1 _0516_ (.Y(_0053_),
    .A(net8));
 sg13g2_inv_1 _0517_ (.Y(_0054_),
    .A(net2));
 sg13g2_inv_1 _0518_ (.Y(_0055_),
    .A(net1));
 sg13g2_nor2_1 _0519_ (.A(_0047_),
    .B(net67),
    .Y(_0056_));
 sg13g2_and2_1 _0520_ (.A(net86),
    .B(net84),
    .X(_0057_));
 sg13g2_nand4_1 _0521_ (.B(net150),
    .C(_0056_),
    .A(net154),
    .Y(_0058_),
    .D(_0057_));
 sg13g2_nor4_1 _0522_ (.A(net151),
    .B(_0450_),
    .C(net147),
    .D(_0058_),
    .Y(_0001_));
 sg13g2_nand2_1 _0523_ (.Y(_0059_),
    .A(\hvsync_gen.hpos[9] ),
    .B(\hvsync_gen.hpos[8] ));
 sg13g2_or3_1 _0524_ (.A(net160),
    .B(net159),
    .C(net157),
    .X(_0060_));
 sg13g2_nand3_1 _0525_ (.B(\hvsync_gen.hpos[9] ),
    .C(_0060_),
    .A(\hvsync_gen.hpos[7] ),
    .Y(_0061_));
 sg13g2_nand4_1 _0526_ (.B(net159),
    .C(net156),
    .A(net160),
    .Y(_0062_),
    .D(net157));
 sg13g2_nor2b_1 _0527_ (.A(\hvsync_gen.hpos[8] ),
    .B_N(\hvsync_gen.hpos[9] ),
    .Y(_0063_));
 sg13g2_a21oi_1 _0528_ (.A1(_0062_),
    .A2(_0063_),
    .Y(_0064_),
    .B1(net60));
 sg13g2_a21oi_1 _0529_ (.A1(_0059_),
    .A2(_0061_),
    .Y(_0000_),
    .B1(net61));
 sg13g2_and2_1 _0530_ (.A(net178),
    .B(net160),
    .X(_0065_));
 sg13g2_nor2_1 _0531_ (.A(net178),
    .B(\hvsync_gen.hpos[4] ),
    .Y(_0066_));
 sg13g2_nor2_1 _0532_ (.A(_0065_),
    .B(_0066_),
    .Y(_0067_));
 sg13g2_a21oi_1 _0533_ (.A1(net177),
    .A2(_0067_),
    .Y(_0068_),
    .B1(_0065_));
 sg13g2_and2_1 _0534_ (.A(net173),
    .B(net159),
    .X(_0069_));
 sg13g2_xor2_1 _0535_ (.B(\hvsync_gen.hpos[5] ),
    .A(net173),
    .X(_0070_));
 sg13g2_xnor2_1 _0536_ (.Y(_0071_),
    .A(net172),
    .B(_0070_));
 sg13g2_nor2_1 _0537_ (.A(_0068_),
    .B(_0071_),
    .Y(_0072_));
 sg13g2_xor2_1 _0538_ (.B(_0071_),
    .A(_0068_),
    .X(_0073_));
 sg13g2_a21oi_1 _0539_ (.A1(net169),
    .A2(_0073_),
    .Y(_0074_),
    .B1(_0072_));
 sg13g2_a21oi_1 _0540_ (.A1(net172),
    .A2(_0070_),
    .Y(_0075_),
    .B1(_0069_));
 sg13g2_xor2_1 _0541_ (.B(net158),
    .A(net170),
    .X(_0076_));
 sg13g2_a21oi_1 _0542_ (.A1(net170),
    .A2(net158),
    .Y(_0077_),
    .B1(net168));
 sg13g2_xnor2_1 _0543_ (.Y(_0078_),
    .A(net168),
    .B(_0076_));
 sg13g2_or2_1 _0544_ (.X(_0079_),
    .B(_0078_),
    .A(_0075_));
 sg13g2_xnor2_1 _0545_ (.Y(_0080_),
    .A(_0075_),
    .B(_0078_));
 sg13g2_xnor2_1 _0546_ (.Y(_0081_),
    .A(_0445_),
    .B(_0080_));
 sg13g2_and2_1 _0547_ (.A(net185),
    .B(\hvsync_gen.hpos[2] ),
    .X(_0082_));
 sg13g2_xor2_1 _0548_ (.B(\hvsync_gen.hpos[2] ),
    .A(net185),
    .X(_0083_));
 sg13g2_a21oi_1 _0549_ (.A1(\counter[1] ),
    .A2(_0083_),
    .Y(_0084_),
    .B1(_0082_));
 sg13g2_and2_1 _0550_ (.A(net182),
    .B(net161),
    .X(_0085_));
 sg13g2_or2_1 _0551_ (.X(_0086_),
    .B(net161),
    .A(net182));
 sg13g2_nor2b_1 _0552_ (.A(_0085_),
    .B_N(_0086_),
    .Y(_0087_));
 sg13g2_xnor2_1 _0553_ (.Y(_0088_),
    .A(net179),
    .B(_0087_));
 sg13g2_nor2_1 _0554_ (.A(_0084_),
    .B(_0088_),
    .Y(_0089_));
 sg13g2_xor2_1 _0555_ (.B(_0088_),
    .A(_0084_),
    .X(_0090_));
 sg13g2_and2_1 _0556_ (.A(net176),
    .B(_0090_),
    .X(_0091_));
 sg13g2_nor2_1 _0557_ (.A(_0089_),
    .B(_0091_),
    .Y(_0092_));
 sg13g2_a21oi_1 _0558_ (.A1(net179),
    .A2(_0086_),
    .Y(_0093_),
    .B1(_0085_));
 sg13g2_xnor2_1 _0559_ (.Y(_0094_),
    .A(net176),
    .B(_0067_));
 sg13g2_nor2_1 _0560_ (.A(_0093_),
    .B(_0094_),
    .Y(_0095_));
 sg13g2_xor2_1 _0561_ (.B(_0094_),
    .A(_0093_),
    .X(_0096_));
 sg13g2_xnor2_1 _0562_ (.Y(_0097_),
    .A(net172),
    .B(_0096_));
 sg13g2_xor2_1 _0563_ (.B(_0083_),
    .A(net182),
    .X(_0098_));
 sg13g2_nand2_1 _0564_ (.Y(_0099_),
    .A(net183),
    .B(net184));
 sg13g2_and4_1 _0565_ (.A(net182),
    .B(net185),
    .C(\hvsync_gen.hpos[0] ),
    .D(net163),
    .X(_0100_));
 sg13g2_nand3_1 _0566_ (.B(_0098_),
    .C(_0100_),
    .A(net179),
    .Y(_0101_));
 sg13g2_nor3_1 _0567_ (.A(net179),
    .B(_0098_),
    .C(_0100_),
    .Y(_0102_));
 sg13g2_o21ai_1 _0568_ (.B1(net184),
    .Y(_0103_),
    .A1(\hvsync_gen.hpos[0] ),
    .A2(net163));
 sg13g2_o21ai_1 _0569_ (.B1(net182),
    .Y(_0104_),
    .A1(net184),
    .A2(net163));
 sg13g2_nand2_1 _0570_ (.Y(_0105_),
    .A(_0103_),
    .B(_0104_));
 sg13g2_a21oi_1 _0571_ (.A1(net179),
    .A2(_0098_),
    .Y(_0106_),
    .B1(_0105_));
 sg13g2_nor3_1 _0572_ (.A(_0091_),
    .B(_0102_),
    .C(_0106_),
    .Y(_0107_));
 sg13g2_o21ai_1 _0573_ (.B1(_0107_),
    .Y(_0108_),
    .A1(net176),
    .A2(_0090_));
 sg13g2_a22oi_1 _0574_ (.Y(_0109_),
    .B1(_0101_),
    .B2(_0108_),
    .A2(_0097_),
    .A1(_0092_));
 sg13g2_a21oi_1 _0575_ (.A1(net172),
    .A2(_0096_),
    .Y(_0110_),
    .B1(_0095_));
 sg13g2_xnor2_1 _0576_ (.Y(_0111_),
    .A(net169),
    .B(_0073_));
 sg13g2_or2_1 _0577_ (.X(_0112_),
    .B(_0111_),
    .A(_0110_));
 sg13g2_o21ai_1 _0578_ (.B1(_0112_),
    .Y(_0113_),
    .A1(_0092_),
    .A2(_0097_));
 sg13g2_a22oi_1 _0579_ (.Y(_0114_),
    .B1(_0110_),
    .B2(_0111_),
    .A2(_0081_),
    .A1(_0074_));
 sg13g2_o21ai_1 _0580_ (.B1(_0114_),
    .Y(_0115_),
    .A1(_0109_),
    .A2(_0113_));
 sg13g2_o21ai_1 _0581_ (.B1(_0115_),
    .Y(_0116_),
    .A1(_0074_),
    .A2(_0081_));
 sg13g2_and2_1 _0582_ (.A(net165),
    .B(net167),
    .X(_0117_));
 sg13g2_xor2_1 _0583_ (.B(net167),
    .A(net165),
    .X(_0118_));
 sg13g2_a21o_1 _0584_ (.A2(_0118_),
    .A1(net146),
    .B1(_0117_),
    .X(_0119_));
 sg13g2_nor2_1 _0585_ (.A(_0444_),
    .B(_0445_),
    .Y(_0120_));
 sg13g2_xor2_1 _0586_ (.B(net165),
    .A(\counter[7] ),
    .X(_0121_));
 sg13g2_xor2_1 _0587_ (.B(_0121_),
    .A(net144),
    .X(_0122_));
 sg13g2_and2_1 _0588_ (.A(net180),
    .B(net182),
    .X(_0123_));
 sg13g2_nor2_1 _0589_ (.A(net180),
    .B(net182),
    .Y(_0124_));
 sg13g2_nor2_1 _0590_ (.A(_0123_),
    .B(_0124_),
    .Y(_0125_));
 sg13g2_a21oi_1 _0591_ (.A1(net153),
    .A2(_0125_),
    .Y(_0126_),
    .B1(_0123_));
 sg13g2_or2_1 _0592_ (.X(_0127_),
    .B(net152),
    .A(net174));
 sg13g2_xor2_1 _0593_ (.B(net152),
    .A(net174),
    .X(_0128_));
 sg13g2_xnor2_1 _0594_ (.Y(_0129_),
    .A(net178),
    .B(_0128_));
 sg13g2_nand2_1 _0595_ (.Y(_0130_),
    .A(_0126_),
    .B(_0129_));
 sg13g2_xor2_1 _0596_ (.B(_0125_),
    .A(net153),
    .X(_0131_));
 sg13g2_nor2_1 _0597_ (.A(net183),
    .B(net184),
    .Y(_0132_));
 sg13g2_a21oi_1 _0598_ (.A1(_0013_),
    .A2(_0099_),
    .Y(_0133_),
    .B1(_0132_));
 sg13g2_nand3_1 _0599_ (.B(_0131_),
    .C(_0133_),
    .A(_0130_),
    .Y(_0134_));
 sg13g2_nand2_1 _0600_ (.Y(_0135_),
    .A(net171),
    .B(net174));
 sg13g2_xor2_1 _0601_ (.B(net174),
    .A(net171),
    .X(_0136_));
 sg13g2_nand2_1 _0602_ (.Y(_0137_),
    .A(net149),
    .B(_0136_));
 sg13g2_xor2_1 _0603_ (.B(_0136_),
    .A(net149),
    .X(_0138_));
 sg13g2_nand2_1 _0604_ (.Y(_0139_),
    .A(net174),
    .B(net178));
 sg13g2_nor2_1 _0605_ (.A(net174),
    .B(net178),
    .Y(_0140_));
 sg13g2_a21oi_1 _0606_ (.A1(_0010_),
    .A2(_0139_),
    .Y(_0141_),
    .B1(_0140_));
 sg13g2_nand2_1 _0607_ (.Y(_0142_),
    .A(_0138_),
    .B(_0141_));
 sg13g2_o21ai_1 _0608_ (.B1(_0142_),
    .Y(_0143_),
    .A1(_0126_),
    .A2(_0129_));
 sg13g2_nand2b_1 _0609_ (.Y(_0144_),
    .B(_0134_),
    .A_N(_0143_));
 sg13g2_nand2_1 _0610_ (.Y(_0145_),
    .A(net167),
    .B(net171));
 sg13g2_xor2_1 _0611_ (.B(net171),
    .A(net167),
    .X(_0146_));
 sg13g2_nand2_1 _0612_ (.Y(_0147_),
    .A(net148),
    .B(_0146_));
 sg13g2_xnor2_1 _0613_ (.Y(_0148_),
    .A(net147),
    .B(_0146_));
 sg13g2_nand3_1 _0614_ (.B(_0137_),
    .C(_0148_),
    .A(_0135_),
    .Y(_0149_));
 sg13g2_o21ai_1 _0615_ (.B1(_0149_),
    .Y(_0150_),
    .A1(_0138_),
    .A2(_0141_));
 sg13g2_nand2b_1 _0616_ (.Y(_0151_),
    .B(_0144_),
    .A_N(_0150_));
 sg13g2_a21oi_1 _0617_ (.A1(_0135_),
    .A2(_0137_),
    .Y(_0152_),
    .B1(_0148_));
 sg13g2_xnor2_1 _0618_ (.Y(_0153_),
    .A(net146),
    .B(_0118_));
 sg13g2_a21oi_1 _0619_ (.A1(_0145_),
    .A2(_0147_),
    .Y(_0154_),
    .B1(_0153_));
 sg13g2_nor2_1 _0620_ (.A(_0152_),
    .B(_0154_),
    .Y(_0155_));
 sg13g2_nand3_1 _0621_ (.B(_0147_),
    .C(_0153_),
    .A(_0145_),
    .Y(_0156_));
 sg13g2_o21ai_1 _0622_ (.B1(_0156_),
    .Y(_0157_),
    .A1(_0119_),
    .A2(_0122_));
 sg13g2_a21oi_1 _0623_ (.A1(_0151_),
    .A2(_0155_),
    .Y(_0158_),
    .B1(_0157_));
 sg13g2_a21oi_1 _0624_ (.A1(_0119_),
    .A2(_0122_),
    .Y(_0159_),
    .B1(_0158_));
 sg13g2_o21ai_1 _0625_ (.B1(_0079_),
    .Y(_0160_),
    .A1(_0445_),
    .A2(_0080_));
 sg13g2_xnor2_1 _0626_ (.Y(_0161_),
    .A(\counter[8] ),
    .B(\counter[7] ));
 sg13g2_xor2_1 _0627_ (.B(_0005_),
    .A(net156),
    .X(_0162_));
 sg13g2_xnor2_1 _0628_ (.Y(_0163_),
    .A(_0161_),
    .B(_0162_));
 sg13g2_xor2_1 _0629_ (.B(\hvsync_gen.vpos[7] ),
    .A(\counter[7] ),
    .X(_0164_));
 sg13g2_a21oi_1 _0630_ (.A1(net144),
    .A2(_0121_),
    .Y(_0165_),
    .B1(_0120_));
 sg13g2_o21ai_1 _0631_ (.B1(net168),
    .Y(_0166_),
    .A1(net170),
    .A2(net158));
 sg13g2_nand2b_1 _0632_ (.Y(_0167_),
    .B(_0166_),
    .A_N(_0077_));
 sg13g2_xnor2_1 _0633_ (.Y(_0168_),
    .A(_0164_),
    .B(_0167_));
 sg13g2_xnor2_1 _0634_ (.Y(_0169_),
    .A(_0163_),
    .B(_0168_));
 sg13g2_xnor2_1 _0635_ (.Y(_0170_),
    .A(_0165_),
    .B(_0169_));
 sg13g2_xnor2_1 _0636_ (.Y(_0171_),
    .A(_0160_),
    .B(_0170_));
 sg13g2_xor2_1 _0637_ (.B(_0171_),
    .A(_0159_),
    .X(_0172_));
 sg13g2_xnor2_1 _0638_ (.Y(_0173_),
    .A(net162),
    .B(\hvsync_gen.vpos[0] ));
 sg13g2_o21ai_1 _0639_ (.B1(_0173_),
    .Y(_0174_),
    .A1(_0116_),
    .A2(_0172_));
 sg13g2_a21oi_2 _0640_ (.B1(_0174_),
    .Y(_0175_),
    .A2(_0172_),
    .A1(_0116_));
 sg13g2_nand2_1 _0641_ (.Y(_0176_),
    .A(net166),
    .B(net146));
 sg13g2_nand3b_1 _0642_ (.B(net155),
    .C(net183),
    .Y(_0177_),
    .A_N(_0131_));
 sg13g2_a22oi_1 _0643_ (.Y(_0178_),
    .B1(net152),
    .B2(net174),
    .A2(net153),
    .A1(net181));
 sg13g2_o21ai_1 _0644_ (.B1(_0127_),
    .Y(_0179_),
    .A1(\counter[4] ),
    .A2(net150));
 sg13g2_a21oi_1 _0645_ (.A1(_0177_),
    .A2(_0178_),
    .Y(_0180_),
    .B1(_0179_));
 sg13g2_a221oi_1 _0646_ (.B2(net169),
    .C1(_0180_),
    .B1(net148),
    .A1(net170),
    .Y(_0181_),
    .A2(net149));
 sg13g2_or2_1 _0647_ (.X(_0182_),
    .B(net147),
    .A(net169));
 sg13g2_o21ai_1 _0648_ (.B1(_0182_),
    .Y(_0183_),
    .A1(net166),
    .A2(net146));
 sg13g2_o21ai_1 _0649_ (.B1(_0176_),
    .Y(_0184_),
    .A1(_0181_),
    .A2(_0183_));
 sg13g2_a21oi_1 _0650_ (.A1(_0082_),
    .A2(_0086_),
    .Y(_0185_),
    .B1(_0085_));
 sg13g2_nor2_1 _0651_ (.A(_0065_),
    .B(_0069_),
    .Y(_0186_));
 sg13g2_o21ai_1 _0652_ (.B1(_0186_),
    .Y(_0187_),
    .A1(_0066_),
    .A2(_0185_));
 sg13g2_o21ai_1 _0653_ (.B1(_0187_),
    .Y(_0188_),
    .A1(net173),
    .A2(\hvsync_gen.hpos[5] ));
 sg13g2_xnor2_1 _0654_ (.Y(_0189_),
    .A(\counter[7] ),
    .B(net170));
 sg13g2_xnor2_1 _0655_ (.Y(_0190_),
    .A(net158),
    .B(net144));
 sg13g2_xnor2_1 _0656_ (.Y(_0191_),
    .A(_0189_),
    .B(_0190_));
 sg13g2_xnor2_1 _0657_ (.Y(_0192_),
    .A(_0188_),
    .B(_0191_));
 sg13g2_xnor2_1 _0658_ (.Y(_0193_),
    .A(_0184_),
    .B(_0192_));
 sg13g2_a21oi_2 _0659_ (.B1(_0175_),
    .Y(_0194_),
    .A2(_0193_),
    .A1(_0053_));
 sg13g2_nand2b_1 _0660_ (.Y(_0195_),
    .B(net164),
    .A_N(net153));
 sg13g2_nand2b_1 _0661_ (.Y(_0196_),
    .B(net153),
    .A_N(net164));
 sg13g2_and2_1 _0662_ (.A(_0195_),
    .B(_0196_),
    .X(_0197_));
 sg13g2_nand2_2 _0663_ (.Y(_0198_),
    .A(\counter[9] ),
    .B(\counter[8] ));
 sg13g2_nor2_1 _0664_ (.A(net172),
    .B(_0198_),
    .Y(_0199_));
 sg13g2_a21o_1 _0665_ (.A2(_0198_),
    .A1(_0008_),
    .B1(_0199_),
    .X(_0200_));
 sg13g2_a21oi_2 _0666_ (.B1(_0199_),
    .Y(_0201_),
    .A2(_0198_),
    .A1(_0008_));
 sg13g2_a21oi_1 _0667_ (.A1(_0005_),
    .A2(_0198_),
    .Y(_0202_),
    .B1(_0004_));
 sg13g2_and3_1 _0668_ (.X(_0203_),
    .A(\counter[7] ),
    .B(_0445_),
    .C(_0198_));
 sg13g2_nor2_1 _0669_ (.A(_0202_),
    .B(_0203_),
    .Y(_0204_));
 sg13g2_nor2b_1 _0670_ (.A(\counter[9] ),
    .B_N(\counter[8] ),
    .Y(_0205_));
 sg13g2_nand2_1 _0671_ (.Y(_0206_),
    .A(_0006_),
    .B(_0205_));
 sg13g2_nand2_1 _0672_ (.Y(_0207_),
    .A(\counter[9] ),
    .B(_0443_));
 sg13g2_o21ai_1 _0673_ (.B1(_0206_),
    .Y(_0208_),
    .A1(_0006_),
    .A2(_0207_));
 sg13g2_nand2b_2 _0674_ (.Y(_0209_),
    .B(_0208_),
    .A_N(_0204_));
 sg13g2_inv_1 _0675_ (.Y(_0210_),
    .A(_0209_));
 sg13g2_o21ai_1 _0676_ (.B1(_0205_),
    .Y(_0211_),
    .A1(_0202_),
    .A2(_0203_));
 sg13g2_and3_1 _0677_ (.X(_0212_),
    .A(_0004_),
    .B(_0207_),
    .C(_0211_));
 sg13g2_a21oi_1 _0678_ (.A1(_0207_),
    .A2(_0211_),
    .Y(_0213_),
    .B1(_0444_));
 sg13g2_or2_1 _0679_ (.X(_0214_),
    .B(_0213_),
    .A(_0212_));
 sg13g2_nor3_2 _0680_ (.A(_0005_),
    .B(_0212_),
    .C(_0213_),
    .Y(_0215_));
 sg13g2_or2_1 _0681_ (.X(_0216_),
    .B(_0214_),
    .A(_0005_));
 sg13g2_a21oi_2 _0682_ (.B1(_0006_),
    .Y(_0217_),
    .A2(\counter[8] ),
    .A1(\counter[9] ));
 sg13g2_a21o_1 _0683_ (.A2(_0211_),
    .A1(_0207_),
    .B1(_0204_),
    .X(_0218_));
 sg13g2_xor2_1 _0684_ (.B(_0218_),
    .A(_0217_),
    .X(_0219_));
 sg13g2_xnor2_1 _0685_ (.Y(_0220_),
    .A(_0217_),
    .B(_0218_));
 sg13g2_nor3_2 _0686_ (.A(_0210_),
    .B(_0215_),
    .C(_0220_),
    .Y(_0221_));
 sg13g2_xnor2_1 _0687_ (.Y(_0222_),
    .A(_0050_),
    .B(_0221_));
 sg13g2_xnor2_1 _0688_ (.Y(_0223_),
    .A(_0005_),
    .B(_0221_));
 sg13g2_nand2_1 _0689_ (.Y(_0224_),
    .A(_0051_),
    .B(_0222_));
 sg13g2_o21ai_1 _0690_ (.B1(_0214_),
    .Y(_0225_),
    .A1(_0005_),
    .A2(_0221_));
 sg13g2_a22oi_1 _0691_ (.Y(_0226_),
    .B1(_0225_),
    .B2(_0216_),
    .A2(_0222_),
    .A1(_0051_));
 sg13g2_nand2_1 _0692_ (.Y(_0227_),
    .A(_0215_),
    .B(_0220_));
 sg13g2_nand2_1 _0693_ (.Y(_0228_),
    .A(_0209_),
    .B(_0227_));
 sg13g2_a221oi_1 _0694_ (.B2(_0216_),
    .C1(_0228_),
    .B1(_0225_),
    .A1(_0051_),
    .Y(_0229_),
    .A2(_0222_));
 sg13g2_xnor2_1 _0695_ (.Y(_0230_),
    .A(_0051_),
    .B(_0229_));
 sg13g2_inv_1 _0696_ (.Y(_0231_),
    .A(_0230_));
 sg13g2_nand2_1 _0697_ (.Y(_0232_),
    .A(_0201_),
    .B(_0230_));
 sg13g2_o21ai_1 _0698_ (.B1(_0223_),
    .Y(_0233_),
    .A1(_0007_),
    .A2(_0229_));
 sg13g2_a22oi_1 _0699_ (.Y(_0234_),
    .B1(_0233_),
    .B2(_0224_),
    .A2(_0230_),
    .A1(_0201_));
 sg13g2_nor4_1 _0700_ (.A(_0050_),
    .B(_0007_),
    .C(_0214_),
    .D(_0221_),
    .Y(_0235_));
 sg13g2_a21oi_1 _0701_ (.A1(_0215_),
    .A2(_0220_),
    .Y(_0236_),
    .B1(_0235_));
 sg13g2_nand2_1 _0702_ (.Y(_0237_),
    .A(_0209_),
    .B(_0236_));
 sg13g2_a221oi_1 _0703_ (.B2(_0224_),
    .C1(_0237_),
    .B1(_0233_),
    .A1(_0201_),
    .Y(_0238_),
    .A2(_0230_));
 sg13g2_xnor2_1 _0704_ (.Y(_0239_),
    .A(_0201_),
    .B(_0238_));
 sg13g2_nand2_1 _0705_ (.Y(_0240_),
    .A(net175),
    .B(_0239_));
 sg13g2_o21ai_1 _0706_ (.B1(_0231_),
    .Y(_0241_),
    .A1(_0200_),
    .A2(_0238_));
 sg13g2_a21oi_1 _0707_ (.A1(_0216_),
    .A2(_0219_),
    .Y(_0242_),
    .B1(_0226_));
 sg13g2_o21ai_1 _0708_ (.B1(_0236_),
    .Y(_0243_),
    .A1(_0209_),
    .A2(_0242_));
 sg13g2_nand2b_1 _0709_ (.Y(_0244_),
    .B(_0234_),
    .A_N(_0243_));
 sg13g2_a21oi_1 _0710_ (.A1(_0216_),
    .A2(_0219_),
    .Y(_0245_),
    .B1(_0209_));
 sg13g2_inv_1 _0711_ (.Y(_0246_),
    .A(_0245_));
 sg13g2_a21oi_1 _0712_ (.A1(_0226_),
    .A2(_0227_),
    .Y(_0247_),
    .B1(_0246_));
 sg13g2_a221oi_1 _0713_ (.B2(_0224_),
    .C1(_0246_),
    .B1(_0233_),
    .A1(_0201_),
    .Y(_0248_),
    .A2(_0230_));
 sg13g2_nor4_1 _0714_ (.A(_0051_),
    .B(_0200_),
    .C(_0223_),
    .D(_0229_),
    .Y(_0249_));
 sg13g2_or3_1 _0715_ (.A(_0243_),
    .B(_0248_),
    .C(_0249_),
    .X(_0250_));
 sg13g2_a221oi_1 _0716_ (.B2(_0247_),
    .C1(_0250_),
    .B1(_0244_),
    .A1(_0232_),
    .Y(_0251_),
    .A2(_0241_));
 sg13g2_nand2_1 _0717_ (.Y(_0252_),
    .A(_0240_),
    .B(_0251_));
 sg13g2_a21o_1 _0718_ (.A2(_0251_),
    .A1(_0240_),
    .B1(_0447_),
    .X(_0253_));
 sg13g2_nand2b_1 _0719_ (.Y(_0254_),
    .B(_0253_),
    .A_N(_0239_));
 sg13g2_and2_1 _0720_ (.A(_0240_),
    .B(_0254_),
    .X(_0255_));
 sg13g2_nand2_1 _0721_ (.Y(_0256_),
    .A(_0447_),
    .B(_0251_));
 sg13g2_nand3_1 _0722_ (.B(_0253_),
    .C(_0256_),
    .A(_0052_),
    .Y(_0257_));
 sg13g2_or2_1 _0723_ (.X(_0258_),
    .B(_0012_),
    .A(net180));
 sg13g2_a21oi_1 _0724_ (.A1(_0253_),
    .A2(_0256_),
    .Y(_0259_),
    .B1(_0123_));
 sg13g2_a221oi_1 _0725_ (.B2(_0011_),
    .C1(_0259_),
    .B1(_0258_),
    .A1(_0013_),
    .Y(_0260_),
    .A2(_0257_));
 sg13g2_a21o_1 _0726_ (.A2(_0256_),
    .A1(_0253_),
    .B1(_0124_),
    .X(_0261_));
 sg13g2_nand2_1 _0727_ (.Y(_0262_),
    .A(net180),
    .B(_0012_));
 sg13g2_nand3_1 _0728_ (.B(_0256_),
    .C(_0262_),
    .A(_0253_),
    .Y(_0263_));
 sg13g2_nand3_1 _0729_ (.B(_0261_),
    .C(_0263_),
    .A(_0011_),
    .Y(_0264_));
 sg13g2_o21ai_1 _0730_ (.B1(_0264_),
    .Y(_0265_),
    .A1(_0255_),
    .A2(_0260_));
 sg13g2_a221oi_1 _0731_ (.B2(_0247_),
    .C1(_0250_),
    .B1(_0244_),
    .A1(net175),
    .Y(_0266_),
    .A2(_0239_));
 sg13g2_or2_1 _0732_ (.X(_0267_),
    .B(_0266_),
    .A(_0251_));
 sg13g2_xnor2_1 _0733_ (.Y(_0268_),
    .A(_0009_),
    .B(_0238_));
 sg13g2_a21oi_1 _0734_ (.A1(_0013_),
    .A2(_0011_),
    .Y(_0269_),
    .B1(_0268_));
 sg13g2_o21ai_1 _0735_ (.B1(_0269_),
    .Y(_0270_),
    .A1(net152),
    .A2(_0252_));
 sg13g2_a221oi_1 _0736_ (.B2(_0267_),
    .C1(_0270_),
    .B1(_0265_),
    .A1(net152),
    .Y(_0271_),
    .A2(_0252_));
 sg13g2_nor2_1 _0737_ (.A(_0010_),
    .B(_0268_),
    .Y(_0272_));
 sg13g2_nand2_1 _0738_ (.Y(_0273_),
    .A(_0252_),
    .B(_0272_));
 sg13g2_o21ai_1 _0739_ (.B1(_0273_),
    .Y(_0274_),
    .A1(_0009_),
    .A2(_0238_));
 sg13g2_o21ai_1 _0740_ (.B1(\counter[1] ),
    .Y(_0275_),
    .A1(net179),
    .A2(net162));
 sg13g2_nand2b_1 _0741_ (.Y(_0276_),
    .B(net164),
    .A_N(_0275_));
 sg13g2_a22oi_1 _0742_ (.Y(_0277_),
    .B1(\hvsync_gen.hpos[2] ),
    .B2(net175),
    .A2(net163),
    .A1(net180));
 sg13g2_or2_1 _0743_ (.X(_0278_),
    .B(net161),
    .A(net172));
 sg13g2_o21ai_1 _0744_ (.B1(_0278_),
    .Y(_0279_),
    .A1(net175),
    .A2(\hvsync_gen.hpos[2] ));
 sg13g2_a21oi_1 _0745_ (.A1(_0276_),
    .A2(_0277_),
    .Y(_0280_),
    .B1(_0279_));
 sg13g2_a21oi_1 _0746_ (.A1(net172),
    .A2(net161),
    .Y(_0281_),
    .B1(_0280_));
 sg13g2_xnor2_1 _0747_ (.Y(_0282_),
    .A(net168),
    .B(net160));
 sg13g2_xnor2_1 _0748_ (.Y(_0283_),
    .A(_0003_),
    .B(_0282_));
 sg13g2_xnor2_1 _0749_ (.Y(_0284_),
    .A(_0281_),
    .B(_0283_));
 sg13g2_xnor2_1 _0750_ (.Y(_0285_),
    .A(_0229_),
    .B(_0284_));
 sg13g2_o21ai_1 _0751_ (.B1(_0285_),
    .Y(_0286_),
    .A1(_0271_),
    .A2(_0274_));
 sg13g2_or3_2 _0752_ (.A(_0271_),
    .B(_0274_),
    .C(_0285_),
    .X(_0287_));
 sg13g2_a21o_1 _0753_ (.A2(_0287_),
    .A1(_0286_),
    .B1(_0197_),
    .X(_0288_));
 sg13g2_nor2_1 _0754_ (.A(net168),
    .B(net150),
    .Y(_0289_));
 sg13g2_o21ai_1 _0755_ (.B1(net181),
    .Y(_0290_),
    .A1(net173),
    .A2(net154));
 sg13g2_a22oi_1 _0756_ (.Y(_0291_),
    .B1(net151),
    .B2(net171),
    .A2(net154),
    .A1(net173));
 sg13g2_o21ai_1 _0757_ (.B1(_0291_),
    .Y(_0292_),
    .A1(_0449_),
    .A2(_0290_));
 sg13g2_o21ai_1 _0758_ (.B1(_0292_),
    .Y(_0293_),
    .A1(net170),
    .A2(net151));
 sg13g2_a22oi_1 _0759_ (.Y(_0294_),
    .B1(net147),
    .B2(net166),
    .A2(net149),
    .A1(net168));
 sg13g2_o21ai_1 _0760_ (.B1(_0294_),
    .Y(_0295_),
    .A1(_0289_),
    .A2(_0293_));
 sg13g2_o21ai_1 _0761_ (.B1(_0295_),
    .Y(_0296_),
    .A1(net166),
    .A2(net148));
 sg13g2_nand3b_1 _0762_ (.B(net162),
    .C(net184),
    .Y(_0297_),
    .A_N(_0098_));
 sg13g2_a22oi_1 _0763_ (.Y(_0298_),
    .B1(\hvsync_gen.hpos[2] ),
    .B2(\counter[1] ),
    .A2(net161),
    .A1(net179));
 sg13g2_or2_1 _0764_ (.X(_0299_),
    .B(net160),
    .A(net175));
 sg13g2_o21ai_1 _0765_ (.B1(_0299_),
    .Y(_0300_),
    .A1(net179),
    .A2(net161));
 sg13g2_a21oi_1 _0766_ (.A1(_0297_),
    .A2(_0298_),
    .Y(_0301_),
    .B1(_0300_));
 sg13g2_a21o_1 _0767_ (.A2(net160),
    .A1(net176),
    .B1(_0301_),
    .X(_0302_));
 sg13g2_xor2_1 _0768_ (.B(net146),
    .A(net159),
    .X(_0303_));
 sg13g2_xnor2_1 _0769_ (.Y(_0304_),
    .A(_0189_),
    .B(_0303_));
 sg13g2_xnor2_1 _0770_ (.Y(_0305_),
    .A(_0296_),
    .B(_0304_));
 sg13g2_or2_1 _0771_ (.X(_0306_),
    .B(_0305_),
    .A(_0302_));
 sg13g2_nand2_1 _0772_ (.Y(_0307_),
    .A(_0302_),
    .B(_0305_));
 sg13g2_and2_1 _0773_ (.A(_0306_),
    .B(_0307_),
    .X(_0308_));
 sg13g2_xor2_1 _0774_ (.B(net6),
    .A(net3),
    .X(_0309_));
 sg13g2_a221oi_1 _0775_ (.B2(_0287_),
    .C1(_0309_),
    .B1(_0286_),
    .A1(_0195_),
    .Y(_0310_),
    .A2(_0196_));
 sg13g2_a221oi_1 _0776_ (.B2(_0307_),
    .C1(_0310_),
    .B1(_0306_),
    .A1(_0053_),
    .Y(_0311_),
    .A2(_0288_));
 sg13g2_a21o_1 _0777_ (.A2(_0308_),
    .A1(net3),
    .B1(_0193_),
    .X(_0312_));
 sg13g2_o21ai_1 _0778_ (.B1(_0194_),
    .Y(_0313_),
    .A1(_0311_),
    .A2(_0312_));
 sg13g2_nor2_1 _0779_ (.A(net168),
    .B(net144),
    .Y(_0314_));
 sg13g2_a22oi_1 _0780_ (.Y(_0315_),
    .B1(net152),
    .B2(net183),
    .A2(net153),
    .A1(net184));
 sg13g2_or2_1 _0781_ (.X(_0316_),
    .B(net149),
    .A(net178));
 sg13g2_o21ai_1 _0782_ (.B1(_0316_),
    .Y(_0317_),
    .A1(net183),
    .A2(net151));
 sg13g2_a22oi_1 _0783_ (.Y(_0318_),
    .B1(net148),
    .B2(net173),
    .A2(net149),
    .A1(net178));
 sg13g2_o21ai_1 _0784_ (.B1(_0318_),
    .Y(_0319_),
    .A1(_0315_),
    .A2(_0317_));
 sg13g2_a22oi_1 _0785_ (.Y(_0320_),
    .B1(_0046_),
    .B2(_0447_),
    .A2(_0450_),
    .A1(_0446_));
 sg13g2_a22oi_1 _0786_ (.Y(_0321_),
    .B1(_0319_),
    .B2(_0320_),
    .A2(net145),
    .A1(net170));
 sg13g2_a22oi_1 _0787_ (.Y(_0322_),
    .B1(net144),
    .B2(net168),
    .A2(\hvsync_gen.vpos[7] ),
    .A1(net165));
 sg13g2_o21ai_1 _0788_ (.B1(_0322_),
    .Y(_0323_),
    .A1(_0314_),
    .A2(_0321_));
 sg13g2_o21ai_1 _0789_ (.B1(_0323_),
    .Y(_0324_),
    .A1(net165),
    .A2(\hvsync_gen.vpos[7] ));
 sg13g2_or2_1 _0790_ (.X(_0325_),
    .B(net159),
    .A(net183));
 sg13g2_nand3_1 _0791_ (.B(net160),
    .C(_0325_),
    .A(net184),
    .Y(_0326_));
 sg13g2_a22oi_1 _0792_ (.Y(_0327_),
    .B1(net157),
    .B2(net178),
    .A2(\hvsync_gen.hpos[5] ),
    .A1(net183));
 sg13g2_or2_1 _0793_ (.X(_0328_),
    .B(net158),
    .A(net181));
 sg13g2_o21ai_1 _0794_ (.B1(_0328_),
    .Y(_0329_),
    .A1(net173),
    .A2(net156));
 sg13g2_a21oi_1 _0795_ (.A1(_0326_),
    .A2(_0327_),
    .Y(_0330_),
    .B1(_0329_));
 sg13g2_a21oi_1 _0796_ (.A1(net173),
    .A2(net156),
    .Y(_0331_),
    .B1(_0330_));
 sg13g2_xnor2_1 _0797_ (.Y(_0332_),
    .A(\hvsync_gen.hpos[8] ),
    .B(\hvsync_gen.vpos[8] ));
 sg13g2_xnor2_1 _0798_ (.Y(_0333_),
    .A(_0189_),
    .B(_0332_));
 sg13g2_xnor2_1 _0799_ (.Y(_0334_),
    .A(_0331_),
    .B(_0333_));
 sg13g2_xnor2_1 _0800_ (.Y(_0335_),
    .A(_0324_),
    .B(_0334_));
 sg13g2_nor2_1 _0801_ (.A(_0197_),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_a21oi_1 _0802_ (.A1(_0049_),
    .A2(net142),
    .Y(_0337_),
    .B1(net143));
 sg13g2_nor2_1 _0803_ (.A(net156),
    .B(\hvsync_gen.hpos[8] ),
    .Y(_0338_));
 sg13g2_and3_1 _0804_ (.X(_0339_),
    .A(net145),
    .B(net75),
    .C(_0057_));
 sg13g2_nor2_1 _0805_ (.A(\hvsync_gen.vpos[9] ),
    .B(_0339_),
    .Y(_0340_));
 sg13g2_o21ai_1 _0806_ (.B1(_0340_),
    .Y(_0341_),
    .A1(_0002_),
    .A2(_0338_));
 sg13g2_a221oi_1 _0807_ (.B2(_0313_),
    .C1(_0341_),
    .B1(_0337_),
    .A1(_0049_),
    .Y(uo_out[6]),
    .A2(_0336_));
 sg13g2_a21o_1 _0808_ (.A2(net143),
    .A1(net7),
    .B1(_0341_),
    .X(_0342_));
 sg13g2_and2_1 _0809_ (.A(_0049_),
    .B(_0193_),
    .X(_0343_));
 sg13g2_nor2_1 _0810_ (.A(net8),
    .B(_0193_),
    .Y(_0344_));
 sg13g2_or3_1 _0811_ (.A(net142),
    .B(_0343_),
    .C(_0344_),
    .X(_0345_));
 sg13g2_a21oi_1 _0812_ (.A1(net142),
    .A2(_0309_),
    .Y(_0346_),
    .B1(net143));
 sg13g2_a21oi_1 _0813_ (.A1(_0345_),
    .A2(_0346_),
    .Y(uo_out[2]),
    .B1(_0342_));
 sg13g2_xor2_1 _0814_ (.B(net5),
    .A(net2),
    .X(_0347_));
 sg13g2_a221oi_1 _0815_ (.B2(_0287_),
    .C1(_0347_),
    .B1(_0286_),
    .A1(_0195_),
    .Y(_0348_),
    .A2(_0196_));
 sg13g2_a221oi_1 _0816_ (.B2(_0307_),
    .C1(_0348_),
    .B1(_0306_),
    .A1(_0053_),
    .Y(_0349_),
    .A2(_0288_));
 sg13g2_a21o_1 _0817_ (.A2(_0308_),
    .A1(net2),
    .B1(_0193_),
    .X(_0350_));
 sg13g2_o21ai_1 _0818_ (.B1(_0194_),
    .Y(_0351_),
    .A1(_0349_),
    .A2(_0350_));
 sg13g2_a21oi_1 _0819_ (.A1(_0054_),
    .A2(net142),
    .Y(_0352_),
    .B1(_0336_));
 sg13g2_a221oi_1 _0820_ (.B2(_0352_),
    .C1(_0341_),
    .B1(_0351_),
    .A1(_0054_),
    .Y(uo_out[5]),
    .A2(net143));
 sg13g2_a21oi_1 _0821_ (.A1(_0054_),
    .A2(_0193_),
    .Y(_0353_),
    .B1(_0344_));
 sg13g2_mux2_1 _0822_ (.A0(_0353_),
    .A1(_0347_),
    .S(net142),
    .X(_0354_));
 sg13g2_nor2_1 _0823_ (.A(net143),
    .B(_0354_),
    .Y(_0355_));
 sg13g2_nor2_1 _0824_ (.A(_0342_),
    .B(_0355_),
    .Y(uo_out[1]));
 sg13g2_xnor2_1 _0825_ (.Y(_0356_),
    .A(net1),
    .B(net4));
 sg13g2_a221oi_1 _0826_ (.B2(_0287_),
    .C1(_0356_),
    .B1(_0286_),
    .A1(_0195_),
    .Y(_0357_),
    .A2(_0196_));
 sg13g2_a221oi_1 _0827_ (.B2(_0307_),
    .C1(_0357_),
    .B1(_0306_),
    .A1(_0053_),
    .Y(_0358_),
    .A2(_0288_));
 sg13g2_a21o_1 _0828_ (.A2(_0308_),
    .A1(_0055_),
    .B1(_0193_),
    .X(_0359_));
 sg13g2_o21ai_1 _0829_ (.B1(_0194_),
    .Y(_0360_),
    .A1(_0358_),
    .A2(_0359_));
 sg13g2_a21oi_1 _0830_ (.A1(net1),
    .A2(net142),
    .Y(_0361_),
    .B1(net143));
 sg13g2_a221oi_1 _0831_ (.B2(_0361_),
    .C1(_0341_),
    .B1(_0360_),
    .A1(net1),
    .Y(uo_out[4]),
    .A2(net143));
 sg13g2_nand2_1 _0832_ (.Y(_0362_),
    .A(net142),
    .B(_0356_));
 sg13g2_and2_1 _0833_ (.A(net1),
    .B(_0193_),
    .X(_0363_));
 sg13g2_nor3_1 _0834_ (.A(net142),
    .B(_0344_),
    .C(_0363_),
    .Y(_0364_));
 sg13g2_nor2_1 _0835_ (.A(net143),
    .B(_0364_),
    .Y(_0365_));
 sg13g2_a21oi_1 _0836_ (.A1(_0362_),
    .A2(_0365_),
    .Y(uo_out[0]),
    .B1(_0342_));
 sg13g2_nor3_1 _0837_ (.A(net145),
    .B(net147),
    .C(net144),
    .Y(_0366_));
 sg13g2_nand3b_1 _0838_ (.B(_0047_),
    .C(_0366_),
    .Y(_0367_),
    .A_N(\hvsync_gen.vpos[7] ));
 sg13g2_nor4_2 _0839_ (.A(net164),
    .B(net162),
    .C(net161),
    .Y(_0368_),
    .D(\hvsync_gen.hpos[2] ));
 sg13g2_nor2_1 _0840_ (.A(net154),
    .B(net155),
    .Y(_0369_));
 sg13g2_nor4_1 _0841_ (.A(\hvsync_gen.hpos[9] ),
    .B(net150),
    .C(net151),
    .D(\hvsync_gen.vpos[9] ),
    .Y(_0370_));
 sg13g2_nor2b_1 _0842_ (.A(_0060_),
    .B_N(_0370_),
    .Y(_0371_));
 sg13g2_nand4_1 _0843_ (.B(_0368_),
    .C(_0369_),
    .A(_0338_),
    .Y(_0372_),
    .D(_0371_));
 sg13g2_nor2_2 _0844_ (.A(_0367_),
    .B(_0372_),
    .Y(_0373_));
 sg13g2_o21ai_1 _0845_ (.B1(net187),
    .Y(_0374_),
    .A1(net185),
    .A2(_0373_));
 sg13g2_a21oi_1 _0846_ (.A1(_0448_),
    .A2(_0373_),
    .Y(_0016_),
    .B1(_0374_));
 sg13g2_a21oi_1 _0847_ (.A1(net184),
    .A2(_0373_),
    .Y(_0375_),
    .B1(net182));
 sg13g2_nor3_2 _0848_ (.A(_0099_),
    .B(_0367_),
    .C(_0372_),
    .Y(_0376_));
 sg13g2_nor3_1 _0849_ (.A(_0048_),
    .B(_0375_),
    .C(_0376_),
    .Y(_0017_));
 sg13g2_xnor2_1 _0850_ (.Y(_0377_),
    .A(net180),
    .B(_0376_));
 sg13g2_nor2_1 _0851_ (.A(_0048_),
    .B(_0377_),
    .Y(_0018_));
 sg13g2_and2_1 _0852_ (.A(_0052_),
    .B(_0376_),
    .X(_0378_));
 sg13g2_o21ai_1 _0853_ (.B1(net187),
    .Y(_0379_),
    .A1(net175),
    .A2(_0378_));
 sg13g2_a21oi_1 _0854_ (.A1(net175),
    .A2(_0378_),
    .Y(_0019_),
    .B1(_0379_));
 sg13g2_nor2b_1 _0855_ (.A(_0139_),
    .B_N(_0376_),
    .Y(_0380_));
 sg13g2_and2_1 _0856_ (.A(net171),
    .B(_0380_),
    .X(_0381_));
 sg13g2_o21ai_1 _0857_ (.B1(net186),
    .Y(_0382_),
    .A1(net171),
    .A2(_0380_));
 sg13g2_nor2_1 _0858_ (.A(_0381_),
    .B(_0382_),
    .Y(_0020_));
 sg13g2_nor2b_1 _0859_ (.A(_0008_),
    .B_N(_0380_),
    .Y(_0383_));
 sg13g2_o21ai_1 _0860_ (.B1(net186),
    .Y(_0384_),
    .A1(net167),
    .A2(_0383_));
 sg13g2_a21oi_1 _0861_ (.A1(net63),
    .A2(_0383_),
    .Y(_0021_),
    .B1(_0384_));
 sg13g2_a21oi_1 _0862_ (.A1(net167),
    .A2(_0381_),
    .Y(_0385_),
    .B1(net165));
 sg13g2_nand3_1 _0863_ (.B(net167),
    .C(_0381_),
    .A(net165),
    .Y(_0386_));
 sg13g2_nand2_1 _0864_ (.Y(_0387_),
    .A(net186),
    .B(_0386_));
 sg13g2_nor2_1 _0865_ (.A(_0385_),
    .B(_0387_),
    .Y(_0022_));
 sg13g2_and3_1 _0866_ (.X(_0388_),
    .A(net167),
    .B(_0050_),
    .C(_0381_));
 sg13g2_o21ai_1 _0867_ (.B1(net186),
    .Y(_0389_),
    .A1(net95),
    .A2(_0388_));
 sg13g2_a21oi_1 _0868_ (.A1(net95),
    .A2(_0388_),
    .Y(_0023_),
    .B1(_0389_));
 sg13g2_or2_1 _0869_ (.X(_0390_),
    .B(_0386_),
    .A(_0444_));
 sg13g2_o21ai_1 _0870_ (.B1(net186),
    .Y(_0391_),
    .A1(_0443_),
    .A2(_0390_));
 sg13g2_a21oi_1 _0871_ (.A1(_0443_),
    .A2(_0390_),
    .Y(_0024_),
    .B1(_0391_));
 sg13g2_nor2_1 _0872_ (.A(_0006_),
    .B(_0390_),
    .Y(_0392_));
 sg13g2_o21ai_1 _0873_ (.B1(net186),
    .Y(_0393_),
    .A1(net72),
    .A2(_0392_));
 sg13g2_a21oi_1 _0874_ (.A1(net72),
    .A2(_0392_),
    .Y(_0025_),
    .B1(_0393_));
 sg13g2_and3_1 _0875_ (.X(_0394_),
    .A(net164),
    .B(net162),
    .C(\hvsync_gen.hpos[2] ));
 sg13g2_and3_2 _0876_ (.X(_0395_),
    .A(net69),
    .B(net99),
    .C(_0394_));
 sg13g2_nor4_1 _0877_ (.A(net159),
    .B(net156),
    .C(net157),
    .D(_0059_),
    .Y(_0396_));
 sg13g2_nand2_1 _0878_ (.Y(_0397_),
    .A(_0395_),
    .B(_0396_));
 sg13g2_and2_2 _0879_ (.A(net187),
    .B(_0397_),
    .X(_0398_));
 sg13g2_nand2_2 _0880_ (.Y(_0399_),
    .A(net187),
    .B(_0397_));
 sg13g2_and2_1 _0881_ (.A(net57),
    .B(_0398_),
    .X(_0026_));
 sg13g2_o21ai_1 _0882_ (.B1(_0398_),
    .Y(_0400_),
    .A1(net164),
    .A2(net162));
 sg13g2_a21oi_1 _0883_ (.A1(net164),
    .A2(net162),
    .Y(_0027_),
    .B1(_0400_));
 sg13g2_a21oi_1 _0884_ (.A1(net164),
    .A2(net162),
    .Y(_0401_),
    .B1(net74));
 sg13g2_nor3_1 _0885_ (.A(_0048_),
    .B(_0394_),
    .C(net80),
    .Y(_0028_));
 sg13g2_o21ai_1 _0886_ (.B1(net187),
    .Y(_0402_),
    .A1(net69),
    .A2(_0394_));
 sg13g2_a21oi_1 _0887_ (.A1(net161),
    .A2(_0394_),
    .Y(_0029_),
    .B1(_0402_));
 sg13g2_a21oi_1 _0888_ (.A1(net69),
    .A2(_0394_),
    .Y(_0403_),
    .B1(net160));
 sg13g2_nor3_1 _0889_ (.A(_0048_),
    .B(_0395_),
    .C(net70),
    .Y(_0030_));
 sg13g2_and2_1 _0890_ (.A(net159),
    .B(_0395_),
    .X(_0404_));
 sg13g2_nor2_1 _0891_ (.A(net159),
    .B(_0395_),
    .Y(_0405_));
 sg13g2_nor3_1 _0892_ (.A(_0399_),
    .B(_0404_),
    .C(net100),
    .Y(_0031_));
 sg13g2_a21oi_1 _0893_ (.A1(net157),
    .A2(_0404_),
    .Y(_0406_),
    .B1(_0399_));
 sg13g2_o21ai_1 _0894_ (.B1(_0406_),
    .Y(_0407_),
    .A1(net157),
    .A2(_0404_));
 sg13g2_inv_1 _0895_ (.Y(_0032_),
    .A(_0407_));
 sg13g2_a21oi_1 _0896_ (.A1(net157),
    .A2(_0404_),
    .Y(_0408_),
    .B1(net156));
 sg13g2_and3_1 _0897_ (.X(_0409_),
    .A(net156),
    .B(net157),
    .C(_0404_));
 sg13g2_nor3_1 _0898_ (.A(_0399_),
    .B(net93),
    .C(_0409_),
    .Y(_0033_));
 sg13g2_nor2_1 _0899_ (.A(net77),
    .B(_0409_),
    .Y(_0410_));
 sg13g2_and2_1 _0900_ (.A(net77),
    .B(_0409_),
    .X(_0411_));
 sg13g2_nor3_1 _0901_ (.A(_0399_),
    .B(_0410_),
    .C(_0411_),
    .Y(_0034_));
 sg13g2_a21oi_1 _0902_ (.A1(net78),
    .A2(_0411_),
    .Y(_0412_),
    .B1(_0399_));
 sg13g2_o21ai_1 _0903_ (.B1(_0412_),
    .Y(_0413_),
    .A1(net78),
    .A2(_0411_));
 sg13g2_inv_1 _0904_ (.Y(_0035_),
    .A(_0413_));
 sg13g2_nand4_1 _0905_ (.B(net151),
    .C(\hvsync_gen.vpos[9] ),
    .A(net150),
    .Y(_0414_),
    .D(_0369_));
 sg13g2_o21ai_1 _0906_ (.B1(net186),
    .Y(_0415_),
    .A1(_0367_),
    .A2(_0414_));
 sg13g2_or2_2 _0907_ (.X(_0416_),
    .B(_0415_),
    .A(_0397_));
 sg13g2_inv_1 _0908_ (.Y(_0417_),
    .A(_0416_));
 sg13g2_a22oi_1 _0909_ (.Y(_0418_),
    .B1(_0417_),
    .B2(net65),
    .A2(_0398_),
    .A1(net155));
 sg13g2_inv_1 _0910_ (.Y(_0036_),
    .A(net66));
 sg13g2_nand2_1 _0911_ (.Y(_0419_),
    .A(net153),
    .B(_0398_));
 sg13g2_xnor2_1 _0912_ (.Y(_0420_),
    .A(net153),
    .B(net155));
 sg13g2_o21ai_1 _0913_ (.B1(_0419_),
    .Y(_0037_),
    .A1(_0416_),
    .A2(_0420_));
 sg13g2_nand3_1 _0914_ (.B(net155),
    .C(_0399_),
    .A(net154),
    .Y(_0421_));
 sg13g2_and2_2 _0915_ (.A(_0399_),
    .B(_0415_),
    .X(_0422_));
 sg13g2_xor2_1 _0916_ (.B(_0421_),
    .A(net151),
    .X(_0423_));
 sg13g2_nor2_1 _0917_ (.A(_0422_),
    .B(_0423_),
    .Y(_0038_));
 sg13g2_nand2_1 _0918_ (.Y(_0424_),
    .A(net149),
    .B(_0398_));
 sg13g2_nand3b_1 _0919_ (.B(net155),
    .C(net154),
    .Y(_0425_),
    .A_N(net103));
 sg13g2_xor2_1 _0920_ (.B(_0425_),
    .A(net149),
    .X(_0426_));
 sg13g2_o21ai_1 _0921_ (.B1(_0424_),
    .Y(_0039_),
    .A1(_0416_),
    .A2(_0426_));
 sg13g2_nand4_1 _0922_ (.B(net155),
    .C(net150),
    .A(net154),
    .Y(_0427_),
    .D(net151));
 sg13g2_nor2_1 _0923_ (.A(_0398_),
    .B(_0427_),
    .Y(_0428_));
 sg13g2_and2_1 _0924_ (.A(net147),
    .B(_0428_),
    .X(_0429_));
 sg13g2_nor2_1 _0925_ (.A(net147),
    .B(_0428_),
    .Y(_0430_));
 sg13g2_nor3_1 _0926_ (.A(_0422_),
    .B(_0429_),
    .C(_0430_),
    .Y(_0040_));
 sg13g2_nand2_1 _0927_ (.Y(_0431_),
    .A(net145),
    .B(_0398_));
 sg13g2_nor2_1 _0928_ (.A(net81),
    .B(_0427_),
    .Y(_0432_));
 sg13g2_xnor2_1 _0929_ (.Y(_0433_),
    .A(net145),
    .B(_0432_));
 sg13g2_o21ai_1 _0930_ (.B1(_0431_),
    .Y(_0041_),
    .A1(_0416_),
    .A2(net82));
 sg13g2_nand3_1 _0931_ (.B(net147),
    .C(net144),
    .A(net145),
    .Y(_0434_));
 sg13g2_nor3_1 _0932_ (.A(_0398_),
    .B(_0427_),
    .C(_0434_),
    .Y(_0435_));
 sg13g2_nor2_1 _0933_ (.A(_0422_),
    .B(_0435_),
    .Y(_0436_));
 sg13g2_a21oi_1 _0934_ (.A1(net145),
    .A2(_0429_),
    .Y(_0437_),
    .B1(net144));
 sg13g2_nor2b_1 _0935_ (.A(net85),
    .B_N(_0436_),
    .Y(_0042_));
 sg13g2_nor4_1 _0936_ (.A(net86),
    .B(_0416_),
    .C(_0427_),
    .D(_0434_),
    .Y(_0438_));
 sg13g2_a21o_1 _0937_ (.A2(_0436_),
    .A1(net86),
    .B1(_0438_),
    .X(_0043_));
 sg13g2_a21oi_1 _0938_ (.A1(_0339_),
    .A2(_0429_),
    .Y(_0439_),
    .B1(_0422_));
 sg13g2_nand3_1 _0939_ (.B(_0057_),
    .C(_0429_),
    .A(net145),
    .Y(_0440_));
 sg13g2_a221oi_1 _0940_ (.B2(_0047_),
    .C1(_0422_),
    .B1(_0440_),
    .A1(_0339_),
    .Y(_0044_),
    .A2(_0429_));
 sg13g2_nand2_1 _0941_ (.Y(_0441_),
    .A(net67),
    .B(_0439_));
 sg13g2_nand2_1 _0942_ (.Y(_0442_),
    .A(net186),
    .B(_0056_));
 sg13g2_o21ai_1 _0943_ (.B1(_0441_),
    .Y(_0045_),
    .A1(_0440_),
    .A2(_0442_));
 sg13g2_dfrbp_1 _0944_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net45),
    .D(net59),
    .Q_N(_0015_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _0945_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net30),
    .D(_0017_),
    .Q_N(_0467_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _0946_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net28),
    .D(_0018_),
    .Q_N(_0012_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _0947_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net26),
    .D(net91),
    .Q_N(_0466_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _0948_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net55),
    .D(_0020_),
    .Q_N(_0008_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _0949_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net53),
    .D(net64),
    .Q_N(_0007_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _0950_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net51),
    .D(_0022_),
    .Q_N(_0005_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _0951_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net49),
    .D(_0023_),
    .Q_N(_0004_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _0952_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net47),
    .D(_0024_),
    .Q_N(_0006_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _0953_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net44),
    .D(net73),
    .Q_N(_0465_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 _0954_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net42),
    .D(_0026_),
    .Q_N(_0014_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 _0955_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net41),
    .D(_0027_),
    .Q_N(_0464_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _0956_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net40),
    .D(_0028_),
    .Q_N(_0463_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _0957_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net39),
    .D(_0029_),
    .Q_N(_0462_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _0958_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net38),
    .D(net71),
    .Q_N(_0461_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _0959_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net37),
    .D(_0031_),
    .Q_N(_0460_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _0960_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net36),
    .D(_0032_),
    .Q_N(_0459_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _0961_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net35),
    .D(_0033_),
    .Q_N(_0458_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _0962_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net34),
    .D(_0034_),
    .Q_N(_0457_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _0963_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net56),
    .D(_0035_),
    .Q_N(_0002_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _0964_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net33),
    .D(net62),
    .Q_N(_0456_),
    .Q(hsync));
 sg13g2_dfrbp_1 _0965_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net32),
    .D(_0036_),
    .Q_N(_0013_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _0966_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net29),
    .D(_0037_),
    .Q_N(_0011_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _0967_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net25),
    .D(_0038_),
    .Q_N(_0010_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _0968_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net52),
    .D(_0039_),
    .Q_N(_0009_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _0969_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net48),
    .D(_0040_),
    .Q_N(_0003_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _0970_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net43),
    .D(net83),
    .Q_N(_0455_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _0971_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net27),
    .D(_0042_),
    .Q_N(_0454_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _0972_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net50),
    .D(_0043_),
    .Q_N(_0453_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _0973_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net31),
    .D(net76),
    .Q_N(_0452_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _0974_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net54),
    .D(net68),
    .Q_N(_0468_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _0975_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net46),
    .D(net89),
    .Q_N(_0451_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_tiehi _0947__26 (.L_HI(net26));
 sg13g2_tiehi _0971__27 (.L_HI(net27));
 sg13g2_tiehi _0946__28 (.L_HI(net28));
 sg13g2_tiehi _0966__29 (.L_HI(net29));
 sg13g2_tiehi _0945__30 (.L_HI(net30));
 sg13g2_tiehi _0973__31 (.L_HI(net31));
 sg13g2_tiehi _0965__32 (.L_HI(net32));
 sg13g2_tiehi _0964__33 (.L_HI(net33));
 sg13g2_tiehi _0962__34 (.L_HI(net34));
 sg13g2_tiehi _0961__35 (.L_HI(net35));
 sg13g2_tiehi _0960__36 (.L_HI(net36));
 sg13g2_tiehi _0959__37 (.L_HI(net37));
 sg13g2_tiehi _0958__38 (.L_HI(net38));
 sg13g2_tiehi _0957__39 (.L_HI(net39));
 sg13g2_tiehi _0956__40 (.L_HI(net40));
 sg13g2_tiehi _0955__41 (.L_HI(net41));
 sg13g2_tiehi _0954__42 (.L_HI(net42));
 sg13g2_tiehi _0970__43 (.L_HI(net43));
 sg13g2_tiehi _0953__44 (.L_HI(net44));
 sg13g2_tiehi _0944__45 (.L_HI(net45));
 sg13g2_tiehi _0975__46 (.L_HI(net46));
 sg13g2_tiehi _0952__47 (.L_HI(net47));
 sg13g2_tiehi _0969__48 (.L_HI(net48));
 sg13g2_tiehi _0951__49 (.L_HI(net49));
 sg13g2_tiehi _0972__50 (.L_HI(net50));
 sg13g2_tiehi _0950__51 (.L_HI(net51));
 sg13g2_tiehi _0968__52 (.L_HI(net52));
 sg13g2_tiehi _0949__53 (.L_HI(net53));
 sg13g2_tiehi _0974__54 (.L_HI(net54));
 sg13g2_tiehi _0948__55 (.L_HI(net55));
 sg13g2_tiehi _0963__56 (.L_HI(net56));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_htfab_checkers_10 (.L_LO(net10));
 sg13g2_tielo tt_um_htfab_checkers_11 (.L_LO(net11));
 sg13g2_tielo tt_um_htfab_checkers_12 (.L_LO(net12));
 sg13g2_tielo tt_um_htfab_checkers_13 (.L_LO(net13));
 sg13g2_tielo tt_um_htfab_checkers_14 (.L_LO(net14));
 sg13g2_tielo tt_um_htfab_checkers_15 (.L_LO(net15));
 sg13g2_tielo tt_um_htfab_checkers_16 (.L_LO(net16));
 sg13g2_tielo tt_um_htfab_checkers_17 (.L_LO(net17));
 sg13g2_tielo tt_um_htfab_checkers_18 (.L_LO(net18));
 sg13g2_tielo tt_um_htfab_checkers_19 (.L_LO(net19));
 sg13g2_tielo tt_um_htfab_checkers_20 (.L_LO(net20));
 sg13g2_tielo tt_um_htfab_checkers_21 (.L_LO(net21));
 sg13g2_tielo tt_um_htfab_checkers_22 (.L_LO(net22));
 sg13g2_tielo tt_um_htfab_checkers_23 (.L_LO(net23));
 sg13g2_tielo tt_um_htfab_checkers_24 (.L_LO(net24));
 sg13g2_tiehi _0967__25 (.L_HI(net25));
 sg13g2_buf_1 _1024_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1025_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout142 (.A(_0175_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_0336_),
    .X(net143));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(net84));
 sg13g2_buf_2 fanout145 (.A(\hvsync_gen.vpos[5] ),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(\hvsync_gen.vpos[5] ),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(net88),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(\hvsync_gen.vpos[4] ),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(\hvsync_gen.vpos[3] ),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(net102),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(\hvsync_gen.vpos[2] ),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(net97),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(net104),
    .X(net155));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(net92));
 sg13g2_buf_2 fanout157 (.A(net101),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(\hvsync_gen.hpos[6] ),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(\hvsync_gen.hpos[5] ),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(\hvsync_gen.hpos[4] ),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(net69),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(net94),
    .X(net162));
 sg13g2_buf_1 fanout163 (.A(\hvsync_gen.hpos[1] ),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(net79),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(net96),
    .X(net165));
 sg13g2_buf_1 fanout166 (.A(\counter[6] ),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(net63),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(\counter[5] ),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(net171),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(\counter[4] ));
 sg13g2_buf_2 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(net177),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(net177),
    .X(net175));
 sg13g2_buf_1 fanout176 (.A(net177),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(\counter[3] ),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(net181),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(net180),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(net181),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(\counter[2] ),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(net183),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(\counter[1] ),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(net98),
    .X(net184));
 sg13g2_buf_1 fanout185 (.A(\counter[0] ),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(net187),
    .X(net186));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_htfab_checkers_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0014_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0015_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0016_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0002_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0064_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0000_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold7 (.A(\counter[5] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0021_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0013_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0418_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold11 (.A(\hvsync_gen.vpos[9] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0045_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold13 (.A(\hvsync_gen.hpos[3] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0403_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0030_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold16 (.A(\counter[9] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0025_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold18 (.A(\hvsync_gen.hpos[2] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold19 (.A(\hvsync_gen.vpos[8] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0044_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold21 (.A(\hvsync_gen.hpos[8] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold22 (.A(\hvsync_gen.hpos[9] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold23 (.A(\hvsync_gen.hpos[0] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0401_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0003_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0433_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0041_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold28 (.A(\hvsync_gen.vpos[6] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0437_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold30 (.A(\hvsync_gen.vpos[7] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold31 (.A(\counter[8] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold32 (.A(\hvsync_gen.vpos[4] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0001_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0012_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0019_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold36 (.A(\hvsync_gen.hpos[7] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0408_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold38 (.A(\hvsync_gen.hpos[1] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold39 (.A(\counter[7] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold40 (.A(\counter[6] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold41 (.A(\hvsync_gen.vpos[1] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold42 (.A(\counter[0] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold43 (.A(\hvsync_gen.hpos[4] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0405_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold45 (.A(\hvsync_gen.hpos[6] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold46 (.A(\hvsync_gen.vpos[2] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0010_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold48 (.A(\hvsync_gen.vpos[0] ),
    .X(net104));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_208 ();
 sg13g2_decap_8 FILLER_16_215 ();
 sg13g2_decap_8 FILLER_16_222 ();
 sg13g2_decap_8 FILLER_16_229 ();
 sg13g2_decap_8 FILLER_16_236 ();
 sg13g2_decap_8 FILLER_16_243 ();
 sg13g2_decap_8 FILLER_16_250 ();
 sg13g2_decap_8 FILLER_16_257 ();
 sg13g2_decap_8 FILLER_16_264 ();
 sg13g2_decap_8 FILLER_16_271 ();
 sg13g2_decap_8 FILLER_16_278 ();
 sg13g2_decap_8 FILLER_16_285 ();
 sg13g2_decap_8 FILLER_16_292 ();
 sg13g2_decap_8 FILLER_16_299 ();
 sg13g2_decap_8 FILLER_16_306 ();
 sg13g2_decap_8 FILLER_16_313 ();
 sg13g2_decap_8 FILLER_16_320 ();
 sg13g2_decap_8 FILLER_16_327 ();
 sg13g2_decap_8 FILLER_16_334 ();
 sg13g2_decap_8 FILLER_16_341 ();
 sg13g2_decap_8 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_355 ();
 sg13g2_decap_8 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_decap_8 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_fill_2 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_191 ();
 sg13g2_decap_4 FILLER_17_201 ();
 sg13g2_fill_2 FILLER_17_214 ();
 sg13g2_decap_8 FILLER_17_220 ();
 sg13g2_decap_4 FILLER_17_227 ();
 sg13g2_decap_8 FILLER_17_235 ();
 sg13g2_decap_4 FILLER_17_242 ();
 sg13g2_decap_8 FILLER_17_250 ();
 sg13g2_decap_8 FILLER_17_257 ();
 sg13g2_decap_8 FILLER_17_264 ();
 sg13g2_decap_8 FILLER_17_271 ();
 sg13g2_decap_8 FILLER_17_278 ();
 sg13g2_decap_8 FILLER_17_285 ();
 sg13g2_decap_8 FILLER_17_292 ();
 sg13g2_decap_8 FILLER_17_299 ();
 sg13g2_decap_8 FILLER_17_306 ();
 sg13g2_decap_8 FILLER_17_313 ();
 sg13g2_decap_8 FILLER_17_320 ();
 sg13g2_decap_8 FILLER_17_327 ();
 sg13g2_decap_8 FILLER_17_334 ();
 sg13g2_decap_8 FILLER_17_341 ();
 sg13g2_decap_8 FILLER_17_348 ();
 sg13g2_decap_8 FILLER_17_355 ();
 sg13g2_decap_8 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_4 FILLER_18_175 ();
 sg13g2_fill_2 FILLER_18_254 ();
 sg13g2_decap_8 FILLER_18_264 ();
 sg13g2_fill_2 FILLER_18_287 ();
 sg13g2_fill_2 FILLER_18_292 ();
 sg13g2_decap_8 FILLER_18_299 ();
 sg13g2_decap_8 FILLER_18_310 ();
 sg13g2_decap_4 FILLER_18_317 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_4 FILLER_19_182 ();
 sg13g2_fill_2 FILLER_19_195 ();
 sg13g2_fill_1 FILLER_19_197 ();
 sg13g2_fill_2 FILLER_19_233 ();
 sg13g2_fill_2 FILLER_19_245 ();
 sg13g2_fill_1 FILLER_19_252 ();
 sg13g2_fill_2 FILLER_19_267 ();
 sg13g2_fill_1 FILLER_19_269 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_4 FILLER_20_182 ();
 sg13g2_fill_1 FILLER_20_186 ();
 sg13g2_fill_1 FILLER_20_213 ();
 sg13g2_decap_4 FILLER_20_222 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_decap_4 FILLER_20_239 ();
 sg13g2_decap_8 FILLER_20_260 ();
 sg13g2_decap_8 FILLER_20_267 ();
 sg13g2_decap_8 FILLER_20_274 ();
 sg13g2_decap_8 FILLER_20_281 ();
 sg13g2_fill_1 FILLER_20_288 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_309 ();
 sg13g2_fill_1 FILLER_20_316 ();
 sg13g2_decap_8 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_345 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_decap_8 FILLER_20_366 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_fill_2 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_fill_2 FILLER_21_208 ();
 sg13g2_decap_4 FILLER_21_218 ();
 sg13g2_fill_1 FILLER_21_222 ();
 sg13g2_fill_2 FILLER_21_236 ();
 sg13g2_decap_4 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_256 ();
 sg13g2_decap_4 FILLER_21_289 ();
 sg13g2_decap_8 FILLER_21_341 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_decap_8 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_172 ();
 sg13g2_fill_1 FILLER_22_179 ();
 sg13g2_decap_4 FILLER_22_206 ();
 sg13g2_fill_2 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_244 ();
 sg13g2_decap_4 FILLER_22_251 ();
 sg13g2_fill_2 FILLER_22_255 ();
 sg13g2_decap_4 FILLER_22_262 ();
 sg13g2_fill_2 FILLER_22_298 ();
 sg13g2_fill_1 FILLER_22_300 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_fill_2 FILLER_23_140 ();
 sg13g2_fill_1 FILLER_23_142 ();
 sg13g2_decap_8 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_23_230 ();
 sg13g2_fill_1 FILLER_23_232 ();
 sg13g2_decap_4 FILLER_23_253 ();
 sg13g2_fill_2 FILLER_23_272 ();
 sg13g2_fill_1 FILLER_23_274 ();
 sg13g2_decap_8 FILLER_23_313 ();
 sg13g2_decap_8 FILLER_23_320 ();
 sg13g2_fill_2 FILLER_23_327 ();
 sg13g2_fill_1 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_346 ();
 sg13g2_fill_1 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_362 ();
 sg13g2_decap_8 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_376 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_4 FILLER_24_126 ();
 sg13g2_fill_2 FILLER_24_130 ();
 sg13g2_decap_4 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_146 ();
 sg13g2_fill_2 FILLER_24_159 ();
 sg13g2_fill_1 FILLER_24_187 ();
 sg13g2_decap_4 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_229 ();
 sg13g2_fill_2 FILLER_24_260 ();
 sg13g2_decap_8 FILLER_24_276 ();
 sg13g2_fill_2 FILLER_24_283 ();
 sg13g2_fill_1 FILLER_24_285 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_4 FILLER_24_308 ();
 sg13g2_fill_2 FILLER_24_333 ();
 sg13g2_fill_1 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_fill_1 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_119 ();
 sg13g2_fill_2 FILLER_25_161 ();
 sg13g2_fill_2 FILLER_25_168 ();
 sg13g2_fill_1 FILLER_25_170 ();
 sg13g2_fill_2 FILLER_25_181 ();
 sg13g2_fill_1 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_201 ();
 sg13g2_decap_8 FILLER_25_208 ();
 sg13g2_fill_2 FILLER_25_215 ();
 sg13g2_decap_4 FILLER_25_222 ();
 sg13g2_fill_1 FILLER_25_226 ();
 sg13g2_decap_4 FILLER_25_236 ();
 sg13g2_fill_1 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_255 ();
 sg13g2_fill_2 FILLER_25_266 ();
 sg13g2_fill_1 FILLER_25_268 ();
 sg13g2_decap_4 FILLER_25_274 ();
 sg13g2_fill_1 FILLER_25_278 ();
 sg13g2_decap_4 FILLER_25_310 ();
 sg13g2_fill_1 FILLER_25_331 ();
 sg13g2_decap_4 FILLER_25_350 ();
 sg13g2_fill_2 FILLER_25_354 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_4 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_fill_2 FILLER_26_126 ();
 sg13g2_fill_1 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_fill_2 FILLER_26_163 ();
 sg13g2_fill_1 FILLER_26_165 ();
 sg13g2_fill_2 FILLER_26_212 ();
 sg13g2_fill_1 FILLER_26_214 ();
 sg13g2_decap_4 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_251 ();
 sg13g2_fill_2 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_decap_8 FILLER_26_306 ();
 sg13g2_decap_4 FILLER_26_313 ();
 sg13g2_fill_2 FILLER_26_317 ();
 sg13g2_fill_2 FILLER_26_324 ();
 sg13g2_decap_4 FILLER_26_330 ();
 sg13g2_decap_8 FILLER_26_338 ();
 sg13g2_decap_4 FILLER_26_345 ();
 sg13g2_fill_2 FILLER_26_349 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_4 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_116 ();
 sg13g2_fill_1 FILLER_27_194 ();
 sg13g2_fill_2 FILLER_27_212 ();
 sg13g2_fill_2 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_fill_1 FILLER_27_249 ();
 sg13g2_fill_1 FILLER_27_265 ();
 sg13g2_fill_2 FILLER_27_274 ();
 sg13g2_decap_4 FILLER_27_285 ();
 sg13g2_fill_1 FILLER_27_289 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_2 FILLER_27_308 ();
 sg13g2_fill_1 FILLER_27_323 ();
 sg13g2_fill_2 FILLER_27_355 ();
 sg13g2_fill_1 FILLER_27_362 ();
 sg13g2_fill_1 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_fill_2 FILLER_27_394 ();
 sg13g2_fill_1 FILLER_27_396 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_4 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_123 ();
 sg13g2_fill_2 FILLER_28_141 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_fill_1 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_191 ();
 sg13g2_fill_2 FILLER_28_245 ();
 sg13g2_fill_1 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_274 ();
 sg13g2_fill_1 FILLER_28_288 ();
 sg13g2_fill_2 FILLER_28_298 ();
 sg13g2_fill_2 FILLER_28_312 ();
 sg13g2_fill_2 FILLER_28_339 ();
 sg13g2_fill_1 FILLER_28_364 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_112 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_163 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_fill_2 FILLER_29_191 ();
 sg13g2_fill_1 FILLER_29_201 ();
 sg13g2_decap_8 FILLER_29_207 ();
 sg13g2_decap_8 FILLER_29_214 ();
 sg13g2_fill_1 FILLER_29_221 ();
 sg13g2_decap_8 FILLER_29_240 ();
 sg13g2_decap_4 FILLER_29_247 ();
 sg13g2_fill_2 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_decap_4 FILLER_29_273 ();
 sg13g2_fill_2 FILLER_29_298 ();
 sg13g2_fill_2 FILLER_29_318 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_367 ();
 sg13g2_fill_1 FILLER_29_374 ();
 sg13g2_decap_4 FILLER_29_389 ();
 sg13g2_fill_1 FILLER_29_397 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_4 FILLER_30_112 ();
 sg13g2_fill_2 FILLER_30_116 ();
 sg13g2_fill_2 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_168 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_fill_1 FILLER_30_194 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_fill_1 FILLER_30_220 ();
 sg13g2_fill_1 FILLER_30_242 ();
 sg13g2_decap_8 FILLER_30_264 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_decap_4 FILLER_30_278 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_4 FILLER_30_294 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_312 ();
 sg13g2_fill_2 FILLER_30_326 ();
 sg13g2_fill_1 FILLER_30_328 ();
 sg13g2_fill_2 FILLER_30_340 ();
 sg13g2_decap_4 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_4 FILLER_31_119 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_fill_1 FILLER_31_150 ();
 sg13g2_fill_2 FILLER_31_161 ();
 sg13g2_fill_1 FILLER_31_176 ();
 sg13g2_fill_2 FILLER_31_183 ();
 sg13g2_fill_1 FILLER_31_185 ();
 sg13g2_fill_2 FILLER_31_192 ();
 sg13g2_fill_2 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_209 ();
 sg13g2_decap_8 FILLER_31_218 ();
 sg13g2_fill_1 FILLER_31_225 ();
 sg13g2_fill_1 FILLER_31_236 ();
 sg13g2_decap_4 FILLER_31_242 ();
 sg13g2_fill_1 FILLER_31_246 ();
 sg13g2_decap_4 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_264 ();
 sg13g2_fill_2 FILLER_31_293 ();
 sg13g2_fill_1 FILLER_31_295 ();
 sg13g2_fill_2 FILLER_31_325 ();
 sg13g2_fill_1 FILLER_31_327 ();
 sg13g2_decap_4 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_368 ();
 sg13g2_fill_1 FILLER_31_374 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_fill_2 FILLER_32_119 ();
 sg13g2_decap_4 FILLER_32_192 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_fill_1 FILLER_32_222 ();
 sg13g2_fill_2 FILLER_32_231 ();
 sg13g2_decap_4 FILLER_32_238 ();
 sg13g2_fill_2 FILLER_32_248 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_fill_1 FILLER_32_279 ();
 sg13g2_decap_4 FILLER_32_285 ();
 sg13g2_fill_1 FILLER_32_289 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_fill_2 FILLER_32_301 ();
 sg13g2_fill_1 FILLER_32_303 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_fill_2 FILLER_32_329 ();
 sg13g2_fill_1 FILLER_32_331 ();
 sg13g2_fill_1 FILLER_32_344 ();
 sg13g2_decap_4 FILLER_32_351 ();
 sg13g2_fill_2 FILLER_32_365 ();
 sg13g2_fill_1 FILLER_32_367 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_119 ();
 sg13g2_fill_1 FILLER_33_146 ();
 sg13g2_fill_2 FILLER_33_169 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_fill_1 FILLER_33_187 ();
 sg13g2_fill_2 FILLER_33_198 ();
 sg13g2_decap_4 FILLER_33_216 ();
 sg13g2_fill_2 FILLER_33_220 ();
 sg13g2_decap_4 FILLER_33_243 ();
 sg13g2_decap_4 FILLER_33_257 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_272 ();
 sg13g2_decap_4 FILLER_33_297 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_314 ();
 sg13g2_fill_2 FILLER_33_331 ();
 sg13g2_fill_1 FILLER_33_333 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_fill_2 FILLER_33_376 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_fill_1 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_167 ();
 sg13g2_fill_1 FILLER_34_169 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_fill_2 FILLER_34_218 ();
 sg13g2_fill_1 FILLER_34_220 ();
 sg13g2_decap_8 FILLER_34_226 ();
 sg13g2_decap_8 FILLER_34_233 ();
 sg13g2_decap_8 FILLER_34_247 ();
 sg13g2_decap_8 FILLER_34_254 ();
 sg13g2_fill_1 FILLER_34_261 ();
 sg13g2_decap_4 FILLER_34_275 ();
 sg13g2_fill_2 FILLER_34_279 ();
 sg13g2_decap_8 FILLER_34_285 ();
 sg13g2_decap_8 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_299 ();
 sg13g2_fill_1 FILLER_34_306 ();
 sg13g2_fill_2 FILLER_34_312 ();
 sg13g2_fill_2 FILLER_34_331 ();
 sg13g2_fill_1 FILLER_34_366 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_4 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_116 ();
 sg13g2_fill_1 FILLER_35_121 ();
 sg13g2_fill_1 FILLER_35_158 ();
 sg13g2_decap_4 FILLER_35_187 ();
 sg13g2_fill_1 FILLER_35_191 ();
 sg13g2_decap_4 FILLER_35_222 ();
 sg13g2_fill_1 FILLER_35_226 ();
 sg13g2_fill_2 FILLER_35_231 ();
 sg13g2_fill_2 FILLER_35_240 ();
 sg13g2_fill_1 FILLER_35_258 ();
 sg13g2_fill_1 FILLER_35_291 ();
 sg13g2_fill_2 FILLER_35_317 ();
 sg13g2_fill_1 FILLER_35_319 ();
 sg13g2_fill_2 FILLER_35_324 ();
 sg13g2_fill_1 FILLER_35_326 ();
 sg13g2_decap_4 FILLER_35_332 ();
 sg13g2_fill_1 FILLER_35_336 ();
 sg13g2_fill_2 FILLER_35_368 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_4 FILLER_36_119 ();
 sg13g2_fill_2 FILLER_36_123 ();
 sg13g2_fill_1 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_decap_8 FILLER_36_220 ();
 sg13g2_decap_8 FILLER_36_227 ();
 sg13g2_fill_1 FILLER_36_234 ();
 sg13g2_fill_1 FILLER_36_251 ();
 sg13g2_decap_8 FILLER_36_257 ();
 sg13g2_fill_1 FILLER_36_264 ();
 sg13g2_fill_2 FILLER_36_273 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_decap_8 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_310 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_330 ();
 sg13g2_fill_1 FILLER_36_344 ();
 sg13g2_fill_1 FILLER_36_361 ();
 sg13g2_fill_1 FILLER_36_371 ();
 sg13g2_fill_2 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_4 FILLER_37_140 ();
 sg13g2_fill_2 FILLER_37_144 ();
 sg13g2_decap_8 FILLER_37_150 ();
 sg13g2_decap_8 FILLER_37_166 ();
 sg13g2_decap_8 FILLER_37_173 ();
 sg13g2_decap_8 FILLER_37_180 ();
 sg13g2_decap_4 FILLER_37_187 ();
 sg13g2_fill_2 FILLER_37_191 ();
 sg13g2_decap_8 FILLER_37_197 ();
 sg13g2_decap_8 FILLER_37_204 ();
 sg13g2_decap_8 FILLER_37_211 ();
 sg13g2_decap_8 FILLER_37_218 ();
 sg13g2_fill_1 FILLER_37_251 ();
 sg13g2_fill_1 FILLER_37_271 ();
 sg13g2_decap_4 FILLER_37_276 ();
 sg13g2_fill_1 FILLER_37_288 ();
 sg13g2_decap_8 FILLER_37_302 ();
 sg13g2_fill_2 FILLER_37_309 ();
 sg13g2_fill_1 FILLER_37_311 ();
 sg13g2_fill_2 FILLER_37_361 ();
 sg13g2_fill_2 FILLER_37_393 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_4 FILLER_38_229 ();
 sg13g2_fill_1 FILLER_38_233 ();
 sg13g2_fill_1 FILLER_38_239 ();
 sg13g2_decap_4 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_265 ();
 sg13g2_fill_2 FILLER_38_272 ();
 sg13g2_fill_1 FILLER_38_274 ();
 sg13g2_fill_2 FILLER_38_282 ();
 sg13g2_fill_1 FILLER_38_284 ();
 sg13g2_decap_8 FILLER_38_304 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_fill_2 FILLER_38_332 ();
 sg13g2_fill_1 FILLER_38_334 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule

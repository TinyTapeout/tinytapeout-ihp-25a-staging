module tt_um_tommythorn_workshop (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire clknet_0_clk;
 wire \pdm_inst.O ;
 wire \pdm_inst.level[0] ;
 wire \pdm_inst.level[10] ;
 wire \pdm_inst.level[11] ;
 wire \pdm_inst.level[12] ;
 wire \pdm_inst.level[13] ;
 wire \pdm_inst.level[14] ;
 wire \pdm_inst.level[15] ;
 wire \pdm_inst.level[1] ;
 wire \pdm_inst.level[2] ;
 wire \pdm_inst.level[3] ;
 wire \pdm_inst.level[4] ;
 wire \pdm_inst.level[5] ;
 wire \pdm_inst.level[6] ;
 wire \pdm_inst.level[7] ;
 wire \pdm_inst.level[8] ;
 wire \pdm_inst.level[9] ;
 wire \pdm_inst.sigma[0] ;
 wire \pdm_inst.sigma[10] ;
 wire \pdm_inst.sigma[11] ;
 wire \pdm_inst.sigma[12] ;
 wire \pdm_inst.sigma[13] ;
 wire \pdm_inst.sigma[14] ;
 wire \pdm_inst.sigma[15] ;
 wire \pdm_inst.sigma[16] ;
 wire \pdm_inst.sigma[17] ;
 wire \pdm_inst.sigma[1] ;
 wire \pdm_inst.sigma[2] ;
 wire \pdm_inst.sigma[3] ;
 wire \pdm_inst.sigma[4] ;
 wire \pdm_inst.sigma[5] ;
 wire \pdm_inst.sigma[6] ;
 wire \pdm_inst.sigma[7] ;
 wire \pdm_inst.sigma[8] ;
 wire \pdm_inst.sigma[9] ;
 wire \rs232in_inst.attention ;
 wire \rs232in_inst.count[0] ;
 wire \rs232in_inst.count[1] ;
 wire \rs232in_inst.count[2] ;
 wire \rs232in_inst.count[3] ;
 wire \rs232in_inst.count[4] ;
 wire \rs232in_inst.received_data[0] ;
 wire \rs232in_inst.received_data[1] ;
 wire \rs232in_inst.received_data[2] ;
 wire \rs232in_inst.received_data[3] ;
 wire \rs232in_inst.received_data[4] ;
 wire \rs232in_inst.received_data[5] ;
 wire \rs232in_inst.received_data[6] ;
 wire \rs232in_inst.received_data[7] ;
 wire \rs232in_inst.rxd ;
 wire \rs232in_inst.rxd2 ;
 wire \rs232in_inst.shift_in[1] ;
 wire \rs232in_inst.shift_in[2] ;
 wire \rs232in_inst.shift_in[3] ;
 wire \rs232in_inst.shift_in[4] ;
 wire \rs232in_inst.shift_in[5] ;
 wire \rs232in_inst.shift_in[6] ;
 wire \rs232in_inst.shift_in[7] ;
 wire \rs232in_inst.ttyclk[0] ;
 wire \rs232in_inst.ttyclk[10] ;
 wire \rs232in_inst.ttyclk[11] ;
 wire \rs232in_inst.ttyclk[12] ;
 wire \rs232in_inst.ttyclk[13] ;
 wire \rs232in_inst.ttyclk[14] ;
 wire \rs232in_inst.ttyclk[15] ;
 wire \rs232in_inst.ttyclk[16] ;
 wire \rs232in_inst.ttyclk[1] ;
 wire \rs232in_inst.ttyclk[2] ;
 wire \rs232in_inst.ttyclk[3] ;
 wire \rs232in_inst.ttyclk[4] ;
 wire \rs232in_inst.ttyclk[5] ;
 wire \rs232in_inst.ttyclk[6] ;
 wire \rs232in_inst.ttyclk[7] ;
 wire \rs232in_inst.ttyclk[8] ;
 wire \rs232in_inst.ttyclk[9] ;
 wire \rs232out_inst.count[0] ;
 wire \rs232out_inst.count[1] ;
 wire \rs232out_inst.count[2] ;
 wire \rs232out_inst.count[3] ;
 wire \rs232out_inst.count[4] ;
 wire \rs232out_inst.serial_out ;
 wire \rs232out_inst.shift_out[1] ;
 wire \rs232out_inst.shift_out[2] ;
 wire \rs232out_inst.shift_out[3] ;
 wire \rs232out_inst.shift_out[4] ;
 wire \rs232out_inst.shift_out[5] ;
 wire \rs232out_inst.shift_out[6] ;
 wire \rs232out_inst.shift_out[7] ;
 wire \rs232out_inst.shift_out[8] ;
 wire \rs232out_inst.transmit_data[0] ;
 wire \rs232out_inst.transmit_data[1] ;
 wire \rs232out_inst.transmit_data[2] ;
 wire \rs232out_inst.transmit_data[3] ;
 wire \rs232out_inst.transmit_data[4] ;
 wire \rs232out_inst.transmit_data[5] ;
 wire \rs232out_inst.transmit_data[6] ;
 wire \rs232out_inst.transmit_data[7] ;
 wire \rs232out_inst.ttyclk[0] ;
 wire \rs232out_inst.ttyclk[10] ;
 wire \rs232out_inst.ttyclk[11] ;
 wire \rs232out_inst.ttyclk[12] ;
 wire \rs232out_inst.ttyclk[13] ;
 wire \rs232out_inst.ttyclk[14] ;
 wire \rs232out_inst.ttyclk[15] ;
 wire \rs232out_inst.ttyclk[16] ;
 wire \rs232out_inst.ttyclk[1] ;
 wire \rs232out_inst.ttyclk[2] ;
 wire \rs232out_inst.ttyclk[3] ;
 wire \rs232out_inst.ttyclk[4] ;
 wire \rs232out_inst.ttyclk[5] ;
 wire \rs232out_inst.ttyclk[6] ;
 wire \rs232out_inst.ttyclk[7] ;
 wire \rs232out_inst.ttyclk[8] ;
 wire \rs232out_inst.ttyclk[9] ;
 wire \rs232out_inst.we ;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;

 sg13g2_inv_1 _0621_ (.Y(_0124_),
    .A(net253));
 sg13g2_inv_1 _0622_ (.Y(_0125_),
    .A(net170));
 sg13g2_inv_1 _0623_ (.Y(_0126_),
    .A(net273));
 sg13g2_inv_1 _0624_ (.Y(_0127_),
    .A(\rs232out_inst.ttyclk[4] ));
 sg13g2_inv_1 _0625_ (.Y(_0128_),
    .A(\rs232out_inst.count[0] ));
 sg13g2_inv_1 _0626_ (.Y(_0129_),
    .A(net168));
 sg13g2_inv_1 _0627_ (.Y(_0130_),
    .A(net212));
 sg13g2_inv_1 _0628_ (.Y(_0131_),
    .A(\rs232in_inst.ttyclk[7] ));
 sg13g2_inv_1 _0629_ (.Y(_0132_),
    .A(\rs232in_inst.received_data[4] ));
 sg13g2_inv_1 _0630_ (.Y(_0133_),
    .A(net322));
 sg13g2_inv_1 _0631_ (.Y(_0134_),
    .A(net1));
 sg13g2_nand2_1 _0632_ (.Y(_0135_),
    .A(net74),
    .B(net68));
 sg13g2_nor2_2 _0633_ (.A(net332),
    .B(_0135_),
    .Y(_0136_));
 sg13g2_nand3b_1 _0634_ (.B(\rs232out_inst.ttyclk[16] ),
    .C(net74),
    .Y(_0137_),
    .A_N(\rs232out_inst.we ));
 sg13g2_or2_1 _0635_ (.X(_0138_),
    .B(\rs232out_inst.ttyclk[2] ),
    .A(\rs232out_inst.ttyclk[1] ));
 sg13g2_nor4_2 _0636_ (.A(net237),
    .B(\rs232out_inst.ttyclk[1] ),
    .C(net222),
    .Y(_0139_),
    .D(net260));
 sg13g2_or2_1 _0637_ (.X(_0140_),
    .B(\rs232out_inst.ttyclk[5] ),
    .A(\rs232out_inst.ttyclk[4] ));
 sg13g2_nor4_2 _0638_ (.A(\rs232out_inst.ttyclk[4] ),
    .B(net233),
    .C(net224),
    .Y(_0141_),
    .D(net292));
 sg13g2_nor4_1 _0639_ (.A(net321),
    .B(net323),
    .C(net263),
    .D(\rs232out_inst.ttyclk[11] ),
    .Y(_0142_));
 sg13g2_nor2_1 _0640_ (.A(\rs232out_inst.ttyclk[16] ),
    .B(\rs232out_inst.ttyclk[12] ),
    .Y(_0143_));
 sg13g2_nand4_1 _0641_ (.B(_0141_),
    .C(_0142_),
    .A(_0139_),
    .Y(_0144_),
    .D(_0143_));
 sg13g2_nor4_1 _0642_ (.A(net319),
    .B(net278),
    .C(net255),
    .D(_0144_),
    .Y(_0145_));
 sg13g2_or2_1 _0643_ (.X(_0001_),
    .B(_0145_),
    .A(_0136_));
 sg13g2_nor2_1 _0644_ (.A(\rs232in_inst.count[0] ),
    .B(\rs232in_inst.count[1] ),
    .Y(_0146_));
 sg13g2_nand2_1 _0645_ (.Y(_0147_),
    .A(_0124_),
    .B(_0125_));
 sg13g2_nor3_2 _0646_ (.A(net267),
    .B(net291),
    .C(net174),
    .Y(_0148_));
 sg13g2_and2_1 _0647_ (.A(_0146_),
    .B(_0148_),
    .X(_0149_));
 sg13g2_nand2_2 _0648_ (.Y(_0150_),
    .A(_0146_),
    .B(_0148_));
 sg13g2_and3_1 _0649_ (.X(_0151_),
    .A(net70),
    .B(\rs232in_inst.rxd2 ),
    .C(_0149_));
 sg13g2_nor2_1 _0650_ (.A(\rs232in_inst.ttyclk[0] ),
    .B(\rs232in_inst.ttyclk[1] ),
    .Y(_0152_));
 sg13g2_nor4_1 _0651_ (.A(\rs232in_inst.ttyclk[0] ),
    .B(\rs232in_inst.ttyclk[1] ),
    .C(\rs232in_inst.ttyclk[2] ),
    .D(net250),
    .Y(_0153_));
 sg13g2_or4_2 _0652_ (.A(\rs232in_inst.ttyclk[0] ),
    .B(\rs232in_inst.ttyclk[1] ),
    .C(\rs232in_inst.ttyclk[2] ),
    .D(net250),
    .X(_0154_));
 sg13g2_nor4_2 _0653_ (.A(\rs232in_inst.ttyclk[4] ),
    .B(\rs232in_inst.ttyclk[5] ),
    .C(net359),
    .Y(_0155_),
    .D(_0154_));
 sg13g2_and2_1 _0654_ (.A(_0131_),
    .B(_0155_),
    .X(_0156_));
 sg13g2_nand2_1 _0655_ (.Y(_0157_),
    .A(_0131_),
    .B(_0155_));
 sg13g2_or2_1 _0656_ (.X(_0158_),
    .B(net305),
    .A(net314));
 sg13g2_nor4_1 _0657_ (.A(net71),
    .B(net330),
    .C(net339),
    .D(net246),
    .Y(_0159_));
 sg13g2_nor3_1 _0658_ (.A(net284),
    .B(net317),
    .C(net234),
    .Y(_0160_));
 sg13g2_nand2_1 _0659_ (.Y(_0161_),
    .A(_0159_),
    .B(_0160_));
 sg13g2_nor3_1 _0660_ (.A(net360),
    .B(_0158_),
    .C(_0161_),
    .Y(_0162_));
 sg13g2_or2_1 _0661_ (.X(_0000_),
    .B(_0162_),
    .A(net57));
 sg13g2_nand2_1 _0662_ (.Y(_0163_),
    .A(net8),
    .B(net2));
 sg13g2_xor2_1 _0663_ (.B(net3),
    .A(net9),
    .X(_0164_));
 sg13g2_nor2b_1 _0664_ (.A(_0163_),
    .B_N(_0164_),
    .Y(_0165_));
 sg13g2_xnor2_1 _0665_ (.Y(uo_out[3]),
    .A(_0163_),
    .B(_0164_));
 sg13g2_a21oi_1 _0666_ (.A1(net9),
    .A2(net3),
    .Y(_0166_),
    .B1(_0165_));
 sg13g2_nand2_1 _0667_ (.Y(_0167_),
    .A(net10),
    .B(net4));
 sg13g2_xnor2_1 _0668_ (.Y(_0168_),
    .A(net10),
    .B(net4));
 sg13g2_xor2_1 _0669_ (.B(_0168_),
    .A(_0166_),
    .X(uo_out[4]));
 sg13g2_o21ai_1 _0670_ (.B1(_0167_),
    .Y(_0169_),
    .A1(_0166_),
    .A2(_0168_));
 sg13g2_inv_1 _0671_ (.Y(_0170_),
    .A(_0169_));
 sg13g2_nand2_1 _0672_ (.Y(_0171_),
    .A(net11),
    .B(net5));
 sg13g2_xnor2_1 _0673_ (.Y(_0172_),
    .A(net11),
    .B(net5));
 sg13g2_xnor2_1 _0674_ (.Y(uo_out[5]),
    .A(_0169_),
    .B(_0172_));
 sg13g2_o21ai_1 _0675_ (.B1(_0171_),
    .Y(_0173_),
    .A1(_0170_),
    .A2(_0172_));
 sg13g2_and2_1 _0676_ (.A(net12),
    .B(net6),
    .X(_0174_));
 sg13g2_or2_1 _0677_ (.X(_0175_),
    .B(net6),
    .A(net12));
 sg13g2_nand2b_1 _0678_ (.Y(_0176_),
    .B(_0175_),
    .A_N(_0174_));
 sg13g2_xnor2_1 _0679_ (.Y(uo_out[6]),
    .A(_0173_),
    .B(_0176_));
 sg13g2_a21oi_1 _0680_ (.A1(_0173_),
    .A2(_0175_),
    .Y(_0177_),
    .B1(_0174_));
 sg13g2_xor2_1 _0681_ (.B(net7),
    .A(net13),
    .X(_0178_));
 sg13g2_xnor2_1 _0682_ (.Y(uo_out[7]),
    .A(_0177_),
    .B(_0178_));
 sg13g2_xor2_1 _0683_ (.B(net2),
    .A(net8),
    .X(uo_out[2]));
 sg13g2_nand2_1 _0684_ (.Y(_0179_),
    .A(net276),
    .B(net182));
 sg13g2_nand2_1 _0685_ (.Y(_0180_),
    .A(net331),
    .B(net324));
 sg13g2_nor2_1 _0686_ (.A(\pdm_inst.level[1] ),
    .B(net357),
    .Y(_0181_));
 sg13g2_xor2_1 _0687_ (.B(net324),
    .A(\pdm_inst.level[1] ),
    .X(_0182_));
 sg13g2_xnor2_1 _0688_ (.Y(_0021_),
    .A(_0179_),
    .B(net325));
 sg13g2_o21ai_1 _0689_ (.B1(_0180_),
    .Y(_0183_),
    .A1(_0179_),
    .A2(_0181_));
 sg13g2_xnor2_1 _0690_ (.Y(_0184_),
    .A(net328),
    .B(net343));
 sg13g2_nor2b_1 _0691_ (.A(_0184_),
    .B_N(_0183_),
    .Y(_0185_));
 sg13g2_xnor2_1 _0692_ (.Y(_0022_),
    .A(_0183_),
    .B(_0184_));
 sg13g2_or2_1 _0693_ (.X(_0186_),
    .B(\pdm_inst.sigma[3] ),
    .A(\pdm_inst.level[3] ));
 sg13g2_xor2_1 _0694_ (.B(\pdm_inst.sigma[3] ),
    .A(\pdm_inst.level[3] ),
    .X(_0187_));
 sg13g2_a21oi_1 _0695_ (.A1(net328),
    .A2(net343),
    .Y(_0188_),
    .B1(_0185_));
 sg13g2_xnor2_1 _0696_ (.Y(_0023_),
    .A(_0187_),
    .B(_0188_));
 sg13g2_nor2b_1 _0697_ (.A(_0184_),
    .B_N(_0187_),
    .Y(_0189_));
 sg13g2_and3_1 _0698_ (.X(_0190_),
    .A(\pdm_inst.level[2] ),
    .B(\pdm_inst.sigma[2] ),
    .C(_0186_));
 sg13g2_a221oi_1 _0699_ (.B2(_0189_),
    .C1(_0190_),
    .B1(_0183_),
    .A1(\pdm_inst.level[3] ),
    .Y(_0191_),
    .A2(\pdm_inst.sigma[3] ));
 sg13g2_xor2_1 _0700_ (.B(net334),
    .A(net280),
    .X(_0192_));
 sg13g2_nor2b_1 _0701_ (.A(_0191_),
    .B_N(_0192_),
    .Y(_0193_));
 sg13g2_xnor2_1 _0702_ (.Y(_0024_),
    .A(_0191_),
    .B(_0192_));
 sg13g2_nor2_1 _0703_ (.A(\pdm_inst.level[5] ),
    .B(\pdm_inst.sigma[5] ),
    .Y(_0194_));
 sg13g2_nand2_1 _0704_ (.Y(_0195_),
    .A(net310),
    .B(\pdm_inst.sigma[5] ));
 sg13g2_nand2b_1 _0705_ (.Y(_0196_),
    .B(_0195_),
    .A_N(_0194_));
 sg13g2_a21oi_1 _0706_ (.A1(net280),
    .A2(net334),
    .Y(_0197_),
    .B1(_0193_));
 sg13g2_xor2_1 _0707_ (.B(_0197_),
    .A(_0196_),
    .X(_0025_));
 sg13g2_nand2_1 _0708_ (.Y(_0198_),
    .A(net308),
    .B(\pdm_inst.sigma[6] ));
 sg13g2_xnor2_1 _0709_ (.Y(_0199_),
    .A(net308),
    .B(net366));
 sg13g2_a22oi_1 _0710_ (.Y(_0200_),
    .B1(\pdm_inst.level[5] ),
    .B2(\pdm_inst.sigma[5] ),
    .A2(\pdm_inst.sigma[4] ),
    .A1(\pdm_inst.level[4] ));
 sg13g2_or2_1 _0711_ (.X(_0201_),
    .B(_0200_),
    .A(_0194_));
 sg13g2_nand3b_1 _0712_ (.B(_0195_),
    .C(_0192_),
    .Y(_0202_),
    .A_N(_0194_));
 sg13g2_o21ai_1 _0713_ (.B1(_0201_),
    .Y(_0203_),
    .A1(_0191_),
    .A2(_0202_));
 sg13g2_nand2b_1 _0714_ (.Y(_0204_),
    .B(_0203_),
    .A_N(_0199_));
 sg13g2_xnor2_1 _0715_ (.Y(_0026_),
    .A(_0199_),
    .B(_0203_));
 sg13g2_nor2_1 _0716_ (.A(\pdm_inst.level[7] ),
    .B(\pdm_inst.sigma[7] ),
    .Y(_0205_));
 sg13g2_nand2_1 _0717_ (.Y(_0206_),
    .A(\pdm_inst.level[7] ),
    .B(\pdm_inst.sigma[7] ));
 sg13g2_xnor2_1 _0718_ (.Y(_0207_),
    .A(net322),
    .B(net364));
 sg13g2_and2_1 _0719_ (.A(_0198_),
    .B(_0204_),
    .X(_0208_));
 sg13g2_xor2_1 _0720_ (.B(_0208_),
    .A(_0207_),
    .X(_0027_));
 sg13g2_or3_1 _0721_ (.A(_0199_),
    .B(_0202_),
    .C(_0207_),
    .X(_0209_));
 sg13g2_o21ai_1 _0722_ (.B1(_0206_),
    .Y(_0210_),
    .A1(_0198_),
    .A2(_0205_));
 sg13g2_nor4_1 _0723_ (.A(_0194_),
    .B(_0199_),
    .C(_0200_),
    .D(_0207_),
    .Y(_0211_));
 sg13g2_nor2_1 _0724_ (.A(_0210_),
    .B(_0211_),
    .Y(_0212_));
 sg13g2_o21ai_1 _0725_ (.B1(_0212_),
    .Y(_0213_),
    .A1(_0191_),
    .A2(_0209_));
 sg13g2_xnor2_1 _0726_ (.Y(_0214_),
    .A(net358),
    .B(net345));
 sg13g2_nor2b_1 _0727_ (.A(_0214_),
    .B_N(_0213_),
    .Y(_0215_));
 sg13g2_xnor2_1 _0728_ (.Y(_0028_),
    .A(_0213_),
    .B(_0214_));
 sg13g2_nor2_1 _0729_ (.A(\pdm_inst.level[9] ),
    .B(\pdm_inst.sigma[9] ),
    .Y(_0216_));
 sg13g2_xor2_1 _0730_ (.B(\pdm_inst.sigma[9] ),
    .A(net326),
    .X(_0217_));
 sg13g2_a21oi_1 _0731_ (.A1(\pdm_inst.level[8] ),
    .A2(net345),
    .Y(_0218_),
    .B1(_0215_));
 sg13g2_xnor2_1 _0732_ (.Y(_0029_),
    .A(_0217_),
    .B(net346));
 sg13g2_nand2_1 _0733_ (.Y(_0219_),
    .A(\pdm_inst.level[10] ),
    .B(net355));
 sg13g2_nor2_1 _0734_ (.A(\pdm_inst.level[10] ),
    .B(net355),
    .Y(_0220_));
 sg13g2_xor2_1 _0735_ (.B(net355),
    .A(\pdm_inst.level[10] ),
    .X(_0221_));
 sg13g2_a22oi_1 _0736_ (.Y(_0222_),
    .B1(\pdm_inst.level[9] ),
    .B2(\pdm_inst.sigma[9] ),
    .A2(\pdm_inst.sigma[8] ),
    .A1(\pdm_inst.level[8] ));
 sg13g2_or2_1 _0737_ (.X(_0223_),
    .B(_0222_),
    .A(_0216_));
 sg13g2_nand2b_1 _0738_ (.Y(_0224_),
    .B(_0217_),
    .A_N(_0214_));
 sg13g2_nand2b_1 _0739_ (.Y(_0225_),
    .B(_0213_),
    .A_N(_0224_));
 sg13g2_and2_1 _0740_ (.A(_0223_),
    .B(_0225_),
    .X(_0226_));
 sg13g2_xnor2_1 _0741_ (.Y(_0013_),
    .A(net356),
    .B(_0226_));
 sg13g2_nor2_1 _0742_ (.A(net298),
    .B(net361),
    .Y(_0227_));
 sg13g2_nand2_1 _0743_ (.Y(_0228_),
    .A(net298),
    .B(net361));
 sg13g2_nand2b_1 _0744_ (.Y(_0229_),
    .B(_0228_),
    .A_N(_0227_));
 sg13g2_o21ai_1 _0745_ (.B1(_0219_),
    .Y(_0230_),
    .A1(_0220_),
    .A2(_0226_));
 sg13g2_xnor2_1 _0746_ (.Y(_0014_),
    .A(_0229_),
    .B(_0230_));
 sg13g2_nand3b_1 _0747_ (.B(_0228_),
    .C(_0221_),
    .Y(_0231_),
    .A_N(_0227_));
 sg13g2_nor2_1 _0748_ (.A(_0224_),
    .B(_0231_),
    .Y(_0232_));
 sg13g2_o21ai_1 _0749_ (.B1(_0228_),
    .Y(_0233_),
    .A1(_0219_),
    .A2(_0227_));
 sg13g2_nor2_1 _0750_ (.A(_0223_),
    .B(_0231_),
    .Y(_0234_));
 sg13g2_or2_1 _0751_ (.X(_0235_),
    .B(_0234_),
    .A(_0233_));
 sg13g2_a21oi_1 _0752_ (.A1(_0213_),
    .A2(_0232_),
    .Y(_0236_),
    .B1(_0235_));
 sg13g2_a21o_1 _0753_ (.A2(_0232_),
    .A1(_0213_),
    .B1(_0235_),
    .X(_0237_));
 sg13g2_nand2_1 _0754_ (.Y(_0238_),
    .A(net300),
    .B(net354));
 sg13g2_xnor2_1 _0755_ (.Y(_0239_),
    .A(net300),
    .B(net354));
 sg13g2_xnor2_1 _0756_ (.Y(_0015_),
    .A(_0237_),
    .B(_0239_));
 sg13g2_nor2_1 _0757_ (.A(net286),
    .B(net363),
    .Y(_0240_));
 sg13g2_nand2_1 _0758_ (.Y(_0241_),
    .A(net286),
    .B(net363));
 sg13g2_nor2b_1 _0759_ (.A(_0240_),
    .B_N(_0241_),
    .Y(_0242_));
 sg13g2_o21ai_1 _0760_ (.B1(_0238_),
    .Y(_0243_),
    .A1(_0236_),
    .A2(_0239_));
 sg13g2_xor2_1 _0761_ (.B(_0243_),
    .A(_0242_),
    .X(_0016_));
 sg13g2_nor2b_1 _0762_ (.A(_0239_),
    .B_N(_0242_),
    .Y(_0244_));
 sg13g2_o21ai_1 _0763_ (.B1(_0241_),
    .Y(_0245_),
    .A1(_0238_),
    .A2(_0240_));
 sg13g2_a21oi_2 _0764_ (.B1(_0245_),
    .Y(_0246_),
    .A2(_0244_),
    .A1(_0237_));
 sg13g2_nand2_1 _0765_ (.Y(_0247_),
    .A(\pdm_inst.level[14] ),
    .B(\pdm_inst.sigma[14] ));
 sg13g2_nor2_1 _0766_ (.A(\pdm_inst.level[14] ),
    .B(\pdm_inst.sigma[14] ),
    .Y(_0248_));
 sg13g2_xor2_1 _0767_ (.B(net350),
    .A(\pdm_inst.level[14] ),
    .X(_0249_));
 sg13g2_xnor2_1 _0768_ (.Y(_0017_),
    .A(_0246_),
    .B(net351));
 sg13g2_nand2_1 _0769_ (.Y(_0250_),
    .A(\pdm_inst.level[15] ),
    .B(\pdm_inst.sigma[15] ));
 sg13g2_nor2_1 _0770_ (.A(\pdm_inst.level[15] ),
    .B(\pdm_inst.sigma[15] ),
    .Y(_0251_));
 sg13g2_xnor2_1 _0771_ (.Y(_0252_),
    .A(net288),
    .B(net348));
 sg13g2_o21ai_1 _0772_ (.B1(_0247_),
    .Y(_0253_),
    .A1(_0246_),
    .A2(_0248_));
 sg13g2_xnor2_1 _0773_ (.Y(_0018_),
    .A(_0252_),
    .B(_0253_));
 sg13g2_nand3b_1 _0774_ (.B(_0249_),
    .C(_0250_),
    .Y(_0254_),
    .A_N(_0251_));
 sg13g2_nor2_1 _0775_ (.A(_0247_),
    .B(_0251_),
    .Y(_0255_));
 sg13g2_a21oi_1 _0776_ (.A1(\pdm_inst.level[15] ),
    .A2(\pdm_inst.sigma[15] ),
    .Y(_0256_),
    .B1(_0255_));
 sg13g2_o21ai_1 _0777_ (.B1(_0256_),
    .Y(_0257_),
    .A1(_0246_),
    .A2(_0254_));
 sg13g2_nor2b_1 _0778_ (.A(net228),
    .B_N(\pdm_inst.sigma[16] ),
    .Y(_0258_));
 sg13g2_xnor2_1 _0779_ (.Y(_0259_),
    .A(net228),
    .B(net337));
 sg13g2_xor2_1 _0780_ (.B(_0259_),
    .A(_0257_),
    .X(_0019_));
 sg13g2_a21oi_1 _0781_ (.A1(_0257_),
    .A2(_0259_),
    .Y(_0020_),
    .B1(net229));
 sg13g2_xor2_1 _0782_ (.B(net182),
    .A(\pdm_inst.level[0] ),
    .X(_0012_));
 sg13g2_nand3_1 _0783_ (.B(net68),
    .C(\rs232in_inst.attention ),
    .A(net73),
    .Y(_0260_));
 sg13g2_mux2_1 _0784_ (.A0(net318),
    .A1(net276),
    .S(net63),
    .X(_0032_));
 sg13g2_mux2_1 _0785_ (.A0(net254),
    .A1(net331),
    .S(net63),
    .X(_0033_));
 sg13g2_mux2_1 _0786_ (.A0(net301),
    .A1(\pdm_inst.level[2] ),
    .S(net63),
    .X(_0034_));
 sg13g2_mux2_1 _0787_ (.A0(net282),
    .A1(\pdm_inst.level[3] ),
    .S(net64),
    .X(_0035_));
 sg13g2_nand2_1 _0788_ (.Y(_0261_),
    .A(net280),
    .B(net66));
 sg13g2_o21ai_1 _0789_ (.B1(_0261_),
    .Y(_0036_),
    .A1(_0132_),
    .A2(net63));
 sg13g2_mux2_1 _0790_ (.A0(net266),
    .A1(net310),
    .S(net66),
    .X(_0037_));
 sg13g2_mux2_1 _0791_ (.A0(net313),
    .A1(net308),
    .S(net66),
    .X(_0038_));
 sg13g2_nor2_2 _0792_ (.A(net220),
    .B(net64),
    .Y(_0262_));
 sg13g2_a21oi_1 _0793_ (.A1(_0133_),
    .A2(net65),
    .Y(_0039_),
    .B1(_0262_));
 sg13g2_mux2_1 _0794_ (.A0(net276),
    .A1(\pdm_inst.level[8] ),
    .S(net63),
    .X(_0040_));
 sg13g2_mux2_1 _0795_ (.A0(\pdm_inst.level[1] ),
    .A1(net326),
    .S(net63),
    .X(_0041_));
 sg13g2_mux2_1 _0796_ (.A0(net328),
    .A1(\pdm_inst.level[10] ),
    .S(net63),
    .X(_0042_));
 sg13g2_mux2_1 _0797_ (.A0(\pdm_inst.level[3] ),
    .A1(net298),
    .S(net66),
    .X(_0043_));
 sg13g2_mux2_1 _0798_ (.A0(net280),
    .A1(net300),
    .S(net66),
    .X(_0044_));
 sg13g2_mux2_1 _0799_ (.A0(\pdm_inst.level[5] ),
    .A1(net286),
    .S(net66),
    .X(_0045_));
 sg13g2_mux2_1 _0800_ (.A0(net308),
    .A1(\pdm_inst.level[14] ),
    .S(net66),
    .X(_0046_));
 sg13g2_nand2_1 _0801_ (.Y(_0263_),
    .A(net288),
    .B(net67));
 sg13g2_o21ai_1 _0802_ (.B1(net289),
    .Y(_0047_),
    .A1(_0133_),
    .A2(net65));
 sg13g2_nand2b_1 _0803_ (.Y(_0264_),
    .B(net68),
    .A_N(net311));
 sg13g2_nor2_1 _0804_ (.A(\rs232out_inst.count[0] ),
    .B(net210),
    .Y(_0265_));
 sg13g2_nand2b_1 _0805_ (.Y(_0266_),
    .B(_0265_),
    .A_N(\rs232out_inst.count[2] ));
 sg13g2_nor2b_2 _0806_ (.A(net73),
    .B_N(net68),
    .Y(_0267_));
 sg13g2_nor2_1 _0807_ (.A(net207),
    .B(_0266_),
    .Y(_0268_));
 sg13g2_a22oi_1 _0808_ (.Y(_0269_),
    .B1(_0267_),
    .B2(_0268_),
    .A2(_0264_),
    .A1(net74));
 sg13g2_inv_1 _0809_ (.Y(_0048_),
    .A(net312));
 sg13g2_mux2_1 _0810_ (.A0(net166),
    .A1(\rs232out_inst.transmit_data[0] ),
    .S(net67),
    .X(_0049_));
 sg13g2_nand2_1 _0811_ (.Y(_0270_),
    .A(net194),
    .B(net64));
 sg13g2_xnor2_1 _0812_ (.Y(_0271_),
    .A(\rs232in_inst.received_data[0] ),
    .B(\rs232in_inst.received_data[1] ));
 sg13g2_o21ai_1 _0813_ (.B1(_0270_),
    .Y(_0050_),
    .A1(net64),
    .A2(_0271_));
 sg13g2_nand3_1 _0814_ (.B(net254),
    .C(\rs232in_inst.received_data[2] ),
    .A(\rs232in_inst.received_data[0] ),
    .Y(_0272_));
 sg13g2_a21o_1 _0815_ (.A2(\rs232in_inst.received_data[1] ),
    .A1(\rs232in_inst.received_data[0] ),
    .B1(\rs232in_inst.received_data[2] ),
    .X(_0273_));
 sg13g2_a21oi_1 _0816_ (.A1(_0272_),
    .A2(_0273_),
    .Y(_0274_),
    .B1(net67));
 sg13g2_a21oi_1 _0817_ (.A1(_0130_),
    .A2(net64),
    .Y(_0051_),
    .B1(_0274_));
 sg13g2_nand4_1 _0818_ (.B(\rs232in_inst.received_data[1] ),
    .C(\rs232in_inst.received_data[2] ),
    .A(\rs232in_inst.received_data[0] ),
    .Y(_0275_),
    .D(\rs232in_inst.received_data[3] ));
 sg13g2_xnor2_1 _0819_ (.Y(_0276_),
    .A(\rs232in_inst.received_data[3] ),
    .B(_0272_));
 sg13g2_mux2_1 _0820_ (.A0(_0276_),
    .A1(net258),
    .S(net64),
    .X(_0052_));
 sg13g2_nand2_1 _0821_ (.Y(_0277_),
    .A(net196),
    .B(net64));
 sg13g2_nor2_1 _0822_ (.A(_0132_),
    .B(_0275_),
    .Y(_0278_));
 sg13g2_a21o_1 _0823_ (.A2(_0275_),
    .A1(_0132_),
    .B1(net63),
    .X(_0279_));
 sg13g2_o21ai_1 _0824_ (.B1(_0277_),
    .Y(_0053_),
    .A1(_0278_),
    .A2(_0279_));
 sg13g2_nor2_1 _0825_ (.A(\rs232in_inst.received_data[5] ),
    .B(_0278_),
    .Y(_0280_));
 sg13g2_and2_1 _0826_ (.A(net266),
    .B(_0278_),
    .X(_0281_));
 sg13g2_nor3_1 _0827_ (.A(net65),
    .B(_0280_),
    .C(_0281_),
    .Y(_0282_));
 sg13g2_a21o_1 _0828_ (.A2(net65),
    .A1(net226),
    .B1(_0282_),
    .X(_0054_));
 sg13g2_nand2_1 _0829_ (.Y(_0283_),
    .A(net184),
    .B(net65));
 sg13g2_nor2_1 _0830_ (.A(\rs232in_inst.received_data[6] ),
    .B(_0281_),
    .Y(_0284_));
 sg13g2_nand2_1 _0831_ (.Y(_0285_),
    .A(\rs232in_inst.received_data[6] ),
    .B(_0281_));
 sg13g2_nand2b_1 _0832_ (.Y(_0286_),
    .B(_0285_),
    .A_N(net65));
 sg13g2_o21ai_1 _0833_ (.B1(_0283_),
    .Y(_0055_),
    .A1(_0284_),
    .A2(_0286_));
 sg13g2_a21oi_1 _0834_ (.A1(net294),
    .A2(net65),
    .Y(_0287_),
    .B1(_0262_));
 sg13g2_a22oi_1 _0835_ (.Y(_0056_),
    .B1(_0286_),
    .B2(_0287_),
    .A2(_0285_),
    .A1(_0262_));
 sg13g2_nor2_1 _0836_ (.A(_0134_),
    .B(net65),
    .Y(_0057_));
 sg13g2_a21oi_1 _0837_ (.A1(\rs232out_inst.we ),
    .A2(net68),
    .Y(_0288_),
    .B1(_0267_));
 sg13g2_inv_1 _0838_ (.Y(_0289_),
    .A(net62));
 sg13g2_nand2b_1 _0839_ (.Y(_0290_),
    .B(\rs232out_inst.count[4] ),
    .A_N(\rs232out_inst.transmit_data[7] ));
 sg13g2_mux2_1 _0840_ (.A0(_0290_),
    .A1(net248),
    .S(net61),
    .X(_0058_));
 sg13g2_nand2_1 _0841_ (.Y(_0291_),
    .A(net237),
    .B(_0136_));
 sg13g2_o21ai_1 _0842_ (.B1(_0291_),
    .Y(_0059_),
    .A1(net68),
    .A2(net237));
 sg13g2_nor2_2 _0843_ (.A(net217),
    .B(_0136_),
    .Y(_0292_));
 sg13g2_nand2b_1 _0844_ (.Y(_0293_),
    .B(_0137_),
    .A_N(\rs232out_inst.ttyclk[0] ));
 sg13g2_nor2_1 _0845_ (.A(\rs232out_inst.ttyclk[1] ),
    .B(_0293_),
    .Y(_0294_));
 sg13g2_xor2_1 _0846_ (.B(_0293_),
    .A(\rs232out_inst.ttyclk[1] ),
    .X(_0295_));
 sg13g2_nor2_1 _0847_ (.A(net218),
    .B(_0295_),
    .Y(_0060_));
 sg13g2_xnor2_1 _0848_ (.Y(_0296_),
    .A(net222),
    .B(_0294_));
 sg13g2_nor2_1 _0849_ (.A(net218),
    .B(net223),
    .Y(_0061_));
 sg13g2_nand2_1 _0850_ (.Y(_0297_),
    .A(_0137_),
    .B(_0139_));
 sg13g2_o21ai_1 _0851_ (.B1(net260),
    .Y(_0298_),
    .A1(_0138_),
    .A2(_0293_));
 sg13g2_a21oi_1 _0852_ (.A1(_0297_),
    .A2(net261),
    .Y(_0062_),
    .B1(net56));
 sg13g2_nand2_1 _0853_ (.Y(_0299_),
    .A(net204),
    .B(_0139_));
 sg13g2_nor2_1 _0854_ (.A(net204),
    .B(_0139_),
    .Y(_0300_));
 sg13g2_nor2_1 _0855_ (.A(net68),
    .B(_0300_),
    .Y(_0301_));
 sg13g2_a22oi_1 _0856_ (.Y(_0063_),
    .B1(net205),
    .B2(_0301_),
    .A2(_0136_),
    .A1(_0127_));
 sg13g2_nor2_1 _0857_ (.A(net68),
    .B(net205),
    .Y(_0302_));
 sg13g2_nor3_1 _0858_ (.A(net233),
    .B(_0289_),
    .C(_0302_),
    .Y(_0303_));
 sg13g2_a21oi_1 _0859_ (.A1(net233),
    .A2(_0302_),
    .Y(_0064_),
    .B1(_0303_));
 sg13g2_or3_1 _0860_ (.A(net224),
    .B(_0140_),
    .C(_0297_),
    .X(_0304_));
 sg13g2_o21ai_1 _0861_ (.B1(net224),
    .Y(_0305_),
    .A1(_0140_),
    .A2(_0297_));
 sg13g2_a21oi_1 _0862_ (.A1(_0304_),
    .A2(_0305_),
    .Y(_0065_),
    .B1(net218));
 sg13g2_nand3_1 _0863_ (.B(_0139_),
    .C(_0141_),
    .A(_0137_),
    .Y(_0306_));
 sg13g2_a21oi_1 _0864_ (.A1(net292),
    .A2(_0304_),
    .Y(_0307_),
    .B1(_0289_));
 sg13g2_nand2_1 _0865_ (.Y(_0066_),
    .A(_0306_),
    .B(_0307_));
 sg13g2_nand2_1 _0866_ (.Y(_0308_),
    .A(net321),
    .B(_0306_));
 sg13g2_or2_1 _0867_ (.X(_0309_),
    .B(_0306_),
    .A(net321));
 sg13g2_nand3_1 _0868_ (.B(_0308_),
    .C(_0309_),
    .A(net61),
    .Y(_0067_));
 sg13g2_nor3_1 _0869_ (.A(net321),
    .B(net323),
    .C(_0306_),
    .Y(_0310_));
 sg13g2_xor2_1 _0870_ (.B(_0309_),
    .A(net323),
    .X(_0311_));
 sg13g2_nor2_1 _0871_ (.A(net56),
    .B(_0311_),
    .Y(_0068_));
 sg13g2_nand2b_2 _0872_ (.Y(_0312_),
    .B(_0310_),
    .A_N(net263));
 sg13g2_nand2b_1 _0873_ (.Y(_0313_),
    .B(net263),
    .A_N(_0310_));
 sg13g2_a21oi_1 _0874_ (.A1(_0312_),
    .A2(net264),
    .Y(_0069_),
    .B1(net56));
 sg13g2_xor2_1 _0875_ (.B(_0312_),
    .A(net336),
    .X(_0314_));
 sg13g2_nor2_1 _0876_ (.A(net56),
    .B(_0314_),
    .Y(_0070_));
 sg13g2_nor3_1 _0877_ (.A(net336),
    .B(net353),
    .C(_0312_),
    .Y(_0315_));
 sg13g2_o21ai_1 _0878_ (.B1(net353),
    .Y(_0316_),
    .A1(net336),
    .A2(_0312_));
 sg13g2_nor2b_1 _0879_ (.A(_0315_),
    .B_N(_0316_),
    .Y(_0317_));
 sg13g2_nor2_1 _0880_ (.A(net56),
    .B(_0317_),
    .Y(_0071_));
 sg13g2_nor4_2 _0881_ (.A(\rs232out_inst.ttyclk[11] ),
    .B(\rs232out_inst.ttyclk[12] ),
    .C(\rs232out_inst.ttyclk[13] ),
    .Y(_0318_),
    .D(_0312_));
 sg13g2_xnor2_1 _0882_ (.Y(_0319_),
    .A(net319),
    .B(_0315_));
 sg13g2_nor2_1 _0883_ (.A(net56),
    .B(net320),
    .Y(_0072_));
 sg13g2_nor2b_1 _0884_ (.A(\rs232out_inst.ttyclk[14] ),
    .B_N(_0318_),
    .Y(_0320_));
 sg13g2_xnor2_1 _0885_ (.Y(_0321_),
    .A(net278),
    .B(_0318_));
 sg13g2_nor2_1 _0886_ (.A(net56),
    .B(net279),
    .Y(_0073_));
 sg13g2_nor2_1 _0887_ (.A(net255),
    .B(_0320_),
    .Y(_0322_));
 sg13g2_a21oi_1 _0888_ (.A1(net255),
    .A2(_0320_),
    .Y(_0323_),
    .B1(net56));
 sg13g2_nor2b_1 _0889_ (.A(net256),
    .B_N(_0323_),
    .Y(_0074_));
 sg13g2_nor2b_1 _0890_ (.A(net73),
    .B_N(net178),
    .Y(_0324_));
 sg13g2_a21oi_1 _0891_ (.A1(net73),
    .A2(\rs232out_inst.transmit_data[0] ),
    .Y(_0325_),
    .B1(_0324_));
 sg13g2_nand2_1 _0892_ (.Y(_0326_),
    .A(net188),
    .B(net60));
 sg13g2_o21ai_1 _0893_ (.B1(_0326_),
    .Y(_0075_),
    .A1(net60),
    .A2(_0325_));
 sg13g2_nor2b_1 _0894_ (.A(net73),
    .B_N(\rs232out_inst.shift_out[3] ),
    .Y(_0327_));
 sg13g2_a21oi_1 _0895_ (.A1(net73),
    .A2(\rs232out_inst.transmit_data[1] ),
    .Y(_0328_),
    .B1(_0327_));
 sg13g2_nand2_1 _0896_ (.Y(_0329_),
    .A(net178),
    .B(net60));
 sg13g2_o21ai_1 _0897_ (.B1(_0329_),
    .Y(_0076_),
    .A1(net60),
    .A2(_0328_));
 sg13g2_nor2b_1 _0898_ (.A(net72),
    .B_N(net172),
    .Y(_0330_));
 sg13g2_a21oi_1 _0899_ (.A1(net72),
    .A2(\rs232out_inst.transmit_data[2] ),
    .Y(_0331_),
    .B1(_0330_));
 sg13g2_nand2_1 _0900_ (.Y(_0332_),
    .A(net180),
    .B(net59));
 sg13g2_o21ai_1 _0901_ (.B1(_0332_),
    .Y(_0077_),
    .A1(net59),
    .A2(_0331_));
 sg13g2_nor2b_1 _0902_ (.A(net72),
    .B_N(\rs232out_inst.shift_out[5] ),
    .Y(_0333_));
 sg13g2_a21oi_1 _0903_ (.A1(net72),
    .A2(\rs232out_inst.transmit_data[3] ),
    .Y(_0334_),
    .B1(_0333_));
 sg13g2_nand2_1 _0904_ (.Y(_0335_),
    .A(net172),
    .B(net59));
 sg13g2_o21ai_1 _0905_ (.B1(_0335_),
    .Y(_0078_),
    .A1(net59),
    .A2(_0334_));
 sg13g2_nor2b_1 _0906_ (.A(net72),
    .B_N(net186),
    .Y(_0336_));
 sg13g2_a21oi_1 _0907_ (.A1(net72),
    .A2(\rs232out_inst.transmit_data[4] ),
    .Y(_0337_),
    .B1(_0336_));
 sg13g2_nand2_1 _0908_ (.Y(_0338_),
    .A(net190),
    .B(net59));
 sg13g2_o21ai_1 _0909_ (.B1(_0338_),
    .Y(_0079_),
    .A1(net59),
    .A2(_0337_));
 sg13g2_nor2b_1 _0910_ (.A(net72),
    .B_N(\rs232out_inst.shift_out[7] ),
    .Y(_0339_));
 sg13g2_a21oi_1 _0911_ (.A1(net72),
    .A2(\rs232out_inst.transmit_data[5] ),
    .Y(_0340_),
    .B1(_0339_));
 sg13g2_nand2_1 _0912_ (.Y(_0341_),
    .A(net186),
    .B(net59));
 sg13g2_o21ai_1 _0913_ (.B1(_0341_),
    .Y(_0080_),
    .A1(net59),
    .A2(_0340_));
 sg13g2_nor2b_1 _0914_ (.A(net74),
    .B_N(\rs232out_inst.shift_out[8] ),
    .Y(_0342_));
 sg13g2_a21oi_1 _0915_ (.A1(net74),
    .A2(net184),
    .Y(_0343_),
    .B1(_0342_));
 sg13g2_nand2_1 _0916_ (.Y(_0344_),
    .A(net192),
    .B(net61));
 sg13g2_o21ai_1 _0917_ (.B1(_0344_),
    .Y(_0081_),
    .A1(net61),
    .A2(_0343_));
 sg13g2_a22oi_1 _0918_ (.Y(_0345_),
    .B1(net60),
    .B2(net176),
    .A2(_0267_),
    .A1(\rs232out_inst.shift_out[1] ));
 sg13g2_inv_1 _0919_ (.Y(_0082_),
    .A(net177));
 sg13g2_a22oi_1 _0920_ (.Y(_0083_),
    .B1(net61),
    .B2(_0128_),
    .A2(_0267_),
    .A1(_0129_));
 sg13g2_nand2_1 _0921_ (.Y(_0346_),
    .A(net202),
    .B(_0289_));
 sg13g2_xor2_1 _0922_ (.B(net210),
    .A(\rs232out_inst.count[0] ),
    .X(_0347_));
 sg13g2_nand2_1 _0923_ (.Y(_0348_),
    .A(net210),
    .B(net61));
 sg13g2_o21ai_1 _0924_ (.B1(_0348_),
    .Y(_0084_),
    .A1(_0346_),
    .A2(_0347_));
 sg13g2_nor2b_1 _0925_ (.A(_0265_),
    .B_N(net202),
    .Y(_0349_));
 sg13g2_o21ai_1 _0926_ (.B1(\rs232out_inst.count[2] ),
    .Y(_0350_),
    .A1(net61),
    .A2(_0349_));
 sg13g2_o21ai_1 _0927_ (.B1(_0350_),
    .Y(_0085_),
    .A1(_0266_),
    .A2(_0346_));
 sg13g2_o21ai_1 _0928_ (.B1(net207),
    .Y(_0351_),
    .A1(_0266_),
    .A2(net61));
 sg13g2_o21ai_1 _0929_ (.B1(_0289_),
    .Y(_0352_),
    .A1(net74),
    .A2(_0268_));
 sg13g2_nand2_1 _0930_ (.Y(_0086_),
    .A(net208),
    .B(_0352_));
 sg13g2_nor2_2 _0931_ (.A(_0002_),
    .B(_0149_),
    .Y(_0353_));
 sg13g2_mux2_1 _0932_ (.A0(net200),
    .A1(net214),
    .S(net242),
    .X(_0087_));
 sg13g2_mux2_1 _0933_ (.A0(net214),
    .A1(net239),
    .S(net242),
    .X(_0088_));
 sg13g2_mux2_1 _0934_ (.A0(net239),
    .A1(net231),
    .S(net242),
    .X(_0089_));
 sg13g2_mux2_1 _0935_ (.A0(net231),
    .A1(net215),
    .S(net242),
    .X(_0090_));
 sg13g2_mux2_1 _0936_ (.A0(net215),
    .A1(net251),
    .S(net242),
    .X(_0091_));
 sg13g2_mux2_1 _0937_ (.A0(net251),
    .A1(\rs232in_inst.shift_in[7] ),
    .S(net242),
    .X(_0092_));
 sg13g2_nor2_1 _0938_ (.A(net271),
    .B(net242),
    .Y(_0354_));
 sg13g2_a21oi_1 _0939_ (.A1(_0126_),
    .A2(net242),
    .Y(_0093_),
    .B1(_0354_));
 sg13g2_nand2_1 _0940_ (.Y(_0355_),
    .A(\rs232in_inst.ttyclk[0] ),
    .B(net57));
 sg13g2_nand2b_1 _0941_ (.Y(_0356_),
    .B(net198),
    .A_N(net69));
 sg13g2_nand4_1 _0942_ (.B(_0126_),
    .C(net243),
    .A(net70),
    .Y(_0357_),
    .D(_0149_));
 sg13g2_nand3_1 _0943_ (.B(_0356_),
    .C(_0357_),
    .A(_0355_),
    .Y(_0094_));
 sg13g2_nand2b_1 _0944_ (.Y(_0358_),
    .B(net241),
    .A_N(net57));
 sg13g2_xor2_1 _0945_ (.B(net303),
    .A(\rs232in_inst.ttyclk[0] ),
    .X(_0359_));
 sg13g2_nand2_1 _0946_ (.Y(_0360_),
    .A(net303),
    .B(net57));
 sg13g2_o21ai_1 _0947_ (.B1(_0360_),
    .Y(_0095_),
    .A1(_0358_),
    .A2(_0359_));
 sg13g2_xnor2_1 _0948_ (.Y(_0361_),
    .A(net269),
    .B(_0152_));
 sg13g2_nand2_1 _0949_ (.Y(_0362_),
    .A(net269),
    .B(net57));
 sg13g2_o21ai_1 _0950_ (.B1(_0362_),
    .Y(_0096_),
    .A1(_0358_),
    .A2(_0361_));
 sg13g2_o21ai_1 _0951_ (.B1(net70),
    .Y(_0363_),
    .A1(_0126_),
    .A2(_0150_));
 sg13g2_or4_1 _0952_ (.A(net69),
    .B(\rs232in_inst.ttyclk[0] ),
    .C(\rs232in_inst.ttyclk[1] ),
    .D(net367),
    .X(_0364_));
 sg13g2_nand3_1 _0953_ (.B(_0363_),
    .C(_0364_),
    .A(net250),
    .Y(_0365_));
 sg13g2_o21ai_1 _0954_ (.B1(_0357_),
    .Y(_0366_),
    .A1(net69),
    .A2(_0154_));
 sg13g2_nand2b_1 _0955_ (.Y(_0097_),
    .B(_0365_),
    .A_N(_0366_));
 sg13g2_nand2_1 _0956_ (.Y(_0367_),
    .A(net69),
    .B(_0150_));
 sg13g2_nand2_1 _0957_ (.Y(_0368_),
    .A(_0010_),
    .B(_0153_));
 sg13g2_xnor2_1 _0958_ (.Y(_0369_),
    .A(_0010_),
    .B(_0154_));
 sg13g2_o21ai_1 _0959_ (.B1(_0367_),
    .Y(_0370_),
    .A1(net71),
    .A2(_0369_));
 sg13g2_a21o_1 _0960_ (.A2(net57),
    .A1(net296),
    .B1(_0370_),
    .X(_0098_));
 sg13g2_o21ai_1 _0961_ (.B1(net71),
    .Y(_0371_),
    .A1(net273),
    .A2(_0150_));
 sg13g2_nor2_1 _0962_ (.A(net340),
    .B(_0150_),
    .Y(_0372_));
 sg13g2_xnor2_1 _0963_ (.Y(_0373_),
    .A(net340),
    .B(_0368_));
 sg13g2_nand2b_1 _0964_ (.Y(_0374_),
    .B(_0373_),
    .A_N(net71));
 sg13g2_o21ai_1 _0965_ (.B1(_0374_),
    .Y(_0099_),
    .A1(_0371_),
    .A2(net341));
 sg13g2_nor2_2 _0966_ (.A(net241),
    .B(_0151_),
    .Y(_0375_));
 sg13g2_nor4_1 _0967_ (.A(\rs232in_inst.ttyclk[4] ),
    .B(\rs232in_inst.ttyclk[5] ),
    .C(net57),
    .D(_0154_),
    .Y(_0376_));
 sg13g2_xnor2_1 _0968_ (.Y(_0377_),
    .A(net274),
    .B(_0376_));
 sg13g2_nor2_1 _0969_ (.A(_0375_),
    .B(net275),
    .Y(_0100_));
 sg13g2_nand2b_1 _0970_ (.Y(_0378_),
    .B(\rs232in_inst.ttyclk[7] ),
    .A_N(_0155_));
 sg13g2_a21oi_1 _0971_ (.A1(_0157_),
    .A2(_0378_),
    .Y(_0379_),
    .B1(net71));
 sg13g2_a21oi_1 _0972_ (.A1(net71),
    .A2(net243),
    .Y(_0380_),
    .B1(_0379_));
 sg13g2_a22oi_1 _0973_ (.Y(_0101_),
    .B1(_0371_),
    .B2(net244),
    .A2(_0151_),
    .A1(_0131_));
 sg13g2_or3_1 _0974_ (.A(net69),
    .B(_0011_),
    .C(_0156_),
    .X(_0381_));
 sg13g2_nand2_1 _0975_ (.Y(_0382_),
    .A(net314),
    .B(_0151_));
 sg13g2_nand3b_1 _0976_ (.B(_0011_),
    .C(_0156_),
    .Y(_0383_),
    .A_N(net69));
 sg13g2_nand4_1 _0977_ (.B(_0381_),
    .C(net315),
    .A(_0367_),
    .Y(_0102_),
    .D(_0383_));
 sg13g2_or2_1 _0978_ (.X(_0384_),
    .B(_0383_),
    .A(net305));
 sg13g2_nand3_1 _0979_ (.B(_0363_),
    .C(_0383_),
    .A(net305),
    .Y(_0385_));
 sg13g2_nand3_1 _0980_ (.B(_0384_),
    .C(net306),
    .A(_0357_),
    .Y(_0103_));
 sg13g2_nor3_2 _0981_ (.A(net57),
    .B(_0157_),
    .C(_0158_),
    .Y(_0386_));
 sg13g2_nand2b_1 _0982_ (.Y(_0387_),
    .B(_0386_),
    .A_N(net284));
 sg13g2_xnor2_1 _0983_ (.Y(_0388_),
    .A(net284),
    .B(_0386_));
 sg13g2_nor2_1 _0984_ (.A(_0375_),
    .B(net285),
    .Y(_0104_));
 sg13g2_xor2_1 _0985_ (.B(_0387_),
    .A(net317),
    .X(_0389_));
 sg13g2_nor2_1 _0986_ (.A(_0375_),
    .B(_0389_),
    .Y(_0105_));
 sg13g2_nand2_2 _0987_ (.Y(_0390_),
    .A(_0160_),
    .B(_0386_));
 sg13g2_o21ai_1 _0988_ (.B1(net234),
    .Y(_0391_),
    .A1(\rs232in_inst.ttyclk[11] ),
    .A2(_0387_));
 sg13g2_a21oi_1 _0989_ (.A1(_0390_),
    .A2(net235),
    .Y(_0106_),
    .B1(_0375_));
 sg13g2_xor2_1 _0990_ (.B(_0390_),
    .A(net330),
    .X(_0392_));
 sg13g2_nor2_1 _0991_ (.A(_0375_),
    .B(_0392_),
    .Y(_0107_));
 sg13g2_nor3_1 _0992_ (.A(net330),
    .B(net339),
    .C(_0390_),
    .Y(_0393_));
 sg13g2_o21ai_1 _0993_ (.B1(net339),
    .Y(_0394_),
    .A1(net330),
    .A2(_0390_));
 sg13g2_nor2b_1 _0994_ (.A(_0393_),
    .B_N(_0394_),
    .Y(_0395_));
 sg13g2_nor2_1 _0995_ (.A(_0375_),
    .B(_0395_),
    .Y(_0108_));
 sg13g2_xnor2_1 _0996_ (.Y(_0396_),
    .A(net246),
    .B(_0393_));
 sg13g2_nor2_1 _0997_ (.A(_0375_),
    .B(net247),
    .Y(_0109_));
 sg13g2_nand2_1 _0998_ (.Y(_0397_),
    .A(\rs232in_inst.count[0] ),
    .B(_0148_));
 sg13g2_nand4_1 _0999_ (.B(_0125_),
    .C(net70),
    .A(net253),
    .Y(_0398_),
    .D(_0148_));
 sg13g2_mux2_1 _1000_ (.A0(net200),
    .A1(\rs232in_inst.received_data[0] ),
    .S(net58),
    .X(_0110_));
 sg13g2_mux2_1 _1001_ (.A0(net214),
    .A1(net254),
    .S(net58),
    .X(_0111_));
 sg13g2_mux2_1 _1002_ (.A0(net239),
    .A1(\rs232in_inst.received_data[2] ),
    .S(net58),
    .X(_0112_));
 sg13g2_mux2_1 _1003_ (.A0(net231),
    .A1(\rs232in_inst.received_data[3] ),
    .S(net58),
    .X(_0113_));
 sg13g2_nor2_1 _1004_ (.A(net215),
    .B(net58),
    .Y(_0399_));
 sg13g2_a21oi_1 _1005_ (.A1(_0132_),
    .A2(net58),
    .Y(_0114_),
    .B1(_0399_));
 sg13g2_mux2_1 _1006_ (.A0(net251),
    .A1(net266),
    .S(net58),
    .X(_0115_));
 sg13g2_mux2_1 _1007_ (.A0(net271),
    .A1(\rs232in_inst.received_data[6] ),
    .S(_0398_),
    .X(_0116_));
 sg13g2_nand2_1 _1008_ (.Y(_0400_),
    .A(net220),
    .B(net58));
 sg13g2_o21ai_1 _1009_ (.B1(_0400_),
    .Y(_0117_),
    .A1(_0126_),
    .A2(_0398_));
 sg13g2_nor3_1 _1010_ (.A(net170),
    .B(_0002_),
    .C(_0397_),
    .Y(_0118_));
 sg13g2_nand3_1 _1011_ (.B(net69),
    .C(_0150_),
    .A(net164),
    .Y(_0401_));
 sg13g2_o21ai_1 _1012_ (.B1(_0401_),
    .Y(_0119_),
    .A1(_0124_),
    .A2(net69));
 sg13g2_o21ai_1 _1013_ (.B1(net170),
    .Y(_0402_),
    .A1(net253),
    .A2(_0363_));
 sg13g2_o21ai_1 _1014_ (.B1(_0402_),
    .Y(_0120_),
    .A1(_0147_),
    .A2(_0367_));
 sg13g2_o21ai_1 _1015_ (.B1(net291),
    .Y(_0403_),
    .A1(_0147_),
    .A2(_0363_));
 sg13g2_or3_1 _1016_ (.A(net291),
    .B(_0147_),
    .C(_0363_),
    .X(_0404_));
 sg13g2_a21oi_1 _1017_ (.A1(_0403_),
    .A2(_0404_),
    .Y(_0121_),
    .B1(_0148_));
 sg13g2_xnor2_1 _1018_ (.Y(_0122_),
    .A(net267),
    .B(_0404_));
 sg13g2_o21ai_1 _1019_ (.B1(net174),
    .Y(_0405_),
    .A1(\rs232in_inst.count[3] ),
    .A2(_0404_));
 sg13g2_inv_1 _1020_ (.Y(_0123_),
    .A(net175));
 sg13g2_dfrbp_1 _1021_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net99),
    .D(_0032_),
    .Q_N(_0485_),
    .Q(\pdm_inst.level[0] ));
 sg13g2_dfrbp_1 _1022_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net31),
    .D(_0033_),
    .Q_N(_0484_),
    .Q(\pdm_inst.level[1] ));
 sg13g2_dfrbp_1 _1023_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net30),
    .D(net302),
    .Q_N(_0483_),
    .Q(\pdm_inst.level[2] ));
 sg13g2_dfrbp_1 _1024_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net144),
    .D(net283),
    .Q_N(_0482_),
    .Q(\pdm_inst.level[3] ));
 sg13g2_dfrbp_1 _1025_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net143),
    .D(net281),
    .Q_N(_0481_),
    .Q(\pdm_inst.level[4] ));
 sg13g2_dfrbp_1 _1026_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net142),
    .D(_0037_),
    .Q_N(_0480_),
    .Q(\pdm_inst.level[5] ));
 sg13g2_dfrbp_1 _1027_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net141),
    .D(_0038_),
    .Q_N(_0479_),
    .Q(\pdm_inst.level[6] ));
 sg13g2_dfrbp_1 _1028_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net140),
    .D(_0039_),
    .Q_N(_0478_),
    .Q(\pdm_inst.level[7] ));
 sg13g2_dfrbp_1 _1029_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net139),
    .D(net277),
    .Q_N(_0477_),
    .Q(\pdm_inst.level[8] ));
 sg13g2_dfrbp_1 _1030_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net138),
    .D(net327),
    .Q_N(_0476_),
    .Q(\pdm_inst.level[9] ));
 sg13g2_dfrbp_1 _1031_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net137),
    .D(net329),
    .Q_N(_0475_),
    .Q(\pdm_inst.level[10] ));
 sg13g2_dfrbp_1 _1032_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net136),
    .D(net299),
    .Q_N(_0474_),
    .Q(\pdm_inst.level[11] ));
 sg13g2_dfrbp_1 _1033_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net135),
    .D(_0044_),
    .Q_N(_0473_),
    .Q(\pdm_inst.level[12] ));
 sg13g2_dfrbp_1 _1034_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net134),
    .D(net287),
    .Q_N(_0472_),
    .Q(\pdm_inst.level[13] ));
 sg13g2_dfrbp_1 _1035_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net133),
    .D(net309),
    .Q_N(_0471_),
    .Q(\pdm_inst.level[14] ));
 sg13g2_dfrbp_1 _1036_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net132),
    .D(net290),
    .Q_N(_0470_),
    .Q(\pdm_inst.level[15] ));
 sg13g2_dfrbp_1 _1037_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net131),
    .D(_0048_),
    .Q_N(_0006_),
    .Q(\rs232out_inst.count[4] ));
 sg13g2_dfrbp_1 _1038_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net130),
    .D(net167),
    .Q_N(_0469_),
    .Q(\rs232out_inst.transmit_data[0] ));
 sg13g2_dfrbp_1 _1039_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net129),
    .D(net195),
    .Q_N(_0468_),
    .Q(\rs232out_inst.transmit_data[1] ));
 sg13g2_dfrbp_1 _1040_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net128),
    .D(net213),
    .Q_N(_0467_),
    .Q(\rs232out_inst.transmit_data[2] ));
 sg13g2_dfrbp_1 _1041_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net127),
    .D(net259),
    .Q_N(_0466_),
    .Q(\rs232out_inst.transmit_data[3] ));
 sg13g2_dfrbp_1 _1042_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net126),
    .D(net197),
    .Q_N(_0465_),
    .Q(\rs232out_inst.transmit_data[4] ));
 sg13g2_dfrbp_1 _1043_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net125),
    .D(net227),
    .Q_N(_0464_),
    .Q(\rs232out_inst.transmit_data[5] ));
 sg13g2_dfrbp_1 _1044_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net124),
    .D(net185),
    .Q_N(_0463_),
    .Q(\rs232out_inst.transmit_data[6] ));
 sg13g2_dfrbp_1 _1045_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net123),
    .D(net295),
    .Q_N(_0462_),
    .Q(\rs232out_inst.transmit_data[7] ));
 sg13g2_dfrbp_1 _1046_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net122),
    .D(_0057_),
    .Q_N(_0007_),
    .Q(\rs232out_inst.we ));
 sg13g2_dfrbp_1 _1047_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net121),
    .D(net249),
    .Q_N(_0461_),
    .Q(\rs232out_inst.shift_out[8] ));
 sg13g2_dfrbp_1 _1048_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net119),
    .D(net238),
    .Q_N(_0460_),
    .Q(\rs232out_inst.ttyclk[0] ));
 sg13g2_dfrbp_1 _1049_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net118),
    .D(net219),
    .Q_N(_0459_),
    .Q(\rs232out_inst.ttyclk[1] ));
 sg13g2_dfrbp_1 _1050_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net117),
    .D(_0061_),
    .Q_N(_0458_),
    .Q(\rs232out_inst.ttyclk[2] ));
 sg13g2_dfrbp_1 _1051_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net116),
    .D(net262),
    .Q_N(_0457_),
    .Q(\rs232out_inst.ttyclk[3] ));
 sg13g2_dfrbp_1 _1052_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net115),
    .D(net206),
    .Q_N(_0004_),
    .Q(\rs232out_inst.ttyclk[4] ));
 sg13g2_dfrbp_1 _1053_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net114),
    .D(_0064_),
    .Q_N(_0456_),
    .Q(\rs232out_inst.ttyclk[5] ));
 sg13g2_dfrbp_1 _1054_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net113),
    .D(net225),
    .Q_N(_0455_),
    .Q(\rs232out_inst.ttyclk[6] ));
 sg13g2_dfrbp_1 _1055_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net112),
    .D(net293),
    .Q_N(_0454_),
    .Q(\rs232out_inst.ttyclk[7] ));
 sg13g2_dfrbp_1 _1056_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net111),
    .D(_0067_),
    .Q_N(_0453_),
    .Q(\rs232out_inst.ttyclk[8] ));
 sg13g2_dfrbp_1 _1057_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net110),
    .D(_0068_),
    .Q_N(_0452_),
    .Q(\rs232out_inst.ttyclk[9] ));
 sg13g2_dfrbp_1 _1058_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net109),
    .D(net265),
    .Q_N(_0451_),
    .Q(\rs232out_inst.ttyclk[10] ));
 sg13g2_dfrbp_1 _1059_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net108),
    .D(_0070_),
    .Q_N(_0450_),
    .Q(\rs232out_inst.ttyclk[11] ));
 sg13g2_dfrbp_1 _1060_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net105),
    .D(_0071_),
    .Q_N(_0449_),
    .Q(\rs232out_inst.ttyclk[12] ));
 sg13g2_dfrbp_1 _1061_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net104),
    .D(_0072_),
    .Q_N(_0448_),
    .Q(\rs232out_inst.ttyclk[13] ));
 sg13g2_dfrbp_1 _1062_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net103),
    .D(_0073_),
    .Q_N(_0447_),
    .Q(\rs232out_inst.ttyclk[14] ));
 sg13g2_dfrbp_1 _1063_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net102),
    .D(net257),
    .Q_N(_0446_),
    .Q(\rs232out_inst.ttyclk[15] ));
 sg13g2_dfrbp_1 _1064_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net100),
    .D(net189),
    .Q_N(_0445_),
    .Q(\rs232out_inst.shift_out[1] ));
 sg13g2_dfrbp_1 _1065_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net98),
    .D(net179),
    .Q_N(_0444_),
    .Q(\rs232out_inst.shift_out[2] ));
 sg13g2_dfrbp_1 _1066_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net97),
    .D(net181),
    .Q_N(_0443_),
    .Q(\rs232out_inst.shift_out[3] ));
 sg13g2_dfrbp_1 _1067_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net96),
    .D(net173),
    .Q_N(_0442_),
    .Q(\rs232out_inst.shift_out[4] ));
 sg13g2_dfrbp_1 _1068_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net95),
    .D(net191),
    .Q_N(_0441_),
    .Q(\rs232out_inst.shift_out[5] ));
 sg13g2_dfrbp_1 _1069_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net94),
    .D(net187),
    .Q_N(_0440_),
    .Q(\rs232out_inst.shift_out[6] ));
 sg13g2_dfrbp_1 _1070_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net101),
    .D(net193),
    .Q_N(_0486_),
    .Q(\rs232out_inst.shift_out[7] ));
 sg13g2_dfrbp_1 _1071_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net93),
    .D(_0000_),
    .Q_N(_0002_),
    .Q(\rs232in_inst.ttyclk[16] ));
 sg13g2_dfrbp_1 _1072_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net106),
    .D(_0082_),
    .Q_N(_0487_),
    .Q(\rs232out_inst.serial_out ));
 sg13g2_dfrbp_1 _1073_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net92),
    .D(net333),
    .Q_N(_0003_),
    .Q(\rs232out_inst.ttyclk[16] ));
 sg13g2_dfrbp_1 _1074_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net90),
    .D(net169),
    .Q_N(_0005_),
    .Q(\rs232out_inst.count[0] ));
 sg13g2_dfrbp_1 _1075_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net89),
    .D(net211),
    .Q_N(_0439_),
    .Q(\rs232out_inst.count[1] ));
 sg13g2_dfrbp_1 _1076_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net88),
    .D(net203),
    .Q_N(_0438_),
    .Q(\rs232out_inst.count[2] ));
 sg13g2_dfrbp_1 _1077_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net107),
    .D(net209),
    .Q_N(_0488_),
    .Q(\rs232out_inst.count[3] ));
 sg13g2_dfrbp_1 _1078_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net145),
    .D(net163),
    .Q_N(_0009_),
    .Q(\rs232in_inst.rxd2 ));
 sg13g2_dfrbp_1 _1079_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net87),
    .D(net2),
    .Q_N(_0437_),
    .Q(\rs232in_inst.rxd ));
 sg13g2_dfrbp_1 _1080_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net86),
    .D(_0087_),
    .Q_N(_0436_),
    .Q(\rs232in_inst.shift_in[1] ));
 sg13g2_dfrbp_1 _1081_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net85),
    .D(_0088_),
    .Q_N(_0435_),
    .Q(\rs232in_inst.shift_in[2] ));
 sg13g2_dfrbp_1 _1082_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net84),
    .D(_0089_),
    .Q_N(_0434_),
    .Q(\rs232in_inst.shift_in[3] ));
 sg13g2_dfrbp_1 _1083_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net83),
    .D(_0090_),
    .Q_N(_0433_),
    .Q(\rs232in_inst.shift_in[4] ));
 sg13g2_dfrbp_1 _1084_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net82),
    .D(_0091_),
    .Q_N(_0432_),
    .Q(\rs232in_inst.shift_in[5] ));
 sg13g2_dfrbp_1 _1085_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net81),
    .D(net252),
    .Q_N(_0431_),
    .Q(\rs232in_inst.shift_in[6] ));
 sg13g2_dfrbp_1 _1086_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net80),
    .D(_0093_),
    .Q_N(_0430_),
    .Q(\rs232in_inst.shift_in[7] ));
 sg13g2_dfrbp_1 _1087_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net79),
    .D(net199),
    .Q_N(_0008_),
    .Q(\rs232in_inst.ttyclk[0] ));
 sg13g2_dfrbp_1 _1088_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net78),
    .D(net304),
    .Q_N(_0429_),
    .Q(\rs232in_inst.ttyclk[1] ));
 sg13g2_dfrbp_1 _1089_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net77),
    .D(net270),
    .Q_N(_0428_),
    .Q(\rs232in_inst.ttyclk[2] ));
 sg13g2_dfrbp_1 _1090_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net76),
    .D(_0097_),
    .Q_N(_0427_),
    .Q(\rs232in_inst.ttyclk[3] ));
 sg13g2_dfrbp_1 _1091_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net75),
    .D(net297),
    .Q_N(_0010_),
    .Q(\rs232in_inst.ttyclk[4] ));
 sg13g2_dfrbp_1 _1092_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net55),
    .D(net342),
    .Q_N(_0426_),
    .Q(\rs232in_inst.ttyclk[5] ));
 sg13g2_dfrbp_1 _1093_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net54),
    .D(_0100_),
    .Q_N(_0425_),
    .Q(\rs232in_inst.ttyclk[6] ));
 sg13g2_dfrbp_1 _1094_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net53),
    .D(net245),
    .Q_N(_0424_),
    .Q(\rs232in_inst.ttyclk[7] ));
 sg13g2_dfrbp_1 _1095_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net52),
    .D(net316),
    .Q_N(_0011_),
    .Q(\rs232in_inst.ttyclk[8] ));
 sg13g2_dfrbp_1 _1096_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net51),
    .D(net307),
    .Q_N(_0423_),
    .Q(\rs232in_inst.ttyclk[9] ));
 sg13g2_dfrbp_1 _1097_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net50),
    .D(_0104_),
    .Q_N(_0422_),
    .Q(\rs232in_inst.ttyclk[10] ));
 sg13g2_dfrbp_1 _1098_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net49),
    .D(_0105_),
    .Q_N(_0421_),
    .Q(\rs232in_inst.ttyclk[11] ));
 sg13g2_dfrbp_1 _1099_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net48),
    .D(net236),
    .Q_N(_0420_),
    .Q(\rs232in_inst.ttyclk[12] ));
 sg13g2_dfrbp_1 _1100_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net47),
    .D(_0107_),
    .Q_N(_0419_),
    .Q(\rs232in_inst.ttyclk[13] ));
 sg13g2_dfrbp_1 _1101_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net46),
    .D(_0108_),
    .Q_N(_0418_),
    .Q(\rs232in_inst.ttyclk[14] ));
 sg13g2_dfrbp_1 _1102_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net45),
    .D(_0109_),
    .Q_N(_0417_),
    .Q(\rs232in_inst.ttyclk[15] ));
 sg13g2_dfrbp_1 _1103_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net44),
    .D(net201),
    .Q_N(_0031_),
    .Q(\rs232in_inst.received_data[0] ));
 sg13g2_dfrbp_1 _1104_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net43),
    .D(_0111_),
    .Q_N(_0416_),
    .Q(\rs232in_inst.received_data[1] ));
 sg13g2_dfrbp_1 _1105_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net42),
    .D(net240),
    .Q_N(_0415_),
    .Q(\rs232in_inst.received_data[2] ));
 sg13g2_dfrbp_1 _1106_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net41),
    .D(net232),
    .Q_N(_0414_),
    .Q(\rs232in_inst.received_data[3] ));
 sg13g2_dfrbp_1 _1107_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net40),
    .D(net216),
    .Q_N(_0413_),
    .Q(\rs232in_inst.received_data[4] ));
 sg13g2_dfrbp_1 _1108_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net39),
    .D(_0115_),
    .Q_N(_0412_),
    .Q(\rs232in_inst.received_data[5] ));
 sg13g2_dfrbp_1 _1109_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net38),
    .D(net272),
    .Q_N(_0411_),
    .Q(\rs232in_inst.received_data[6] ));
 sg13g2_dfrbp_1 _1110_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net37),
    .D(net221),
    .Q_N(_0410_),
    .Q(\rs232in_inst.received_data[7] ));
 sg13g2_dfrbp_1 _1111_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net36),
    .D(net171),
    .Q_N(_0409_),
    .Q(\rs232in_inst.attention ));
 sg13g2_dfrbp_1 _1112_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net35),
    .D(net165),
    .Q_N(_0030_),
    .Q(\rs232in_inst.count[0] ));
 sg13g2_dfrbp_1 _1113_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net33),
    .D(_0120_),
    .Q_N(_0408_),
    .Q(\rs232in_inst.count[1] ));
 sg13g2_dfrbp_1 _1114_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net120),
    .D(_0121_),
    .Q_N(_0407_),
    .Q(\rs232in_inst.count[2] ));
 sg13g2_dfrbp_1 _1115_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net34),
    .D(net268),
    .Q_N(_0406_),
    .Q(\rs232in_inst.count[3] ));
 sg13g2_dfrbp_1 _1116_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net146),
    .D(_0123_),
    .Q_N(_0489_),
    .Q(\rs232in_inst.count[4] ));
 sg13g2_dfrbp_1 _1117_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net147),
    .D(net183),
    .Q_N(_0490_),
    .Q(\pdm_inst.sigma[0] ));
 sg13g2_dfrbp_1 _1118_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net148),
    .D(_0021_),
    .Q_N(_0491_),
    .Q(\pdm_inst.sigma[1] ));
 sg13g2_dfrbp_1 _1119_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net149),
    .D(_0022_),
    .Q_N(_0492_),
    .Q(\pdm_inst.sigma[2] ));
 sg13g2_dfrbp_1 _1120_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net150),
    .D(net344),
    .Q_N(_0493_),
    .Q(\pdm_inst.sigma[3] ));
 sg13g2_dfrbp_1 _1121_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net151),
    .D(_0024_),
    .Q_N(_0494_),
    .Q(\pdm_inst.sigma[4] ));
 sg13g2_dfrbp_1 _1122_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net152),
    .D(net335),
    .Q_N(_0495_),
    .Q(\pdm_inst.sigma[5] ));
 sg13g2_dfrbp_1 _1123_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net153),
    .D(_0026_),
    .Q_N(_0496_),
    .Q(\pdm_inst.sigma[6] ));
 sg13g2_dfrbp_1 _1124_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net154),
    .D(net365),
    .Q_N(_0497_),
    .Q(\pdm_inst.sigma[7] ));
 sg13g2_dfrbp_1 _1125_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net155),
    .D(_0028_),
    .Q_N(_0498_),
    .Q(\pdm_inst.sigma[8] ));
 sg13g2_dfrbp_1 _1126_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net156),
    .D(net347),
    .Q_N(_0499_),
    .Q(\pdm_inst.sigma[9] ));
 sg13g2_dfrbp_1 _1127_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net157),
    .D(_0013_),
    .Q_N(_0500_),
    .Q(\pdm_inst.sigma[10] ));
 sg13g2_dfrbp_1 _1128_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net158),
    .D(net362),
    .Q_N(_0501_),
    .Q(\pdm_inst.sigma[11] ));
 sg13g2_dfrbp_1 _1129_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net159),
    .D(_0015_),
    .Q_N(_0502_),
    .Q(\pdm_inst.sigma[12] ));
 sg13g2_dfrbp_1 _1130_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net160),
    .D(_0016_),
    .Q_N(_0503_),
    .Q(\pdm_inst.sigma[13] ));
 sg13g2_dfrbp_1 _1131_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net161),
    .D(net352),
    .Q_N(_0504_),
    .Q(\pdm_inst.sigma[14] ));
 sg13g2_dfrbp_1 _1132_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net162),
    .D(net349),
    .Q_N(_0505_),
    .Q(\pdm_inst.sigma[15] ));
 sg13g2_dfrbp_1 _1133_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net32),
    .D(net338),
    .Q_N(_0506_),
    .Q(\pdm_inst.sigma[16] ));
 sg13g2_dfrbp_1 _1134_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net91),
    .D(net230),
    .Q_N(\pdm_inst.O ),
    .Q(\pdm_inst.sigma[17] ));
 sg13g2_tiehi _1022__31 (.L_HI(net31));
 sg13g2_tiehi _1133__32 (.L_HI(net32));
 sg13g2_tiehi _1113__33 (.L_HI(net33));
 sg13g2_tiehi _1115__34 (.L_HI(net34));
 sg13g2_tiehi _1112__35 (.L_HI(net35));
 sg13g2_tiehi _1111__36 (.L_HI(net36));
 sg13g2_tiehi _1110__37 (.L_HI(net37));
 sg13g2_tiehi _1109__38 (.L_HI(net38));
 sg13g2_tiehi _1108__39 (.L_HI(net39));
 sg13g2_tiehi _1107__40 (.L_HI(net40));
 sg13g2_tiehi _1106__41 (.L_HI(net41));
 sg13g2_tiehi _1105__42 (.L_HI(net42));
 sg13g2_tiehi _1104__43 (.L_HI(net43));
 sg13g2_tiehi _1103__44 (.L_HI(net44));
 sg13g2_tiehi _1102__45 (.L_HI(net45));
 sg13g2_tiehi _1101__46 (.L_HI(net46));
 sg13g2_tiehi _1100__47 (.L_HI(net47));
 sg13g2_tiehi _1099__48 (.L_HI(net48));
 sg13g2_tiehi _1098__49 (.L_HI(net49));
 sg13g2_tiehi _1097__50 (.L_HI(net50));
 sg13g2_tiehi _1096__51 (.L_HI(net51));
 sg13g2_tiehi _1095__52 (.L_HI(net52));
 sg13g2_tiehi _1094__53 (.L_HI(net53));
 sg13g2_tiehi _1093__54 (.L_HI(net54));
 sg13g2_tiehi _1092__55 (.L_HI(net55));
 sg13g2_tiehi _1091__56 (.L_HI(net75));
 sg13g2_tiehi _1090__57 (.L_HI(net76));
 sg13g2_tiehi _1089__58 (.L_HI(net77));
 sg13g2_tiehi _1088__59 (.L_HI(net78));
 sg13g2_tiehi _1087__60 (.L_HI(net79));
 sg13g2_tiehi _1086__61 (.L_HI(net80));
 sg13g2_tiehi _1085__62 (.L_HI(net81));
 sg13g2_tiehi _1084__63 (.L_HI(net82));
 sg13g2_tiehi _1083__64 (.L_HI(net83));
 sg13g2_tiehi _1082__65 (.L_HI(net84));
 sg13g2_tiehi _1081__66 (.L_HI(net85));
 sg13g2_tiehi _1080__67 (.L_HI(net86));
 sg13g2_tiehi _1079__68 (.L_HI(net87));
 sg13g2_tiehi _1076__69 (.L_HI(net88));
 sg13g2_tiehi _1075__70 (.L_HI(net89));
 sg13g2_tiehi _1074__71 (.L_HI(net90));
 sg13g2_tiehi _1134__72 (.L_HI(net91));
 sg13g2_tiehi _1073__73 (.L_HI(net92));
 sg13g2_tiehi _1071__74 (.L_HI(net93));
 sg13g2_tiehi _1069__75 (.L_HI(net94));
 sg13g2_tiehi _1068__76 (.L_HI(net95));
 sg13g2_tiehi _1067__77 (.L_HI(net96));
 sg13g2_tiehi _1066__78 (.L_HI(net97));
 sg13g2_tiehi _1065__79 (.L_HI(net98));
 sg13g2_tiehi _1021__80 (.L_HI(net99));
 sg13g2_tiehi _1064__81 (.L_HI(net100));
 sg13g2_tiehi _1070__82 (.L_HI(net101));
 sg13g2_tiehi _1063__83 (.L_HI(net102));
 sg13g2_tiehi _1062__84 (.L_HI(net103));
 sg13g2_tiehi _1061__85 (.L_HI(net104));
 sg13g2_tiehi _1060__86 (.L_HI(net105));
 sg13g2_tiehi _1072__87 (.L_HI(net106));
 sg13g2_tiehi _1077__88 (.L_HI(net107));
 sg13g2_tiehi _1059__89 (.L_HI(net108));
 sg13g2_tiehi _1058__90 (.L_HI(net109));
 sg13g2_tiehi _1057__91 (.L_HI(net110));
 sg13g2_tiehi _1056__92 (.L_HI(net111));
 sg13g2_tiehi _1055__93 (.L_HI(net112));
 sg13g2_tiehi _1054__94 (.L_HI(net113));
 sg13g2_tiehi _1053__95 (.L_HI(net114));
 sg13g2_tiehi _1052__96 (.L_HI(net115));
 sg13g2_tiehi _1051__97 (.L_HI(net116));
 sg13g2_tiehi _1050__98 (.L_HI(net117));
 sg13g2_tiehi _1049__99 (.L_HI(net118));
 sg13g2_tiehi _1048__100 (.L_HI(net119));
 sg13g2_tiehi _1114__101 (.L_HI(net120));
 sg13g2_tiehi _1047__102 (.L_HI(net121));
 sg13g2_tiehi _1046__103 (.L_HI(net122));
 sg13g2_tiehi _1045__104 (.L_HI(net123));
 sg13g2_tiehi _1044__105 (.L_HI(net124));
 sg13g2_tiehi _1043__106 (.L_HI(net125));
 sg13g2_tiehi _1042__107 (.L_HI(net126));
 sg13g2_tiehi _1041__108 (.L_HI(net127));
 sg13g2_tiehi _1040__109 (.L_HI(net128));
 sg13g2_tiehi _1039__110 (.L_HI(net129));
 sg13g2_tiehi _1038__111 (.L_HI(net130));
 sg13g2_tiehi _1037__112 (.L_HI(net131));
 sg13g2_tiehi _1036__113 (.L_HI(net132));
 sg13g2_tiehi _1035__114 (.L_HI(net133));
 sg13g2_tiehi _1034__115 (.L_HI(net134));
 sg13g2_tiehi _1033__116 (.L_HI(net135));
 sg13g2_tiehi _1032__117 (.L_HI(net136));
 sg13g2_tiehi _1031__118 (.L_HI(net137));
 sg13g2_tiehi _1030__119 (.L_HI(net138));
 sg13g2_tiehi _1029__120 (.L_HI(net139));
 sg13g2_tiehi _1028__121 (.L_HI(net140));
 sg13g2_tiehi _1027__122 (.L_HI(net141));
 sg13g2_tiehi _1026__123 (.L_HI(net142));
 sg13g2_tiehi _1025__124 (.L_HI(net143));
 sg13g2_tiehi _1024__125 (.L_HI(net144));
 sg13g2_tiehi _1078__126 (.L_HI(net145));
 sg13g2_tiehi _1116__127 (.L_HI(net146));
 sg13g2_tiehi _1117__128 (.L_HI(net147));
 sg13g2_tiehi _1118__129 (.L_HI(net148));
 sg13g2_tiehi _1119__130 (.L_HI(net149));
 sg13g2_tiehi _1120__131 (.L_HI(net150));
 sg13g2_tiehi _1121__132 (.L_HI(net151));
 sg13g2_tiehi _1122__133 (.L_HI(net152));
 sg13g2_tiehi _1123__134 (.L_HI(net153));
 sg13g2_tiehi _1124__135 (.L_HI(net154));
 sg13g2_tiehi _1125__136 (.L_HI(net155));
 sg13g2_tiehi _1126__137 (.L_HI(net156));
 sg13g2_tiehi _1127__138 (.L_HI(net157));
 sg13g2_tiehi _1128__139 (.L_HI(net158));
 sg13g2_tiehi _1129__140 (.L_HI(net159));
 sg13g2_tiehi _1130__141 (.L_HI(net160));
 sg13g2_tiehi _1131__142 (.L_HI(net161));
 sg13g2_tiehi _1132__143 (.L_HI(net162));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_tommythorn_workshop_15 (.L_LO(net15));
 sg13g2_tielo tt_um_tommythorn_workshop_16 (.L_LO(net16));
 sg13g2_tielo tt_um_tommythorn_workshop_17 (.L_LO(net17));
 sg13g2_tielo tt_um_tommythorn_workshop_18 (.L_LO(net18));
 sg13g2_tielo tt_um_tommythorn_workshop_19 (.L_LO(net19));
 sg13g2_tielo tt_um_tommythorn_workshop_20 (.L_LO(net20));
 sg13g2_tielo tt_um_tommythorn_workshop_21 (.L_LO(net21));
 sg13g2_tielo tt_um_tommythorn_workshop_22 (.L_LO(net22));
 sg13g2_tielo tt_um_tommythorn_workshop_23 (.L_LO(net23));
 sg13g2_tielo tt_um_tommythorn_workshop_24 (.L_LO(net24));
 sg13g2_tielo tt_um_tommythorn_workshop_25 (.L_LO(net25));
 sg13g2_tielo tt_um_tommythorn_workshop_26 (.L_LO(net26));
 sg13g2_tielo tt_um_tommythorn_workshop_27 (.L_LO(net27));
 sg13g2_tielo tt_um_tommythorn_workshop_28 (.L_LO(net28));
 sg13g2_tielo tt_um_tommythorn_workshop_29 (.L_LO(net29));
 sg13g2_tiehi _1023__30 (.L_HI(net30));
 sg13g2_buf_1 _1265_ (.A(\rs232out_inst.serial_out ),
    .X(uo_out[0]));
 sg13g2_buf_1 _1266_ (.A(\pdm_inst.O ),
    .X(uo_out[1]));
 sg13g2_buf_2 fanout56 (.A(_0292_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0151_),
    .X(net57));
 sg13g2_buf_4 fanout58 (.X(net58),
    .A(_0398_));
 sg13g2_buf_2 fanout59 (.A(net62),
    .X(net59));
 sg13g2_buf_1 fanout60 (.A(net62),
    .X(net60));
 sg13g2_buf_4 fanout61 (.X(net61),
    .A(net62));
 sg13g2_buf_1 fanout62 (.A(_0288_),
    .X(net62));
 sg13g2_buf_4 fanout63 (.X(net63),
    .A(net64));
 sg13g2_buf_2 fanout64 (.A(net67),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(net66),
    .X(net65));
 sg13g2_buf_4 fanout66 (.X(net66),
    .A(net67));
 sg13g2_buf_2 fanout67 (.A(_0260_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(\rs232out_inst.ttyclk[16] ),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(net71),
    .X(net69));
 sg13g2_buf_1 fanout70 (.A(net71),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(\rs232in_inst.ttyclk[16] ),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(net74),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(\rs232out_inst.count[4] ),
    .X(net74));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[0]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[3]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[4]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_tielo tt_um_tommythorn_workshop_14 (.L_LO(net14));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\rs232in_inst.rxd ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0030_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0119_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0031_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0049_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0005_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0083_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold8 (.A(\rs232in_inst.count[1] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0118_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold10 (.A(\rs232out_inst.shift_out[4] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0078_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold12 (.A(\rs232in_inst.count[4] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0405_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold14 (.A(\rs232out_inst.serial_out ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0345_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold16 (.A(\rs232out_inst.shift_out[2] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0076_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold18 (.A(\rs232out_inst.shift_out[3] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0077_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold20 (.A(\pdm_inst.sigma[0] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0012_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold22 (.A(\rs232out_inst.transmit_data[6] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0055_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold24 (.A(\rs232out_inst.shift_out[6] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0080_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold26 (.A(\rs232out_inst.shift_out[1] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0075_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold28 (.A(\rs232out_inst.shift_out[5] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0079_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold30 (.A(\rs232out_inst.shift_out[7] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0081_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold32 (.A(\rs232out_inst.transmit_data[1] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0050_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold34 (.A(\rs232out_inst.transmit_data[4] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0053_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0008_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0094_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold38 (.A(\rs232in_inst.shift_in[1] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0110_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0006_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0085_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0004_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0299_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0063_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold45 (.A(\rs232out_inst.count[3] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0351_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0086_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold48 (.A(\rs232out_inst.count[1] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0084_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold50 (.A(\rs232out_inst.transmit_data[2] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0051_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold52 (.A(\rs232in_inst.shift_in[2] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold53 (.A(\rs232in_inst.shift_in[5] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0114_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0003_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0292_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0060_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold58 (.A(\rs232in_inst.received_data[7] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0117_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold60 (.A(\rs232out_inst.ttyclk[2] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0296_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold62 (.A(\rs232out_inst.ttyclk[6] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0065_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold64 (.A(\rs232out_inst.transmit_data[5] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0054_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold66 (.A(\pdm_inst.sigma[17] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0258_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0020_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold69 (.A(\rs232in_inst.shift_in[4] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0113_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold71 (.A(\rs232out_inst.ttyclk[5] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold72 (.A(\rs232in_inst.ttyclk[12] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0391_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0106_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold75 (.A(\rs232out_inst.ttyclk[0] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0059_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold77 (.A(\rs232in_inst.shift_in[3] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0112_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0002_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0353_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0009_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0380_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0101_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold84 (.A(\rs232in_inst.ttyclk[15] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0396_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold86 (.A(\rs232out_inst.shift_out[8] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0058_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold88 (.A(\rs232in_inst.ttyclk[3] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold89 (.A(\rs232in_inst.shift_in[6] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0092_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold91 (.A(\rs232in_inst.count[0] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold92 (.A(\rs232in_inst.received_data[1] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold93 (.A(\rs232out_inst.ttyclk[15] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0322_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0074_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold96 (.A(\rs232out_inst.transmit_data[3] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0052_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold98 (.A(\rs232out_inst.ttyclk[3] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0298_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0062_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold101 (.A(\rs232out_inst.ttyclk[10] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0313_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0069_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold104 (.A(\rs232in_inst.received_data[5] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold105 (.A(\rs232in_inst.count[3] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0122_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold107 (.A(\rs232in_inst.ttyclk[2] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0096_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold109 (.A(\rs232in_inst.shift_in[7] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0116_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold111 (.A(\rs232in_inst.rxd2 ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold112 (.A(\rs232in_inst.ttyclk[6] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0377_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold114 (.A(\pdm_inst.level[0] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0040_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold116 (.A(\rs232out_inst.ttyclk[14] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0321_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold118 (.A(\pdm_inst.level[4] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0036_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold120 (.A(\rs232in_inst.received_data[3] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0035_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold122 (.A(\rs232in_inst.ttyclk[10] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0388_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold124 (.A(\pdm_inst.level[13] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0045_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold126 (.A(\pdm_inst.level[15] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0263_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0047_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold129 (.A(\rs232in_inst.count[2] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold130 (.A(\rs232out_inst.ttyclk[7] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0066_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold132 (.A(\rs232out_inst.transmit_data[7] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0056_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold134 (.A(\rs232in_inst.ttyclk[4] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0098_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold136 (.A(\pdm_inst.level[11] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0043_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold138 (.A(\pdm_inst.level[12] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold139 (.A(\rs232in_inst.received_data[2] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0034_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold141 (.A(\rs232in_inst.ttyclk[1] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0095_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold143 (.A(\rs232in_inst.ttyclk[9] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0385_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0103_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold146 (.A(\pdm_inst.level[6] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0046_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold148 (.A(\pdm_inst.level[5] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0007_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0269_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold151 (.A(\rs232in_inst.received_data[6] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold152 (.A(\rs232in_inst.ttyclk[8] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0382_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0102_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold155 (.A(\rs232in_inst.ttyclk[11] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold156 (.A(\rs232in_inst.received_data[0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold157 (.A(\rs232out_inst.ttyclk[13] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0319_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold159 (.A(\rs232out_inst.ttyclk[8] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold160 (.A(\pdm_inst.level[7] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold161 (.A(\rs232out_inst.ttyclk[9] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold162 (.A(\pdm_inst.sigma[1] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0182_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold164 (.A(\pdm_inst.level[9] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0041_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold166 (.A(\pdm_inst.level[2] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0042_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold168 (.A(\rs232in_inst.ttyclk[13] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold169 (.A(\pdm_inst.level[1] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold170 (.A(\rs232out_inst.we ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0001_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold172 (.A(\pdm_inst.sigma[4] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0025_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold174 (.A(\rs232out_inst.ttyclk[11] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold175 (.A(\pdm_inst.sigma[16] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0019_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold177 (.A(\rs232in_inst.ttyclk[14] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold178 (.A(\rs232in_inst.ttyclk[5] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0372_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0099_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold181 (.A(\pdm_inst.sigma[2] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0023_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold183 (.A(\pdm_inst.sigma[8] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0218_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0029_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold186 (.A(\pdm_inst.sigma[15] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0018_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold188 (.A(\pdm_inst.sigma[14] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0249_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0017_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold191 (.A(\rs232out_inst.ttyclk[12] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold192 (.A(\pdm_inst.sigma[12] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold193 (.A(\pdm_inst.sigma[10] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0221_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold195 (.A(\pdm_inst.sigma[1] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold196 (.A(\pdm_inst.level[8] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold197 (.A(\rs232in_inst.ttyclk[6] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0157_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold199 (.A(\pdm_inst.sigma[11] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0014_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold201 (.A(\pdm_inst.sigma[13] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold202 (.A(\pdm_inst.sigma[7] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0027_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold204 (.A(\pdm_inst.sigma[6] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold205 (.A(\rs232in_inst.ttyclk[2] ),
    .X(net367));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_4 FILLER_8_294 ();
 sg13g2_fill_1 FILLER_8_298 ();
 sg13g2_decap_8 FILLER_8_303 ();
 sg13g2_decap_8 FILLER_8_310 ();
 sg13g2_decap_8 FILLER_8_317 ();
 sg13g2_decap_8 FILLER_8_345 ();
 sg13g2_decap_8 FILLER_8_352 ();
 sg13g2_decap_8 FILLER_8_359 ();
 sg13g2_decap_8 FILLER_8_366 ();
 sg13g2_decap_8 FILLER_8_373 ();
 sg13g2_decap_8 FILLER_8_380 ();
 sg13g2_decap_8 FILLER_8_387 ();
 sg13g2_decap_8 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_4 FILLER_9_217 ();
 sg13g2_fill_2 FILLER_9_221 ();
 sg13g2_decap_4 FILLER_9_231 ();
 sg13g2_fill_2 FILLER_9_235 ();
 sg13g2_decap_8 FILLER_9_242 ();
 sg13g2_decap_8 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_260 ();
 sg13g2_decap_4 FILLER_9_267 ();
 sg13g2_fill_2 FILLER_9_271 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_fill_2 FILLER_10_189 ();
 sg13g2_fill_1 FILLER_10_191 ();
 sg13g2_decap_4 FILLER_10_204 ();
 sg13g2_fill_2 FILLER_10_208 ();
 sg13g2_fill_2 FILLER_10_257 ();
 sg13g2_fill_1 FILLER_10_269 ();
 sg13g2_decap_8 FILLER_10_274 ();
 sg13g2_fill_2 FILLER_10_281 ();
 sg13g2_fill_1 FILLER_10_304 ();
 sg13g2_fill_2 FILLER_10_314 ();
 sg13g2_fill_2 FILLER_10_333 ();
 sg13g2_fill_1 FILLER_10_335 ();
 sg13g2_fill_1 FILLER_10_341 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_4 FILLER_10_403 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_fill_1 FILLER_11_221 ();
 sg13g2_fill_2 FILLER_11_257 ();
 sg13g2_fill_1 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_286 ();
 sg13g2_fill_1 FILLER_11_293 ();
 sg13g2_fill_2 FILLER_11_309 ();
 sg13g2_fill_2 FILLER_11_320 ();
 sg13g2_fill_2 FILLER_11_327 ();
 sg13g2_fill_1 FILLER_11_336 ();
 sg13g2_fill_2 FILLER_11_358 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_fill_2 FILLER_12_161 ();
 sg13g2_fill_1 FILLER_12_163 ();
 sg13g2_fill_2 FILLER_12_195 ();
 sg13g2_fill_1 FILLER_12_197 ();
 sg13g2_fill_2 FILLER_12_265 ();
 sg13g2_fill_1 FILLER_12_267 ();
 sg13g2_decap_4 FILLER_12_294 ();
 sg13g2_fill_1 FILLER_12_298 ();
 sg13g2_fill_2 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_fill_2 FILLER_12_357 ();
 sg13g2_fill_2 FILLER_12_367 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_4 FILLER_13_147 ();
 sg13g2_fill_2 FILLER_13_151 ();
 sg13g2_fill_2 FILLER_13_179 ();
 sg13g2_fill_1 FILLER_13_181 ();
 sg13g2_fill_2 FILLER_13_230 ();
 sg13g2_fill_2 FILLER_13_257 ();
 sg13g2_fill_1 FILLER_13_291 ();
 sg13g2_fill_2 FILLER_13_359 ();
 sg13g2_fill_1 FILLER_13_361 ();
 sg13g2_decap_4 FILLER_13_389 ();
 sg13g2_fill_2 FILLER_13_393 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_4 FILLER_14_154 ();
 sg13g2_fill_1 FILLER_14_158 ();
 sg13g2_fill_1 FILLER_14_186 ();
 sg13g2_fill_2 FILLER_14_217 ();
 sg13g2_fill_1 FILLER_14_250 ();
 sg13g2_fill_2 FILLER_14_259 ();
 sg13g2_fill_1 FILLER_14_261 ();
 sg13g2_decap_4 FILLER_14_292 ();
 sg13g2_fill_2 FILLER_14_330 ();
 sg13g2_fill_1 FILLER_14_332 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_4 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_4 FILLER_15_154 ();
 sg13g2_fill_1 FILLER_15_158 ();
 sg13g2_fill_1 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_222 ();
 sg13g2_decap_4 FILLER_15_232 ();
 sg13g2_fill_2 FILLER_15_315 ();
 sg13g2_fill_1 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_fill_2 FILLER_16_140 ();
 sg13g2_fill_2 FILLER_16_156 ();
 sg13g2_decap_4 FILLER_16_162 ();
 sg13g2_fill_2 FILLER_16_166 ();
 sg13g2_fill_2 FILLER_16_186 ();
 sg13g2_fill_1 FILLER_16_188 ();
 sg13g2_fill_1 FILLER_16_212 ();
 sg13g2_fill_2 FILLER_16_254 ();
 sg13g2_fill_1 FILLER_16_269 ();
 sg13g2_fill_1 FILLER_16_304 ();
 sg13g2_fill_1 FILLER_16_329 ();
 sg13g2_fill_2 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_fill_2 FILLER_17_133 ();
 sg13g2_fill_1 FILLER_17_135 ();
 sg13g2_fill_2 FILLER_17_145 ();
 sg13g2_fill_2 FILLER_17_238 ();
 sg13g2_fill_2 FILLER_17_296 ();
 sg13g2_fill_1 FILLER_17_298 ();
 sg13g2_fill_2 FILLER_17_341 ();
 sg13g2_fill_1 FILLER_17_343 ();
 sg13g2_fill_2 FILLER_17_349 ();
 sg13g2_fill_1 FILLER_17_351 ();
 sg13g2_fill_2 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_fill_2 FILLER_17_394 ();
 sg13g2_fill_1 FILLER_17_396 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_fill_1 FILLER_18_119 ();
 sg13g2_decap_4 FILLER_18_156 ();
 sg13g2_fill_1 FILLER_18_160 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_1 FILLER_18_230 ();
 sg13g2_fill_2 FILLER_18_286 ();
 sg13g2_fill_2 FILLER_18_298 ();
 sg13g2_fill_1 FILLER_18_352 ();
 sg13g2_decap_4 FILLER_18_382 ();
 sg13g2_fill_2 FILLER_18_386 ();
 sg13g2_fill_2 FILLER_18_392 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_4 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_134 ();
 sg13g2_fill_2 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_167 ();
 sg13g2_fill_2 FILLER_19_176 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_1 FILLER_19_216 ();
 sg13g2_fill_1 FILLER_19_232 ();
 sg13g2_fill_1 FILLER_19_246 ();
 sg13g2_fill_1 FILLER_19_261 ();
 sg13g2_fill_2 FILLER_19_312 ();
 sg13g2_fill_1 FILLER_19_392 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_fill_2 FILLER_20_119 ();
 sg13g2_fill_1 FILLER_20_121 ();
 sg13g2_decap_4 FILLER_20_148 ();
 sg13g2_fill_1 FILLER_20_152 ();
 sg13g2_fill_2 FILLER_20_182 ();
 sg13g2_fill_1 FILLER_20_184 ();
 sg13g2_fill_1 FILLER_20_215 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_fill_2 FILLER_20_268 ();
 sg13g2_fill_1 FILLER_20_270 ();
 sg13g2_fill_2 FILLER_20_289 ();
 sg13g2_fill_1 FILLER_20_308 ();
 sg13g2_fill_1 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_150 ();
 sg13g2_decap_4 FILLER_21_157 ();
 sg13g2_fill_1 FILLER_21_161 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_fill_1 FILLER_21_186 ();
 sg13g2_decap_4 FILLER_21_238 ();
 sg13g2_fill_2 FILLER_21_242 ();
 sg13g2_fill_2 FILLER_21_252 ();
 sg13g2_fill_2 FILLER_21_273 ();
 sg13g2_fill_1 FILLER_21_275 ();
 sg13g2_fill_2 FILLER_21_302 ();
 sg13g2_fill_2 FILLER_21_330 ();
 sg13g2_fill_1 FILLER_21_332 ();
 sg13g2_fill_2 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_fill_2 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_135 ();
 sg13g2_fill_1 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_152 ();
 sg13g2_fill_1 FILLER_22_186 ();
 sg13g2_fill_2 FILLER_22_196 ();
 sg13g2_fill_1 FILLER_22_198 ();
 sg13g2_fill_2 FILLER_22_216 ();
 sg13g2_fill_2 FILLER_22_298 ();
 sg13g2_fill_2 FILLER_22_353 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_4 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_110 ();
 sg13g2_decap_8 FILLER_23_117 ();
 sg13g2_decap_8 FILLER_23_124 ();
 sg13g2_fill_1 FILLER_23_157 ();
 sg13g2_decap_4 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_249 ();
 sg13g2_fill_2 FILLER_23_300 ();
 sg13g2_fill_1 FILLER_23_302 ();
 sg13g2_fill_2 FILLER_23_320 ();
 sg13g2_fill_1 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_4 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_88 ();
 sg13g2_fill_2 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_129 ();
 sg13g2_decap_4 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_172 ();
 sg13g2_fill_2 FILLER_24_187 ();
 sg13g2_decap_4 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_fill_2 FILLER_24_276 ();
 sg13g2_fill_1 FILLER_24_292 ();
 sg13g2_fill_2 FILLER_24_320 ();
 sg13g2_fill_2 FILLER_24_333 ();
 sg13g2_fill_1 FILLER_24_390 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_4 FILLER_25_77 ();
 sg13g2_fill_1 FILLER_25_81 ();
 sg13g2_fill_1 FILLER_25_108 ();
 sg13g2_fill_1 FILLER_25_166 ();
 sg13g2_fill_1 FILLER_25_212 ();
 sg13g2_fill_2 FILLER_25_222 ();
 sg13g2_fill_2 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_339 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_95 ();
 sg13g2_fill_2 FILLER_26_102 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_fill_2 FILLER_26_197 ();
 sg13g2_fill_2 FILLER_26_208 ();
 sg13g2_fill_1 FILLER_26_210 ();
 sg13g2_decap_4 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_decap_4 FILLER_26_239 ();
 sg13g2_fill_1 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_300 ();
 sg13g2_fill_2 FILLER_26_311 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_fill_2 FILLER_26_354 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_fill_2 FILLER_27_77 ();
 sg13g2_fill_1 FILLER_27_79 ();
 sg13g2_fill_1 FILLER_27_156 ();
 sg13g2_fill_2 FILLER_27_282 ();
 sg13g2_fill_1 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_315 ();
 sg13g2_fill_2 FILLER_27_320 ();
 sg13g2_fill_2 FILLER_27_342 ();
 sg13g2_fill_1 FILLER_27_363 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_4 FILLER_28_101 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_2 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_169 ();
 sg13g2_fill_2 FILLER_28_221 ();
 sg13g2_fill_1 FILLER_28_223 ();
 sg13g2_fill_2 FILLER_28_232 ();
 sg13g2_fill_2 FILLER_28_255 ();
 sg13g2_fill_1 FILLER_28_262 ();
 sg13g2_fill_2 FILLER_28_370 ();
 sg13g2_fill_2 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_4 FILLER_29_56 ();
 sg13g2_fill_1 FILLER_29_60 ();
 sg13g2_fill_2 FILLER_29_92 ();
 sg13g2_fill_1 FILLER_29_94 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_fill_1 FILLER_29_168 ();
 sg13g2_fill_2 FILLER_29_217 ();
 sg13g2_fill_2 FILLER_29_261 ();
 sg13g2_fill_2 FILLER_29_267 ();
 sg13g2_fill_1 FILLER_29_269 ();
 sg13g2_fill_1 FILLER_29_301 ();
 sg13g2_fill_1 FILLER_29_325 ();
 sg13g2_fill_1 FILLER_29_392 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_4 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_110 ();
 sg13g2_fill_1 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_fill_2 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_90 ();
 sg13g2_fill_1 FILLER_31_92 ();
 sg13g2_fill_1 FILLER_31_131 ();
 sg13g2_fill_1 FILLER_31_150 ();
 sg13g2_fill_1 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_218 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_326 ();
 sg13g2_fill_1 FILLER_31_339 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_fill_2 FILLER_32_63 ();
 sg13g2_fill_2 FILLER_32_122 ();
 sg13g2_fill_2 FILLER_32_153 ();
 sg13g2_fill_2 FILLER_32_185 ();
 sg13g2_fill_1 FILLER_32_250 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_fill_1 FILLER_32_279 ();
 sg13g2_fill_2 FILLER_32_289 ();
 sg13g2_fill_1 FILLER_32_326 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_4 FILLER_33_63 ();
 sg13g2_fill_2 FILLER_33_67 ();
 sg13g2_fill_1 FILLER_33_95 ();
 sg13g2_fill_1 FILLER_33_135 ();
 sg13g2_fill_1 FILLER_33_190 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_fill_2 FILLER_33_339 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_4 FILLER_34_77 ();
 sg13g2_fill_2 FILLER_34_81 ();
 sg13g2_fill_2 FILLER_34_114 ();
 sg13g2_fill_1 FILLER_34_116 ();
 sg13g2_fill_2 FILLER_34_247 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_fill_2 FILLER_34_306 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_104 ();
 sg13g2_fill_1 FILLER_35_106 ();
 sg13g2_fill_1 FILLER_35_124 ();
 sg13g2_fill_1 FILLER_35_138 ();
 sg13g2_fill_2 FILLER_35_166 ();
 sg13g2_fill_2 FILLER_35_205 ();
 sg13g2_fill_1 FILLER_35_224 ();
 sg13g2_fill_2 FILLER_35_275 ();
 sg13g2_fill_1 FILLER_35_304 ();
 sg13g2_fill_1 FILLER_35_340 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_fill_2 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_108 ();
 sg13g2_fill_1 FILLER_36_176 ();
 sg13g2_fill_2 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_203 ();
 sg13g2_fill_2 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_273 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_fill_2 FILLER_36_350 ();
 sg13g2_fill_2 FILLER_36_378 ();
 sg13g2_fill_1 FILLER_36_380 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_fill_2 FILLER_37_98 ();
 sg13g2_fill_1 FILLER_37_100 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_fill_2 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_223 ();
 sg13g2_fill_1 FILLER_37_225 ();
 sg13g2_fill_2 FILLER_37_273 ();
 sg13g2_fill_2 FILLER_37_301 ();
 sg13g2_fill_1 FILLER_37_303 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_92 ();
 sg13g2_fill_1 FILLER_38_94 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_fill_1 FILLER_38_168 ();
 sg13g2_fill_2 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_245 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_358 ();
 sg13g2_fill_1 FILLER_38_373 ();
 sg13g2_fill_2 FILLER_38_392 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net19;
 assign uio_oe[6] = net20;
 assign uio_oe[7] = net21;
 assign uio_out[0] = net22;
 assign uio_out[1] = net23;
 assign uio_out[2] = net24;
 assign uio_out[3] = net25;
 assign uio_out[4] = net26;
 assign uio_out[5] = net27;
 assign uio_out[6] = net28;
 assign uio_out[7] = net29;
endmodule

module tt_um_lif_network_MR (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire \lif_net.input_current_output[0] ;
 wire \lif_net.input_current_output[1] ;
 wire \lif_net.input_current_output[2] ;
 wire \lif_net.input_current_output[3] ;
 wire \lif_net.neuron1.spike ;
 wire \lif_net.neuron1.state[1] ;
 wire \lif_net.neuron1.state[2] ;
 wire \lif_net.neuron1.state[3] ;
 wire \lif_net.neuron2.spike ;
 wire \lif_net.neuron2.state[1] ;
 wire \lif_net.neuron2.state[2] ;
 wire \lif_net.neuron2.state[3] ;
 wire \lif_net.neuron3.spike ;
 wire \lif_net.neuron3.state[1] ;
 wire \lif_net.neuron3.state[2] ;
 wire \lif_net.neuron3.state[3] ;
 wire \lif_net.output_neuron.spike ;
 wire \lif_net.output_neuron.state[1] ;
 wire \lif_net.output_neuron.state[2] ;
 wire \lif_net.output_neuron.state[3] ;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net43;
 wire net44;
 wire net45;
 wire clknet_0_clk;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;

 sg13g2_inv_1 _100_ (.Y(_038_),
    .A(net54));
 sg13g2_inv_1 _101_ (.Y(_039_),
    .A(net1));
 sg13g2_nand2b_1 _102_ (.Y(_040_),
    .B(net1),
    .A_N(net56));
 sg13g2_nand2_1 _103_ (.Y(_041_),
    .A(\lif_net.output_neuron.state[1] ),
    .B(\lif_net.input_current_output[0] ));
 sg13g2_nand2_1 _104_ (.Y(_042_),
    .A(\lif_net.output_neuron.state[2] ),
    .B(\lif_net.input_current_output[1] ));
 sg13g2_xnor2_1 _105_ (.Y(_043_),
    .A(\lif_net.output_neuron.state[2] ),
    .B(\lif_net.input_current_output[1] ));
 sg13g2_xnor2_1 _106_ (.Y(_044_),
    .A(_041_),
    .B(_043_));
 sg13g2_nor2_1 _107_ (.A(_040_),
    .B(_044_),
    .Y(_000_));
 sg13g2_o21ai_1 _108_ (.B1(_042_),
    .Y(_045_),
    .A1(_041_),
    .A2(_043_));
 sg13g2_xnor2_1 _109_ (.Y(_046_),
    .A(\lif_net.output_neuron.state[3] ),
    .B(net49));
 sg13g2_inv_1 _110_ (.Y(_047_),
    .A(_046_));
 sg13g2_and2_1 _111_ (.A(_045_),
    .B(_047_),
    .X(_048_));
 sg13g2_nor2_1 _112_ (.A(net49),
    .B(_045_),
    .Y(_049_));
 sg13g2_nor3_1 _113_ (.A(_040_),
    .B(_048_),
    .C(net50),
    .Y(_001_));
 sg13g2_a21oi_1 _114_ (.A1(_045_),
    .A2(_047_),
    .Y(_050_),
    .B1(net46));
 sg13g2_and3_1 _115_ (.X(_051_),
    .A(net46),
    .B(_045_),
    .C(_047_));
 sg13g2_nor3_1 _116_ (.A(_040_),
    .B(net47),
    .C(_051_),
    .Y(_002_));
 sg13g2_nand2_1 _117_ (.Y(_052_),
    .A(_038_),
    .B(net1));
 sg13g2_nand2_1 _118_ (.Y(_053_),
    .A(net58),
    .B(net2));
 sg13g2_nand2_1 _119_ (.Y(_054_),
    .A(net66),
    .B(net3));
 sg13g2_xnor2_1 _120_ (.Y(_055_),
    .A(\lif_net.neuron3.state[2] ),
    .B(net3));
 sg13g2_xnor2_1 _121_ (.Y(_056_),
    .A(_053_),
    .B(_055_));
 sg13g2_nor2_1 _122_ (.A(_052_),
    .B(net59),
    .Y(_003_));
 sg13g2_o21ai_1 _123_ (.B1(_054_),
    .Y(_057_),
    .A1(_053_),
    .A2(_055_));
 sg13g2_xnor2_1 _124_ (.Y(_058_),
    .A(\lif_net.neuron3.state[3] ),
    .B(net4));
 sg13g2_inv_1 _125_ (.Y(_059_),
    .A(_058_));
 sg13g2_and2_1 _126_ (.A(_057_),
    .B(_059_),
    .X(_060_));
 sg13g2_nor2_1 _127_ (.A(net4),
    .B(_057_),
    .Y(_061_));
 sg13g2_nor3_1 _128_ (.A(_052_),
    .B(_060_),
    .C(_061_),
    .Y(_004_));
 sg13g2_a21oi_1 _129_ (.A1(_057_),
    .A2(_059_),
    .Y(_062_),
    .B1(net5));
 sg13g2_and3_1 _130_ (.X(_063_),
    .A(net5),
    .B(_057_),
    .C(_059_));
 sg13g2_nor3_1 _131_ (.A(_052_),
    .B(net67),
    .C(_063_),
    .Y(_005_));
 sg13g2_nand2b_1 _132_ (.Y(_064_),
    .B(net1),
    .A_N(net55));
 sg13g2_inv_1 _133_ (.Y(_065_),
    .A(_064_));
 sg13g2_nand2_1 _134_ (.Y(_066_),
    .A(net62),
    .B(net6));
 sg13g2_nand2_1 _135_ (.Y(_067_),
    .A(net64),
    .B(net7));
 sg13g2_xnor2_1 _136_ (.Y(_016_),
    .A(\lif_net.neuron2.state[2] ),
    .B(net7));
 sg13g2_xnor2_1 _137_ (.Y(_017_),
    .A(_066_),
    .B(_016_));
 sg13g2_nor2_1 _138_ (.A(_064_),
    .B(net63),
    .Y(_006_));
 sg13g2_o21ai_1 _139_ (.B1(_067_),
    .Y(_018_),
    .A1(_066_),
    .A2(_016_));
 sg13g2_xor2_1 _140_ (.B(net8),
    .A(net55),
    .X(_019_));
 sg13g2_o21ai_1 _141_ (.B1(_065_),
    .Y(_020_),
    .A1(net8),
    .A2(_018_));
 sg13g2_a21oi_1 _142_ (.A1(_018_),
    .A2(_019_),
    .Y(_007_),
    .B1(_020_));
 sg13g2_a21oi_1 _143_ (.A1(_018_),
    .A2(_019_),
    .Y(_021_),
    .B1(net9));
 sg13g2_and3_1 _144_ (.X(_022_),
    .A(net9),
    .B(_018_),
    .C(_019_));
 sg13g2_nor3_1 _145_ (.A(_064_),
    .B(_021_),
    .C(_022_),
    .Y(_008_));
 sg13g2_nand2b_2 _146_ (.Y(_023_),
    .B(net1),
    .A_N(net52));
 sg13g2_nand2_1 _147_ (.Y(_024_),
    .A(net60),
    .B(net10));
 sg13g2_nand2_1 _148_ (.Y(_025_),
    .A(net65),
    .B(net11));
 sg13g2_xnor2_1 _149_ (.Y(_026_),
    .A(\lif_net.neuron1.state[2] ),
    .B(net11));
 sg13g2_xnor2_1 _150_ (.Y(_027_),
    .A(_024_),
    .B(_026_));
 sg13g2_nor2_1 _151_ (.A(_023_),
    .B(net61),
    .Y(_009_));
 sg13g2_o21ai_1 _152_ (.B1(_025_),
    .Y(_028_),
    .A1(_024_),
    .A2(_026_));
 sg13g2_xnor2_1 _153_ (.Y(_029_),
    .A(net52),
    .B(net12));
 sg13g2_inv_1 _154_ (.Y(_030_),
    .A(_029_));
 sg13g2_and2_1 _155_ (.A(_028_),
    .B(_030_),
    .X(_031_));
 sg13g2_nor2_1 _156_ (.A(net12),
    .B(_028_),
    .Y(_032_));
 sg13g2_nor3_1 _157_ (.A(_023_),
    .B(_031_),
    .C(_032_),
    .Y(_010_));
 sg13g2_a21oi_1 _158_ (.A1(_028_),
    .A2(_030_),
    .Y(_033_),
    .B1(net13));
 sg13g2_and3_1 _159_ (.X(_034_),
    .A(net13),
    .B(_028_),
    .C(_030_));
 sg13g2_nor3_1 _160_ (.A(_023_),
    .B(_033_),
    .C(_034_),
    .Y(_011_));
 sg13g2_nor2_1 _161_ (.A(_038_),
    .B(_023_),
    .Y(_013_));
 sg13g2_nor2b_1 _162_ (.A(net54),
    .B_N(net52),
    .Y(_035_));
 sg13g2_a21o_1 _163_ (.A2(_035_),
    .A1(net1),
    .B1(_013_),
    .X(_012_));
 sg13g2_xnor2_1 _164_ (.Y(_036_),
    .A(net55),
    .B(_035_));
 sg13g2_nor2_1 _165_ (.A(_039_),
    .B(_036_),
    .Y(_014_));
 sg13g2_o21ai_1 _166_ (.B1(net52),
    .Y(_037_),
    .A1(\lif_net.neuron2.state[3] ),
    .A2(\lif_net.neuron3.state[3] ));
 sg13g2_nor2_1 _167_ (.A(_039_),
    .B(net53),
    .Y(_015_));
 sg13g2_buf_1 _168_ (.A(\lif_net.neuron2.state[3] ),
    .X(\lif_net.neuron2.spike ));
 sg13g2_buf_1 _169_ (.A(\lif_net.neuron1.state[3] ),
    .X(\lif_net.neuron1.spike ));
 sg13g2_buf_1 _170_ (.A(\lif_net.neuron3.state[3] ),
    .X(\lif_net.neuron3.spike ));
 sg13g2_buf_1 _171_ (.A(\lif_net.output_neuron.state[3] ),
    .X(\lif_net.output_neuron.spike ));
 sg13g2_dfrbp_1 _172_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net36),
    .D(net57),
    .Q_N(_083_),
    .Q(\lif_net.output_neuron.state[1] ));
 sg13g2_dfrbp_1 _173_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net35),
    .D(net51),
    .Q_N(_082_),
    .Q(\lif_net.output_neuron.state[2] ));
 sg13g2_dfrbp_1 _174_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net34),
    .D(net48),
    .Q_N(_081_),
    .Q(\lif_net.output_neuron.state[3] ));
 sg13g2_dfrbp_1 _175_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net33),
    .D(_003_),
    .Q_N(_080_),
    .Q(\lif_net.neuron3.state[1] ));
 sg13g2_dfrbp_1 _176_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net32),
    .D(_004_),
    .Q_N(_079_),
    .Q(\lif_net.neuron3.state[2] ));
 sg13g2_dfrbp_1 _177_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net31),
    .D(_005_),
    .Q_N(_078_),
    .Q(\lif_net.neuron3.state[3] ));
 sg13g2_dfrbp_1 _178_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net30),
    .D(_006_),
    .Q_N(_077_),
    .Q(\lif_net.neuron2.state[1] ));
 sg13g2_dfrbp_1 _179_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net29),
    .D(_007_),
    .Q_N(_076_),
    .Q(\lif_net.neuron2.state[2] ));
 sg13g2_dfrbp_1 _180_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net28),
    .D(_008_),
    .Q_N(_075_),
    .Q(\lif_net.neuron2.state[3] ));
 sg13g2_dfrbp_1 _181_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net27),
    .D(_009_),
    .Q_N(_074_),
    .Q(\lif_net.neuron1.state[1] ));
 sg13g2_dfrbp_1 _182_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net26),
    .D(_010_),
    .Q_N(_073_),
    .Q(\lif_net.neuron1.state[2] ));
 sg13g2_dfrbp_1 _183_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net41),
    .D(_011_),
    .Q_N(_072_),
    .Q(\lif_net.neuron1.state[3] ));
 sg13g2_dfrbp_1 _184_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net40),
    .D(_012_),
    .Q_N(_071_),
    .Q(\lif_net.input_current_output[0] ));
 sg13g2_dfrbp_1 _185_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net39),
    .D(_013_),
    .Q_N(_070_),
    .Q(\lif_net.input_current_output[1] ));
 sg13g2_dfrbp_1 _186_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net38),
    .D(_014_),
    .Q_N(_069_),
    .Q(\lif_net.input_current_output[2] ));
 sg13g2_dfrbp_1 _187_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net37),
    .D(_015_),
    .Q_N(_068_),
    .Q(\lif_net.input_current_output[3] ));
 sg13g2_tiehi _181__27 (.L_HI(net27));
 sg13g2_tiehi _180__28 (.L_HI(net28));
 sg13g2_tiehi _179__29 (.L_HI(net29));
 sg13g2_tiehi _178__30 (.L_HI(net30));
 sg13g2_tiehi _177__31 (.L_HI(net31));
 sg13g2_tiehi _176__32 (.L_HI(net32));
 sg13g2_tiehi _175__33 (.L_HI(net33));
 sg13g2_tiehi _174__34 (.L_HI(net34));
 sg13g2_tiehi _173__35 (.L_HI(net35));
 sg13g2_tiehi _172__36 (.L_HI(net36));
 sg13g2_tiehi _187__37 (.L_HI(net37));
 sg13g2_tiehi _186__38 (.L_HI(net38));
 sg13g2_tiehi _185__39 (.L_HI(net39));
 sg13g2_tiehi _184__40 (.L_HI(net40));
 sg13g2_tiehi _183__41 (.L_HI(net41));
 sg13g2_tiehi tt_um_lif_network_MR_42 (.L_HI(net42));
 sg13g2_tiehi tt_um_lif_network_MR_43 (.L_HI(net43));
 sg13g2_tiehi tt_um_lif_network_MR_44 (.L_HI(net44));
 sg13g2_tiehi tt_um_lif_network_MR_45 (.L_HI(net45));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_lif_network_MR_15 (.L_LO(net15));
 sg13g2_tielo tt_um_lif_network_MR_16 (.L_LO(net16));
 sg13g2_tielo tt_um_lif_network_MR_17 (.L_LO(net17));
 sg13g2_tielo tt_um_lif_network_MR_18 (.L_LO(net18));
 sg13g2_tielo tt_um_lif_network_MR_19 (.L_LO(net19));
 sg13g2_tielo tt_um_lif_network_MR_20 (.L_LO(net20));
 sg13g2_tielo tt_um_lif_network_MR_21 (.L_LO(net21));
 sg13g2_tielo tt_um_lif_network_MR_22 (.L_LO(net22));
 sg13g2_tielo tt_um_lif_network_MR_23 (.L_LO(net23));
 sg13g2_tielo tt_um_lif_network_MR_24 (.L_LO(net24));
 sg13g2_tielo tt_um_lif_network_MR_25 (.L_LO(net25));
 sg13g2_tiehi _182__26 (.L_HI(net26));
 sg13g2_buf_1 _220_ (.A(\lif_net.neuron1.spike ),
    .X(uio_out[4]));
 sg13g2_buf_1 _221_ (.A(\lif_net.neuron2.spike ),
    .X(uio_out[5]));
 sg13g2_buf_2 _222_ (.A(\lif_net.neuron3.spike ),
    .X(uio_out[6]));
 sg13g2_buf_2 _223_ (.A(\lif_net.output_neuron.spike ),
    .X(uio_out[7]));
 sg13g2_buf_1 _224_ (.A(\lif_net.output_neuron.spike ),
    .X(uo_out[0]));
 sg13g2_buf_1 _225_ (.A(\lif_net.neuron1.spike ),
    .X(uo_out[1]));
 sg13g2_buf_1 _226_ (.A(\lif_net.neuron2.spike ),
    .X(uo_out[2]));
 sg13g2_buf_1 _227_ (.A(\lif_net.neuron3.spike ),
    .X(uo_out[3]));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[1]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[2]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[3]),
    .X(net13));
 sg13g2_tielo tt_um_lif_network_MR_14 (.L_LO(net14));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\lif_net.input_current_output[3] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold2 (.A(_050_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold3 (.A(_002_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold4 (.A(\lif_net.input_current_output[2] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold5 (.A(_049_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold6 (.A(_001_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold7 (.A(\lif_net.neuron1.state[3] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold8 (.A(_037_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold9 (.A(\lif_net.neuron3.state[3] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold10 (.A(\lif_net.neuron2.state[3] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold11 (.A(\lif_net.output_neuron.state[3] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold12 (.A(_000_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold13 (.A(\lif_net.neuron3.state[1] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold14 (.A(_056_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold15 (.A(\lif_net.neuron1.state[1] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold16 (.A(_027_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold17 (.A(\lif_net.neuron2.state[1] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold18 (.A(_017_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold19 (.A(\lif_net.neuron2.state[2] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold20 (.A(\lif_net.neuron1.state[2] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold21 (.A(\lif_net.neuron3.state[2] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold22 (.A(_062_),
    .X(net67));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_fill_2 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_4 FILLER_27_280 ();
 sg13g2_fill_1 FILLER_27_284 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_decap_8 FILLER_27_330 ();
 sg13g2_decap_8 FILLER_27_337 ();
 sg13g2_decap_8 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_280 ();
 sg13g2_fill_1 FILLER_28_282 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_fill_2 FILLER_28_294 ();
 sg13g2_fill_2 FILLER_28_300 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_decap_8 FILLER_28_349 ();
 sg13g2_decap_8 FILLER_28_356 ();
 sg13g2_decap_8 FILLER_28_363 ();
 sg13g2_decap_8 FILLER_28_370 ();
 sg13g2_decap_8 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_decap_4 FILLER_29_268 ();
 sg13g2_fill_1 FILLER_29_307 ();
 sg13g2_fill_1 FILLER_29_324 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_4 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_234 ();
 sg13g2_fill_1 FILLER_30_265 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_367 ();
 sg13g2_decap_8 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_fill_1 FILLER_31_224 ();
 sg13g2_decap_4 FILLER_31_248 ();
 sg13g2_fill_2 FILLER_31_252 ();
 sg13g2_decap_4 FILLER_31_296 ();
 sg13g2_decap_8 FILLER_31_352 ();
 sg13g2_decap_8 FILLER_31_359 ();
 sg13g2_decap_8 FILLER_31_366 ();
 sg13g2_decap_8 FILLER_31_373 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_fill_2 FILLER_32_236 ();
 sg13g2_fill_2 FILLER_32_243 ();
 sg13g2_fill_1 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_decap_8 FILLER_32_351 ();
 sg13g2_decap_8 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_4 FILLER_33_217 ();
 sg13g2_fill_1 FILLER_33_221 ();
 sg13g2_fill_2 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_273 ();
 sg13g2_fill_2 FILLER_33_293 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_decap_4 FILLER_33_317 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_4 FILLER_34_217 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_decap_4 FILLER_34_238 ();
 sg13g2_fill_2 FILLER_34_242 ();
 sg13g2_fill_2 FILLER_34_260 ();
 sg13g2_fill_1 FILLER_34_287 ();
 sg13g2_fill_1 FILLER_34_293 ();
 sg13g2_fill_2 FILLER_34_320 ();
 sg13g2_fill_1 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_337 ();
 sg13g2_decap_8 FILLER_34_344 ();
 sg13g2_decap_8 FILLER_34_351 ();
 sg13g2_decap_8 FILLER_34_358 ();
 sg13g2_decap_8 FILLER_34_365 ();
 sg13g2_decap_8 FILLER_34_372 ();
 sg13g2_decap_8 FILLER_34_379 ();
 sg13g2_decap_8 FILLER_34_386 ();
 sg13g2_decap_8 FILLER_34_393 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_4 FILLER_35_217 ();
 sg13g2_fill_2 FILLER_35_221 ();
 sg13g2_fill_1 FILLER_35_231 ();
 sg13g2_fill_2 FILLER_35_237 ();
 sg13g2_fill_2 FILLER_35_265 ();
 sg13g2_fill_2 FILLER_35_279 ();
 sg13g2_decap_8 FILLER_35_310 ();
 sg13g2_fill_1 FILLER_35_317 ();
 sg13g2_decap_8 FILLER_35_331 ();
 sg13g2_decap_8 FILLER_35_338 ();
 sg13g2_decap_8 FILLER_35_345 ();
 sg13g2_decap_8 FILLER_35_352 ();
 sg13g2_decap_8 FILLER_35_359 ();
 sg13g2_decap_8 FILLER_35_366 ();
 sg13g2_decap_8 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_380 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_fill_2 FILLER_36_217 ();
 sg13g2_fill_1 FILLER_36_219 ();
 sg13g2_decap_4 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_fill_1 FILLER_36_284 ();
 sg13g2_decap_8 FILLER_36_333 ();
 sg13g2_decap_8 FILLER_36_340 ();
 sg13g2_decap_8 FILLER_36_347 ();
 sg13g2_decap_8 FILLER_36_354 ();
 sg13g2_decap_8 FILLER_36_361 ();
 sg13g2_decap_8 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_decap_8 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_389 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_fill_2 FILLER_37_224 ();
 sg13g2_fill_1 FILLER_37_226 ();
 sg13g2_fill_2 FILLER_37_253 ();
 sg13g2_fill_1 FILLER_37_277 ();
 sg13g2_decap_8 FILLER_37_324 ();
 sg13g2_decap_8 FILLER_37_331 ();
 sg13g2_decap_8 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_37_345 ();
 sg13g2_decap_8 FILLER_37_352 ();
 sg13g2_decap_8 FILLER_37_359 ();
 sg13g2_decap_8 FILLER_37_366 ();
 sg13g2_decap_8 FILLER_37_373 ();
 sg13g2_decap_8 FILLER_37_380 ();
 sg13g2_decap_8 FILLER_37_387 ();
 sg13g2_decap_8 FILLER_37_394 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_123 ();
 sg13g2_decap_8 FILLER_38_130 ();
 sg13g2_decap_8 FILLER_38_137 ();
 sg13g2_decap_8 FILLER_38_144 ();
 sg13g2_fill_1 FILLER_38_151 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_decap_8 FILLER_38_212 ();
 sg13g2_decap_8 FILLER_38_219 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_decap_4 FILLER_38_233 ();
 sg13g2_fill_1 FILLER_38_237 ();
 sg13g2_decap_4 FILLER_38_242 ();
 sg13g2_fill_1 FILLER_38_246 ();
 sg13g2_fill_2 FILLER_38_259 ();
 sg13g2_fill_1 FILLER_38_275 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_decap_4 FILLER_38_340 ();
 sg13g2_decap_4 FILLER_38_348 ();
 sg13g2_decap_4 FILLER_38_356 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_decap_4 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net42;
 assign uio_oe[5] = net43;
 assign uio_oe[6] = net44;
 assign uio_oe[7] = net45;
 assign uio_out[0] = net18;
 assign uio_out[1] = net19;
 assign uio_out[2] = net20;
 assign uio_out[3] = net21;
 assign uo_out[4] = net22;
 assign uo_out[5] = net23;
 assign uo_out[6] = net24;
 assign uo_out[7] = net25;
endmodule

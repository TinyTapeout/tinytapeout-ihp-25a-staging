module tt_um_wokwi_group_13 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire \proj_10.net11 ;
 wire \proj_10.net12 ;
 wire \proj_10.net13 ;
 wire \proj_10.net14 ;
 wire \proj_10.net15 ;
 wire \proj_10.net16 ;
 wire \proj_10.net17 ;
 wire \proj_10.net18 ;
 wire \proj_10.net24 ;
 wire \proj_10.net25 ;
 wire \proj_10.net26 ;
 wire \proj_10.net27 ;
 wire \proj_10.net28 ;
 wire \proj_10.net29 ;
 wire \proj_10.net30 ;
 wire \proj_10.net31 ;
 wire \proj_10.net32 ;
 wire \proj_10.net33 ;
 wire \proj_10.net34 ;
 wire \proj_10.net35 ;
 wire \proj_10.net36 ;
 wire \proj_10.net37 ;
 wire \proj_10.net38 ;
 wire \proj_10.net39 ;
 wire \proj_10.net40 ;
 wire \proj_10.net41 ;
 wire \proj_10.net42 ;
 wire \proj_10.net43 ;
 wire \proj_10.net44 ;
 wire \proj_10.net45 ;
 wire \proj_10.net46 ;
 wire \proj_10.net47 ;
 wire \proj_10.net48 ;
 wire \proj_10.net49 ;
 wire \proj_10.net50 ;
 wire \proj_10.net51 ;
 wire \proj_10.net52 ;
 wire \proj_10.net53 ;
 wire \proj_10.net54 ;
 wire \proj_10.net55 ;
 wire \proj_10.net56 ;
 wire \proj_10.net57 ;
 wire \proj_10.net59 ;
 wire \proj_10.net60 ;
 wire \proj_10.net61 ;
 wire \proj_10.net62 ;
 wire \proj_10.net63 ;
 wire \proj_10.net64 ;
 wire \proj_10.net66 ;
 wire \proj_10.net69 ;
 wire \proj_10.net71 ;
 wire \proj_10.net72 ;
 wire \proj_10.net73 ;
 wire \proj_10.net74 ;
 wire \proj_10.net75 ;
 wire \proj_10.net76 ;
 wire \proj_10.net77 ;
 wire \proj_10.net78 ;
 wire \proj_10.net79 ;
 wire \proj_10.net80 ;
 wire \proj_10.net82 ;
 wire \proj_10.net83 ;
 wire \proj_10.net85 ;
 wire \proj_10.net87 ;
 wire \proj_10.net89 ;
 wire \proj_10.net92 ;
 wire \proj_10.net93 ;
 wire \proj_10.net94 ;
 wire \proj_10.net95 ;
 wire \proj_10.net96 ;
 wire \proj_11.net10 ;
 wire \proj_11.net11 ;
 wire \proj_11.net12 ;
 wire \proj_11.net9 ;
 wire \proj_12.net10 ;
 wire \proj_12.net11 ;
 wire \proj_12.net17 ;
 wire \proj_12.net19 ;
 wire \proj_12.net20 ;
 wire \proj_12.net7 ;
 wire \proj_12.net8 ;
 wire \proj_12.net9 ;
 wire \proj_13.net10 ;
 wire \proj_13.net11 ;
 wire \proj_13.net12 ;
 wire \proj_13.net13 ;
 wire \proj_13.net14 ;
 wire \proj_13.net15 ;
 wire \proj_13.net16 ;
 wire \proj_13.net22 ;
 wire \proj_13.net23 ;
 wire \proj_13.net24 ;
 wire \proj_13.net25 ;
 wire \proj_13.net26 ;
 wire \proj_13.net27 ;
 wire \proj_13.net28 ;
 wire \proj_13.net29 ;
 wire \proj_13.net30 ;
 wire \proj_13.net31 ;
 wire \proj_13.net32 ;
 wire \proj_13.net33 ;
 wire \proj_13.net34 ;
 wire \proj_13.net35 ;
 wire \proj_13.net36 ;
 wire \proj_13.net37 ;
 wire \proj_13.net38 ;
 wire \proj_13.net39 ;
 wire \proj_13.net40 ;
 wire \proj_13.net41 ;
 wire \proj_13.net42 ;
 wire \proj_13.net43 ;
 wire \proj_13.net44 ;
 wire \proj_14.net3 ;
 wire \proj_15.net10 ;
 wire \proj_15.net11 ;
 wire \proj_15.net12 ;
 wire \proj_15.net9 ;
 wire \proj__0.net10 ;
 wire \proj__0.net11 ;
 wire \proj__1.net10 ;
 wire \proj__1.net11 ;
 wire \proj__1.net12 ;
 wire \proj__1.net13 ;
 wire \proj__2.net12 ;
 wire \proj__2.net13 ;
 wire \proj__2.net14 ;
 wire \proj__2.net6 ;
 wire \proj__3.net14 ;
 wire \proj__3.net15 ;
 wire \proj__3.net16 ;
 wire \proj__3.net17 ;
 wire \proj__3.net18 ;
 wire \proj__3.net19 ;
 wire \proj__3.net2 ;
 wire \proj__3.net20 ;
 wire \proj__3.net21 ;
 wire \proj__3.net22 ;
 wire \proj__3.net23 ;
 wire \proj__3.net24 ;
 wire \proj__3.net25 ;
 wire \proj__3.net26 ;
 wire \proj__3.net27 ;
 wire \proj__3.net28 ;
 wire \proj__3.net29 ;
 wire \proj__3.net3 ;
 wire \proj__3.net4 ;
 wire \proj__3.net5 ;
 wire \proj__3.net6 ;
 wire \proj__3.net7 ;
 wire \proj__3.net8 ;
 wire \proj__4.net100 ;
 wire \proj__4.net101 ;
 wire \proj__4.net102 ;
 wire \proj__4.net103 ;
 wire \proj__4.net104 ;
 wire \proj__4.net105 ;
 wire \proj__4.net106 ;
 wire \proj__4.net109 ;
 wire \proj__4.net110 ;
 wire \proj__4.net111 ;
 wire \proj__4.net112 ;
 wire \proj__4.net113 ;
 wire \proj__4.net114 ;
 wire \proj__4.net115 ;
 wire \proj__4.net116 ;
 wire \proj__4.net117 ;
 wire \proj__4.net118 ;
 wire \proj__4.net119 ;
 wire \proj__4.net120 ;
 wire \proj__4.net121 ;
 wire \proj__4.net122 ;
 wire \proj__4.net125 ;
 wire \proj__4.net126 ;
 wire \proj__4.net127 ;
 wire \proj__4.net128 ;
 wire \proj__4.net129 ;
 wire \proj__4.net130 ;
 wire \proj__4.net131 ;
 wire \proj__4.net132 ;
 wire \proj__4.net133 ;
 wire \proj__4.net134 ;
 wire \proj__4.net135 ;
 wire \proj__4.net136 ;
 wire \proj__4.net137 ;
 wire \proj__4.net138 ;
 wire \proj__4.net139 ;
 wire \proj__4.net140 ;
 wire \proj__4.net16 ;
 wire \proj__4.net17 ;
 wire \proj__4.net18 ;
 wire \proj__4.net2 ;
 wire \proj__4.net20 ;
 wire \proj__4.net21 ;
 wire \proj__4.net22 ;
 wire \proj__4.net23 ;
 wire \proj__4.net24 ;
 wire \proj__4.net25 ;
 wire \proj__4.net26 ;
 wire \proj__4.net27 ;
 wire \proj__4.net28 ;
 wire \proj__4.net29 ;
 wire \proj__4.net3 ;
 wire \proj__4.net30 ;
 wire \proj__4.net31 ;
 wire \proj__4.net32 ;
 wire \proj__4.net33 ;
 wire \proj__4.net34 ;
 wire \proj__4.net35 ;
 wire \proj__4.net36 ;
 wire \proj__4.net37 ;
 wire \proj__4.net38 ;
 wire \proj__4.net4 ;
 wire \proj__4.net40 ;
 wire \proj__4.net41 ;
 wire \proj__4.net42 ;
 wire \proj__4.net44 ;
 wire \proj__4.net46 ;
 wire \proj__4.net47 ;
 wire \proj__4.net48 ;
 wire \proj__4.net49 ;
 wire \proj__4.net5 ;
 wire \proj__4.net50 ;
 wire \proj__4.net51 ;
 wire \proj__4.net52 ;
 wire \proj__4.net53 ;
 wire \proj__4.net54 ;
 wire \proj__4.net55 ;
 wire \proj__4.net56 ;
 wire \proj__4.net57 ;
 wire \proj__4.net58 ;
 wire \proj__4.net6 ;
 wire \proj__4.net60 ;
 wire \proj__4.net62 ;
 wire \proj__4.net63 ;
 wire \proj__4.net64 ;
 wire \proj__4.net65 ;
 wire \proj__4.net66 ;
 wire \proj__4.net67 ;
 wire \proj__4.net68 ;
 wire \proj__4.net69 ;
 wire \proj__4.net7 ;
 wire \proj__4.net70 ;
 wire \proj__4.net71 ;
 wire \proj__4.net72 ;
 wire \proj__4.net73 ;
 wire \proj__4.net74 ;
 wire \proj__4.net77 ;
 wire \proj__4.net78 ;
 wire \proj__4.net79 ;
 wire \proj__4.net8 ;
 wire \proj__4.net80 ;
 wire \proj__4.net81 ;
 wire \proj__4.net82 ;
 wire \proj__4.net83 ;
 wire \proj__4.net84 ;
 wire \proj__4.net85 ;
 wire \proj__4.net86 ;
 wire \proj__4.net87 ;
 wire \proj__4.net88 ;
 wire \proj__4.net89 ;
 wire \proj__4.net9 ;
 wire \proj__4.net90 ;
 wire \proj__4.net92 ;
 wire \proj__4.net94 ;
 wire \proj__4.net95 ;
 wire \proj__4.net96 ;
 wire \proj__4.net97 ;
 wire \proj__4.net98 ;
 wire \proj__4.net99 ;
 wire \proj__5.net12 ;
 wire \proj__5.net13 ;
 wire \proj__5.net14 ;
 wire \proj__5.net6 ;
 wire \proj__6.net10 ;
 wire \proj__6.net100 ;
 wire \proj__6.net101 ;
 wire \proj__6.net102 ;
 wire \proj__6.net103 ;
 wire \proj__6.net104 ;
 wire \proj__6.net105 ;
 wire \proj__6.net106 ;
 wire \proj__6.net107 ;
 wire \proj__6.net11 ;
 wire \proj__6.net12 ;
 wire \proj__6.net13 ;
 wire \proj__6.net14 ;
 wire \proj__6.net15 ;
 wire \proj__6.net16 ;
 wire \proj__6.net17 ;
 wire \proj__6.net20 ;
 wire \proj__6.net21 ;
 wire \proj__6.net23 ;
 wire \proj__6.net24 ;
 wire \proj__6.net25 ;
 wire \proj__6.net26 ;
 wire \proj__6.net27 ;
 wire \proj__6.net28 ;
 wire \proj__6.net29 ;
 wire \proj__6.net30 ;
 wire \proj__6.net31 ;
 wire \proj__6.net32 ;
 wire \proj__6.net33 ;
 wire \proj__6.net34 ;
 wire \proj__6.net35 ;
 wire \proj__6.net36 ;
 wire \proj__6.net37 ;
 wire \proj__6.net38 ;
 wire \proj__6.net39 ;
 wire \proj__6.net40 ;
 wire \proj__6.net41 ;
 wire \proj__6.net42 ;
 wire \proj__6.net43 ;
 wire \proj__6.net44 ;
 wire \proj__6.net45 ;
 wire \proj__6.net46 ;
 wire \proj__6.net47 ;
 wire \proj__6.net48 ;
 wire \proj__6.net49 ;
 wire \proj__6.net50 ;
 wire \proj__6.net51 ;
 wire \proj__6.net52 ;
 wire \proj__6.net53 ;
 wire \proj__6.net54 ;
 wire \proj__6.net55 ;
 wire \proj__6.net56 ;
 wire \proj__6.net57 ;
 wire \proj__6.net58 ;
 wire \proj__6.net59 ;
 wire \proj__6.net60 ;
 wire \proj__6.net61 ;
 wire \proj__6.net62 ;
 wire \proj__6.net63 ;
 wire \proj__6.net64 ;
 wire \proj__6.net65 ;
 wire \proj__6.net66 ;
 wire \proj__6.net72 ;
 wire \proj__6.net74 ;
 wire \proj__6.net75 ;
 wire \proj__6.net76 ;
 wire \proj__6.net77 ;
 wire \proj__6.net78 ;
 wire \proj__6.net79 ;
 wire \proj__6.net80 ;
 wire \proj__6.net81 ;
 wire \proj__6.net82 ;
 wire \proj__6.net83 ;
 wire \proj__6.net84 ;
 wire \proj__6.net85 ;
 wire \proj__6.net86 ;
 wire \proj__6.net87 ;
 wire \proj__6.net88 ;
 wire \proj__6.net90 ;
 wire \proj__6.net91 ;
 wire \proj__6.net92 ;
 wire \proj__6.net93 ;
 wire \proj__6.net94 ;
 wire \proj__6.net95 ;
 wire \proj__6.net96 ;
 wire \proj__6.net97 ;
 wire \proj__6.net98 ;
 wire \proj__6.net99 ;
 wire \proj__7.net11 ;
 wire \proj__7.net12 ;
 wire \proj__7.net4 ;
 wire \proj__7.net5 ;
 wire \proj__9.net15 ;
 wire \proj__9.net16 ;
 wire \proj__9.net18 ;
 wire \proj__9.net19 ;
 wire \proj__9.net20 ;
 wire \proj__9.net5 ;
 wire \proj__9.net6 ;
 wire \proj__9.net7 ;
 wire \proj__9.net8 ;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire \proj_10.flop1/_0_ ;
 wire \proj_10.flop1/_1_ ;
 wire net266;
 wire net267;
 wire \proj_10.flop1/notq ;
 wire \proj_10.flop10/_0_ ;
 wire \proj_10.flop10/_1_ ;
 wire net268;
 wire net269;
 wire \proj_10.flop10/notq ;
 wire \proj_10.flop11/_0_ ;
 wire \proj_10.flop11/_1_ ;
 wire net270;
 wire net271;
 wire \proj_10.flop11/notq ;
 wire \proj_10.flop12/_0_ ;
 wire \proj_10.flop12/_1_ ;
 wire net272;
 wire net273;
 wire \proj_10.flop12/notq ;
 wire \proj_10.flop13/_0_ ;
 wire \proj_10.flop13/_1_ ;
 wire net274;
 wire net275;
 wire \proj_10.flop13/notq ;
 wire \proj_10.flop14/_0_ ;
 wire \proj_10.flop14/_1_ ;
 wire net276;
 wire net277;
 wire \proj_10.flop14/notq ;
 wire \proj_10.flop2/_0_ ;
 wire \proj_10.flop2/_1_ ;
 wire net278;
 wire net279;
 wire \proj_10.flop2/notq ;
 wire \proj_10.flop3/_0_ ;
 wire \proj_10.flop3/_1_ ;
 wire net280;
 wire net281;
 wire \proj_10.flop3/notq ;
 wire \proj_10.flop4/_0_ ;
 wire \proj_10.flop4/_1_ ;
 wire net282;
 wire net283;
 wire \proj_10.flop4/notq ;
 wire \proj_10.flop5/_0_ ;
 wire \proj_10.flop5/_1_ ;
 wire net284;
 wire net285;
 wire \proj_10.flop5/notq ;
 wire \proj_10.flop6/_0_ ;
 wire \proj_10.flop6/_1_ ;
 wire net286;
 wire net287;
 wire \proj_10.flop6/notq ;
 wire \proj_10.flop7/_0_ ;
 wire \proj_10.flop7/_1_ ;
 wire net288;
 wire net289;
 wire \proj_10.flop7/notq ;
 wire \proj_10.flop8/_0_ ;
 wire \proj_10.flop8/_1_ ;
 wire net290;
 wire net291;
 wire \proj_10.flop8/notq ;
 wire \proj_10.flop9/_0_ ;
 wire \proj_10.flop9/_1_ ;
 wire net292;
 wire net293;
 wire \proj_10.flop9/notq ;
 wire \proj_12.flop1/_0_ ;
 wire \proj_12.flop1/_1_ ;
 wire net294;
 wire net295;
 wire \proj_12.flop2/_0_ ;
 wire \proj_12.flop2/_1_ ;
 wire net296;
 wire net297;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire \proj__4.flop1/notq ;
 wire net458;
 wire \proj__4.flop2/notq ;
 wire net459;
 wire \proj__4.flop3/notq ;
 wire \proj__4.flop4/notq ;
 wire \proj__6.flop0/_0_ ;
 wire \proj__6.flop0/_1_ ;
 wire net298;
 wire net299;
 wire \proj__6.flop0/notq ;
 wire \proj__6.flop1/_0_ ;
 wire \proj__6.flop1/_1_ ;
 wire net300;
 wire net301;
 wire \proj__6.flop1/notq ;
 wire \proj__6.flop10/_0_ ;
 wire \proj__6.flop10/_1_ ;
 wire net302;
 wire net303;
 wire \proj__6.flop10/notq ;
 wire \proj__6.flop11/_0_ ;
 wire \proj__6.flop11/_1_ ;
 wire net304;
 wire net305;
 wire \proj__6.flop11/notq ;
 wire \proj__6.flop12/_0_ ;
 wire \proj__6.flop12/_1_ ;
 wire net306;
 wire net307;
 wire \proj__6.flop12/notq ;
 wire \proj__6.flop13/_0_ ;
 wire \proj__6.flop13/_1_ ;
 wire net308;
 wire net309;
 wire \proj__6.flop13/notq ;
 wire \proj__6.flop14/_0_ ;
 wire \proj__6.flop14/_1_ ;
 wire net310;
 wire net311;
 wire \proj__6.flop14/notq ;
 wire \proj__6.flop15/_0_ ;
 wire \proj__6.flop15/_1_ ;
 wire net312;
 wire net313;
 wire \proj__6.flop15/notq ;
 wire \proj__6.flop16/_0_ ;
 wire \proj__6.flop16/_1_ ;
 wire net314;
 wire net315;
 wire \proj__6.flop16/notq ;
 wire \proj__6.flop17/_0_ ;
 wire \proj__6.flop17/_1_ ;
 wire net316;
 wire net317;
 wire \proj__6.flop17/notq ;
 wire \proj__6.flop18/_0_ ;
 wire \proj__6.flop18/_1_ ;
 wire net318;
 wire net319;
 wire \proj__6.flop18/notq ;
 wire \proj__6.flop19/_0_ ;
 wire \proj__6.flop19/_1_ ;
 wire net320;
 wire net321;
 wire \proj__6.flop19/notq ;
 wire \proj__6.flop2/_0_ ;
 wire \proj__6.flop2/_1_ ;
 wire net322;
 wire net323;
 wire \proj__6.flop2/notq ;
 wire \proj__6.flop20/_0_ ;
 wire \proj__6.flop20/_1_ ;
 wire net324;
 wire net325;
 wire \proj__6.flop20/notq ;
 wire \proj__6.flop21/_0_ ;
 wire \proj__6.flop21/_1_ ;
 wire net326;
 wire net327;
 wire \proj__6.flop21/notq ;
 wire \proj__6.flop22/_0_ ;
 wire \proj__6.flop22/_1_ ;
 wire net328;
 wire net329;
 wire \proj__6.flop22/notq ;
 wire \proj__6.flop23/_0_ ;
 wire \proj__6.flop23/_1_ ;
 wire net330;
 wire net331;
 wire \proj__6.flop23/notq ;
 wire \proj__6.flop24/_0_ ;
 wire \proj__6.flop24/_1_ ;
 wire net332;
 wire net333;
 wire \proj__6.flop24/notq ;
 wire \proj__6.flop25/_0_ ;
 wire \proj__6.flop25/_1_ ;
 wire net334;
 wire net335;
 wire \proj__6.flop25/notq ;
 wire \proj__6.flop26/_0_ ;
 wire \proj__6.flop26/_1_ ;
 wire net336;
 wire net337;
 wire \proj__6.flop26/notq ;
 wire \proj__6.flop27/_0_ ;
 wire \proj__6.flop27/_1_ ;
 wire net338;
 wire net339;
 wire \proj__6.flop27/notq ;
 wire \proj__6.flop28/_0_ ;
 wire \proj__6.flop28/_1_ ;
 wire net340;
 wire net341;
 wire \proj__6.flop28/notq ;
 wire \proj__6.flop29/_0_ ;
 wire \proj__6.flop29/_1_ ;
 wire net342;
 wire net343;
 wire \proj__6.flop29/notq ;
 wire \proj__6.flop3/_0_ ;
 wire \proj__6.flop3/_1_ ;
 wire net344;
 wire net345;
 wire \proj__6.flop3/notq ;
 wire \proj__6.flop30/_0_ ;
 wire \proj__6.flop30/_1_ ;
 wire net346;
 wire net347;
 wire \proj__6.flop30/notq ;
 wire \proj__6.flop31/_0_ ;
 wire \proj__6.flop31/_1_ ;
 wire net348;
 wire net349;
 wire \proj__6.flop31/notq ;
 wire \proj__6.flop33/_0_ ;
 wire \proj__6.flop33/_1_ ;
 wire net350;
 wire net351;
 wire \proj__6.flop33/notq ;
 wire \proj__6.flop34/_0_ ;
 wire \proj__6.flop34/_1_ ;
 wire net352;
 wire net353;
 wire \proj__6.flop34/notq ;
 wire \proj__6.flop35/_0_ ;
 wire \proj__6.flop35/_1_ ;
 wire net354;
 wire net355;
 wire \proj__6.flop35/notq ;
 wire \proj__6.flop36/_0_ ;
 wire \proj__6.flop36/_1_ ;
 wire net356;
 wire net357;
 wire \proj__6.flop36/notq ;
 wire \proj__6.flop37/_0_ ;
 wire \proj__6.flop37/_1_ ;
 wire net358;
 wire net359;
 wire \proj__6.flop37/notq ;
 wire \proj__6.flop38/_0_ ;
 wire \proj__6.flop38/_1_ ;
 wire net360;
 wire net361;
 wire \proj__6.flop38/notq ;
 wire \proj__6.flop39/_0_ ;
 wire \proj__6.flop39/_1_ ;
 wire net362;
 wire net363;
 wire \proj__6.flop39/notq ;
 wire \proj__6.flop4/_0_ ;
 wire \proj__6.flop4/_1_ ;
 wire net364;
 wire net365;
 wire \proj__6.flop4/notq ;
 wire \proj__6.flop40/_0_ ;
 wire \proj__6.flop40/_1_ ;
 wire net366;
 wire net367;
 wire \proj__6.flop40/notq ;
 wire \proj__6.flop5/_0_ ;
 wire \proj__6.flop5/_1_ ;
 wire net368;
 wire net369;
 wire \proj__6.flop5/notq ;
 wire \proj__6.flop6/_0_ ;
 wire \proj__6.flop6/_1_ ;
 wire net370;
 wire net371;
 wire \proj__6.flop6/notq ;
 wire \proj__6.flop7/_0_ ;
 wire \proj__6.flop7/_1_ ;
 wire net372;
 wire net373;
 wire \proj__6.flop7/notq ;
 wire \proj__6.flop8/_0_ ;
 wire \proj__6.flop8/_1_ ;
 wire net374;
 wire net375;
 wire \proj__6.flop8/notq ;
 wire \proj__6.flop9/_0_ ;
 wire \proj__6.flop9/_1_ ;
 wire net376;
 wire net377;
 wire \proj__6.flop9/notq ;
 wire \proj__9.flop1/_0_ ;
 wire \proj__9.flop1/_1_ ;
 wire net378;
 wire net379;
 wire \proj__9.flop1/notq ;
 wire \proj__9.flop2/_0_ ;
 wire \proj__9.flop2/_1_ ;
 wire net380;
 wire net381;
 wire \proj__9.flop2/notq ;
 wire \proj__9.flop3/_0_ ;
 wire \proj__9.flop3/_1_ ;
 wire net382;
 wire net383;
 wire \proj__9.flop3/notq ;
 wire \proj__9.flop4/_0_ ;
 wire \proj__9.flop4/_1_ ;
 wire net384;
 wire net385;
 wire \proj__9.flop4/notq ;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;

 sg13g2_inv_1 _339_ (.Y(_059_),
    .A(net143));
 sg13g2_inv_1 _340_ (.Y(_060_),
    .A(\proj__0.net10 ));
 sg13g2_inv_1 _341_ (.Y(_061_),
    .A(\proj__0.net11 ));
 sg13g2_and2_2 _342_ (.A(net6),
    .B(net7),
    .X(_062_));
 sg13g2_nor2b_2 _343_ (.A(net9),
    .B_N(net8),
    .Y(_063_));
 sg13g2_nand3_1 _344_ (.B(_062_),
    .C(_063_),
    .A(\proj__7.net5 ),
    .Y(_064_));
 sg13g2_nand2_2 _345_ (.Y(_065_),
    .A(net8),
    .B(net9));
 sg13g2_nor2_1 _346_ (.A(net6),
    .B(net7),
    .Y(_066_));
 sg13g2_nor2b_2 _347_ (.A(_065_),
    .B_N(_066_),
    .Y(_067_));
 sg13g2_nand2_1 _348_ (.Y(_068_),
    .A(\proj_12.net11 ),
    .B(_067_));
 sg13g2_nor2b_1 _349_ (.A(net6),
    .B_N(net7),
    .Y(_069_));
 sg13g2_nor2b_1 _350_ (.A(net8),
    .B_N(net9),
    .Y(_070_));
 sg13g2_and2_2 _351_ (.A(_069_),
    .B(_070_),
    .X(_071_));
 sg13g2_nor2_1 _352_ (.A(net8),
    .B(net9),
    .Y(_072_));
 sg13g2_or2_1 _353_ (.X(_073_),
    .B(net9),
    .A(net8));
 sg13g2_nand2_1 _354_ (.Y(_074_),
    .A(net9),
    .B(_062_));
 sg13g2_o21ai_1 _355_ (.B1(_074_),
    .Y(_000_),
    .A1(_062_),
    .A2(_073_));
 sg13g2_and2_2 _356_ (.A(_063_),
    .B(_069_),
    .X(_001_));
 sg13g2_and2_2 _357_ (.A(_063_),
    .B(_066_),
    .X(_002_));
 sg13g2_a22oi_1 _358_ (.Y(_003_),
    .B1(_002_),
    .B2(\proj__4.net9 ),
    .A2(_000_),
    .A1(net131));
 sg13g2_a22oi_1 _359_ (.Y(_004_),
    .B1(_001_),
    .B2(\proj__6.net17 ),
    .A2(_071_),
    .A1(\proj_10.net18 ));
 sg13g2_nand4_1 _360_ (.B(_068_),
    .C(_003_),
    .A(_064_),
    .Y(uo_out[7]),
    .D(_004_));
 sg13g2_and2_1 _361_ (.A(_062_),
    .B(_070_),
    .X(_005_));
 sg13g2_a22oi_1 _362_ (.Y(_006_),
    .B1(_005_),
    .B2(\proj_11.net9 ),
    .A2(_001_),
    .A1(\proj__6.net10 ));
 sg13g2_nand3_1 _363_ (.B(_062_),
    .C(_063_),
    .A(\proj__7.net4 ),
    .Y(_007_));
 sg13g2_nor2b_2 _364_ (.A(net7),
    .B_N(net6),
    .Y(_008_));
 sg13g2_nand3_1 _365_ (.B(_063_),
    .C(_008_),
    .A(\proj__5.net6 ),
    .Y(_009_));
 sg13g2_and2_2 _366_ (.A(_062_),
    .B(_072_),
    .X(_010_));
 sg13g2_and2_2 _367_ (.A(_072_),
    .B(_008_),
    .X(_011_));
 sg13g2_a22oi_1 _368_ (.Y(_012_),
    .B1(_011_),
    .B2(\proj__1.net10 ),
    .A2(_010_),
    .A1(\proj__3.net2 ));
 sg13g2_nand4_1 _369_ (.B(_007_),
    .C(_009_),
    .A(_006_),
    .Y(_013_),
    .D(_012_));
 sg13g2_nor2b_2 _370_ (.A(_065_),
    .B_N(_008_),
    .Y(_014_));
 sg13g2_a22oi_1 _371_ (.Y(_015_),
    .B1(_014_),
    .B2(\proj_13.net10 ),
    .A2(_071_),
    .A1(\proj_10.net11 ));
 sg13g2_nand3b_1 _372_ (.B(net7),
    .C(\proj_14.net3 ),
    .Y(_016_),
    .A_N(net6));
 sg13g2_nor2_1 _373_ (.A(_065_),
    .B(_016_),
    .Y(_017_));
 sg13g2_a21oi_1 _374_ (.A1(\proj_12.net7 ),
    .A2(_067_),
    .Y(_018_),
    .B1(_017_));
 sg13g2_and3_2 _375_ (.X(_019_),
    .A(net8),
    .B(net9),
    .C(_062_));
 sg13g2_and2_2 _376_ (.A(_070_),
    .B(_008_),
    .X(_020_));
 sg13g2_a22oi_1 _377_ (.Y(_021_),
    .B1(_020_),
    .B2(\proj__9.net5 ),
    .A2(_019_),
    .A1(\proj_15.net9 ));
 sg13g2_and2_1 _378_ (.A(_069_),
    .B(_072_),
    .X(_022_));
 sg13g2_a22oi_1 _379_ (.Y(_023_),
    .B1(_022_),
    .B2(\proj__2.net6 ),
    .A2(_002_),
    .A1(\proj__4.net2 ));
 sg13g2_nand4_1 _380_ (.B(_018_),
    .C(_021_),
    .A(_015_),
    .Y(_024_),
    .D(_023_));
 sg13g2_or2_1 _381_ (.X(uo_out[0]),
    .B(_024_),
    .A(_013_));
 sg13g2_and2_1 _382_ (.A(_066_),
    .B(_072_),
    .X(_025_));
 sg13g2_or4_1 _383_ (.A(net6),
    .B(net7),
    .C(net8),
    .D(net9),
    .X(_026_));
 sg13g2_o21ai_1 _384_ (.B1(_026_),
    .Y(_027_),
    .A1(_065_),
    .A2(_016_));
 sg13g2_a221oi_1 _385_ (.B2(\proj__4.net3 ),
    .C1(_027_),
    .B1(_002_),
    .A1(\proj__6.net11 ),
    .Y(_028_),
    .A2(_001_));
 sg13g2_a22oi_1 _386_ (.Y(_029_),
    .B1(_020_),
    .B2(\proj__9.net6 ),
    .A2(_014_),
    .A1(\proj_13.net11 ));
 sg13g2_a22oi_1 _387_ (.Y(_030_),
    .B1(_019_),
    .B2(\proj_15.net10 ),
    .A2(_071_),
    .A1(\proj_10.net12 ));
 sg13g2_a22oi_1 _388_ (.Y(_031_),
    .B1(_010_),
    .B2(\proj__3.net3 ),
    .A2(_067_),
    .A1(\proj_12.net8 ));
 sg13g2_and2_1 _389_ (.A(_030_),
    .B(_031_),
    .X(_032_));
 sg13g2_a22oi_1 _390_ (.Y(_033_),
    .B1(_011_),
    .B2(\proj__1.net11 ),
    .A2(_005_),
    .A1(\proj_11.net10 ));
 sg13g2_and3_1 _391_ (.X(_034_),
    .A(_028_),
    .B(_029_),
    .C(_033_));
 sg13g2_a22oi_1 _392_ (.Y(uo_out[1]),
    .B1(_032_),
    .B2(_034_),
    .A2(_025_),
    .A1(_059_));
 sg13g2_nand2_1 _393_ (.Y(_035_),
    .A(\proj_15.net11 ),
    .B(_019_));
 sg13g2_a221oi_1 _394_ (.B2(\proj__4.net4 ),
    .C1(_027_),
    .B1(_002_),
    .A1(\proj__6.net12 ),
    .Y(_036_),
    .A2(_001_));
 sg13g2_a22oi_1 _395_ (.Y(_037_),
    .B1(_010_),
    .B2(\proj__3.net4 ),
    .A2(_067_),
    .A1(\proj_12.net9 ));
 sg13g2_a22oi_1 _396_ (.Y(_038_),
    .B1(_020_),
    .B2(\proj__9.net7 ),
    .A2(_005_),
    .A1(\proj_11.net11 ));
 sg13g2_a22oi_1 _397_ (.Y(_039_),
    .B1(_014_),
    .B2(\proj_13.net12 ),
    .A2(_071_),
    .A1(\proj_10.net13 ));
 sg13g2_and4_1 _398_ (.A(_035_),
    .B(_037_),
    .C(_038_),
    .D(_039_),
    .X(_040_));
 sg13g2_a22oi_1 _399_ (.Y(uo_out[2]),
    .B1(_036_),
    .B2(_040_),
    .A2(_025_),
    .A1(_060_));
 sg13g2_and2_1 _400_ (.A(\proj_11.net12 ),
    .B(_005_),
    .X(_041_));
 sg13g2_a221oi_1 _401_ (.B2(\proj__3.net5 ),
    .C1(_041_),
    .B1(_010_),
    .A1(\proj__6.net13 ),
    .Y(_042_),
    .A2(_001_));
 sg13g2_a22oi_1 _402_ (.Y(_043_),
    .B1(_014_),
    .B2(\proj_13.net13 ),
    .A2(_002_),
    .A1(\proj__4.net5 ));
 sg13g2_a22oi_1 _403_ (.Y(_044_),
    .B1(_020_),
    .B2(\proj__9.net8 ),
    .A2(_067_),
    .A1(\proj_12.net10 ));
 sg13g2_a21oi_1 _404_ (.A1(\proj_10.net14 ),
    .A2(_071_),
    .Y(_045_),
    .B1(_025_));
 sg13g2_a22oi_1 _405_ (.Y(_046_),
    .B1(_019_),
    .B2(\proj_15.net12 ),
    .A2(_011_),
    .A1(\proj__1.net12 ));
 sg13g2_and4_1 _406_ (.A(_043_),
    .B(_044_),
    .C(_045_),
    .D(_046_),
    .X(_047_));
 sg13g2_a22oi_1 _407_ (.Y(uo_out[3]),
    .B1(_042_),
    .B2(_047_),
    .A2(_025_),
    .A1(_061_));
 sg13g2_o21ai_1 _408_ (.B1(_074_),
    .Y(_048_),
    .A1(net6),
    .A2(_073_));
 sg13g2_o21ai_1 _409_ (.B1(net136),
    .Y(_049_),
    .A1(_067_),
    .A2(_048_));
 sg13g2_a22oi_1 _410_ (.Y(_050_),
    .B1(_011_),
    .B2(\proj__1.net13 ),
    .A2(_071_),
    .A1(\proj_10.net15 ));
 sg13g2_a22oi_1 _411_ (.Y(_051_),
    .B1(_010_),
    .B2(\proj__3.net6 ),
    .A2(_002_),
    .A1(\proj__4.net6 ));
 sg13g2_a22oi_1 _412_ (.Y(_052_),
    .B1(_014_),
    .B2(\proj_13.net14 ),
    .A2(_001_),
    .A1(\proj__6.net14 ));
 sg13g2_nand4_1 _413_ (.B(_050_),
    .C(_051_),
    .A(_049_),
    .Y(uo_out[4]),
    .D(_052_));
 sg13g2_a22oi_1 _414_ (.Y(_053_),
    .B1(_048_),
    .B2(net134),
    .A2(_001_),
    .A1(\proj__6.net15 ));
 sg13g2_a22oi_1 _415_ (.Y(_054_),
    .B1(_014_),
    .B2(\proj_13.net15 ),
    .A2(_010_),
    .A1(\proj__3.net7 ));
 sg13g2_a22oi_1 _416_ (.Y(_055_),
    .B1(_002_),
    .B2(\proj__4.net7 ),
    .A2(_071_),
    .A1(\proj_10.net16 ));
 sg13g2_nand3_1 _417_ (.B(_054_),
    .C(_055_),
    .A(_053_),
    .Y(uo_out[5]));
 sg13g2_a22oi_1 _418_ (.Y(_056_),
    .B1(_002_),
    .B2(\proj__4.net8 ),
    .A2(_000_),
    .A1(net132));
 sg13g2_a22oi_1 _419_ (.Y(_057_),
    .B1(_010_),
    .B2(\proj__3.net8 ),
    .A2(_071_),
    .A1(\proj_10.net17 ));
 sg13g2_a22oi_1 _420_ (.Y(_058_),
    .B1(_014_),
    .B2(\proj_13.net16 ),
    .A2(_001_),
    .A1(\proj__6.net16 ));
 sg13g2_nand3_1 _421_ (.B(_057_),
    .C(_058_),
    .A(_056_),
    .Y(uo_out[6]));
 sg13g2_tiehi \proj__4.mux106/_0__345  (.L_HI(net386));
 sg13g2_tiehi \proj__4.mux107/_0__346  (.L_HI(net387));
 sg13g2_tiehi \proj__4.mux107/_0__347  (.L_HI(net388));
 sg13g2_tiehi \proj__4.mux108/_0__348  (.L_HI(net389));
 sg13g2_tiehi \proj__4.mux108/_0__349  (.L_HI(net390));
 sg13g2_tiehi \proj__4.mux109/_0__350  (.L_HI(net391));
 sg13g2_tiehi \proj__4.mux109/_0__351  (.L_HI(net392));
 sg13g2_tiehi \proj__4.mux110/_0__352  (.L_HI(net393));
 sg13g2_tiehi \proj__4.mux111/_0__353  (.L_HI(net394));
 sg13g2_tiehi \proj__4.mux111/_0__354  (.L_HI(net395));
 sg13g2_tiehi \proj__4.mux112/_0__355  (.L_HI(net396));
 sg13g2_tiehi \proj__4.mux112/_0__356  (.L_HI(net397));
 sg13g2_tiehi \proj__4.mux113/_0__357  (.L_HI(net398));
 sg13g2_tiehi \proj__4.mux113/_0__358  (.L_HI(net399));
 sg13g2_tiehi \proj__4.mux3/_0__359  (.L_HI(net400));
 sg13g2_tiehi \proj__4.mux32/_0__360  (.L_HI(net401));
 sg13g2_tiehi \proj__4.mux33/_0__361  (.L_HI(net402));
 sg13g2_tiehi \proj__4.mux34/_0__362  (.L_HI(net403));
 sg13g2_tiehi \proj__4.mux34/_0__363  (.L_HI(net404));
 sg13g2_tiehi \proj__4.mux38/_0__364  (.L_HI(net405));
 sg13g2_tiehi \proj__4.mux4/_0__365  (.L_HI(net406));
 sg13g2_tiehi \proj__4.mux4/_0__366  (.L_HI(net407));
 sg13g2_tiehi \proj__4.mux47/_0__367  (.L_HI(net408));
 sg13g2_tiehi \proj__4.mux47/_0__368  (.L_HI(net409));
 sg13g2_tiehi \proj__4.mux48/_0__369  (.L_HI(net410));
 sg13g2_tiehi \proj__4.mux50/_0__370  (.L_HI(net411));
 sg13g2_tiehi \proj__4.mux50/_0__371  (.L_HI(net412));
 sg13g2_tiehi \proj__4.mux52/_0__372  (.L_HI(net413));
 sg13g2_tiehi \proj__4.mux53/_0__373  (.L_HI(net414));
 sg13g2_tiehi \proj__4.mux53/_0__374  (.L_HI(net415));
 sg13g2_tiehi \proj__4.mux61/_0__375  (.L_HI(net416));
 sg13g2_tiehi \proj__4.mux62/_0__376  (.L_HI(net417));
 sg13g2_tiehi \proj__4.mux63/_0__377  (.L_HI(net418));
 sg13g2_tiehi \proj__4.mux63/_0__378  (.L_HI(net419));
 sg13g2_tiehi \proj__4.mux64/_0__379  (.L_HI(net420));
 sg13g2_tiehi \proj__4.mux65/_0__380  (.L_HI(net421));
 sg13g2_tiehi \proj__4.mux65/_0__381  (.L_HI(net422));
 sg13g2_tiehi \proj__4.mux66/_0__382  (.L_HI(net423));
 sg13g2_tiehi \proj__4.mux67/_0__383  (.L_HI(net424));
 sg13g2_tiehi \proj__4.mux67/_0__384  (.L_HI(net425));
 sg13g2_tiehi \proj__4.mux68/_0__385  (.L_HI(net426));
 sg13g2_tiehi \proj__4.mux76/_0__386  (.L_HI(net427));
 sg13g2_tiehi \proj__4.mux76/_0__387  (.L_HI(net428));
 sg13g2_tiehi \proj__4.mux77/_0__388  (.L_HI(net429));
 sg13g2_tiehi \proj__4.mux78/_0__389  (.L_HI(net430));
 sg13g2_tiehi \proj__4.mux78/_0__390  (.L_HI(net431));
 sg13g2_tiehi \proj__4.mux79/_0__391  (.L_HI(net432));
 sg13g2_tiehi \proj__4.mux79/_0__392  (.L_HI(net433));
 sg13g2_tiehi \proj__4.mux8/_0__393  (.L_HI(net434));
 sg13g2_tiehi \proj__4.mux80/_0__394  (.L_HI(net435));
 sg13g2_tiehi \proj__4.mux80/_0__395  (.L_HI(net436));
 sg13g2_tiehi \proj__4.mux81/_0__396  (.L_HI(net437));
 sg13g2_tiehi \proj__4.mux81/_0__397  (.L_HI(net438));
 sg13g2_tiehi \proj__4.mux82/_0__398  (.L_HI(net439));
 sg13g2_tiehi \proj__4.mux82/_0__399  (.L_HI(net440));
 sg13g2_tiehi \proj__4.mux83/_0__400  (.L_HI(net441));
 sg13g2_tiehi \proj__4.mux91/_0__401  (.L_HI(net442));
 sg13g2_tiehi \proj__4.mux92/_0__402  (.L_HI(net443));
 sg13g2_tiehi \proj__4.mux93/_0__403  (.L_HI(net444));
 sg13g2_tiehi \proj__4.mux94/_0__404  (.L_HI(net445));
 sg13g2_tiehi \proj__4.mux94/_0__405  (.L_HI(net446));
 sg13g2_tiehi \proj__4.mux96/_0__406  (.L_HI(net447));
 sg13g2_tiehi \proj__4.mux98/_0__407  (.L_HI(net448));
 sg13g2_tiehi \proj__4.mux98/_0__408  (.L_HI(net449));
 sg13g2_tiehi \proj__4.xor1/_0__409  (.L_HI(net450));
 sg13g2_tiehi \proj__2.flop1/_1__410  (.L_HI(net451));
 sg13g2_tielo \proj_10.flop10/dffsr_11  (.L_LO(net11));
 sg13g2_tielo \proj_10.flop10/_5__12  (.L_LO(net12));
 sg13g2_tielo \proj_10.flop11/dffsr_13  (.L_LO(net13));
 sg13g2_tielo \proj_10.flop11/_5__14  (.L_LO(net14));
 sg13g2_tielo \proj_10.flop12/dffsr_15  (.L_LO(net15));
 sg13g2_tielo \proj_10.flop12/_5__16  (.L_LO(net16));
 sg13g2_tielo \proj_10.flop13/dffsr_17  (.L_LO(net17));
 sg13g2_tielo \proj_10.flop13/_5__18  (.L_LO(net18));
 sg13g2_tielo \proj_10.flop14/dffsr_19  (.L_LO(net19));
 sg13g2_tielo \proj_10.flop14/_5__20  (.L_LO(net20));
 sg13g2_tielo \proj_10.flop2/dffsr_21  (.L_LO(net21));
 sg13g2_tielo \proj_10.flop3/dffsr_22  (.L_LO(net22));
 sg13g2_tielo \proj_10.flop4/dffsr_23  (.L_LO(net23));
 sg13g2_tielo \proj_10.flop5/dffsr_24  (.L_LO(net24));
 sg13g2_tielo \proj_10.flop6/dffsr_25  (.L_LO(net25));
 sg13g2_tielo \proj_10.flop7/dffsr_26  (.L_LO(net26));
 sg13g2_tielo \proj_10.flop8/dffsr_27  (.L_LO(net27));
 sg13g2_tielo \proj_10.flop9/dffsr_28  (.L_LO(net28));
 sg13g2_tielo \proj_10.mux11/_0__29  (.L_LO(net29));
 sg13g2_tielo \proj_10.mux12/_0__30  (.L_LO(net30));
 sg13g2_tielo \proj_10.mux13/_0__31  (.L_LO(net31));
 sg13g2_tielo \proj_10.mux14/_0__32  (.L_LO(net32));
 sg13g2_tielo \proj_10.mux15/_0__33  (.L_LO(net33));
 sg13g2_tielo \proj_10.mux16/_0__34  (.L_LO(net34));
 sg13g2_tielo \proj_10.mux17/_0__35  (.L_LO(net35));
 sg13g2_tielo \proj_10.mux18/_0__36  (.L_LO(net36));
 sg13g2_tielo \proj_10.mux19/_0__37  (.L_LO(net37));
 sg13g2_tielo \proj_10.mux20/_0__38  (.L_LO(net38));
 sg13g2_tielo \proj_10.mux21/_0__39  (.L_LO(net39));
 sg13g2_tielo \proj_10.mux21/_0__40  (.L_LO(net40));
 sg13g2_tielo \proj_10.mux22/_0__41  (.L_LO(net41));
 sg13g2_tielo \proj_10.mux23/_0__42  (.L_LO(net42));
 sg13g2_tielo \proj_10.mux23/_0__43  (.L_LO(net43));
 sg13g2_tielo \proj_10.mux25/_0__44  (.L_LO(net44));
 sg13g2_tielo \proj_10.mux26/_0__45  (.L_LO(net45));
 sg13g2_tielo \proj_10.mux27/_0__46  (.L_LO(net46));
 sg13g2_tielo \proj_10.mux29/_0__47  (.L_LO(net47));
 sg13g2_tielo \proj_10.mux30/_0__48  (.L_LO(net48));
 sg13g2_tielo \proj_10.mux31/_0__49  (.L_LO(net49));
 sg13g2_tielo \proj_10.mux32/_0__50  (.L_LO(net50));
 sg13g2_tielo \proj_10.mux33/_0__51  (.L_LO(net51));
 sg13g2_tielo \proj_10.mux34/_0__52  (.L_LO(net52));
 sg13g2_tielo \proj_10.mux35/_0__53  (.L_LO(net53));
 sg13g2_tielo \proj_10.mux36/_0__54  (.L_LO(net54));
 sg13g2_tielo \proj_10.not16/_0__55  (.L_LO(net55));
 sg13g2_tielo \proj_10.not6/_0__56  (.L_LO(net56));
 sg13g2_tielo \proj_10.not7/_0__57  (.L_LO(net57));
 sg13g2_tielo \proj_12.flop1/dffsr_58  (.L_LO(net58));
 sg13g2_tielo \proj_12.flop1/_4__59  (.L_LO(net59));
 sg13g2_tielo \proj_12.flop1/_5__60  (.L_LO(net60));
 sg13g2_tielo \proj_12.flop2/_4__61  (.L_LO(net61));
 sg13g2_tielo \proj_12.flop2/_5__62  (.L_LO(net62));
 sg13g2_tielo \proj_14.and1/_0__63  (.L_LO(net63));
 sg13g2_tielo \proj__1.xor1/_0__64  (.L_LO(net64));
 sg13g2_tielo \proj__2.flop1/_1__65  (.L_LO(net65));
 sg13g2_tielo \proj__3.flop1/_1__66  (.L_LO(net66));
 sg13g2_tielo \proj__4.flop1/_1__67  (.L_LO(net67));
 sg13g2_tielo \proj__4.flop2/_1__68  (.L_LO(net68));
 sg13g2_tielo \proj__4.flop3/_1__69  (.L_LO(net69));
 sg13g2_tielo \proj__4.flop4/_1__70  (.L_LO(net70));
 sg13g2_tielo \proj__4.mux1/_0__71  (.L_LO(net71));
 sg13g2_tielo \proj__4.mux1/_0__72  (.L_LO(net72));
 sg13g2_tielo \proj__4.mux106/_0__73  (.L_LO(net73));
 sg13g2_tielo \proj__4.mux110/_0__74  (.L_LO(net74));
 sg13g2_tielo \proj__4.mux2/_0__75  (.L_LO(net75));
 sg13g2_tielo \proj__4.mux2/_0__76  (.L_LO(net76));
 sg13g2_tielo \proj__4.mux3/_0__77  (.L_LO(net77));
 sg13g2_tielo \proj__4.mux31/_0__78  (.L_LO(net78));
 sg13g2_tielo \proj__4.mux31/_0__79  (.L_LO(net79));
 sg13g2_tielo \proj__4.mux32/_0__80  (.L_LO(net80));
 sg13g2_tielo \proj__4.mux33/_0__81  (.L_LO(net81));
 sg13g2_tielo \proj__4.mux35/_0__82  (.L_LO(net82));
 sg13g2_tielo \proj__4.mux35/_0__83  (.L_LO(net83));
 sg13g2_tielo \proj__4.mux36/_0__84  (.L_LO(net84));
 sg13g2_tielo \proj__4.mux36/_0__85  (.L_LO(net85));
 sg13g2_tielo \proj__4.mux37/_0__86  (.L_LO(net86));
 sg13g2_tielo \proj__4.mux37/_0__87  (.L_LO(net87));
 sg13g2_tielo \proj__4.mux38/_0__88  (.L_LO(net88));
 sg13g2_tielo \proj__4.mux46/_0__89  (.L_LO(net89));
 sg13g2_tielo \proj__4.mux46/_0__90  (.L_LO(net90));
 sg13g2_tielo \proj__4.mux48/_0__91  (.L_LO(net91));
 sg13g2_tielo \proj__4.mux49/_0__92  (.L_LO(net92));
 sg13g2_tielo \proj__4.mux49/_0__93  (.L_LO(net93));
 sg13g2_tielo \proj__4.mux5/_0__94  (.L_LO(net94));
 sg13g2_tielo \proj__4.mux5/_0__95  (.L_LO(net95));
 sg13g2_tielo \proj__4.mux51/_0__96  (.L_LO(net96));
 sg13g2_tielo \proj__4.mux51/_0__97  (.L_LO(net97));
 sg13g2_tielo \proj__4.mux52/_0__98  (.L_LO(net98));
 sg13g2_tielo \proj__4.mux6/_0__99  (.L_LO(net99));
 sg13g2_tielo \proj__4.mux6/_0__100  (.L_LO(net100));
 sg13g2_tielo \proj__4.mux61/_0__101  (.L_LO(net101));
 sg13g2_tielo \proj__4.mux62/_0__102  (.L_LO(net102));
 sg13g2_tielo \proj__4.mux64/_0__103  (.L_LO(net103));
 sg13g2_tielo \proj__4.mux66/_0__104  (.L_LO(net104));
 sg13g2_tielo \proj__4.mux68/_0__105  (.L_LO(net105));
 sg13g2_tielo \proj__4.mux7/_0__106  (.L_LO(net106));
 sg13g2_tielo \proj__4.mux7/_0__107  (.L_LO(net107));
 sg13g2_tielo \proj__4.mux77/_0__108  (.L_LO(net108));
 sg13g2_tielo \proj__4.mux8/_0__109  (.L_LO(net109));
 sg13g2_tielo \proj__4.mux83/_0__110  (.L_LO(net110));
 sg13g2_tielo \proj__4.mux91/_0__111  (.L_LO(net111));
 sg13g2_tielo \proj__4.mux92/_0__112  (.L_LO(net112));
 sg13g2_tielo \proj__4.mux93/_0__113  (.L_LO(net113));
 sg13g2_tielo \proj__4.mux95/_0__114  (.L_LO(net114));
 sg13g2_tielo \proj__4.mux95/_0__115  (.L_LO(net115));
 sg13g2_tielo \proj__4.mux96/_0__116  (.L_LO(net116));
 sg13g2_tielo \proj__4.mux97/_0__117  (.L_LO(net117));
 sg13g2_tielo \proj__4.mux97/_0__118  (.L_LO(net118));
 sg13g2_tielo \proj__6.flop0/_4__119  (.L_LO(net119));
 sg13g2_tielo \proj__6.flop0/_5__120  (.L_LO(net120));
 sg13g2_tielo \proj__6.flop1/_4__121  (.L_LO(net121));
 sg13g2_tielo \proj__6.flop1/_5__122  (.L_LO(net122));
 sg13g2_tielo \proj__6.flop10/_4__123  (.L_LO(net123));
 sg13g2_tielo \proj__6.flop10/_5__124  (.L_LO(net124));
 sg13g2_tielo \proj__6.flop11/_4__125  (.L_LO(net125));
 sg13g2_tielo \proj__6.flop11/_5__126  (.L_LO(net126));
 sg13g2_tielo \proj__6.flop12/_4__127  (.L_LO(net168));
 sg13g2_tielo \proj__6.flop12/_5__128  (.L_LO(net169));
 sg13g2_tielo \proj__6.flop13/_4__129  (.L_LO(net170));
 sg13g2_tielo \proj__6.flop13/_5__130  (.L_LO(net171));
 sg13g2_tielo \proj__6.flop14/_4__131  (.L_LO(net172));
 sg13g2_tielo \proj__6.flop14/_5__132  (.L_LO(net173));
 sg13g2_tielo \proj__6.flop15/_4__133  (.L_LO(net174));
 sg13g2_tielo \proj__6.flop15/_5__134  (.L_LO(net175));
 sg13g2_tielo \proj__6.flop16/_4__135  (.L_LO(net176));
 sg13g2_tielo \proj__6.flop16/_5__136  (.L_LO(net177));
 sg13g2_tielo \proj__6.flop17/_4__137  (.L_LO(net178));
 sg13g2_tielo \proj__6.flop17/_5__138  (.L_LO(net179));
 sg13g2_tielo \proj__6.flop18/_4__139  (.L_LO(net180));
 sg13g2_tielo \proj__6.flop18/_5__140  (.L_LO(net181));
 sg13g2_tielo \proj__6.flop19/_4__141  (.L_LO(net182));
 sg13g2_tielo \proj__6.flop19/_5__142  (.L_LO(net183));
 sg13g2_tielo \proj__6.flop2/_4__143  (.L_LO(net184));
 sg13g2_tielo \proj__6.flop2/_5__144  (.L_LO(net185));
 sg13g2_tielo \proj__6.flop20/_4__145  (.L_LO(net186));
 sg13g2_tielo \proj__6.flop20/_5__146  (.L_LO(net187));
 sg13g2_tielo \proj__6.flop21/_4__147  (.L_LO(net188));
 sg13g2_tielo \proj__6.flop21/_5__148  (.L_LO(net189));
 sg13g2_tielo \proj__6.flop22/_4__149  (.L_LO(net190));
 sg13g2_tielo \proj__6.flop22/_5__150  (.L_LO(net191));
 sg13g2_tielo \proj__6.flop23/_4__151  (.L_LO(net192));
 sg13g2_tielo \proj__6.flop23/_5__152  (.L_LO(net193));
 sg13g2_tielo \proj__6.flop24/_4__153  (.L_LO(net194));
 sg13g2_tielo \proj__6.flop24/_5__154  (.L_LO(net195));
 sg13g2_tielo \proj__6.flop25/_4__155  (.L_LO(net196));
 sg13g2_tielo \proj__6.flop25/_5__156  (.L_LO(net197));
 sg13g2_tielo \proj__6.flop26/_4__157  (.L_LO(net198));
 sg13g2_tielo \proj__6.flop26/_5__158  (.L_LO(net199));
 sg13g2_tielo \proj__6.flop27/_4__159  (.L_LO(net200));
 sg13g2_tielo \proj__6.flop27/_5__160  (.L_LO(net201));
 sg13g2_tielo \proj__6.flop28/_4__161  (.L_LO(net202));
 sg13g2_tielo \proj__6.flop28/_5__162  (.L_LO(net203));
 sg13g2_tielo \proj__6.flop29/_4__163  (.L_LO(net204));
 sg13g2_tielo \proj__6.flop29/_5__164  (.L_LO(net205));
 sg13g2_tielo \proj__6.flop3/_4__165  (.L_LO(net206));
 sg13g2_tielo \proj__6.flop3/_5__166  (.L_LO(net207));
 sg13g2_tielo \proj__6.flop30/_4__167  (.L_LO(net208));
 sg13g2_tielo \proj__6.flop30/_5__168  (.L_LO(net209));
 sg13g2_tielo \proj__6.flop31/_4__169  (.L_LO(net210));
 sg13g2_tielo \proj__6.flop31/_5__170  (.L_LO(net211));
 sg13g2_tielo \proj__6.flop33/_4__171  (.L_LO(net212));
 sg13g2_tielo \proj__6.flop33/_5__172  (.L_LO(net213));
 sg13g2_tielo \proj__6.flop34/_4__173  (.L_LO(net214));
 sg13g2_tielo \proj__6.flop34/_5__174  (.L_LO(net215));
 sg13g2_tielo \proj__6.flop35/_4__175  (.L_LO(net216));
 sg13g2_tielo \proj__6.flop35/_5__176  (.L_LO(net217));
 sg13g2_tielo \proj__6.flop36/_4__177  (.L_LO(net218));
 sg13g2_tielo \proj__6.flop36/_5__178  (.L_LO(net219));
 sg13g2_tielo \proj__6.flop37/_4__179  (.L_LO(net220));
 sg13g2_tielo \proj__6.flop37/_5__180  (.L_LO(net221));
 sg13g2_tielo \proj__6.flop38/_4__181  (.L_LO(net222));
 sg13g2_tielo \proj__6.flop38/_5__182  (.L_LO(net223));
 sg13g2_tielo \proj__6.flop39/_4__183  (.L_LO(net224));
 sg13g2_tielo \proj__6.flop39/_5__184  (.L_LO(net225));
 sg13g2_tielo \proj__6.flop4/_4__185  (.L_LO(net226));
 sg13g2_tielo \proj__6.flop4/_5__186  (.L_LO(net227));
 sg13g2_tielo \proj__6.flop40/_4__187  (.L_LO(net228));
 sg13g2_tielo \proj__6.flop40/_5__188  (.L_LO(net229));
 sg13g2_tielo \proj__6.flop5/_4__189  (.L_LO(net230));
 sg13g2_tielo \proj__6.flop5/_5__190  (.L_LO(net231));
 sg13g2_tielo \proj__6.flop6/_4__191  (.L_LO(net232));
 sg13g2_tielo \proj__6.flop6/_5__192  (.L_LO(net233));
 sg13g2_tielo \proj__6.flop7/_4__193  (.L_LO(net234));
 sg13g2_tielo \proj__6.flop7/_5__194  (.L_LO(net235));
 sg13g2_tielo \proj__6.flop8/_4__195  (.L_LO(net236));
 sg13g2_tielo \proj__6.flop8/_5__196  (.L_LO(net237));
 sg13g2_tielo \proj__6.flop9/_4__197  (.L_LO(net238));
 sg13g2_tielo \proj__6.flop9/_5__198  (.L_LO(net239));
 sg13g2_tielo \proj__9.flop1/dffsr_199  (.L_LO(net240));
 sg13g2_tielo \proj__9.flop1/_5__200  (.L_LO(net241));
 sg13g2_tielo \proj__9.flop2/dffsr_201  (.L_LO(net242));
 sg13g2_tielo \proj__9.flop2/_5__202  (.L_LO(net243));
 sg13g2_tielo \proj__9.flop3/dffsr_203  (.L_LO(net244));
 sg13g2_tielo \proj__9.flop3/_5__204  (.L_LO(net245));
 sg13g2_tielo \proj__9.flop4/dffsr_205  (.L_LO(net246));
 sg13g2_tielo \proj__9.flop4/_5__206  (.L_LO(net247));
 sg13g2_tielo \proj__9.not1/_0__207  (.L_LO(net248));
 sg13g2_tielo tt_um_wokwi_group_13_208 (.L_LO(net249));
 sg13g2_tielo tt_um_wokwi_group_13_209 (.L_LO(net250));
 sg13g2_tielo tt_um_wokwi_group_13_210 (.L_LO(net251));
 sg13g2_tielo tt_um_wokwi_group_13_211 (.L_LO(net252));
 sg13g2_tielo tt_um_wokwi_group_13_212 (.L_LO(net253));
 sg13g2_tielo tt_um_wokwi_group_13_213 (.L_LO(net254));
 sg13g2_tielo tt_um_wokwi_group_13_214 (.L_LO(net255));
 sg13g2_tielo tt_um_wokwi_group_13_215 (.L_LO(net256));
 sg13g2_tielo tt_um_wokwi_group_13_216 (.L_LO(net257));
 sg13g2_tielo tt_um_wokwi_group_13_217 (.L_LO(net258));
 sg13g2_tielo tt_um_wokwi_group_13_218 (.L_LO(net259));
 sg13g2_tielo tt_um_wokwi_group_13_219 (.L_LO(net260));
 sg13g2_tielo tt_um_wokwi_group_13_220 (.L_LO(net261));
 sg13g2_tielo tt_um_wokwi_group_13_221 (.L_LO(net262));
 sg13g2_tielo tt_um_wokwi_group_13_222 (.L_LO(net263));
 sg13g2_tielo tt_um_wokwi_group_13_223 (.L_LO(net264));
 sg13g2_tielo \proj_10.flop1/dffsr_224  (.L_LO(net265));
 sg13g2_and2_2 \proj_10.and1/_0_  (.A(net4),
    .B(net3),
    .X(\proj_10.net96 ));
 sg13g2_inv_1 \proj_10.flop1/_4_  (.Y(\proj_10.flop1/_0_ ),
    .A(\proj_10.net43 ));
 sg13g2_inv_1 \proj_10.flop1/_5_  (.Y(\proj_10.flop1/_1_ ),
    .A(\proj_10.net42 ));
 sg13g2_tielo \proj_10.flop1/dffsr_225  (.L_LO(net266));
 sg13g2_tielo \proj_10.flop10/dffsr_226  (.L_LO(net267));
 sg13g2_sdfbbp_1 \proj_10.flop1/dffsr  (.Q(\proj_10.net28 ),
    .Q_N(\proj_10.flop1/notq ),
    .RESET_B(\proj_10.flop1/_0_ ),
    .SET_B(\proj_10.flop1/_1_ ),
    .D(\proj_10.net41 ),
    .SCE(net266),
    .SCD(net265),
    .CLK(net10));
 sg13g2_inv_1 \proj_10.flop10/_4_  (.Y(\proj_10.flop10/_0_ ),
    .A(\proj_10.net82 ));
 sg13g2_inv_1 \proj_10.flop10/_5_  (.Y(\proj_10.flop10/_1_ ),
    .A(net12));
 sg13g2_tielo \proj_10.flop10/dffsr_227  (.L_LO(net268));
 sg13g2_tielo \proj_10.flop11/dffsr_228  (.L_LO(net269));
 sg13g2_sdfbbp_1 \proj_10.flop10/dffsr  (.Q(\proj_10.net83 ),
    .Q_N(\proj_10.flop10/notq ),
    .RESET_B(\proj_10.flop10/_0_ ),
    .SET_B(\proj_10.flop10/_1_ ),
    .D(\proj_10.net80 ),
    .SCE(net268),
    .SCD(net267),
    .CLK(net11));
 sg13g2_inv_1 \proj_10.flop11/_4_  (.Y(\proj_10.flop11/_0_ ),
    .A(\proj_10.net82 ));
 sg13g2_inv_1 \proj_10.flop11/_5_  (.Y(\proj_10.flop11/_1_ ),
    .A(net14));
 sg13g2_tielo \proj_10.flop11/dffsr_229  (.L_LO(net270));
 sg13g2_tielo \proj_10.flop12/dffsr_230  (.L_LO(net271));
 sg13g2_sdfbbp_1 \proj_10.flop11/dffsr  (.Q(\proj_10.net85 ),
    .Q_N(\proj_10.flop11/notq ),
    .RESET_B(\proj_10.flop11/_0_ ),
    .SET_B(\proj_10.flop11/_1_ ),
    .D(\proj_10.net83 ),
    .SCE(net270),
    .SCD(net269),
    .CLK(net13));
 sg13g2_inv_1 \proj_10.flop12/_4_  (.Y(\proj_10.flop12/_0_ ),
    .A(\proj_10.net82 ));
 sg13g2_inv_1 \proj_10.flop12/_5_  (.Y(\proj_10.flop12/_1_ ),
    .A(net16));
 sg13g2_tielo \proj_10.flop12/dffsr_231  (.L_LO(net272));
 sg13g2_tielo \proj_10.flop13/dffsr_232  (.L_LO(net273));
 sg13g2_sdfbbp_1 \proj_10.flop12/dffsr  (.Q(\proj_10.net87 ),
    .Q_N(\proj_10.flop12/notq ),
    .RESET_B(\proj_10.flop12/_0_ ),
    .SET_B(\proj_10.flop12/_1_ ),
    .D(\proj_10.net85 ),
    .SCE(net272),
    .SCD(net271),
    .CLK(net15));
 sg13g2_inv_1 \proj_10.flop13/_4_  (.Y(\proj_10.flop13/_0_ ),
    .A(\proj_10.net82 ));
 sg13g2_inv_1 \proj_10.flop13/_5_  (.Y(\proj_10.flop13/_1_ ),
    .A(net18));
 sg13g2_tielo \proj_10.flop13/dffsr_233  (.L_LO(net274));
 sg13g2_tielo \proj_10.flop14/dffsr_234  (.L_LO(net275));
 sg13g2_sdfbbp_1 \proj_10.flop13/dffsr  (.Q(\proj_10.net89 ),
    .Q_N(\proj_10.flop13/notq ),
    .RESET_B(\proj_10.flop13/_0_ ),
    .SET_B(\proj_10.flop13/_1_ ),
    .D(\proj_10.net87 ),
    .SCE(net274),
    .SCD(net273),
    .CLK(net17));
 sg13g2_inv_1 \proj_10.flop14/_4_  (.Y(\proj_10.flop14/_0_ ),
    .A(\proj_10.net82 ));
 sg13g2_inv_1 \proj_10.flop14/_5_  (.Y(\proj_10.flop14/_1_ ),
    .A(net20));
 sg13g2_tielo \proj_10.flop14/dffsr_235  (.L_LO(net276));
 sg13g2_tielo \proj_10.flop2/dffsr_236  (.L_LO(net277));
 sg13g2_sdfbbp_1 \proj_10.flop14/dffsr  (.Q(\proj_10.net71 ),
    .Q_N(\proj_10.flop14/notq ),
    .RESET_B(\proj_10.flop14/_0_ ),
    .SET_B(\proj_10.flop14/_1_ ),
    .D(\proj_10.net89 ),
    .SCE(net276),
    .SCD(net275),
    .CLK(net19));
 sg13g2_inv_1 \proj_10.flop2/_4_  (.Y(\proj_10.flop2/_0_ ),
    .A(\proj_10.net45 ));
 sg13g2_inv_1 \proj_10.flop2/_5_  (.Y(\proj_10.flop2/_1_ ),
    .A(\proj_10.net44 ));
 sg13g2_tielo \proj_10.flop2/dffsr_237  (.L_LO(net278));
 sg13g2_tielo \proj_10.flop3/dffsr_238  (.L_LO(net279));
 sg13g2_sdfbbp_1 \proj_10.flop2/dffsr  (.Q(\proj_10.net33 ),
    .Q_N(\proj_10.flop2/notq ),
    .RESET_B(\proj_10.flop2/_0_ ),
    .SET_B(\proj_10.flop2/_1_ ),
    .D(\proj_10.net28 ),
    .SCE(net278),
    .SCD(net277),
    .CLK(net21));
 sg13g2_inv_1 \proj_10.flop3/_4_  (.Y(\proj_10.flop3/_0_ ),
    .A(\proj_10.net47 ));
 sg13g2_inv_1 \proj_10.flop3/_5_  (.Y(\proj_10.flop3/_1_ ),
    .A(\proj_10.net46 ));
 sg13g2_tielo \proj_10.flop3/dffsr_239  (.L_LO(net280));
 sg13g2_tielo \proj_10.flop4/dffsr_240  (.L_LO(net281));
 sg13g2_sdfbbp_1 \proj_10.flop3/dffsr  (.Q(\proj_10.net48 ),
    .Q_N(\proj_10.flop3/notq ),
    .RESET_B(\proj_10.flop3/_0_ ),
    .SET_B(\proj_10.flop3/_1_ ),
    .D(\proj_10.net33 ),
    .SCE(net280),
    .SCD(net279),
    .CLK(net22));
 sg13g2_inv_1 \proj_10.flop4/_4_  (.Y(\proj_10.flop4/_0_ ),
    .A(\proj_10.net50 ));
 sg13g2_inv_1 \proj_10.flop4/_5_  (.Y(\proj_10.flop4/_1_ ),
    .A(\proj_10.net49 ));
 sg13g2_tielo \proj_10.flop4/dffsr_241  (.L_LO(net282));
 sg13g2_tielo \proj_10.flop5/dffsr_242  (.L_LO(net283));
 sg13g2_sdfbbp_1 \proj_10.flop4/dffsr  (.Q(\proj_10.net51 ),
    .Q_N(\proj_10.flop4/notq ),
    .RESET_B(\proj_10.flop4/_0_ ),
    .SET_B(\proj_10.flop4/_1_ ),
    .D(\proj_10.net48 ),
    .SCE(net282),
    .SCD(net281),
    .CLK(net23));
 sg13g2_inv_1 \proj_10.flop5/_4_  (.Y(\proj_10.flop5/_0_ ),
    .A(\proj_10.net53 ));
 sg13g2_inv_1 \proj_10.flop5/_5_  (.Y(\proj_10.flop5/_1_ ),
    .A(\proj_10.net52 ));
 sg13g2_tielo \proj_10.flop5/dffsr_243  (.L_LO(net284));
 sg13g2_tielo \proj_10.flop6/dffsr_244  (.L_LO(net285));
 sg13g2_sdfbbp_1 \proj_10.flop5/dffsr  (.Q(\proj_10.net54 ),
    .Q_N(\proj_10.flop5/notq ),
    .RESET_B(\proj_10.flop5/_0_ ),
    .SET_B(\proj_10.flop5/_1_ ),
    .D(\proj_10.net51 ),
    .SCE(net284),
    .SCD(net283),
    .CLK(net24));
 sg13g2_inv_1 \proj_10.flop6/_4_  (.Y(\proj_10.flop6/_0_ ),
    .A(\proj_10.net56 ));
 sg13g2_inv_1 \proj_10.flop6/_5_  (.Y(\proj_10.flop6/_1_ ),
    .A(\proj_10.net55 ));
 sg13g2_tielo \proj_10.flop6/dffsr_245  (.L_LO(net286));
 sg13g2_tielo \proj_10.flop7/dffsr_246  (.L_LO(net287));
 sg13g2_sdfbbp_1 \proj_10.flop6/dffsr  (.Q(\proj_10.net57 ),
    .Q_N(\proj_10.flop6/notq ),
    .RESET_B(\proj_10.flop6/_0_ ),
    .SET_B(\proj_10.flop6/_1_ ),
    .D(\proj_10.net54 ),
    .SCE(net286),
    .SCD(net285),
    .CLK(net25));
 sg13g2_inv_1 \proj_10.flop7/_4_  (.Y(\proj_10.flop7/_0_ ),
    .A(\proj_10.net73 ));
 sg13g2_inv_1 \proj_10.flop7/_5_  (.Y(\proj_10.flop7/_1_ ),
    .A(\proj_10.net72 ));
 sg13g2_tielo \proj_10.flop7/dffsr_247  (.L_LO(net288));
 sg13g2_tielo \proj_10.flop8/dffsr_248  (.L_LO(net289));
 sg13g2_sdfbbp_1 \proj_10.flop7/dffsr  (.Q(\proj_10.net74 ),
    .Q_N(\proj_10.flop7/notq ),
    .RESET_B(\proj_10.flop7/_0_ ),
    .SET_B(\proj_10.flop7/_1_ ),
    .D(\proj_10.net71 ),
    .SCE(net288),
    .SCD(net287),
    .CLK(net26));
 sg13g2_inv_1 \proj_10.flop8/_4_  (.Y(\proj_10.flop8/_0_ ),
    .A(\proj_10.net76 ));
 sg13g2_inv_1 \proj_10.flop8/_5_  (.Y(\proj_10.flop8/_1_ ),
    .A(\proj_10.net75 ));
 sg13g2_tielo \proj_10.flop8/dffsr_249  (.L_LO(net290));
 sg13g2_tielo \proj_10.flop9/dffsr_250  (.L_LO(net291));
 sg13g2_sdfbbp_1 \proj_10.flop8/dffsr  (.Q(\proj_10.net77 ),
    .Q_N(\proj_10.flop8/notq ),
    .RESET_B(\proj_10.flop8/_0_ ),
    .SET_B(\proj_10.flop8/_1_ ),
    .D(\proj_10.net74 ),
    .SCE(net290),
    .SCD(net289),
    .CLK(net27));
 sg13g2_inv_1 \proj_10.flop9/_4_  (.Y(\proj_10.flop9/_0_ ),
    .A(\proj_10.net79 ));
 sg13g2_inv_1 \proj_10.flop9/_5_  (.Y(\proj_10.flop9/_1_ ),
    .A(\proj_10.net78 ));
 sg13g2_tielo \proj_10.flop9/dffsr_251  (.L_LO(net292));
 sg13g2_tielo \proj_12.flop1/dffsr_252  (.L_LO(net293));
 sg13g2_sdfbbp_1 \proj_10.flop9/dffsr  (.Q(\proj_10.net80 ),
    .Q_N(\proj_10.flop9/notq ),
    .RESET_B(\proj_10.flop9/_0_ ),
    .SET_B(\proj_10.flop9/_1_ ),
    .D(\proj_10.net77 ),
    .SCE(net292),
    .SCD(net291),
    .CLK(net28));
 sg13g2_mux2_1 \proj_10.mux1/_0_  (.A0(\proj_10.net24 ),
    .A1(\proj_10.net25 ),
    .S(net5),
    .X(\proj_10.net12 ));
 sg13g2_mux2_1 \proj_10.mux10/_0_  (.A0(\proj_10.net38 ),
    .A1(\proj_10.net37 ),
    .S(\proj_10.net30 ),
    .X(\proj_10.net40 ));
 sg13g2_mux2_1 \proj_10.mux11/_0_  (.A0(net29),
    .A1(net148),
    .S(\proj_10.net59 ),
    .X(\proj_10.net42 ));
 sg13g2_mux2_1 \proj_10.mux12/_0_  (.A0(net30),
    .A1(\proj_10.net60 ),
    .S(\proj_10.net59 ),
    .X(\proj_10.net43 ));
 sg13g2_mux2_1 \proj_10.mux13/_0_  (.A0(net31),
    .A1(net146),
    .S(\proj_10.net59 ),
    .X(\proj_10.net44 ));
 sg13g2_mux2_1 \proj_10.mux14/_0_  (.A0(net32),
    .A1(\proj_10.net61 ),
    .S(\proj_10.net59 ),
    .X(\proj_10.net45 ));
 sg13g2_mux2_1 \proj_10.mux15/_0_  (.A0(net33),
    .A1(net142),
    .S(\proj_10.net59 ),
    .X(\proj_10.net46 ));
 sg13g2_mux2_1 \proj_10.mux16/_0_  (.A0(net34),
    .A1(\proj_10.net62 ),
    .S(\proj_10.net59 ),
    .X(\proj_10.net47 ));
 sg13g2_mux2_1 \proj_10.mux17/_0_  (.A0(net35),
    .A1(net139),
    .S(\proj_10.net59 ),
    .X(\proj_10.net49 ));
 sg13g2_mux2_1 \proj_10.mux18/_0_  (.A0(net36),
    .A1(\proj_10.net63 ),
    .S(\proj_10.net59 ),
    .X(\proj_10.net50 ));
 sg13g2_mux2_1 \proj_10.mux19/_0_  (.A0(net37),
    .A1(net137),
    .S(\proj_10.net59 ),
    .X(\proj_10.net52 ));
 sg13g2_mux2_1 \proj_10.mux2/_0_  (.A0(\proj_10.net25 ),
    .A1(\proj_10.net24 ),
    .S(net5),
    .X(\proj_10.net16 ));
 sg13g2_mux2_1 \proj_10.mux20/_0_  (.A0(net38),
    .A1(\proj_10.net64 ),
    .S(\proj_10.net59 ),
    .X(\proj_10.net53 ));
 sg13g2_mux2_1 \proj_10.mux21/_0_  (.A0(net39),
    .A1(net40),
    .S(\proj_10.net59 ),
    .X(\proj_10.net55 ));
 sg13g2_mux2_1 \proj_10.mux22/_0_  (.A0(net41),
    .A1(\proj_10.net66 ),
    .S(\proj_10.net59 ),
    .X(\proj_10.net56 ));
 sg13g2_mux2_1 \proj_10.mux23/_0_  (.A0(net42),
    .A1(net43),
    .S(net129),
    .X(\proj_10.net18 ));
 sg13g2_mux2_1 \proj_10.mux24/_0_  (.A0(\proj_10.net57 ),
    .A1(\proj_10.net51 ),
    .S(net133),
    .X(\proj_10.net41 ));
 sg13g2_mux2_1 \proj_10.mux25/_0_  (.A0(\proj_10.net48 ),
    .A1(net44),
    .S(net133),
    .X(\proj_10.net34 ));
 sg13g2_mux2_1 \proj_10.mux26/_0_  (.A0(\proj_10.net51 ),
    .A1(net45),
    .S(net133),
    .X(\proj_10.net29 ));
 sg13g2_mux2_1 \proj_10.mux27/_0_  (.A0(\proj_10.net54 ),
    .A1(net46),
    .S(net133),
    .X(\proj_10.net37 ));
 sg13g2_mux2_1 \proj_10.mux28/_0_  (.A0(\proj_10.net57 ),
    .A1(\proj_10.net51 ),
    .S(net133),
    .X(\proj_10.net38 ));
 sg13g2_mux2_1 \proj_10.mux29/_0_  (.A0(net47),
    .A1(\proj_10.net48 ),
    .S(net133),
    .X(\proj_10.net69 ));
 sg13g2_mux2_1 \proj_10.mux3/_0_  (.A0(\proj_10.net26 ),
    .A1(\proj_10.net27 ),
    .S(net132),
    .X(\proj_10.net13 ));
 sg13g2_mux2_2 \proj_10.mux30/_0_  (.A0(net48),
    .A1(net137),
    .S(net133),
    .X(\proj_10.net30 ));
 sg13g2_mux2_1 \proj_10.mux31/_0_  (.A0(net49),
    .A1(net1),
    .S(\proj_10.net82 ),
    .X(\proj_10.net72 ));
 sg13g2_mux2_1 \proj_10.mux32/_0_  (.A0(net50),
    .A1(\proj_10.net92 ),
    .S(\proj_10.net82 ),
    .X(\proj_10.net73 ));
 sg13g2_mux2_1 \proj_10.mux33/_0_  (.A0(net51),
    .A1(net146),
    .S(\proj_10.net82 ),
    .X(\proj_10.net75 ));
 sg13g2_mux2_1 \proj_10.mux34/_0_  (.A0(net52),
    .A1(\proj_10.net93 ),
    .S(\proj_10.net82 ),
    .X(\proj_10.net76 ));
 sg13g2_mux2_1 \proj_10.mux35/_0_  (.A0(net53),
    .A1(net142),
    .S(\proj_10.net82 ),
    .X(\proj_10.net78 ));
 sg13g2_mux2_1 \proj_10.mux36/_0_  (.A0(net54),
    .A1(\proj_10.net94 ),
    .S(\proj_10.net82 ),
    .X(\proj_10.net79 ));
 sg13g2_mux2_1 \proj_10.mux37/_0_  (.A0(\proj_10.net31 ),
    .A1(\proj_10.net74 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net11 ));
 sg13g2_mux2_1 \proj_10.mux38/_0_  (.A0(\proj_10.net35 ),
    .A1(\proj_10.net77 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net24 ));
 sg13g2_mux2_1 \proj_10.mux39/_0_  (.A0(\proj_10.net36 ),
    .A1(\proj_10.net87 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net26 ));
 sg13g2_mux2_1 \proj_10.mux4/_0_  (.A0(\proj_10.net27 ),
    .A1(\proj_10.net26 ),
    .S(net132),
    .X(\proj_10.net15 ));
 sg13g2_mux2_1 \proj_10.mux40/_0_  (.A0(\proj_10.net32 ),
    .A1(\proj_10.net85 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net14 ));
 sg13g2_mux2_1 \proj_10.mux41/_0_  (.A0(\proj_10.net39 ),
    .A1(\proj_10.net83 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net27 ));
 sg13g2_mux2_1 \proj_10.mux42/_0_  (.A0(\proj_10.net40 ),
    .A1(\proj_10.net71 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net25 ));
 sg13g2_mux2_1 \proj_10.mux43/_0_  (.A0(\proj_10.net69 ),
    .A1(\proj_10.net95 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net17 ));
 sg13g2_mux2_1 \proj_10.mux5/_0_  (.A0(\proj_10.net28 ),
    .A1(\proj_10.net29 ),
    .S(\proj_10.net30 ),
    .X(\proj_10.net31 ));
 sg13g2_mux2_1 \proj_10.mux6/_0_  (.A0(\proj_10.net29 ),
    .A1(\proj_10.net28 ),
    .S(\proj_10.net30 ),
    .X(\proj_10.net32 ));
 sg13g2_mux2_1 \proj_10.mux7/_0_  (.A0(\proj_10.net33 ),
    .A1(\proj_10.net34 ),
    .S(\proj_10.net30 ),
    .X(\proj_10.net35 ));
 sg13g2_mux2_1 \proj_10.mux8/_0_  (.A0(\proj_10.net34 ),
    .A1(\proj_10.net33 ),
    .S(\proj_10.net30 ),
    .X(\proj_10.net36 ));
 sg13g2_mux2_1 \proj_10.mux9/_0_  (.A0(\proj_10.net37 ),
    .A1(\proj_10.net38 ),
    .S(\proj_10.net30 ),
    .X(\proj_10.net39 ));
 sg13g2_inv_1 \proj_10.not1/_0_  (.Y(\proj_10.net60 ),
    .A(net148));
 sg13g2_inv_1 \proj_10.not10/_0_  (.Y(\proj_10.net94 ),
    .A(net142));
 sg13g2_inv_1 \proj_10.not16/_0_  (.Y(\proj_10.net82 ),
    .A(net55));
 sg13g2_inv_1 \proj_10.not2/_0_  (.Y(\proj_10.net61 ),
    .A(net146));
 sg13g2_inv_1 \proj_10.not3/_0_  (.Y(\proj_10.net62 ),
    .A(net142));
 sg13g2_inv_1 \proj_10.not4/_0_  (.Y(\proj_10.net63 ),
    .A(net139));
 sg13g2_inv_1 \proj_10.not5/_0_  (.Y(\proj_10.net64 ),
    .A(net137));
 sg13g2_inv_1 \proj_10.not6/_0_  (.Y(\proj_10.net66 ),
    .A(net56));
 sg13g2_inv_1 \proj_10.not7/_0_  (.Y(\proj_10.net59 ),
    .A(net57));
 sg13g2_inv_1 \proj_10.not8/_0_  (.Y(\proj_10.net92 ),
    .A(net148));
 sg13g2_inv_1 \proj_10.not9/_0_  (.Y(\proj_10.net93 ),
    .A(net146));
 sg13g2_or2_1 \proj_10.or1/_0_  (.X(\proj_10.net95 ),
    .B(\proj_10.net80 ),
    .A(\proj_10.net89 ));
 sg13g2_inv_1 \proj_11.not1/_0_  (.Y(\proj_11.net9 ),
    .A(net147));
 sg13g2_inv_1 \proj_11.not2/_0_  (.Y(\proj_11.net10 ),
    .A(net143));
 sg13g2_inv_1 \proj_11.not3/_0_  (.Y(\proj_11.net11 ),
    .A(net141));
 sg13g2_inv_1 \proj_11.not4/_0_  (.Y(\proj_11.net12 ),
    .A(net138));
 sg13g2_inv_1 \proj_12.flop1/_4_  (.Y(\proj_12.flop1/_0_ ),
    .A(net59));
 sg13g2_inv_1 \proj_12.flop1/_5_  (.Y(\proj_12.flop1/_1_ ),
    .A(net60));
 sg13g2_tielo \proj_12.flop1/dffsr_253  (.L_LO(net294));
 sg13g2_tielo \proj_12.flop2/dffsr_254  (.L_LO(net295));
 sg13g2_sdfbbp_1 \proj_12.flop1/dffsr  (.Q(\proj_12.net19 ),
    .Q_N(\proj_12.net17 ),
    .RESET_B(\proj_12.flop1/_0_ ),
    .SET_B(\proj_12.flop1/_1_ ),
    .D(\proj_12.net17 ),
    .SCE(net294),
    .SCD(net293),
    .CLK(net58));
 sg13g2_inv_1 \proj_12.flop2/_4_  (.Y(\proj_12.flop2/_0_ ),
    .A(net61));
 sg13g2_inv_1 \proj_12.flop2/_5_  (.Y(\proj_12.flop2/_1_ ),
    .A(net62));
 sg13g2_tielo \proj_12.flop2/dffsr_255  (.L_LO(net296));
 sg13g2_tielo \proj__6.flop0/dffsr_256  (.L_LO(net297));
 sg13g2_sdfbbp_1 \proj_12.flop2/dffsr  (.Q(\proj_12.net11 ),
    .Q_N(\proj_12.net20 ),
    .RESET_B(\proj_12.flop2/_0_ ),
    .SET_B(\proj_12.flop2/_1_ ),
    .D(\proj_12.net20 ),
    .SCE(net296),
    .SCD(net295),
    .CLK(\proj_12.net19 ));
 sg13g2_inv_1 \proj_12.not1/_0_  (.Y(\proj_12.net7 ),
    .A(net148));
 sg13g2_inv_1 \proj_12.not2/_0_  (.Y(\proj_12.net8 ),
    .A(net143));
 sg13g2_inv_1 \proj_12.not3/_0_  (.Y(\proj_12.net9 ),
    .A(net141));
 sg13g2_inv_1 \proj_12.not4/_0_  (.Y(\proj_12.net10 ),
    .A(net138));
 sg13g2_or2_1 \proj_13.or1/_0_  (.X(\proj_13.net22 ),
    .B(net132),
    .A(net130));
 sg13g2_or2_1 \proj_13.or10/_0_  (.X(\proj_13.net30 ),
    .B(net148),
    .A(net2));
 sg13g2_or2_1 \proj_13.or11/_0_  (.X(\proj_13.net31 ),
    .B(\proj_13.net30 ),
    .A(net137));
 sg13g2_or2_1 \proj_13.or12/_0_  (.X(\proj_13.net32 ),
    .B(\proj_13.net31 ),
    .A(net138));
 sg13g2_or2_1 \proj_13.or13/_0_  (.X(\proj_13.net33 ),
    .B(\proj_13.net32 ),
    .A(net134));
 sg13g2_or2_1 \proj_13.or14/_0_  (.X(\proj_13.net34 ),
    .B(\proj_13.net33 ),
    .A(net132));
 sg13g2_or2_1 \proj_13.or15/_0_  (.X(\proj_13.net12 ),
    .B(\proj_13.net34 ),
    .A(net131));
 sg13g2_or2_1 \proj_13.or16/_0_  (.X(\proj_13.net35 ),
    .B(net145),
    .A(net140));
 sg13g2_or2_1 \proj_13.or17/_0_  (.X(\proj_13.net27 ),
    .B(\proj_13.net26 ),
    .A(net147));
 sg13g2_or2_1 \proj_13.or18/_0_  (.X(\proj_13.net36 ),
    .B(net135),
    .A(\proj_13.net35 ));
 sg13g2_or2_1 \proj_13.or19/_0_  (.X(\proj_13.net37 ),
    .B(net134),
    .A(\proj_13.net36 ));
 sg13g2_or2_1 \proj_13.or2/_0_  (.X(\proj_13.net23 ),
    .B(net134),
    .A(\proj_13.net22 ));
 sg13g2_or2_1 \proj_13.or20/_0_  (.X(\proj_13.net13 ),
    .B(net129),
    .A(\proj_13.net37 ));
 sg13g2_or2_1 \proj_13.or21/_0_  (.X(\proj_13.net38 ),
    .B(net145),
    .A(net134));
 sg13g2_or2_1 \proj_13.or22/_0_  (.X(\proj_13.net14 ),
    .B(net130),
    .A(\proj_13.net38 ));
 sg13g2_or2_1 \proj_13.or23/_0_  (.X(\proj_13.net39 ),
    .B(net134),
    .A(net136));
 sg13g2_or2_1 \proj_13.or24/_0_  (.X(\proj_13.net40 ),
    .B(net138),
    .A(\proj_13.net39 ));
 sg13g2_or2_1 \proj_13.or25/_0_  (.X(\proj_13.net15 ),
    .B(net129),
    .A(\proj_13.net40 ));
 sg13g2_or2_1 \proj_13.or26/_0_  (.X(\proj_13.net41 ),
    .B(net140),
    .A(net145));
 sg13g2_or2_1 \proj_13.or27/_0_  (.X(\proj_13.net42 ),
    .B(net139),
    .A(\proj_13.net41 ));
 sg13g2_or2_1 \proj_13.or28/_0_  (.X(\proj_13.net43 ),
    .B(net135),
    .A(\proj_13.net42 ));
 sg13g2_or2_1 \proj_13.or29/_0_  (.X(\proj_13.net44 ),
    .B(net134),
    .A(\proj_13.net43 ));
 sg13g2_or2_1 \proj_13.or3/_0_  (.X(\proj_13.net24 ),
    .B(net137),
    .A(\proj_13.net23 ));
 sg13g2_or2_1 \proj_13.or30/_0_  (.X(\proj_13.net16 ),
    .B(net129),
    .A(\proj_13.net44 ));
 sg13g2_or2_1 \proj_13.or4/_0_  (.X(\proj_13.net25 ),
    .B(net2),
    .A(\proj_13.net24 ));
 sg13g2_or2_1 \proj_13.or5/_0_  (.X(\proj_13.net10 ),
    .B(net144),
    .A(\proj_13.net25 ));
 sg13g2_or2_1 \proj_13.or6/_0_  (.X(\proj_13.net26 ),
    .B(net143),
    .A(net141));
 sg13g2_or2_1 \proj_13.or7/_0_  (.X(\proj_13.net28 ),
    .B(\proj_13.net27 ),
    .A(net138));
 sg13g2_or2_1 \proj_13.or8/_0_  (.X(\proj_13.net29 ),
    .B(\proj_13.net28 ),
    .A(net132));
 sg13g2_or2_1 \proj_13.or9/_0_  (.X(\proj_13.net11 ),
    .B(\proj_13.net29 ),
    .A(net131));
 sg13g2_and2_1 \proj_14.and1/_0_  (.A(net132),
    .B(net63),
    .X(\proj_14.net3 ));
 sg13g2_inv_1 \proj_15.not2/_0_  (.Y(\proj_15.net10 ),
    .A(net144));
 sg13g2_inv_1 \proj_15.not3/_0_  (.Y(\proj_15.net11 ),
    .A(net141));
 sg13g2_inv_1 \proj_15.not4/_0_  (.Y(\proj_15.net12 ),
    .A(net138));
 sg13g2_xor2_1 \proj_15.xor1/_0_  (.B(net147),
    .A(net143),
    .X(\proj_15.net9 ));
 sg13g2_inv_1 \proj__0.not1/_0_  (.Y(\proj__0.net10 ),
    .A(net147));
 sg13g2_or2_1 \proj__0.or1/_0_  (.X(\proj__0.net11 ),
    .B(net140),
    .A(net138));
 sg13g2_nand2_1 \proj__1.nand1/_0_  (.Y(\proj__1.net10 ),
    .A(net143),
    .B(net147));
 sg13g2_inv_1 \proj__1.not1/_0_  (.Y(\proj__1.net12 ),
    .A(net136));
 sg13g2_or2_1 \proj__1.or1/_0_  (.X(\proj__1.net11 ),
    .B(net140),
    .A(net138));
 sg13g2_xor2_1 \proj__1.xor1/_0_  (.B(net64),
    .A(net134),
    .X(\proj__1.net13 ));
 sg13g2_dfrbp_1 \proj__2.flop1/_1_  (.CLK(net65),
    .RESET_B(net451),
    .D(\proj__2.net12 ),
    .Q_N(\proj__2.net12 ),
    .Q(\proj__2.net13 ));
 sg13g2_tiehi \proj__2.flop2/_1__411  (.L_HI(net452));
 sg13g2_dfrbp_1 \proj__2.flop2/_1_  (.CLK(\proj__2.net13 ),
    .RESET_B(net452),
    .D(\proj__2.net14 ),
    .Q_N(\proj__2.net14 ),
    .Q(\proj__2.net6 ));
 sg13g2_tiehi \proj__3.flop1/_1__412  (.L_HI(net453));
 sg13g2_and2_1 \proj__3.and10/_0_  (.A(\proj__3.net14 ),
    .B(\proj__3.net24 ),
    .X(\proj__3.net6 ));
 sg13g2_and2_1 \proj__3.and11/_0_  (.A(\proj__3.net17 ),
    .B(\proj__3.net18 ),
    .X(\proj__3.net25 ));
 sg13g2_and2_1 \proj__3.and12/_0_  (.A(\proj__3.net15 ),
    .B(\proj__3.net25 ),
    .X(\proj__3.net5 ));
 sg13g2_and2_1 \proj__3.and13/_0_  (.A(\proj__3.net17 ),
    .B(\proj__3.net18 ),
    .X(\proj__3.net26 ));
 sg13g2_and2_1 \proj__3.and14/_0_  (.A(\proj__3.net14 ),
    .B(\proj__3.net26 ),
    .X(\proj__3.net4 ));
 sg13g2_and2_1 \proj__3.and15/_0_  (.A(\proj__3.net16 ),
    .B(\proj__3.net18 ),
    .X(\proj__3.net27 ));
 sg13g2_and2_1 \proj__3.and16/_0_  (.A(\proj__3.net15 ),
    .B(\proj__3.net27 ),
    .X(\proj__3.net28 ));
 sg13g2_and2_1 \proj__3.and17/_0_  (.A(\proj__3.net16 ),
    .B(\proj__3.net18 ),
    .X(\proj__3.net29 ));
 sg13g2_and2_1 \proj__3.and18/_0_  (.A(\proj__3.net14 ),
    .B(\proj__3.net29 ),
    .X(\proj__3.net7 ));
 sg13g2_and2_1 \proj__3.and3/_0_  (.A(\proj__3.net17 ),
    .B(\proj__3.net15 ),
    .X(\proj__3.net20 ));
 sg13g2_and2_1 \proj__3.and4/_0_  (.A(\proj__3.net19 ),
    .B(\proj__3.net20 ),
    .X(\proj__3.net2 ));
 sg13g2_and2_1 \proj__3.and5/_0_  (.A(\proj__3.net17 ),
    .B(\proj__3.net19 ),
    .X(\proj__3.net21 ));
 sg13g2_and2_1 \proj__3.and6/_0_  (.A(\proj__3.net14 ),
    .B(\proj__3.net21 ),
    .X(\proj__3.net3 ));
 sg13g2_and2_1 \proj__3.and7/_0_  (.A(\proj__3.net16 ),
    .B(\proj__3.net19 ),
    .X(\proj__3.net22 ));
 sg13g2_and2_1 \proj__3.and8/_0_  (.A(\proj__3.net15 ),
    .B(\proj__3.net22 ),
    .X(\proj__3.net23 ));
 sg13g2_and2_1 \proj__3.and9/_0_  (.A(\proj__3.net16 ),
    .B(\proj__3.net19 ),
    .X(\proj__3.net24 ));
 sg13g2_dfrbp_1 \proj__3.flop1/_1_  (.CLK(net66),
    .RESET_B(net453),
    .D(\proj__3.net14 ),
    .Q_N(\proj__3.net14 ),
    .Q(\proj__3.net15 ));
 sg13g2_tiehi \proj__3.flop2/_1__413  (.L_HI(net454));
 sg13g2_dfrbp_1 \proj__3.flop2/_1_  (.CLK(\proj__3.net15 ),
    .RESET_B(net454),
    .D(\proj__3.net16 ),
    .Q_N(\proj__3.net16 ),
    .Q(\proj__3.net17 ));
 sg13g2_tiehi \proj__3.flop3/_1__414  (.L_HI(net455));
 sg13g2_dfrbp_1 \proj__3.flop3/_1_  (.CLK(\proj__3.net17 ),
    .RESET_B(net455),
    .D(\proj__3.net18 ),
    .Q_N(\proj__3.net18 ),
    .Q(\proj__3.net19 ));
 sg13g2_tiehi \proj__4.flop1/_1__415  (.L_HI(net456));
 sg13g2_or2_1 \proj__3.or1/_0_  (.X(\proj__3.net8 ),
    .B(\proj__3.net23 ),
    .A(\proj__3.net28 ));
 sg13g2_and2_1 \proj__4.and1/_0_  (.A(net385),
    .B(net157),
    .X(\proj__4.net40 ));
 sg13g2_and2_1 \proj__4.and2/_0_  (.A(\proj__4.net40 ),
    .B(net152),
    .X(\proj__4.net41 ));
 sg13g2_and2_1 \proj__4.and3/_0_  (.A(\proj__4.net41 ),
    .B(net150),
    .X(\proj__4.net42 ));
 sg13g2_and2_1 \proj__4.and5/_0_  (.A(net154),
    .B(net166),
    .X(\proj__4.net139 ));
 sg13g2_and2_1 \proj__4.and6/_0_  (.A(\proj__4.net34 ),
    .B(net151),
    .X(\proj__4.net140 ));
 sg13g2_and2_1 \proj__4.and7/_0_  (.A(\proj__4.net140 ),
    .B(\proj__4.net139 ),
    .X(\proj__4.net9 ));
 sg13g2_dfrbp_1 \proj__4.flop1/_1_  (.CLK(net67),
    .RESET_B(net456),
    .D(\proj__4.net35 ),
    .Q_N(\proj__4.flop1/notq ),
    .Q(\proj__4.net16 ));
 sg13g2_tiehi \proj__4.flop2/_1__416  (.L_HI(net457));
 sg13g2_dfrbp_1 \proj__4.flop2/_1_  (.CLK(net68),
    .RESET_B(net457),
    .D(\proj__4.net36 ),
    .Q_N(\proj__4.flop2/notq ),
    .Q(\proj__4.net26 ));
 sg13g2_tiehi \proj__4.flop3/_1__417  (.L_HI(net458));
 sg13g2_dfrbp_1 \proj__4.flop3/_1_  (.CLK(net69),
    .RESET_B(net458),
    .D(\proj__4.net37 ),
    .Q_N(\proj__4.flop3/notq ),
    .Q(\proj__4.net31 ));
 sg13g2_tiehi \proj__4.flop4/_1__418  (.L_HI(net459));
 sg13g2_dfrbp_1 \proj__4.flop4/_1_  (.CLK(net70),
    .RESET_B(net459),
    .D(\proj__4.net38 ),
    .Q_N(\proj__4.flop4/notq ),
    .Q(\proj__4.net34 ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_mux2_1 \proj__4.mux1/_0_  (.A0(net71),
    .A1(net72),
    .S(net163),
    .X(\proj__4.net17 ));
 sg13g2_mux2_1 \proj__4.mux10/_0_  (.A0(\proj__4.net20 ),
    .A1(\proj__4.net21 ),
    .S(net153),
    .X(\proj__4.net28 ));
 sg13g2_mux2_1 \proj__4.mux100/_0_  (.A0(\proj__4.net111 ),
    .A1(\proj__4.net112 ),
    .S(net155),
    .X(\proj__4.net118 ));
 sg13g2_mux2_1 \proj__4.mux101/_0_  (.A0(\proj__4.net113 ),
    .A1(\proj__4.net114 ),
    .S(net155),
    .X(\proj__4.net119 ));
 sg13g2_mux2_1 \proj__4.mux102/_0_  (.A0(\proj__4.net115 ),
    .A1(\proj__4.net116 ),
    .S(net155),
    .X(\proj__4.net120 ));
 sg13g2_mux2_1 \proj__4.mux103/_0_  (.A0(\proj__4.net119 ),
    .A1(\proj__4.net120 ),
    .S(\proj__4.net31 ),
    .X(\proj__4.net121 ));
 sg13g2_mux2_1 \proj__4.mux104/_0_  (.A0(\proj__4.net117 ),
    .A1(\proj__4.net118 ),
    .S(\proj__4.net31 ),
    .X(\proj__4.net122 ));
 sg13g2_mux2_1 \proj__4.mux105/_0_  (.A0(\proj__4.net122 ),
    .A1(\proj__4.net121 ),
    .S(net149),
    .X(\proj__4.net7 ));
 sg13g2_mux2_1 \proj__4.mux106/_0_  (.A0(net386),
    .A1(net73),
    .S(net162),
    .X(\proj__4.net125 ));
 sg13g2_mux2_1 \proj__4.mux107/_0_  (.A0(net387),
    .A1(net388),
    .S(net162),
    .X(\proj__4.net126 ));
 sg13g2_mux2_1 \proj__4.mux108/_0_  (.A0(net389),
    .A1(net390),
    .S(net162),
    .X(\proj__4.net127 ));
 sg13g2_mux2_1 \proj__4.mux109/_0_  (.A0(net391),
    .A1(net392),
    .S(net162),
    .X(\proj__4.net128 ));
 sg13g2_mux2_1 \proj__4.mux11/_0_  (.A0(\proj__4.net22 ),
    .A1(\proj__4.net23 ),
    .S(net153),
    .X(\proj__4.net29 ));
 sg13g2_mux2_1 \proj__4.mux110/_0_  (.A0(net393),
    .A1(net74),
    .S(net164),
    .X(\proj__4.net129 ));
 sg13g2_mux2_1 \proj__4.mux111/_0_  (.A0(net394),
    .A1(net395),
    .S(net164),
    .X(\proj__4.net130 ));
 sg13g2_mux2_1 \proj__4.mux112/_0_  (.A0(net396),
    .A1(net397),
    .S(net164),
    .X(\proj__4.net131 ));
 sg13g2_mux2_1 \proj__4.mux113/_0_  (.A0(net398),
    .A1(net399),
    .S(net164),
    .X(\proj__4.net132 ));
 sg13g2_mux2_1 \proj__4.mux114/_0_  (.A0(\proj__4.net125 ),
    .A1(\proj__4.net126 ),
    .S(net156),
    .X(\proj__4.net133 ));
 sg13g2_mux2_1 \proj__4.mux115/_0_  (.A0(\proj__4.net127 ),
    .A1(\proj__4.net128 ),
    .S(net156),
    .X(\proj__4.net134 ));
 sg13g2_mux2_1 \proj__4.mux116/_0_  (.A0(\proj__4.net129 ),
    .A1(\proj__4.net130 ),
    .S(net156),
    .X(\proj__4.net135 ));
 sg13g2_mux2_1 \proj__4.mux117/_0_  (.A0(\proj__4.net131 ),
    .A1(\proj__4.net132 ),
    .S(net153),
    .X(\proj__4.net136 ));
 sg13g2_mux2_1 \proj__4.mux118/_0_  (.A0(\proj__4.net135 ),
    .A1(\proj__4.net136 ),
    .S(net151),
    .X(\proj__4.net137 ));
 sg13g2_mux2_1 \proj__4.mux119/_0_  (.A0(\proj__4.net133 ),
    .A1(\proj__4.net134 ),
    .S(net151),
    .X(\proj__4.net138 ));
 sg13g2_mux2_1 \proj__4.mux12/_0_  (.A0(\proj__4.net24 ),
    .A1(\proj__4.net25 ),
    .S(net153),
    .X(\proj__4.net30 ));
 sg13g2_mux2_1 \proj__4.mux120/_0_  (.A0(\proj__4.net138 ),
    .A1(\proj__4.net137 ),
    .S(net149),
    .X(\proj__4.net8 ));
 sg13g2_mux2_1 \proj__4.mux13/_0_  (.A0(\proj__4.net29 ),
    .A1(\proj__4.net30 ),
    .S(net150),
    .X(\proj__4.net32 ));
 sg13g2_mux2_1 \proj__4.mux14/_0_  (.A0(\proj__4.net27 ),
    .A1(\proj__4.net28 ),
    .S(net150),
    .X(\proj__4.net33 ));
 sg13g2_mux2_1 \proj__4.mux15/_0_  (.A0(\proj__4.net33 ),
    .A1(\proj__4.net32 ),
    .S(net149),
    .X(\proj__4.net2 ));
 sg13g2_mux2_1 \proj__4.mux2/_0_  (.A0(net75),
    .A1(net76),
    .S(net163),
    .X(\proj__4.net18 ));
 sg13g2_mux2_1 \proj__4.mux3/_0_  (.A0(net77),
    .A1(net400),
    .S(net163),
    .X(\proj__4.net20 ));
 sg13g2_mux2_1 \proj__4.mux31/_0_  (.A0(net78),
    .A1(net79),
    .S(net160),
    .X(\proj__4.net44 ));
 sg13g2_mux2_1 \proj__4.mux32/_0_  (.A0(net80),
    .A1(net401),
    .S(net160),
    .X(\proj__4.net46 ));
 sg13g2_mux2_1 \proj__4.mux33/_0_  (.A0(net81),
    .A1(net402),
    .S(net159),
    .X(\proj__4.net47 ));
 sg13g2_mux2_1 \proj__4.mux34/_0_  (.A0(net403),
    .A1(net404),
    .S(net159),
    .X(\proj__4.net48 ));
 sg13g2_mux2_1 \proj__4.mux35/_0_  (.A0(net82),
    .A1(net83),
    .S(net160),
    .X(\proj__4.net49 ));
 sg13g2_mux2_1 \proj__4.mux36/_0_  (.A0(net84),
    .A1(net85),
    .S(net160),
    .X(\proj__4.net50 ));
 sg13g2_mux2_1 \proj__4.mux37/_0_  (.A0(net86),
    .A1(net87),
    .S(net159),
    .X(\proj__4.net51 ));
 sg13g2_mux2_1 \proj__4.mux38/_0_  (.A0(net405),
    .A1(net88),
    .S(net159),
    .X(\proj__4.net52 ));
 sg13g2_mux2_1 \proj__4.mux39/_0_  (.A0(\proj__4.net44 ),
    .A1(\proj__4.net46 ),
    .S(net154),
    .X(\proj__4.net53 ));
 sg13g2_mux2_1 \proj__4.mux4/_0_  (.A0(net406),
    .A1(net407),
    .S(net163),
    .X(\proj__4.net21 ));
 sg13g2_mux2_1 \proj__4.mux40/_0_  (.A0(\proj__4.net47 ),
    .A1(\proj__4.net48 ),
    .S(net154),
    .X(\proj__4.net54 ));
 sg13g2_mux2_1 \proj__4.mux41/_0_  (.A0(\proj__4.net49 ),
    .A1(\proj__4.net50 ),
    .S(net154),
    .X(\proj__4.net55 ));
 sg13g2_mux2_1 \proj__4.mux42/_0_  (.A0(\proj__4.net51 ),
    .A1(\proj__4.net52 ),
    .S(net154),
    .X(\proj__4.net56 ));
 sg13g2_mux2_1 \proj__4.mux43/_0_  (.A0(\proj__4.net55 ),
    .A1(\proj__4.net56 ),
    .S(net151),
    .X(\proj__4.net57 ));
 sg13g2_mux2_1 \proj__4.mux44/_0_  (.A0(\proj__4.net53 ),
    .A1(\proj__4.net54 ),
    .S(net151),
    .X(\proj__4.net58 ));
 sg13g2_mux2_1 \proj__4.mux45/_0_  (.A0(\proj__4.net58 ),
    .A1(\proj__4.net57 ),
    .S(net149),
    .X(\proj__4.net3 ));
 sg13g2_mux2_1 \proj__4.mux46/_0_  (.A0(net89),
    .A1(net90),
    .S(net165),
    .X(\proj__4.net60 ));
 sg13g2_mux2_1 \proj__4.mux47/_0_  (.A0(net408),
    .A1(net409),
    .S(net165),
    .X(\proj__4.net62 ));
 sg13g2_mux2_1 \proj__4.mux48/_0_  (.A0(net91),
    .A1(net410),
    .S(net165),
    .X(\proj__4.net63 ));
 sg13g2_mux2_1 \proj__4.mux49/_0_  (.A0(net92),
    .A1(net93),
    .S(net165),
    .X(\proj__4.net64 ));
 sg13g2_mux2_1 \proj__4.mux5/_0_  (.A0(net94),
    .A1(net95),
    .S(net162),
    .X(\proj__4.net22 ));
 sg13g2_mux2_1 \proj__4.mux50/_0_  (.A0(net411),
    .A1(net412),
    .S(net161),
    .X(\proj__4.net65 ));
 sg13g2_mux2_1 \proj__4.mux51/_0_  (.A0(net96),
    .A1(net97),
    .S(net160),
    .X(\proj__4.net66 ));
 sg13g2_mux2_1 \proj__4.mux52/_0_  (.A0(net413),
    .A1(net98),
    .S(net160),
    .X(\proj__4.net67 ));
 sg13g2_mux2_1 \proj__4.mux53/_0_  (.A0(net414),
    .A1(net415),
    .S(net160),
    .X(\proj__4.net68 ));
 sg13g2_mux2_1 \proj__4.mux54/_0_  (.A0(\proj__4.net60 ),
    .A1(\proj__4.net62 ),
    .S(net155),
    .X(\proj__4.net69 ));
 sg13g2_mux2_1 \proj__4.mux55/_0_  (.A0(\proj__4.net63 ),
    .A1(\proj__4.net64 ),
    .S(net155),
    .X(\proj__4.net70 ));
 sg13g2_mux2_1 \proj__4.mux56/_0_  (.A0(\proj__4.net65 ),
    .A1(\proj__4.net66 ),
    .S(net154),
    .X(\proj__4.net71 ));
 sg13g2_mux2_1 \proj__4.mux57/_0_  (.A0(\proj__4.net67 ),
    .A1(\proj__4.net68 ),
    .S(net154),
    .X(\proj__4.net72 ));
 sg13g2_mux2_1 \proj__4.mux58/_0_  (.A0(\proj__4.net71 ),
    .A1(\proj__4.net72 ),
    .S(net151),
    .X(\proj__4.net73 ));
 sg13g2_mux2_1 \proj__4.mux59/_0_  (.A0(\proj__4.net69 ),
    .A1(\proj__4.net70 ),
    .S(net151),
    .X(\proj__4.net74 ));
 sg13g2_mux2_1 \proj__4.mux6/_0_  (.A0(net99),
    .A1(net100),
    .S(net162),
    .X(\proj__4.net23 ));
 sg13g2_mux2_1 \proj__4.mux60/_0_  (.A0(\proj__4.net74 ),
    .A1(\proj__4.net73 ),
    .S(net149),
    .X(\proj__4.net4 ));
 sg13g2_mux2_1 \proj__4.mux61/_0_  (.A0(net416),
    .A1(net101),
    .S(net159),
    .X(\proj__4.net77 ));
 sg13g2_mux2_1 \proj__4.mux62/_0_  (.A0(net102),
    .A1(net417),
    .S(net159),
    .X(\proj__4.net78 ));
 sg13g2_mux2_1 \proj__4.mux63/_0_  (.A0(net418),
    .A1(net419),
    .S(net157),
    .X(\proj__4.net79 ));
 sg13g2_mux2_1 \proj__4.mux64/_0_  (.A0(net103),
    .A1(net420),
    .S(net157),
    .X(\proj__4.net80 ));
 sg13g2_mux2_1 \proj__4.mux65/_0_  (.A0(net421),
    .A1(net422),
    .S(net159),
    .X(\proj__4.net81 ));
 sg13g2_mux2_1 \proj__4.mux66/_0_  (.A0(net423),
    .A1(net104),
    .S(net159),
    .X(\proj__4.net82 ));
 sg13g2_mux2_1 \proj__4.mux67/_0_  (.A0(net424),
    .A1(net425),
    .S(net157),
    .X(\proj__4.net83 ));
 sg13g2_mux2_1 \proj__4.mux68/_0_  (.A0(net105),
    .A1(net426),
    .S(net157),
    .X(\proj__4.net84 ));
 sg13g2_mux2_1 \proj__4.mux69/_0_  (.A0(\proj__4.net77 ),
    .A1(\proj__4.net78 ),
    .S(net153),
    .X(\proj__4.net85 ));
 sg13g2_mux2_1 \proj__4.mux7/_0_  (.A0(net106),
    .A1(net107),
    .S(net162),
    .X(\proj__4.net24 ));
 sg13g2_mux2_1 \proj__4.mux70/_0_  (.A0(\proj__4.net79 ),
    .A1(\proj__4.net80 ),
    .S(net153),
    .X(\proj__4.net86 ));
 sg13g2_mux2_1 \proj__4.mux71/_0_  (.A0(\proj__4.net81 ),
    .A1(\proj__4.net82 ),
    .S(net152),
    .X(\proj__4.net87 ));
 sg13g2_mux2_1 \proj__4.mux72/_0_  (.A0(\proj__4.net83 ),
    .A1(\proj__4.net84 ),
    .S(net152),
    .X(\proj__4.net88 ));
 sg13g2_mux2_1 \proj__4.mux73/_0_  (.A0(\proj__4.net87 ),
    .A1(\proj__4.net88 ),
    .S(net150),
    .X(\proj__4.net89 ));
 sg13g2_mux2_1 \proj__4.mux74/_0_  (.A0(\proj__4.net85 ),
    .A1(\proj__4.net86 ),
    .S(net150),
    .X(\proj__4.net90 ));
 sg13g2_mux2_1 \proj__4.mux75/_0_  (.A0(\proj__4.net90 ),
    .A1(\proj__4.net89 ),
    .S(net149),
    .X(\proj__4.net5 ));
 sg13g2_mux2_1 \proj__4.mux76/_0_  (.A0(net427),
    .A1(net428),
    .S(net157),
    .X(\proj__4.net92 ));
 sg13g2_mux2_1 \proj__4.mux77/_0_  (.A0(net429),
    .A1(net108),
    .S(net157),
    .X(\proj__4.net94 ));
 sg13g2_mux2_1 \proj__4.mux78/_0_  (.A0(net430),
    .A1(net431),
    .S(net158),
    .X(\proj__4.net95 ));
 sg13g2_mux2_1 \proj__4.mux79/_0_  (.A0(net432),
    .A1(net433),
    .S(net158),
    .X(\proj__4.net96 ));
 sg13g2_mux2_1 \proj__4.mux8/_0_  (.A0(net109),
    .A1(net434),
    .S(net162),
    .X(\proj__4.net25 ));
 sg13g2_mux2_1 \proj__4.mux80/_0_  (.A0(net435),
    .A1(net436),
    .S(net158),
    .X(\proj__4.net97 ));
 sg13g2_mux2_1 \proj__4.mux81/_0_  (.A0(net437),
    .A1(net438),
    .S(net158),
    .X(\proj__4.net98 ));
 sg13g2_mux2_1 \proj__4.mux82/_0_  (.A0(net439),
    .A1(net440),
    .S(net158),
    .X(\proj__4.net99 ));
 sg13g2_mux2_1 \proj__4.mux83/_0_  (.A0(net441),
    .A1(net110),
    .S(net158),
    .X(\proj__4.net100 ));
 sg13g2_mux2_1 \proj__4.mux84/_0_  (.A0(\proj__4.net92 ),
    .A1(\proj__4.net94 ),
    .S(net152),
    .X(\proj__4.net101 ));
 sg13g2_mux2_1 \proj__4.mux85/_0_  (.A0(\proj__4.net95 ),
    .A1(\proj__4.net96 ),
    .S(net152),
    .X(\proj__4.net102 ));
 sg13g2_mux2_1 \proj__4.mux86/_0_  (.A0(\proj__4.net97 ),
    .A1(\proj__4.net98 ),
    .S(net152),
    .X(\proj__4.net103 ));
 sg13g2_mux2_1 \proj__4.mux87/_0_  (.A0(\proj__4.net99 ),
    .A1(\proj__4.net100 ),
    .S(net152),
    .X(\proj__4.net104 ));
 sg13g2_mux2_1 \proj__4.mux88/_0_  (.A0(\proj__4.net103 ),
    .A1(\proj__4.net104 ),
    .S(net150),
    .X(\proj__4.net105 ));
 sg13g2_mux2_1 \proj__4.mux89/_0_  (.A0(\proj__4.net101 ),
    .A1(\proj__4.net102 ),
    .S(net150),
    .X(\proj__4.net106 ));
 sg13g2_mux2_1 \proj__4.mux9/_0_  (.A0(\proj__4.net17 ),
    .A1(\proj__4.net18 ),
    .S(net153),
    .X(\proj__4.net27 ));
 sg13g2_mux2_1 \proj__4.mux90/_0_  (.A0(\proj__4.net106 ),
    .A1(\proj__4.net105 ),
    .S(net149),
    .X(\proj__4.net6 ));
 sg13g2_mux2_1 \proj__4.mux91/_0_  (.A0(net442),
    .A1(net111),
    .S(net165),
    .X(\proj__4.net109 ));
 sg13g2_mux2_1 \proj__4.mux92/_0_  (.A0(net112),
    .A1(net443),
    .S(net165),
    .X(\proj__4.net110 ));
 sg13g2_mux2_1 \proj__4.mux93/_0_  (.A0(net444),
    .A1(net113),
    .S(net165),
    .X(\proj__4.net111 ));
 sg13g2_mux2_1 \proj__4.mux94/_0_  (.A0(net445),
    .A1(net446),
    .S(net165),
    .X(\proj__4.net112 ));
 sg13g2_mux2_1 \proj__4.mux95/_0_  (.A0(net114),
    .A1(net115),
    .S(net166),
    .X(\proj__4.net113 ));
 sg13g2_mux2_1 \proj__4.mux96/_0_  (.A0(net447),
    .A1(net116),
    .S(net166),
    .X(\proj__4.net114 ));
 sg13g2_mux2_1 \proj__4.mux97/_0_  (.A0(net117),
    .A1(net118),
    .S(net166),
    .X(\proj__4.net115 ));
 sg13g2_mux2_1 \proj__4.mux98/_0_  (.A0(net448),
    .A1(net449),
    .S(net166),
    .X(\proj__4.net116 ));
 sg13g2_mux2_1 \proj__4.mux99/_0_  (.A0(\proj__4.net109 ),
    .A1(\proj__4.net110 ),
    .S(net154),
    .X(\proj__4.net117 ));
 sg13g2_xor2_1 \proj__4.xor1/_0_  (.B(net157),
    .A(net450),
    .X(\proj__4.net35 ));
 sg13g2_xor2_1 \proj__4.xor2/_0_  (.B(net152),
    .A(\proj__4.net40 ),
    .X(\proj__4.net36 ));
 sg13g2_xor2_1 \proj__4.xor3/_0_  (.B(net150),
    .A(\proj__4.net41 ),
    .X(\proj__4.net37 ));
 sg13g2_xor2_1 \proj__4.xor4/_0_  (.B(net149),
    .A(\proj__4.net42 ),
    .X(\proj__4.net38 ));
 sg13g2_and2_1 \proj__5.and1/_0_  (.A(net144),
    .B(net1),
    .X(\proj__5.net12 ));
 sg13g2_and2_1 \proj__5.and2/_0_  (.A(net3),
    .B(net142),
    .X(\proj__5.net13 ));
 sg13g2_and2_1 \proj__5.and3/_0_  (.A(net131),
    .B(\proj__5.net13 ),
    .X(\proj__5.net14 ));
 sg13g2_and2_1 \proj__5.and4/_0_  (.A(\proj__5.net14 ),
    .B(\proj__5.net12 ),
    .X(\proj__5.net6 ));
 sg13g2_and2_1 \proj__6.and1/_0_  (.A(\proj__6.net61 ),
    .B(\proj__6.net62 ),
    .X(\proj__6.net63 ));
 sg13g2_and2_2 \proj__6.and10/_0_  (.A(\proj__6.net64 ),
    .B(net139),
    .X(\proj__6.net32 ));
 sg13g2_and2_2 \proj__6.and11/_0_  (.A(\proj__6.net65 ),
    .B(net139),
    .X(\proj__6.net42 ));
 sg13g2_and2_2 \proj__6.and12/_0_  (.A(\proj__6.net66 ),
    .B(net139),
    .X(\proj__6.net52 ));
 sg13g2_and2_1 \proj__6.and13/_0_  (.A(net129),
    .B(\proj__6.net74 ),
    .X(\proj__6.net10 ));
 sg13g2_and2_1 \proj__6.and14/_0_  (.A(net129),
    .B(\proj__6.net76 ),
    .X(\proj__6.net11 ));
 sg13g2_and2_1 \proj__6.and15/_0_  (.A(net129),
    .B(\proj__6.net78 ),
    .X(\proj__6.net12 ));
 sg13g2_and2_1 \proj__6.and16/_0_  (.A(net129),
    .B(\proj__6.net80 ),
    .X(\proj__6.net13 ));
 sg13g2_and2_1 \proj__6.and17/_0_  (.A(net130),
    .B(\proj__6.net82 ),
    .X(\proj__6.net14 ));
 sg13g2_and2_1 \proj__6.and18/_0_  (.A(net130),
    .B(\proj__6.net84 ),
    .X(\proj__6.net15 ));
 sg13g2_and2_1 \proj__6.and19/_0_  (.A(net130),
    .B(\proj__6.net86 ),
    .X(\proj__6.net16 ));
 sg13g2_and2_1 \proj__6.and2/_0_  (.A(net148),
    .B(net146),
    .X(\proj__6.net66 ));
 sg13g2_and2_1 \proj__6.and20/_0_  (.A(net130),
    .B(\proj__6.net88 ),
    .X(\proj__6.net17 ));
 sg13g2_and2_1 \proj__6.and3/_0_  (.A(net140),
    .B(\proj__6.net63 ),
    .X(\proj__6.net20 ));
 sg13g2_and2_1 \proj__6.and4/_0_  (.A(net147),
    .B(\proj__6.net62 ),
    .X(\proj__6.net64 ));
 sg13g2_and2_1 \proj__6.and5/_0_  (.A(net142),
    .B(\proj__6.net66 ),
    .X(\proj__6.net51 ));
 sg13g2_and2_1 \proj__6.and6/_0_  (.A(net140),
    .B(\proj__6.net64 ),
    .X(\proj__6.net31 ));
 sg13g2_and2_1 \proj__6.and7/_0_  (.A(\proj__6.net61 ),
    .B(net145),
    .X(\proj__6.net65 ));
 sg13g2_and2_2 \proj__6.and8/_0_  (.A(\proj__6.net63 ),
    .B(net139),
    .X(\proj__6.net21 ));
 sg13g2_and2_1 \proj__6.and9/_0_  (.A(net140),
    .B(\proj__6.net65 ),
    .X(\proj__6.net41 ));
 sg13g2_inv_1 \proj__6.flop0/_4_  (.Y(\proj__6.flop0/_0_ ),
    .A(net119));
 sg13g2_inv_1 \proj__6.flop0/_5_  (.Y(\proj__6.flop0/_1_ ),
    .A(net120));
 sg13g2_tielo \proj__6.flop0/dffsr_257  (.L_LO(net298));
 sg13g2_tielo \proj__6.flop1/dffsr_258  (.L_LO(net299));
 sg13g2_sdfbbp_1 \proj__6.flop0/dffsr  (.Q(\proj__6.net23 ),
    .Q_N(\proj__6.flop0/notq ),
    .RESET_B(\proj__6.flop0/_0_ ),
    .SET_B(\proj__6.flop0/_1_ ),
    .D(\proj__6.net20 ),
    .SCE(net298),
    .SCD(net297),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop1/_4_  (.Y(\proj__6.flop1/_0_ ),
    .A(net121));
 sg13g2_inv_1 \proj__6.flop1/_5_  (.Y(\proj__6.flop1/_1_ ),
    .A(net122));
 sg13g2_tielo \proj__6.flop1/dffsr_259  (.L_LO(net300));
 sg13g2_tielo \proj__6.flop10/dffsr_260  (.L_LO(net301));
 sg13g2_sdfbbp_1 \proj__6.flop1/dffsr  (.Q(\proj__6.net24 ),
    .Q_N(\proj__6.flop1/notq ),
    .RESET_B(\proj__6.flop1/_0_ ),
    .SET_B(\proj__6.flop1/_1_ ),
    .D(\proj__6.net23 ),
    .SCE(net300),
    .SCD(net299),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop10/_4_  (.Y(\proj__6.flop10/_0_ ),
    .A(net123));
 sg13g2_inv_1 \proj__6.flop10/_5_  (.Y(\proj__6.flop10/_1_ ),
    .A(net124));
 sg13g2_tielo \proj__6.flop10/dffsr_261  (.L_LO(net302));
 sg13g2_tielo \proj__6.flop11/dffsr_262  (.L_LO(net303));
 sg13g2_sdfbbp_1 \proj__6.flop10/dffsr  (.Q(\proj__6.net36 ),
    .Q_N(\proj__6.flop10/notq ),
    .RESET_B(\proj__6.flop10/_0_ ),
    .SET_B(\proj__6.flop10/_1_ ),
    .D(\proj__6.net35 ),
    .SCE(net302),
    .SCD(net301),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop11/_4_  (.Y(\proj__6.flop11/_0_ ),
    .A(net125));
 sg13g2_inv_1 \proj__6.flop11/_5_  (.Y(\proj__6.flop11/_1_ ),
    .A(net126));
 sg13g2_tielo \proj__6.flop11/dffsr_263  (.L_LO(net304));
 sg13g2_tielo \proj__6.flop12/dffsr_264  (.L_LO(net305));
 sg13g2_sdfbbp_1 \proj__6.flop11/dffsr  (.Q(\proj__6.net35 ),
    .Q_N(\proj__6.flop11/notq ),
    .RESET_B(\proj__6.flop11/_0_ ),
    .SET_B(\proj__6.flop11/_1_ ),
    .D(\proj__6.net37 ),
    .SCE(net304),
    .SCD(net303),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop12/_4_  (.Y(\proj__6.flop12/_0_ ),
    .A(net168));
 sg13g2_inv_1 \proj__6.flop12/_5_  (.Y(\proj__6.flop12/_1_ ),
    .A(net169));
 sg13g2_tielo \proj__6.flop12/dffsr_265  (.L_LO(net306));
 sg13g2_tielo \proj__6.flop13/dffsr_266  (.L_LO(net307));
 sg13g2_sdfbbp_1 \proj__6.flop12/dffsr  (.Q(\proj__6.net38 ),
    .Q_N(\proj__6.flop12/notq ),
    .RESET_B(\proj__6.flop12/_0_ ),
    .SET_B(\proj__6.flop12/_1_ ),
    .D(\proj__6.net34 ),
    .SCE(net306),
    .SCD(net305),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop13/_4_  (.Y(\proj__6.flop13/_0_ ),
    .A(net170));
 sg13g2_inv_1 \proj__6.flop13/_5_  (.Y(\proj__6.flop13/_1_ ),
    .A(net171));
 sg13g2_tielo \proj__6.flop13/dffsr_267  (.L_LO(net308));
 sg13g2_tielo \proj__6.flop14/dffsr_268  (.L_LO(net309));
 sg13g2_sdfbbp_1 \proj__6.flop13/dffsr  (.Q(\proj__6.net39 ),
    .Q_N(\proj__6.flop13/notq ),
    .RESET_B(\proj__6.flop13/_0_ ),
    .SET_B(\proj__6.flop13/_1_ ),
    .D(\proj__6.net38 ),
    .SCE(net308),
    .SCD(net307),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop14/_4_  (.Y(\proj__6.flop14/_0_ ),
    .A(net172));
 sg13g2_inv_1 \proj__6.flop14/_5_  (.Y(\proj__6.flop14/_1_ ),
    .A(net173));
 sg13g2_tielo \proj__6.flop14/dffsr_269  (.L_LO(net310));
 sg13g2_tielo \proj__6.flop15/dffsr_270  (.L_LO(net311));
 sg13g2_sdfbbp_1 \proj__6.flop14/dffsr  (.Q(\proj__6.net40 ),
    .Q_N(\proj__6.flop14/notq ),
    .RESET_B(\proj__6.flop14/_0_ ),
    .SET_B(\proj__6.flop14/_1_ ),
    .D(\proj__6.net39 ),
    .SCE(net310),
    .SCD(net309),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop15/_4_  (.Y(\proj__6.flop15/_0_ ),
    .A(net174));
 sg13g2_inv_1 \proj__6.flop15/_5_  (.Y(\proj__6.flop15/_1_ ),
    .A(net175));
 sg13g2_tielo \proj__6.flop15/dffsr_271  (.L_LO(net312));
 sg13g2_tielo \proj__6.flop16/dffsr_272  (.L_LO(net313));
 sg13g2_sdfbbp_1 \proj__6.flop15/dffsr  (.Q(\proj__6.net37 ),
    .Q_N(\proj__6.flop15/notq ),
    .RESET_B(\proj__6.flop15/_0_ ),
    .SET_B(\proj__6.flop15/_1_ ),
    .D(\proj__6.net40 ),
    .SCE(net312),
    .SCD(net311),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop16/_4_  (.Y(\proj__6.flop16/_0_ ),
    .A(net176));
 sg13g2_inv_1 \proj__6.flop16/_5_  (.Y(\proj__6.flop16/_1_ ),
    .A(net177));
 sg13g2_tielo \proj__6.flop16/dffsr_273  (.L_LO(net314));
 sg13g2_tielo \proj__6.flop17/dffsr_274  (.L_LO(net315));
 sg13g2_sdfbbp_1 \proj__6.flop16/dffsr  (.Q(\proj__6.net43 ),
    .Q_N(\proj__6.flop16/notq ),
    .RESET_B(\proj__6.flop16/_0_ ),
    .SET_B(\proj__6.flop16/_1_ ),
    .D(\proj__6.net41 ),
    .SCE(net314),
    .SCD(net313),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop17/_4_  (.Y(\proj__6.flop17/_0_ ),
    .A(net178));
 sg13g2_inv_1 \proj__6.flop17/_5_  (.Y(\proj__6.flop17/_1_ ),
    .A(net179));
 sg13g2_tielo \proj__6.flop17/dffsr_275  (.L_LO(net316));
 sg13g2_tielo \proj__6.flop18/dffsr_276  (.L_LO(net317));
 sg13g2_sdfbbp_1 \proj__6.flop17/dffsr  (.Q(\proj__6.net44 ),
    .Q_N(\proj__6.flop17/notq ),
    .RESET_B(\proj__6.flop17/_0_ ),
    .SET_B(\proj__6.flop17/_1_ ),
    .D(\proj__6.net43 ),
    .SCE(net316),
    .SCD(net315),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop18/_4_  (.Y(\proj__6.flop18/_0_ ),
    .A(net180));
 sg13g2_inv_1 \proj__6.flop18/_5_  (.Y(\proj__6.flop18/_1_ ),
    .A(net181));
 sg13g2_tielo \proj__6.flop18/dffsr_277  (.L_LO(net318));
 sg13g2_tielo \proj__6.flop19/dffsr_278  (.L_LO(net319));
 sg13g2_sdfbbp_1 \proj__6.flop18/dffsr  (.Q(\proj__6.net46 ),
    .Q_N(\proj__6.flop18/notq ),
    .RESET_B(\proj__6.flop18/_0_ ),
    .SET_B(\proj__6.flop18/_1_ ),
    .D(\proj__6.net45 ),
    .SCE(net318),
    .SCD(net317),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop19/_4_  (.Y(\proj__6.flop19/_0_ ),
    .A(net182));
 sg13g2_inv_1 \proj__6.flop19/_5_  (.Y(\proj__6.flop19/_1_ ),
    .A(net183));
 sg13g2_tielo \proj__6.flop19/dffsr_279  (.L_LO(net320));
 sg13g2_tielo \proj__6.flop2/dffsr_280  (.L_LO(net321));
 sg13g2_sdfbbp_1 \proj__6.flop19/dffsr  (.Q(\proj__6.net45 ),
    .Q_N(\proj__6.flop19/notq ),
    .RESET_B(\proj__6.flop19/_0_ ),
    .SET_B(\proj__6.flop19/_1_ ),
    .D(\proj__6.net47 ),
    .SCE(net320),
    .SCD(net319),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop2/_4_  (.Y(\proj__6.flop2/_0_ ),
    .A(net184));
 sg13g2_inv_1 \proj__6.flop2/_5_  (.Y(\proj__6.flop2/_1_ ),
    .A(net185));
 sg13g2_tielo \proj__6.flop2/dffsr_281  (.L_LO(net322));
 sg13g2_tielo \proj__6.flop20/dffsr_282  (.L_LO(net323));
 sg13g2_sdfbbp_1 \proj__6.flop2/dffsr  (.Q(\proj__6.net26 ),
    .Q_N(\proj__6.flop2/notq ),
    .RESET_B(\proj__6.flop2/_0_ ),
    .SET_B(\proj__6.flop2/_1_ ),
    .D(\proj__6.net25 ),
    .SCE(net322),
    .SCD(net321),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop20/_4_  (.Y(\proj__6.flop20/_0_ ),
    .A(net186));
 sg13g2_inv_1 \proj__6.flop20/_5_  (.Y(\proj__6.flop20/_1_ ),
    .A(net187));
 sg13g2_tielo \proj__6.flop20/dffsr_283  (.L_LO(net324));
 sg13g2_tielo \proj__6.flop21/dffsr_284  (.L_LO(net325));
 sg13g2_sdfbbp_1 \proj__6.flop20/dffsr  (.Q(\proj__6.net48 ),
    .Q_N(\proj__6.flop20/notq ),
    .RESET_B(\proj__6.flop20/_0_ ),
    .SET_B(\proj__6.flop20/_1_ ),
    .D(\proj__6.net44 ),
    .SCE(net324),
    .SCD(net323),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop21/_4_  (.Y(\proj__6.flop21/_0_ ),
    .A(net188));
 sg13g2_inv_1 \proj__6.flop21/_5_  (.Y(\proj__6.flop21/_1_ ),
    .A(net189));
 sg13g2_tielo \proj__6.flop21/dffsr_285  (.L_LO(net326));
 sg13g2_tielo \proj__6.flop22/dffsr_286  (.L_LO(net327));
 sg13g2_sdfbbp_1 \proj__6.flop21/dffsr  (.Q(\proj__6.net49 ),
    .Q_N(\proj__6.flop21/notq ),
    .RESET_B(\proj__6.flop21/_0_ ),
    .SET_B(\proj__6.flop21/_1_ ),
    .D(\proj__6.net48 ),
    .SCE(net326),
    .SCD(net325),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop22/_4_  (.Y(\proj__6.flop22/_0_ ),
    .A(net190));
 sg13g2_inv_1 \proj__6.flop22/_5_  (.Y(\proj__6.flop22/_1_ ),
    .A(net191));
 sg13g2_tielo \proj__6.flop22/dffsr_287  (.L_LO(net328));
 sg13g2_tielo \proj__6.flop23/dffsr_288  (.L_LO(net329));
 sg13g2_sdfbbp_1 \proj__6.flop22/dffsr  (.Q(\proj__6.net50 ),
    .Q_N(\proj__6.flop22/notq ),
    .RESET_B(\proj__6.flop22/_0_ ),
    .SET_B(\proj__6.flop22/_1_ ),
    .D(\proj__6.net49 ),
    .SCE(net328),
    .SCD(net327),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop23/_4_  (.Y(\proj__6.flop23/_0_ ),
    .A(net192));
 sg13g2_inv_1 \proj__6.flop23/_5_  (.Y(\proj__6.flop23/_1_ ),
    .A(net193));
 sg13g2_tielo \proj__6.flop23/dffsr_289  (.L_LO(net330));
 sg13g2_tielo \proj__6.flop24/dffsr_290  (.L_LO(net331));
 sg13g2_sdfbbp_1 \proj__6.flop23/dffsr  (.Q(\proj__6.net47 ),
    .Q_N(\proj__6.flop23/notq ),
    .RESET_B(\proj__6.flop23/_0_ ),
    .SET_B(\proj__6.flop23/_1_ ),
    .D(\proj__6.net50 ),
    .SCE(net330),
    .SCD(net329),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop24/_4_  (.Y(\proj__6.flop24/_0_ ),
    .A(net194));
 sg13g2_inv_1 \proj__6.flop24/_5_  (.Y(\proj__6.flop24/_1_ ),
    .A(net195));
 sg13g2_tielo \proj__6.flop24/dffsr_291  (.L_LO(net332));
 sg13g2_tielo \proj__6.flop25/dffsr_292  (.L_LO(net333));
 sg13g2_sdfbbp_1 \proj__6.flop24/dffsr  (.Q(\proj__6.net53 ),
    .Q_N(\proj__6.flop24/notq ),
    .RESET_B(\proj__6.flop24/_0_ ),
    .SET_B(\proj__6.flop24/_1_ ),
    .D(\proj__6.net51 ),
    .SCE(net332),
    .SCD(net331),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop25/_4_  (.Y(\proj__6.flop25/_0_ ),
    .A(net196));
 sg13g2_inv_1 \proj__6.flop25/_5_  (.Y(\proj__6.flop25/_1_ ),
    .A(net197));
 sg13g2_tielo \proj__6.flop25/dffsr_293  (.L_LO(net334));
 sg13g2_tielo \proj__6.flop26/dffsr_294  (.L_LO(net335));
 sg13g2_sdfbbp_1 \proj__6.flop25/dffsr  (.Q(\proj__6.net54 ),
    .Q_N(\proj__6.flop25/notq ),
    .RESET_B(\proj__6.flop25/_0_ ),
    .SET_B(\proj__6.flop25/_1_ ),
    .D(\proj__6.net53 ),
    .SCE(net334),
    .SCD(net333),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop26/_4_  (.Y(\proj__6.flop26/_0_ ),
    .A(net198));
 sg13g2_inv_1 \proj__6.flop26/_5_  (.Y(\proj__6.flop26/_1_ ),
    .A(net199));
 sg13g2_tielo \proj__6.flop26/dffsr_295  (.L_LO(net336));
 sg13g2_tielo \proj__6.flop27/dffsr_296  (.L_LO(net337));
 sg13g2_sdfbbp_1 \proj__6.flop26/dffsr  (.Q(\proj__6.net56 ),
    .Q_N(\proj__6.flop26/notq ),
    .RESET_B(\proj__6.flop26/_0_ ),
    .SET_B(\proj__6.flop26/_1_ ),
    .D(\proj__6.net55 ),
    .SCE(net336),
    .SCD(net335),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop27/_4_  (.Y(\proj__6.flop27/_0_ ),
    .A(net200));
 sg13g2_inv_1 \proj__6.flop27/_5_  (.Y(\proj__6.flop27/_1_ ),
    .A(net201));
 sg13g2_tielo \proj__6.flop27/dffsr_297  (.L_LO(net338));
 sg13g2_tielo \proj__6.flop28/dffsr_298  (.L_LO(net339));
 sg13g2_sdfbbp_1 \proj__6.flop27/dffsr  (.Q(\proj__6.net55 ),
    .Q_N(\proj__6.flop27/notq ),
    .RESET_B(\proj__6.flop27/_0_ ),
    .SET_B(\proj__6.flop27/_1_ ),
    .D(\proj__6.net57 ),
    .SCE(net338),
    .SCD(net337),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop28/_4_  (.Y(\proj__6.flop28/_0_ ),
    .A(net202));
 sg13g2_inv_1 \proj__6.flop28/_5_  (.Y(\proj__6.flop28/_1_ ),
    .A(net203));
 sg13g2_tielo \proj__6.flop28/dffsr_299  (.L_LO(net340));
 sg13g2_tielo \proj__6.flop29/dffsr_300  (.L_LO(net341));
 sg13g2_sdfbbp_1 \proj__6.flop28/dffsr  (.Q(\proj__6.net58 ),
    .Q_N(\proj__6.flop28/notq ),
    .RESET_B(\proj__6.flop28/_0_ ),
    .SET_B(\proj__6.flop28/_1_ ),
    .D(\proj__6.net54 ),
    .SCE(net340),
    .SCD(net339),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop29/_4_  (.Y(\proj__6.flop29/_0_ ),
    .A(net204));
 sg13g2_inv_1 \proj__6.flop29/_5_  (.Y(\proj__6.flop29/_1_ ),
    .A(net205));
 sg13g2_tielo \proj__6.flop29/dffsr_301  (.L_LO(net342));
 sg13g2_tielo \proj__6.flop3/dffsr_302  (.L_LO(net343));
 sg13g2_sdfbbp_1 \proj__6.flop29/dffsr  (.Q(\proj__6.net59 ),
    .Q_N(\proj__6.flop29/notq ),
    .RESET_B(\proj__6.flop29/_0_ ),
    .SET_B(\proj__6.flop29/_1_ ),
    .D(\proj__6.net58 ),
    .SCE(net342),
    .SCD(net341),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop3/_4_  (.Y(\proj__6.flop3/_0_ ),
    .A(net206));
 sg13g2_inv_1 \proj__6.flop3/_5_  (.Y(\proj__6.flop3/_1_ ),
    .A(net207));
 sg13g2_tielo \proj__6.flop3/dffsr_303  (.L_LO(net344));
 sg13g2_tielo \proj__6.flop30/dffsr_304  (.L_LO(net345));
 sg13g2_sdfbbp_1 \proj__6.flop3/dffsr  (.Q(\proj__6.net25 ),
    .Q_N(\proj__6.flop3/notq ),
    .RESET_B(\proj__6.flop3/_0_ ),
    .SET_B(\proj__6.flop3/_1_ ),
    .D(\proj__6.net27 ),
    .SCE(net344),
    .SCD(net343),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop30/_4_  (.Y(\proj__6.flop30/_0_ ),
    .A(net208));
 sg13g2_inv_1 \proj__6.flop30/_5_  (.Y(\proj__6.flop30/_1_ ),
    .A(net209));
 sg13g2_tielo \proj__6.flop30/dffsr_305  (.L_LO(net346));
 sg13g2_tielo \proj__6.flop31/dffsr_306  (.L_LO(net347));
 sg13g2_sdfbbp_1 \proj__6.flop30/dffsr  (.Q(\proj__6.net60 ),
    .Q_N(\proj__6.flop30/notq ),
    .RESET_B(\proj__6.flop30/_0_ ),
    .SET_B(\proj__6.flop30/_1_ ),
    .D(\proj__6.net59 ),
    .SCE(net346),
    .SCD(net345),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop31/_4_  (.Y(\proj__6.flop31/_0_ ),
    .A(net210));
 sg13g2_inv_1 \proj__6.flop31/_5_  (.Y(\proj__6.flop31/_1_ ),
    .A(net211));
 sg13g2_tielo \proj__6.flop31/dffsr_307  (.L_LO(net348));
 sg13g2_tielo \proj__6.flop33/dffsr_308  (.L_LO(net349));
 sg13g2_sdfbbp_1 \proj__6.flop31/dffsr  (.Q(\proj__6.net57 ),
    .Q_N(\proj__6.flop31/notq ),
    .RESET_B(\proj__6.flop31/_0_ ),
    .SET_B(\proj__6.flop31/_1_ ),
    .D(\proj__6.net60 ),
    .SCE(net348),
    .SCD(net347),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop33/_4_  (.Y(\proj__6.flop33/_0_ ),
    .A(net212));
 sg13g2_inv_1 \proj__6.flop33/_5_  (.Y(\proj__6.flop33/_1_ ),
    .A(net213));
 sg13g2_tielo \proj__6.flop33/dffsr_309  (.L_LO(net350));
 sg13g2_tielo \proj__6.flop34/dffsr_310  (.L_LO(net351));
 sg13g2_sdfbbp_1 \proj__6.flop33/dffsr  (.Q(\proj__6.net74 ),
    .Q_N(\proj__6.flop33/notq ),
    .RESET_B(\proj__6.flop33/_0_ ),
    .SET_B(\proj__6.flop33/_1_ ),
    .D(\proj__6.net72 ),
    .SCE(net350),
    .SCD(net349),
    .CLK(net135));
 sg13g2_inv_1 \proj__6.flop34/_4_  (.Y(\proj__6.flop34/_0_ ),
    .A(net214));
 sg13g2_inv_1 \proj__6.flop34/_5_  (.Y(\proj__6.flop34/_1_ ),
    .A(net215));
 sg13g2_tielo \proj__6.flop34/dffsr_311  (.L_LO(net352));
 sg13g2_tielo \proj__6.flop35/dffsr_312  (.L_LO(net353));
 sg13g2_sdfbbp_1 \proj__6.flop34/dffsr  (.Q(\proj__6.net76 ),
    .Q_N(\proj__6.flop34/notq ),
    .RESET_B(\proj__6.flop34/_0_ ),
    .SET_B(\proj__6.flop34/_1_ ),
    .D(\proj__6.net75 ),
    .SCE(net352),
    .SCD(net351),
    .CLK(net135));
 sg13g2_inv_1 \proj__6.flop35/_4_  (.Y(\proj__6.flop35/_0_ ),
    .A(net216));
 sg13g2_inv_1 \proj__6.flop35/_5_  (.Y(\proj__6.flop35/_1_ ),
    .A(net217));
 sg13g2_tielo \proj__6.flop35/dffsr_313  (.L_LO(net354));
 sg13g2_tielo \proj__6.flop36/dffsr_314  (.L_LO(net355));
 sg13g2_sdfbbp_1 \proj__6.flop35/dffsr  (.Q(\proj__6.net78 ),
    .Q_N(\proj__6.flop35/notq ),
    .RESET_B(\proj__6.flop35/_0_ ),
    .SET_B(\proj__6.flop35/_1_ ),
    .D(\proj__6.net77 ),
    .SCE(net354),
    .SCD(net353),
    .CLK(net135));
 sg13g2_inv_1 \proj__6.flop36/_4_  (.Y(\proj__6.flop36/_0_ ),
    .A(net218));
 sg13g2_inv_1 \proj__6.flop36/_5_  (.Y(\proj__6.flop36/_1_ ),
    .A(net219));
 sg13g2_tielo \proj__6.flop36/dffsr_315  (.L_LO(net356));
 sg13g2_tielo \proj__6.flop37/dffsr_316  (.L_LO(net357));
 sg13g2_sdfbbp_1 \proj__6.flop36/dffsr  (.Q(\proj__6.net80 ),
    .Q_N(\proj__6.flop36/notq ),
    .RESET_B(\proj__6.flop36/_0_ ),
    .SET_B(\proj__6.flop36/_1_ ),
    .D(\proj__6.net79 ),
    .SCE(net356),
    .SCD(net355),
    .CLK(net135));
 sg13g2_inv_1 \proj__6.flop37/_4_  (.Y(\proj__6.flop37/_0_ ),
    .A(net220));
 sg13g2_inv_1 \proj__6.flop37/_5_  (.Y(\proj__6.flop37/_1_ ),
    .A(net221));
 sg13g2_tielo \proj__6.flop37/dffsr_317  (.L_LO(net358));
 sg13g2_tielo \proj__6.flop38/dffsr_318  (.L_LO(net359));
 sg13g2_sdfbbp_1 \proj__6.flop37/dffsr  (.Q(\proj__6.net82 ),
    .Q_N(\proj__6.flop37/notq ),
    .RESET_B(\proj__6.flop37/_0_ ),
    .SET_B(\proj__6.flop37/_1_ ),
    .D(\proj__6.net81 ),
    .SCE(net358),
    .SCD(net357),
    .CLK(net136));
 sg13g2_inv_1 \proj__6.flop38/_4_  (.Y(\proj__6.flop38/_0_ ),
    .A(net222));
 sg13g2_inv_1 \proj__6.flop38/_5_  (.Y(\proj__6.flop38/_1_ ),
    .A(net223));
 sg13g2_tielo \proj__6.flop38/dffsr_319  (.L_LO(net360));
 sg13g2_tielo \proj__6.flop39/dffsr_320  (.L_LO(net361));
 sg13g2_sdfbbp_1 \proj__6.flop38/dffsr  (.Q(\proj__6.net84 ),
    .Q_N(\proj__6.flop38/notq ),
    .RESET_B(\proj__6.flop38/_0_ ),
    .SET_B(\proj__6.flop38/_1_ ),
    .D(\proj__6.net83 ),
    .SCE(net360),
    .SCD(net359),
    .CLK(net135));
 sg13g2_inv_1 \proj__6.flop39/_4_  (.Y(\proj__6.flop39/_0_ ),
    .A(net224));
 sg13g2_inv_1 \proj__6.flop39/_5_  (.Y(\proj__6.flop39/_1_ ),
    .A(net225));
 sg13g2_tielo \proj__6.flop39/dffsr_321  (.L_LO(net362));
 sg13g2_tielo \proj__6.flop4/dffsr_322  (.L_LO(net363));
 sg13g2_sdfbbp_1 \proj__6.flop39/dffsr  (.Q(\proj__6.net86 ),
    .Q_N(\proj__6.flop39/notq ),
    .RESET_B(\proj__6.flop39/_0_ ),
    .SET_B(\proj__6.flop39/_1_ ),
    .D(\proj__6.net85 ),
    .SCE(net362),
    .SCD(net361),
    .CLK(net135));
 sg13g2_inv_1 \proj__6.flop4/_4_  (.Y(\proj__6.flop4/_0_ ),
    .A(net226));
 sg13g2_inv_1 \proj__6.flop4/_5_  (.Y(\proj__6.flop4/_1_ ),
    .A(net227));
 sg13g2_tielo \proj__6.flop4/dffsr_323  (.L_LO(net364));
 sg13g2_tielo \proj__6.flop40/dffsr_324  (.L_LO(net365));
 sg13g2_sdfbbp_1 \proj__6.flop4/dffsr  (.Q(\proj__6.net28 ),
    .Q_N(\proj__6.flop4/notq ),
    .RESET_B(\proj__6.flop4/_0_ ),
    .SET_B(\proj__6.flop4/_1_ ),
    .D(\proj__6.net24 ),
    .SCE(net364),
    .SCD(net363),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop40/_4_  (.Y(\proj__6.flop40/_0_ ),
    .A(net228));
 sg13g2_inv_1 \proj__6.flop40/_5_  (.Y(\proj__6.flop40/_1_ ),
    .A(net229));
 sg13g2_tielo \proj__6.flop40/dffsr_325  (.L_LO(net366));
 sg13g2_tielo \proj__6.flop5/dffsr_326  (.L_LO(net367));
 sg13g2_sdfbbp_1 \proj__6.flop40/dffsr  (.Q(\proj__6.net88 ),
    .Q_N(\proj__6.flop40/notq ),
    .RESET_B(\proj__6.flop40/_0_ ),
    .SET_B(\proj__6.flop40/_1_ ),
    .D(\proj__6.net87 ),
    .SCE(net366),
    .SCD(net365),
    .CLK(net137));
 sg13g2_inv_1 \proj__6.flop5/_4_  (.Y(\proj__6.flop5/_0_ ),
    .A(net230));
 sg13g2_inv_1 \proj__6.flop5/_5_  (.Y(\proj__6.flop5/_1_ ),
    .A(net231));
 sg13g2_tielo \proj__6.flop5/dffsr_327  (.L_LO(net368));
 sg13g2_tielo \proj__6.flop6/dffsr_328  (.L_LO(net369));
 sg13g2_sdfbbp_1 \proj__6.flop5/dffsr  (.Q(\proj__6.net29 ),
    .Q_N(\proj__6.flop5/notq ),
    .RESET_B(\proj__6.flop5/_0_ ),
    .SET_B(\proj__6.flop5/_1_ ),
    .D(\proj__6.net28 ),
    .SCE(net368),
    .SCD(net367),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop6/_4_  (.Y(\proj__6.flop6/_0_ ),
    .A(net232));
 sg13g2_inv_1 \proj__6.flop6/_5_  (.Y(\proj__6.flop6/_1_ ),
    .A(net233));
 sg13g2_tielo \proj__6.flop6/dffsr_329  (.L_LO(net370));
 sg13g2_tielo \proj__6.flop7/dffsr_330  (.L_LO(net371));
 sg13g2_sdfbbp_1 \proj__6.flop6/dffsr  (.Q(\proj__6.net30 ),
    .Q_N(\proj__6.flop6/notq ),
    .RESET_B(\proj__6.flop6/_0_ ),
    .SET_B(\proj__6.flop6/_1_ ),
    .D(\proj__6.net29 ),
    .SCE(net370),
    .SCD(net369),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop7/_4_  (.Y(\proj__6.flop7/_0_ ),
    .A(net234));
 sg13g2_inv_1 \proj__6.flop7/_5_  (.Y(\proj__6.flop7/_1_ ),
    .A(net235));
 sg13g2_tielo \proj__6.flop7/dffsr_331  (.L_LO(net372));
 sg13g2_tielo \proj__6.flop8/dffsr_332  (.L_LO(net373));
 sg13g2_sdfbbp_1 \proj__6.flop7/dffsr  (.Q(\proj__6.net27 ),
    .Q_N(\proj__6.flop7/notq ),
    .RESET_B(\proj__6.flop7/_0_ ),
    .SET_B(\proj__6.flop7/_1_ ),
    .D(\proj__6.net30 ),
    .SCE(net372),
    .SCD(net371),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop8/_4_  (.Y(\proj__6.flop8/_0_ ),
    .A(net236));
 sg13g2_inv_1 \proj__6.flop8/_5_  (.Y(\proj__6.flop8/_1_ ),
    .A(net237));
 sg13g2_tielo \proj__6.flop8/dffsr_333  (.L_LO(net374));
 sg13g2_tielo \proj__6.flop9/dffsr_334  (.L_LO(net375));
 sg13g2_sdfbbp_1 \proj__6.flop8/dffsr  (.Q(\proj__6.net33 ),
    .Q_N(\proj__6.flop8/notq ),
    .RESET_B(\proj__6.flop8/_0_ ),
    .SET_B(\proj__6.flop8/_1_ ),
    .D(\proj__6.net31 ),
    .SCE(net374),
    .SCD(net373),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop9/_4_  (.Y(\proj__6.flop9/_0_ ),
    .A(net238));
 sg13g2_inv_1 \proj__6.flop9/_5_  (.Y(\proj__6.flop9/_1_ ),
    .A(net239));
 sg13g2_tielo \proj__6.flop9/dffsr_335  (.L_LO(net376));
 sg13g2_tielo \proj__9.flop1/dffsr_336  (.L_LO(net377));
 sg13g2_sdfbbp_1 \proj__6.flop9/dffsr  (.Q(\proj__6.net34 ),
    .Q_N(\proj__6.flop9/notq ),
    .RESET_B(\proj__6.flop9/_0_ ),
    .SET_B(\proj__6.flop9/_1_ ),
    .D(\proj__6.net33 ),
    .SCE(net376),
    .SCD(net375),
    .CLK(\proj__6.net32 ));
 sg13g2_mux2_1 \proj__6.mux1/_0_  (.A0(\proj__6.net53 ),
    .A1(\proj__6.net43 ),
    .S(net127),
    .X(\proj__6.net91 ));
 sg13g2_mux2_1 \proj__6.mux10/_0_  (.A0(\proj__6.net59 ),
    .A1(\proj__6.net49 ),
    .S(net128),
    .X(\proj__6.net98 ));
 sg13g2_mux2_1 \proj__6.mux11/_0_  (.A0(\proj__6.net39 ),
    .A1(\proj__6.net29 ),
    .S(net127),
    .X(\proj__6.net99 ));
 sg13g2_mux2_1 \proj__6.mux12/_0_  (.A0(\proj__6.net98 ),
    .A1(\proj__6.net99 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net79 ));
 sg13g2_mux2_1 \proj__6.mux13/_0_  (.A0(\proj__6.net60 ),
    .A1(\proj__6.net50 ),
    .S(\proj__6.net90 ),
    .X(\proj__6.net100 ));
 sg13g2_mux2_1 \proj__6.mux14/_0_  (.A0(\proj__6.net40 ),
    .A1(\proj__6.net30 ),
    .S(net127),
    .X(\proj__6.net101 ));
 sg13g2_mux2_1 \proj__6.mux15/_0_  (.A0(\proj__6.net100 ),
    .A1(\proj__6.net101 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net81 ));
 sg13g2_mux2_1 \proj__6.mux16/_0_  (.A0(\proj__6.net57 ),
    .A1(\proj__6.net47 ),
    .S(net128),
    .X(\proj__6.net102 ));
 sg13g2_mux2_1 \proj__6.mux17/_0_  (.A0(\proj__6.net37 ),
    .A1(\proj__6.net27 ),
    .S(net127),
    .X(\proj__6.net103 ));
 sg13g2_mux2_1 \proj__6.mux18/_0_  (.A0(\proj__6.net102 ),
    .A1(\proj__6.net103 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net83 ));
 sg13g2_mux2_1 \proj__6.mux19/_0_  (.A0(\proj__6.net55 ),
    .A1(\proj__6.net45 ),
    .S(net128),
    .X(\proj__6.net104 ));
 sg13g2_mux2_1 \proj__6.mux2/_0_  (.A0(\proj__6.net54 ),
    .A1(\proj__6.net44 ),
    .S(net128),
    .X(\proj__6.net94 ));
 sg13g2_mux2_1 \proj__6.mux20/_0_  (.A0(\proj__6.net35 ),
    .A1(\proj__6.net25 ),
    .S(net128),
    .X(\proj__6.net105 ));
 sg13g2_mux2_1 \proj__6.mux21/_0_  (.A0(\proj__6.net104 ),
    .A1(\proj__6.net105 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net85 ));
 sg13g2_mux2_1 \proj__6.mux22/_0_  (.A0(\proj__6.net56 ),
    .A1(\proj__6.net46 ),
    .S(net128),
    .X(\proj__6.net106 ));
 sg13g2_mux2_1 \proj__6.mux23/_0_  (.A0(\proj__6.net36 ),
    .A1(\proj__6.net26 ),
    .S(net128),
    .X(\proj__6.net107 ));
 sg13g2_mux2_1 \proj__6.mux24/_0_  (.A0(\proj__6.net106 ),
    .A1(\proj__6.net107 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net87 ));
 sg13g2_mux2_1 \proj__6.mux3/_0_  (.A0(\proj__6.net34 ),
    .A1(\proj__6.net24 ),
    .S(net127),
    .X(\proj__6.net95 ));
 sg13g2_mux2_1 \proj__6.mux4/_0_  (.A0(\proj__6.net94 ),
    .A1(\proj__6.net95 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net75 ));
 sg13g2_mux2_1 \proj__6.mux5/_0_  (.A0(\proj__6.net33 ),
    .A1(\proj__6.net23 ),
    .S(net127),
    .X(\proj__6.net92 ));
 sg13g2_mux2_1 \proj__6.mux6/_0_  (.A0(\proj__6.net58 ),
    .A1(\proj__6.net48 ),
    .S(net127),
    .X(\proj__6.net96 ));
 sg13g2_mux2_1 \proj__6.mux7/_0_  (.A0(\proj__6.net38 ),
    .A1(\proj__6.net28 ),
    .S(net127),
    .X(\proj__6.net97 ));
 sg13g2_mux2_1 \proj__6.mux8/_0_  (.A0(\proj__6.net96 ),
    .A1(\proj__6.net97 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net77 ));
 sg13g2_mux2_1 \proj__6.mux9/_0_  (.A0(\proj__6.net91 ),
    .A1(\proj__6.net92 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net72 ));
 sg13g2_inv_1 \proj__6.not1/_0_  (.Y(\proj__6.net61 ),
    .A(net147));
 sg13g2_inv_1 \proj__6.not2/_0_  (.Y(\proj__6.net62 ),
    .A(net145));
 sg13g2_inv_1 \proj__6.not3/_0_  (.Y(\proj__6.net90 ),
    .A(net133));
 sg13g2_inv_4 \proj__6.not4/_0_  (.A(net132),
    .Y(\proj__6.net93 ));
 sg13g2_nand2_1 \proj__7.nand1/_0_  (.Y(\proj__7.net11 ),
    .A(net144),
    .B(net147));
 sg13g2_nand2_1 \proj__7.nand2/_0_  (.Y(\proj__7.net12 ),
    .A(net140),
    .B(net144));
 sg13g2_nand2_1 \proj__7.nand3/_0_  (.Y(\proj__7.net4 ),
    .A(\proj__7.net5 ),
    .B(\proj__7.net11 ));
 sg13g2_nand2_1 \proj__7.nand4/_0_  (.Y(\proj__7.net5 ),
    .A(\proj__7.net12 ),
    .B(\proj__7.net4 ));
 sg13g2_and2_1 \proj__9.and1/_0_  (.A(net143),
    .B(\proj__9.net16 ),
    .X(\proj__9.net5 ));
 sg13g2_and2_1 \proj__9.and2/_0_  (.A(net143),
    .B(\proj__9.net18 ),
    .X(\proj__9.net6 ));
 sg13g2_and2_1 \proj__9.and3/_0_  (.A(net144),
    .B(\proj__9.net19 ),
    .X(\proj__9.net7 ));
 sg13g2_and2_1 \proj__9.and4/_0_  (.A(net144),
    .B(\proj__9.net20 ),
    .X(\proj__9.net8 ));
 sg13g2_inv_1 \proj__9.flop1/_4_  (.Y(\proj__9.flop1/_0_ ),
    .A(\proj__9.net15 ));
 sg13g2_inv_1 \proj__9.flop1/_5_  (.Y(\proj__9.flop1/_1_ ),
    .A(net241));
 sg13g2_tielo \proj__9.flop1/dffsr_337  (.L_LO(net378));
 sg13g2_tielo \proj__9.flop2/dffsr_338  (.L_LO(net379));
 sg13g2_sdfbbp_1 \proj__9.flop1/dffsr  (.Q(\proj__9.net16 ),
    .Q_N(\proj__9.flop1/notq ),
    .RESET_B(\proj__9.flop1/_0_ ),
    .SET_B(\proj__9.flop1/_1_ ),
    .D(net148),
    .SCE(net378),
    .SCD(net377),
    .CLK(net240));
 sg13g2_inv_1 \proj__9.flop2/_4_  (.Y(\proj__9.flop2/_0_ ),
    .A(\proj__9.net15 ));
 sg13g2_inv_1 \proj__9.flop2/_5_  (.Y(\proj__9.flop2/_1_ ),
    .A(net243));
 sg13g2_tielo \proj__9.flop2/dffsr_339  (.L_LO(net380));
 sg13g2_tielo \proj__9.flop3/dffsr_340  (.L_LO(net381));
 sg13g2_sdfbbp_1 \proj__9.flop2/dffsr  (.Q(\proj__9.net18 ),
    .Q_N(\proj__9.flop2/notq ),
    .RESET_B(\proj__9.flop2/_0_ ),
    .SET_B(\proj__9.flop2/_1_ ),
    .D(\proj__9.net16 ),
    .SCE(net380),
    .SCD(net379),
    .CLK(net242));
 sg13g2_inv_1 \proj__9.flop3/_4_  (.Y(\proj__9.flop3/_0_ ),
    .A(\proj__9.net15 ));
 sg13g2_inv_1 \proj__9.flop3/_5_  (.Y(\proj__9.flop3/_1_ ),
    .A(net245));
 sg13g2_tielo \proj__9.flop3/dffsr_341  (.L_LO(net382));
 sg13g2_tielo \proj__9.flop4/dffsr_342  (.L_LO(net383));
 sg13g2_sdfbbp_1 \proj__9.flop3/dffsr  (.Q(\proj__9.net19 ),
    .Q_N(\proj__9.flop3/notq ),
    .RESET_B(\proj__9.flop3/_0_ ),
    .SET_B(\proj__9.flop3/_1_ ),
    .D(\proj__9.net18 ),
    .SCE(net382),
    .SCD(net381),
    .CLK(net244));
 sg13g2_inv_1 \proj__9.flop4/_4_  (.Y(\proj__9.flop4/_0_ ),
    .A(\proj__9.net15 ));
 sg13g2_inv_1 \proj__9.flop4/_5_  (.Y(\proj__9.flop4/_1_ ),
    .A(net247));
 sg13g2_tielo \proj__9.flop4/dffsr_343  (.L_LO(net384));
 sg13g2_tiehi \proj__4.and1/_0__344  (.L_HI(net385));
 sg13g2_sdfbbp_1 \proj__9.flop4/dffsr  (.Q(\proj__9.net20 ),
    .Q_N(\proj__9.flop4/notq ),
    .RESET_B(\proj__9.flop4/_0_ ),
    .SET_B(\proj__9.flop4/_1_ ),
    .D(\proj__9.net19 ),
    .SCE(net384),
    .SCD(net383),
    .CLK(net246));
 sg13g2_inv_1 \proj__9.not1/_0_  (.Y(\proj__9.net15 ),
    .A(net248));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(net128));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(\proj__6.net90 ));
 sg13g2_buf_2 fanout129 (.A(net131),
    .X(net129));
 sg13g2_buf_1 fanout130 (.A(net131),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(ui_in[7]),
    .X(net131));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(net5));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(net4));
 sg13g2_buf_2 fanout134 (.A(net4),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(ui_in[4]),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(net3),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(net142),
    .X(net140));
 sg13g2_buf_1 fanout141 (.A(net142),
    .X(net141));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(net2));
 sg13g2_buf_2 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(net145),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(net146),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(ui_in[1]),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(net1));
 sg13g2_buf_4 fanout149 (.X(net149),
    .A(\proj__4.net34 ));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(net151));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(\proj__4.net31 ));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(net153));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(net156));
 sg13g2_buf_4 fanout154 (.X(net154),
    .A(net156));
 sg13g2_buf_2 fanout155 (.A(net156),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(\proj__4.net26 ),
    .X(net156));
 sg13g2_buf_4 fanout157 (.X(net157),
    .A(net161));
 sg13g2_buf_2 fanout158 (.A(net161),
    .X(net158));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(net160));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(net161));
 sg13g2_buf_2 fanout161 (.A(net167),
    .X(net161));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(net164));
 sg13g2_buf_2 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(net167),
    .X(net164));
 sg13g2_buf_4 fanout165 (.X(net165),
    .A(net167));
 sg13g2_buf_2 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(\proj__4.net16 ),
    .X(net167));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_tielo \proj_10.flop1/dffsr_10  (.L_LO(net10));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_4 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_193 ();
 sg13g2_decap_8 FILLER_9_198 ();
 sg13g2_decap_8 FILLER_9_209 ();
 sg13g2_decap_8 FILLER_9_216 ();
 sg13g2_decap_8 FILLER_9_223 ();
 sg13g2_fill_2 FILLER_9_230 ();
 sg13g2_decap_4 FILLER_9_236 ();
 sg13g2_fill_1 FILLER_9_240 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_4 FILLER_9_259 ();
 sg13g2_fill_2 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_268 ();
 sg13g2_fill_1 FILLER_9_275 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_fill_2 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_306 ();
 sg13g2_decap_8 FILLER_9_313 ();
 sg13g2_decap_8 FILLER_9_320 ();
 sg13g2_decap_8 FILLER_9_327 ();
 sg13g2_decap_8 FILLER_9_334 ();
 sg13g2_decap_8 FILLER_9_341 ();
 sg13g2_decap_8 FILLER_9_348 ();
 sg13g2_decap_8 FILLER_9_355 ();
 sg13g2_decap_8 FILLER_9_362 ();
 sg13g2_decap_8 FILLER_9_369 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_fill_2 FILLER_10_154 ();
 sg13g2_fill_1 FILLER_10_156 ();
 sg13g2_decap_8 FILLER_10_160 ();
 sg13g2_decap_8 FILLER_10_170 ();
 sg13g2_fill_1 FILLER_10_177 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_fill_2 FILLER_11_179 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_4 FILLER_11_200 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_decap_8 FILLER_11_222 ();
 sg13g2_fill_2 FILLER_11_229 ();
 sg13g2_decap_4 FILLER_11_234 ();
 sg13g2_fill_2 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_243 ();
 sg13g2_decap_8 FILLER_11_258 ();
 sg13g2_fill_1 FILLER_11_265 ();
 sg13g2_decap_4 FILLER_11_270 ();
 sg13g2_fill_1 FILLER_11_274 ();
 sg13g2_decap_8 FILLER_11_278 ();
 sg13g2_fill_1 FILLER_11_285 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_fill_2 FILLER_11_301 ();
 sg13g2_fill_1 FILLER_11_303 ();
 sg13g2_decap_4 FILLER_11_308 ();
 sg13g2_fill_1 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_317 ();
 sg13g2_decap_8 FILLER_11_324 ();
 sg13g2_decap_8 FILLER_11_331 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_decap_8 FILLER_11_345 ();
 sg13g2_decap_8 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_fill_2 FILLER_12_119 ();
 sg13g2_fill_1 FILLER_12_121 ();
 sg13g2_decap_4 FILLER_12_125 ();
 sg13g2_fill_2 FILLER_12_129 ();
 sg13g2_decap_8 FILLER_12_135 ();
 sg13g2_fill_1 FILLER_12_142 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_4 FILLER_12_162 ();
 sg13g2_decap_8 FILLER_12_169 ();
 sg13g2_fill_2 FILLER_12_176 ();
 sg13g2_decap_8 FILLER_12_188 ();
 sg13g2_decap_4 FILLER_12_195 ();
 sg13g2_fill_2 FILLER_12_203 ();
 sg13g2_fill_1 FILLER_12_205 ();
 sg13g2_decap_4 FILLER_12_213 ();
 sg13g2_fill_1 FILLER_12_255 ();
 sg13g2_decap_8 FILLER_12_260 ();
 sg13g2_decap_4 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_271 ();
 sg13g2_fill_1 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_295 ();
 sg13g2_decap_8 FILLER_12_302 ();
 sg13g2_fill_1 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_327 ();
 sg13g2_decap_8 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_341 ();
 sg13g2_decap_8 FILLER_12_348 ();
 sg13g2_decap_8 FILLER_12_355 ();
 sg13g2_decap_8 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_369 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_4 FILLER_13_232 ();
 sg13g2_fill_1 FILLER_13_253 ();
 sg13g2_decap_8 FILLER_13_328 ();
 sg13g2_decap_8 FILLER_13_335 ();
 sg13g2_decap_8 FILLER_13_342 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_fill_2 FILLER_14_105 ();
 sg13g2_fill_1 FILLER_14_107 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_fill_2 FILLER_14_127 ();
 sg13g2_fill_1 FILLER_14_129 ();
 sg13g2_fill_2 FILLER_14_136 ();
 sg13g2_fill_1 FILLER_14_138 ();
 sg13g2_fill_1 FILLER_14_142 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_fill_2 FILLER_14_158 ();
 sg13g2_decap_4 FILLER_14_171 ();
 sg13g2_fill_2 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_fill_2 FILLER_14_196 ();
 sg13g2_decap_4 FILLER_14_205 ();
 sg13g2_decap_8 FILLER_14_212 ();
 sg13g2_decap_4 FILLER_14_219 ();
 sg13g2_fill_2 FILLER_14_223 ();
 sg13g2_decap_8 FILLER_14_229 ();
 sg13g2_decap_4 FILLER_14_236 ();
 sg13g2_fill_1 FILLER_14_240 ();
 sg13g2_fill_2 FILLER_14_249 ();
 sg13g2_fill_1 FILLER_14_251 ();
 sg13g2_fill_1 FILLER_14_256 ();
 sg13g2_decap_8 FILLER_14_261 ();
 sg13g2_decap_4 FILLER_14_268 ();
 sg13g2_decap_8 FILLER_14_275 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_fill_2 FILLER_14_290 ();
 sg13g2_fill_2 FILLER_14_296 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_1 FILLER_14_307 ();
 sg13g2_fill_2 FILLER_14_311 ();
 sg13g2_fill_1 FILLER_14_313 ();
 sg13g2_decap_8 FILLER_14_317 ();
 sg13g2_fill_1 FILLER_14_324 ();
 sg13g2_fill_2 FILLER_14_332 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_decap_8 FILLER_14_345 ();
 sg13g2_decap_4 FILLER_14_356 ();
 sg13g2_fill_1 FILLER_14_360 ();
 sg13g2_fill_2 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_4 FILLER_14_385 ();
 sg13g2_decap_4 FILLER_14_393 ();
 sg13g2_fill_1 FILLER_14_397 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_fill_1 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_decap_4 FILLER_15_172 ();
 sg13g2_fill_2 FILLER_15_176 ();
 sg13g2_fill_2 FILLER_15_221 ();
 sg13g2_fill_1 FILLER_15_296 ();
 sg13g2_fill_1 FILLER_15_332 ();
 sg13g2_fill_1 FILLER_15_368 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_fill_2 FILLER_16_77 ();
 sg13g2_fill_1 FILLER_16_114 ();
 sg13g2_decap_8 FILLER_16_123 ();
 sg13g2_fill_1 FILLER_16_130 ();
 sg13g2_decap_4 FILLER_16_135 ();
 sg13g2_fill_1 FILLER_16_139 ();
 sg13g2_decap_8 FILLER_16_144 ();
 sg13g2_fill_1 FILLER_16_151 ();
 sg13g2_decap_4 FILLER_16_166 ();
 sg13g2_fill_1 FILLER_16_170 ();
 sg13g2_decap_4 FILLER_16_175 ();
 sg13g2_fill_2 FILLER_16_190 ();
 sg13g2_decap_8 FILLER_16_205 ();
 sg13g2_decap_4 FILLER_16_212 ();
 sg13g2_fill_2 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_232 ();
 sg13g2_fill_1 FILLER_16_239 ();
 sg13g2_fill_2 FILLER_16_243 ();
 sg13g2_decap_4 FILLER_16_255 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_fill_1 FILLER_16_287 ();
 sg13g2_decap_4 FILLER_16_292 ();
 sg13g2_fill_1 FILLER_16_296 ();
 sg13g2_decap_8 FILLER_16_305 ();
 sg13g2_fill_2 FILLER_16_312 ();
 sg13g2_fill_1 FILLER_16_314 ();
 sg13g2_decap_4 FILLER_16_319 ();
 sg13g2_fill_2 FILLER_16_323 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_fill_2 FILLER_16_349 ();
 sg13g2_fill_1 FILLER_16_354 ();
 sg13g2_fill_2 FILLER_16_358 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_4 FILLER_16_382 ();
 sg13g2_fill_1 FILLER_16_386 ();
 sg13g2_fill_2 FILLER_16_393 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_4 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_89 ();
 sg13g2_decap_4 FILLER_17_103 ();
 sg13g2_decap_8 FILLER_17_111 ();
 sg13g2_decap_4 FILLER_17_118 ();
 sg13g2_decap_4 FILLER_17_126 ();
 sg13g2_fill_1 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_134 ();
 sg13g2_fill_1 FILLER_17_136 ();
 sg13g2_fill_1 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_201 ();
 sg13g2_decap_4 FILLER_17_208 ();
 sg13g2_fill_2 FILLER_17_216 ();
 sg13g2_fill_1 FILLER_17_218 ();
 sg13g2_decap_8 FILLER_17_240 ();
 sg13g2_decap_4 FILLER_17_247 ();
 sg13g2_fill_1 FILLER_17_251 ();
 sg13g2_decap_8 FILLER_17_256 ();
 sg13g2_decap_8 FILLER_17_270 ();
 sg13g2_decap_4 FILLER_17_277 ();
 sg13g2_fill_2 FILLER_17_281 ();
 sg13g2_fill_2 FILLER_17_293 ();
 sg13g2_fill_1 FILLER_17_295 ();
 sg13g2_fill_2 FILLER_17_306 ();
 sg13g2_decap_8 FILLER_17_318 ();
 sg13g2_decap_4 FILLER_17_325 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_4 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_145 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_decap_8 FILLER_18_163 ();
 sg13g2_decap_4 FILLER_18_176 ();
 sg13g2_fill_1 FILLER_18_180 ();
 sg13g2_decap_4 FILLER_18_185 ();
 sg13g2_fill_2 FILLER_18_189 ();
 sg13g2_fill_2 FILLER_18_230 ();
 sg13g2_fill_1 FILLER_18_232 ();
 sg13g2_decap_8 FILLER_18_276 ();
 sg13g2_decap_4 FILLER_18_287 ();
 sg13g2_fill_1 FILLER_18_291 ();
 sg13g2_fill_2 FILLER_18_299 ();
 sg13g2_decap_8 FILLER_18_309 ();
 sg13g2_fill_2 FILLER_18_316 ();
 sg13g2_fill_1 FILLER_18_318 ();
 sg13g2_decap_4 FILLER_18_323 ();
 sg13g2_decap_8 FILLER_18_339 ();
 sg13g2_fill_1 FILLER_18_346 ();
 sg13g2_decap_4 FILLER_18_351 ();
 sg13g2_fill_1 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_18_370 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_4 FILLER_18_384 ();
 sg13g2_decap_4 FILLER_18_392 ();
 sg13g2_fill_2 FILLER_18_396 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_fill_2 FILLER_19_49 ();
 sg13g2_fill_1 FILLER_19_51 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_fill_1 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_82 ();
 sg13g2_decap_4 FILLER_19_89 ();
 sg13g2_decap_4 FILLER_19_97 ();
 sg13g2_fill_1 FILLER_19_101 ();
 sg13g2_decap_4 FILLER_19_109 ();
 sg13g2_fill_1 FILLER_19_113 ();
 sg13g2_fill_2 FILLER_19_118 ();
 sg13g2_fill_1 FILLER_19_120 ();
 sg13g2_decap_4 FILLER_19_124 ();
 sg13g2_fill_2 FILLER_19_128 ();
 sg13g2_fill_2 FILLER_19_137 ();
 sg13g2_fill_1 FILLER_19_139 ();
 sg13g2_decap_4 FILLER_19_150 ();
 sg13g2_decap_4 FILLER_19_199 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_fill_2 FILLER_19_224 ();
 sg13g2_fill_1 FILLER_19_226 ();
 sg13g2_decap_4 FILLER_19_231 ();
 sg13g2_fill_2 FILLER_19_239 ();
 sg13g2_fill_2 FILLER_19_248 ();
 sg13g2_fill_1 FILLER_19_250 ();
 sg13g2_decap_4 FILLER_19_257 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_fill_2 FILLER_20_35 ();
 sg13g2_fill_1 FILLER_20_37 ();
 sg13g2_fill_1 FILLER_20_46 ();
 sg13g2_fill_2 FILLER_20_73 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_fill_2 FILLER_20_150 ();
 sg13g2_decap_8 FILLER_20_166 ();
 sg13g2_fill_1 FILLER_20_173 ();
 sg13g2_fill_2 FILLER_20_178 ();
 sg13g2_decap_8 FILLER_20_183 ();
 sg13g2_decap_4 FILLER_20_190 ();
 sg13g2_fill_2 FILLER_20_194 ();
 sg13g2_fill_2 FILLER_20_218 ();
 sg13g2_fill_2 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_271 ();
 sg13g2_fill_1 FILLER_20_278 ();
 sg13g2_decap_8 FILLER_20_286 ();
 sg13g2_fill_2 FILLER_20_293 ();
 sg13g2_fill_1 FILLER_20_295 ();
 sg13g2_fill_2 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_310 ();
 sg13g2_fill_1 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_321 ();
 sg13g2_decap_8 FILLER_20_328 ();
 sg13g2_decap_4 FILLER_20_354 ();
 sg13g2_fill_1 FILLER_20_358 ();
 sg13g2_decap_4 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_25 ();
 sg13g2_decap_4 FILLER_21_32 ();
 sg13g2_fill_1 FILLER_21_36 ();
 sg13g2_decap_8 FILLER_21_51 ();
 sg13g2_fill_2 FILLER_21_62 ();
 sg13g2_fill_2 FILLER_21_73 ();
 sg13g2_fill_1 FILLER_21_75 ();
 sg13g2_decap_4 FILLER_21_80 ();
 sg13g2_fill_1 FILLER_21_84 ();
 sg13g2_fill_2 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_95 ();
 sg13g2_fill_1 FILLER_21_102 ();
 sg13g2_decap_8 FILLER_21_117 ();
 sg13g2_decap_8 FILLER_21_124 ();
 sg13g2_decap_8 FILLER_21_144 ();
 sg13g2_decap_4 FILLER_21_151 ();
 sg13g2_fill_1 FILLER_21_155 ();
 sg13g2_decap_8 FILLER_21_160 ();
 sg13g2_decap_4 FILLER_21_167 ();
 sg13g2_fill_2 FILLER_21_171 ();
 sg13g2_decap_8 FILLER_21_183 ();
 sg13g2_decap_4 FILLER_21_190 ();
 sg13g2_decap_8 FILLER_21_218 ();
 sg13g2_fill_2 FILLER_21_225 ();
 sg13g2_decap_8 FILLER_21_232 ();
 sg13g2_fill_1 FILLER_21_239 ();
 sg13g2_fill_2 FILLER_21_275 ();
 sg13g2_decap_4 FILLER_21_316 ();
 sg13g2_fill_2 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_356 ();
 sg13g2_decap_8 FILLER_21_363 ();
 sg13g2_decap_8 FILLER_21_370 ();
 sg13g2_decap_8 FILLER_21_377 ();
 sg13g2_decap_8 FILLER_21_384 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_30 ();
 sg13g2_fill_1 FILLER_22_55 ();
 sg13g2_fill_1 FILLER_22_80 ();
 sg13g2_decap_4 FILLER_22_99 ();
 sg13g2_decap_8 FILLER_22_121 ();
 sg13g2_fill_2 FILLER_22_128 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_decap_4 FILLER_22_145 ();
 sg13g2_fill_2 FILLER_22_149 ();
 sg13g2_fill_2 FILLER_22_194 ();
 sg13g2_fill_1 FILLER_22_196 ();
 sg13g2_decap_4 FILLER_22_236 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_decap_4 FILLER_22_253 ();
 sg13g2_fill_2 FILLER_22_257 ();
 sg13g2_decap_4 FILLER_22_263 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_4 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_295 ();
 sg13g2_decap_4 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_4 FILLER_22_315 ();
 sg13g2_fill_2 FILLER_22_319 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_26 ();
 sg13g2_decap_8 FILLER_23_33 ();
 sg13g2_fill_1 FILLER_23_40 ();
 sg13g2_decap_8 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_60 ();
 sg13g2_fill_1 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_78 ();
 sg13g2_decap_8 FILLER_23_89 ();
 sg13g2_decap_4 FILLER_23_96 ();
 sg13g2_fill_2 FILLER_23_100 ();
 sg13g2_decap_8 FILLER_23_120 ();
 sg13g2_decap_8 FILLER_23_149 ();
 sg13g2_fill_1 FILLER_23_160 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_fill_1 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_229 ();
 sg13g2_fill_1 FILLER_23_269 ();
 sg13g2_decap_4 FILLER_23_317 ();
 sg13g2_fill_1 FILLER_23_321 ();
 sg13g2_fill_1 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_338 ();
 sg13g2_decap_8 FILLER_23_345 ();
 sg13g2_fill_2 FILLER_23_352 ();
 sg13g2_fill_2 FILLER_23_358 ();
 sg13g2_fill_1 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_fill_2 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_48 ();
 sg13g2_decap_4 FILLER_24_55 ();
 sg13g2_fill_2 FILLER_24_59 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_fill_1 FILLER_24_88 ();
 sg13g2_fill_2 FILLER_24_99 ();
 sg13g2_decap_4 FILLER_24_109 ();
 sg13g2_fill_2 FILLER_24_113 ();
 sg13g2_fill_2 FILLER_24_125 ();
 sg13g2_fill_1 FILLER_24_127 ();
 sg13g2_decap_8 FILLER_24_148 ();
 sg13g2_decap_8 FILLER_24_155 ();
 sg13g2_fill_1 FILLER_24_162 ();
 sg13g2_fill_1 FILLER_24_171 ();
 sg13g2_decap_4 FILLER_24_175 ();
 sg13g2_fill_1 FILLER_24_179 ();
 sg13g2_fill_2 FILLER_24_187 ();
 sg13g2_fill_1 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_194 ();
 sg13g2_decap_8 FILLER_24_226 ();
 sg13g2_decap_8 FILLER_24_241 ();
 sg13g2_fill_2 FILLER_24_248 ();
 sg13g2_fill_1 FILLER_24_250 ();
 sg13g2_decap_4 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_259 ();
 sg13g2_decap_4 FILLER_24_264 ();
 sg13g2_fill_2 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_decap_4 FILLER_24_292 ();
 sg13g2_fill_2 FILLER_24_307 ();
 sg13g2_decap_4 FILLER_24_313 ();
 sg13g2_fill_1 FILLER_24_317 ();
 sg13g2_fill_1 FILLER_24_328 ();
 sg13g2_fill_2 FILLER_24_346 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_fill_1 FILLER_24_389 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_17 ();
 sg13g2_decap_8 FILLER_25_24 ();
 sg13g2_decap_4 FILLER_25_31 ();
 sg13g2_fill_2 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_55 ();
 sg13g2_fill_1 FILLER_25_83 ();
 sg13g2_fill_2 FILLER_25_112 ();
 sg13g2_fill_1 FILLER_25_114 ();
 sg13g2_fill_2 FILLER_25_123 ();
 sg13g2_decap_8 FILLER_25_149 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_decap_8 FILLER_25_200 ();
 sg13g2_decap_4 FILLER_25_207 ();
 sg13g2_fill_2 FILLER_25_211 ();
 sg13g2_decap_8 FILLER_25_233 ();
 sg13g2_decap_8 FILLER_25_250 ();
 sg13g2_decap_4 FILLER_25_257 ();
 sg13g2_fill_2 FILLER_25_261 ();
 sg13g2_fill_1 FILLER_25_293 ();
 sg13g2_decap_8 FILLER_25_339 ();
 sg13g2_decap_8 FILLER_25_346 ();
 sg13g2_decap_4 FILLER_25_353 ();
 sg13g2_decap_8 FILLER_25_362 ();
 sg13g2_fill_1 FILLER_25_369 ();
 sg13g2_fill_1 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_fill_2 FILLER_25_389 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_4 ();
 sg13g2_decap_4 FILLER_26_26 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_4 FILLER_26_63 ();
 sg13g2_fill_2 FILLER_26_67 ();
 sg13g2_fill_2 FILLER_26_97 ();
 sg13g2_decap_4 FILLER_26_109 ();
 sg13g2_fill_2 FILLER_26_113 ();
 sg13g2_fill_2 FILLER_26_133 ();
 sg13g2_fill_1 FILLER_26_135 ();
 sg13g2_fill_2 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_152 ();
 sg13g2_decap_4 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_171 ();
 sg13g2_decap_4 FILLER_26_177 ();
 sg13g2_fill_2 FILLER_26_181 ();
 sg13g2_decap_4 FILLER_26_187 ();
 sg13g2_fill_1 FILLER_26_209 ();
 sg13g2_fill_2 FILLER_26_231 ();
 sg13g2_decap_4 FILLER_26_239 ();
 sg13g2_fill_1 FILLER_26_243 ();
 sg13g2_fill_2 FILLER_26_258 ();
 sg13g2_fill_1 FILLER_26_260 ();
 sg13g2_fill_2 FILLER_26_267 ();
 sg13g2_fill_1 FILLER_26_269 ();
 sg13g2_fill_2 FILLER_26_274 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_fill_2 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_330 ();
 sg13g2_decap_4 FILLER_26_337 ();
 sg13g2_fill_1 FILLER_26_341 ();
 sg13g2_decap_4 FILLER_26_362 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_4 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_4 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_fill_2 FILLER_27_50 ();
 sg13g2_fill_1 FILLER_27_52 ();
 sg13g2_decap_4 FILLER_27_78 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_93 ();
 sg13g2_decap_8 FILLER_27_137 ();
 sg13g2_decap_4 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_148 ();
 sg13g2_decap_4 FILLER_27_153 ();
 sg13g2_fill_2 FILLER_27_167 ();
 sg13g2_decap_8 FILLER_27_179 ();
 sg13g2_fill_2 FILLER_27_186 ();
 sg13g2_decap_8 FILLER_27_194 ();
 sg13g2_decap_4 FILLER_27_201 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_fill_2 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_254 ();
 sg13g2_fill_1 FILLER_27_261 ();
 sg13g2_decap_8 FILLER_27_276 ();
 sg13g2_fill_1 FILLER_27_283 ();
 sg13g2_decap_4 FILLER_27_289 ();
 sg13g2_fill_1 FILLER_27_312 ();
 sg13g2_fill_1 FILLER_27_341 ();
 sg13g2_fill_2 FILLER_27_370 ();
 sg13g2_decap_8 FILLER_27_376 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_decap_4 FILLER_27_390 ();
 sg13g2_fill_1 FILLER_27_394 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_4 ();
 sg13g2_fill_2 FILLER_28_9 ();
 sg13g2_fill_1 FILLER_28_31 ();
 sg13g2_fill_2 FILLER_28_37 ();
 sg13g2_decap_8 FILLER_28_57 ();
 sg13g2_fill_1 FILLER_28_64 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_101 ();
 sg13g2_decap_8 FILLER_28_108 ();
 sg13g2_decap_4 FILLER_28_115 ();
 sg13g2_fill_1 FILLER_28_119 ();
 sg13g2_fill_2 FILLER_28_124 ();
 sg13g2_fill_1 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_137 ();
 sg13g2_decap_4 FILLER_28_164 ();
 sg13g2_fill_2 FILLER_28_178 ();
 sg13g2_decap_4 FILLER_28_190 ();
 sg13g2_fill_2 FILLER_28_194 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_fill_1 FILLER_28_233 ();
 sg13g2_decap_4 FILLER_28_250 ();
 sg13g2_fill_2 FILLER_28_254 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_295 ();
 sg13g2_decap_4 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_306 ();
 sg13g2_decap_4 FILLER_28_322 ();
 sg13g2_fill_2 FILLER_28_326 ();
 sg13g2_decap_4 FILLER_28_338 ();
 sg13g2_decap_8 FILLER_28_352 ();
 sg13g2_fill_2 FILLER_28_359 ();
 sg13g2_fill_1 FILLER_28_361 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_2 FILLER_29_31 ();
 sg13g2_fill_1 FILLER_29_37 ();
 sg13g2_decap_4 FILLER_29_57 ();
 sg13g2_decap_4 FILLER_29_95 ();
 sg13g2_fill_2 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_decap_8 FILLER_29_146 ();
 sg13g2_decap_8 FILLER_29_153 ();
 sg13g2_decap_4 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_164 ();
 sg13g2_decap_4 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_fill_1 FILLER_29_196 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_decap_8 FILLER_29_215 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_231 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_fill_2 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_276 ();
 sg13g2_decap_8 FILLER_29_293 ();
 sg13g2_decap_8 FILLER_29_310 ();
 sg13g2_fill_1 FILLER_29_317 ();
 sg13g2_fill_2 FILLER_29_338 ();
 sg13g2_fill_1 FILLER_29_340 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_4 FILLER_29_358 ();
 sg13g2_fill_1 FILLER_29_362 ();
 sg13g2_decap_4 FILLER_29_375 ();
 sg13g2_fill_1 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_19 ();
 sg13g2_decap_8 FILLER_30_26 ();
 sg13g2_decap_4 FILLER_30_33 ();
 sg13g2_decap_8 FILLER_30_51 ();
 sg13g2_decap_8 FILLER_30_58 ();
 sg13g2_fill_1 FILLER_30_73 ();
 sg13g2_fill_2 FILLER_30_78 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_fill_1 FILLER_30_93 ();
 sg13g2_fill_2 FILLER_30_108 ();
 sg13g2_decap_4 FILLER_30_114 ();
 sg13g2_fill_1 FILLER_30_118 ();
 sg13g2_fill_2 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_178 ();
 sg13g2_fill_1 FILLER_30_189 ();
 sg13g2_decap_4 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_197 ();
 sg13g2_fill_1 FILLER_30_234 ();
 sg13g2_decap_4 FILLER_30_247 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_decap_8 FILLER_30_267 ();
 sg13g2_decap_4 FILLER_30_274 ();
 sg13g2_fill_1 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_297 ();
 sg13g2_fill_2 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_351 ();
 sg13g2_decap_8 FILLER_30_358 ();
 sg13g2_decap_8 FILLER_30_386 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_28 ();
 sg13g2_fill_1 FILLER_31_30 ();
 sg13g2_fill_1 FILLER_31_55 ();
 sg13g2_decap_4 FILLER_31_71 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_fill_2 FILLER_31_89 ();
 sg13g2_fill_1 FILLER_31_99 ();
 sg13g2_decap_4 FILLER_31_120 ();
 sg13g2_fill_1 FILLER_31_124 ();
 sg13g2_fill_1 FILLER_31_130 ();
 sg13g2_fill_2 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_146 ();
 sg13g2_decap_8 FILLER_31_153 ();
 sg13g2_fill_1 FILLER_31_160 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_fill_2 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_207 ();
 sg13g2_fill_2 FILLER_31_220 ();
 sg13g2_fill_1 FILLER_31_222 ();
 sg13g2_fill_2 FILLER_31_229 ();
 sg13g2_fill_1 FILLER_31_231 ();
 sg13g2_fill_2 FILLER_31_238 ();
 sg13g2_fill_1 FILLER_31_240 ();
 sg13g2_decap_8 FILLER_31_247 ();
 sg13g2_decap_8 FILLER_31_254 ();
 sg13g2_decap_8 FILLER_31_261 ();
 sg13g2_decap_4 FILLER_31_288 ();
 sg13g2_fill_1 FILLER_31_297 ();
 sg13g2_decap_4 FILLER_31_316 ();
 sg13g2_fill_2 FILLER_31_320 ();
 sg13g2_decap_4 FILLER_31_337 ();
 sg13g2_fill_2 FILLER_31_361 ();
 sg13g2_fill_1 FILLER_31_363 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_26 ();
 sg13g2_decap_4 FILLER_32_33 ();
 sg13g2_fill_1 FILLER_32_37 ();
 sg13g2_decap_8 FILLER_32_54 ();
 sg13g2_decap_4 FILLER_32_61 ();
 sg13g2_decap_4 FILLER_32_83 ();
 sg13g2_decap_4 FILLER_32_99 ();
 sg13g2_decap_4 FILLER_32_111 ();
 sg13g2_decap_4 FILLER_32_123 ();
 sg13g2_fill_1 FILLER_32_127 ();
 sg13g2_decap_8 FILLER_32_138 ();
 sg13g2_fill_1 FILLER_32_145 ();
 sg13g2_fill_2 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_174 ();
 sg13g2_decap_8 FILLER_32_179 ();
 sg13g2_decap_4 FILLER_32_186 ();
 sg13g2_fill_2 FILLER_32_190 ();
 sg13g2_fill_2 FILLER_32_215 ();
 sg13g2_decap_8 FILLER_32_233 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_279 ();
 sg13g2_fill_2 FILLER_32_286 ();
 sg13g2_fill_1 FILLER_32_288 ();
 sg13g2_decap_8 FILLER_32_299 ();
 sg13g2_fill_2 FILLER_32_320 ();
 sg13g2_decap_8 FILLER_32_326 ();
 sg13g2_fill_2 FILLER_32_333 ();
 sg13g2_fill_1 FILLER_32_335 ();
 sg13g2_decap_8 FILLER_32_349 ();
 sg13g2_decap_8 FILLER_32_356 ();
 sg13g2_fill_2 FILLER_32_363 ();
 sg13g2_fill_1 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_32_384 ();
 sg13g2_decap_4 FILLER_32_391 ();
 sg13g2_fill_2 FILLER_32_395 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_9 ();
 sg13g2_decap_4 FILLER_33_30 ();
 sg13g2_fill_2 FILLER_33_54 ();
 sg13g2_decap_8 FILLER_33_66 ();
 sg13g2_decap_8 FILLER_33_73 ();
 sg13g2_fill_2 FILLER_33_80 ();
 sg13g2_decap_4 FILLER_33_97 ();
 sg13g2_decap_8 FILLER_33_111 ();
 sg13g2_fill_2 FILLER_33_118 ();
 sg13g2_fill_1 FILLER_33_120 ();
 sg13g2_fill_2 FILLER_33_149 ();
 sg13g2_fill_2 FILLER_33_155 ();
 sg13g2_fill_2 FILLER_33_161 ();
 sg13g2_fill_1 FILLER_33_163 ();
 sg13g2_fill_1 FILLER_33_190 ();
 sg13g2_decap_8 FILLER_33_202 ();
 sg13g2_decap_4 FILLER_33_209 ();
 sg13g2_fill_1 FILLER_33_218 ();
 sg13g2_fill_2 FILLER_33_227 ();
 sg13g2_fill_1 FILLER_33_229 ();
 sg13g2_fill_2 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_253 ();
 sg13g2_fill_1 FILLER_33_269 ();
 sg13g2_decap_4 FILLER_33_287 ();
 sg13g2_decap_4 FILLER_33_355 ();
 sg13g2_fill_1 FILLER_33_359 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_24 ();
 sg13g2_fill_1 FILLER_34_26 ();
 sg13g2_fill_1 FILLER_34_49 ();
 sg13g2_fill_1 FILLER_34_79 ();
 sg13g2_fill_2 FILLER_34_100 ();
 sg13g2_fill_1 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_127 ();
 sg13g2_decap_8 FILLER_34_142 ();
 sg13g2_decap_4 FILLER_34_149 ();
 sg13g2_fill_1 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_158 ();
 sg13g2_fill_1 FILLER_34_160 ();
 sg13g2_decap_4 FILLER_34_165 ();
 sg13g2_decap_8 FILLER_34_173 ();
 sg13g2_fill_2 FILLER_34_180 ();
 sg13g2_fill_1 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_186 ();
 sg13g2_fill_1 FILLER_34_210 ();
 sg13g2_fill_2 FILLER_34_223 ();
 sg13g2_fill_2 FILLER_34_233 ();
 sg13g2_fill_1 FILLER_34_235 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_4 FILLER_34_259 ();
 sg13g2_fill_1 FILLER_34_263 ();
 sg13g2_decap_8 FILLER_34_278 ();
 sg13g2_decap_4 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_302 ();
 sg13g2_decap_8 FILLER_34_307 ();
 sg13g2_decap_4 FILLER_34_317 ();
 sg13g2_decap_4 FILLER_34_325 ();
 sg13g2_fill_1 FILLER_34_329 ();
 sg13g2_decap_4 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_337 ();
 sg13g2_fill_1 FILLER_34_348 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_fill_2 FILLER_34_364 ();
 sg13g2_fill_1 FILLER_34_370 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_4 FILLER_34_389 ();
 sg13g2_fill_1 FILLER_34_396 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_43 ();
 sg13g2_fill_1 FILLER_35_45 ();
 sg13g2_decap_8 FILLER_35_76 ();
 sg13g2_decap_4 FILLER_35_83 ();
 sg13g2_fill_2 FILLER_35_99 ();
 sg13g2_fill_1 FILLER_35_101 ();
 sg13g2_decap_4 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_116 ();
 sg13g2_fill_1 FILLER_35_122 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_fill_2 FILLER_35_191 ();
 sg13g2_decap_4 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_201 ();
 sg13g2_fill_2 FILLER_35_206 ();
 sg13g2_fill_1 FILLER_35_208 ();
 sg13g2_decap_8 FILLER_35_219 ();
 sg13g2_decap_4 FILLER_35_226 ();
 sg13g2_fill_1 FILLER_35_251 ();
 sg13g2_fill_1 FILLER_35_279 ();
 sg13g2_fill_1 FILLER_35_315 ();
 sg13g2_fill_2 FILLER_35_326 ();
 sg13g2_fill_1 FILLER_35_363 ();
 sg13g2_fill_2 FILLER_35_369 ();
 sg13g2_fill_1 FILLER_35_371 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_30 ();
 sg13g2_decap_8 FILLER_36_41 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_77 ();
 sg13g2_fill_1 FILLER_36_79 ();
 sg13g2_decap_8 FILLER_36_100 ();
 sg13g2_fill_1 FILLER_36_107 ();
 sg13g2_decap_8 FILLER_36_122 ();
 sg13g2_fill_2 FILLER_36_129 ();
 sg13g2_fill_2 FILLER_36_135 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_decap_4 FILLER_36_145 ();
 sg13g2_decap_8 FILLER_36_152 ();
 sg13g2_decap_8 FILLER_36_159 ();
 sg13g2_fill_2 FILLER_36_166 ();
 sg13g2_fill_2 FILLER_36_171 ();
 sg13g2_fill_1 FILLER_36_173 ();
 sg13g2_fill_2 FILLER_36_177 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_fill_2 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_228 ();
 sg13g2_decap_4 FILLER_36_235 ();
 sg13g2_decap_8 FILLER_36_248 ();
 sg13g2_decap_8 FILLER_36_255 ();
 sg13g2_decap_4 FILLER_36_262 ();
 sg13g2_fill_2 FILLER_36_266 ();
 sg13g2_decap_4 FILLER_36_276 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_decap_4 FILLER_36_293 ();
 sg13g2_fill_2 FILLER_36_297 ();
 sg13g2_fill_2 FILLER_36_303 ();
 sg13g2_fill_1 FILLER_36_305 ();
 sg13g2_fill_2 FILLER_36_309 ();
 sg13g2_decap_8 FILLER_36_314 ();
 sg13g2_decap_8 FILLER_36_321 ();
 sg13g2_fill_1 FILLER_36_328 ();
 sg13g2_fill_2 FILLER_36_357 ();
 sg13g2_fill_1 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_363 ();
 sg13g2_decap_4 FILLER_36_370 ();
 sg13g2_fill_2 FILLER_36_386 ();
 sg13g2_fill_1 FILLER_36_388 ();
 sg13g2_fill_2 FILLER_36_392 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_4 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_19 ();
 sg13g2_fill_1 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_51 ();
 sg13g2_decap_8 FILLER_37_72 ();
 sg13g2_fill_1 FILLER_37_79 ();
 sg13g2_fill_2 FILLER_37_96 ();
 sg13g2_fill_2 FILLER_37_120 ();
 sg13g2_decap_8 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_244 ();
 sg13g2_decap_8 FILLER_37_284 ();
 sg13g2_fill_2 FILLER_37_291 ();
 sg13g2_fill_1 FILLER_37_293 ();
 sg13g2_fill_1 FILLER_37_332 ();
 sg13g2_fill_2 FILLER_37_368 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_4 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_25 ();
 sg13g2_fill_1 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_68 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_fill_1 FILLER_38_154 ();
 sg13g2_fill_1 FILLER_38_167 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_fill_2 FILLER_38_184 ();
 sg13g2_decap_8 FILLER_38_190 ();
 sg13g2_decap_8 FILLER_38_197 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_fill_1 FILLER_38_208 ();
 sg13g2_decap_4 FILLER_38_221 ();
 sg13g2_fill_1 FILLER_38_225 ();
 sg13g2_decap_8 FILLER_38_230 ();
 sg13g2_decap_8 FILLER_38_237 ();
 sg13g2_fill_2 FILLER_38_244 ();
 sg13g2_fill_1 FILLER_38_246 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_fill_2 FILLER_38_277 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_333 ();
 sg13g2_fill_2 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_360 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_decap_4 FILLER_38_384 ();
 sg13g2_fill_2 FILLER_38_388 ();
 sg13g2_decap_4 FILLER_38_394 ();
 sg13g2_fill_1 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net249;
 assign uio_oe[1] = net250;
 assign uio_oe[2] = net251;
 assign uio_oe[3] = net252;
 assign uio_oe[4] = net253;
 assign uio_oe[5] = net254;
 assign uio_oe[6] = net255;
 assign uio_oe[7] = net256;
 assign uio_out[0] = net257;
 assign uio_out[1] = net258;
 assign uio_out[2] = net259;
 assign uio_out[3] = net260;
 assign uio_out[4] = net261;
 assign uio_out[5] = net262;
 assign uio_out[6] = net263;
 assign uio_out[7] = net264;
endmodule

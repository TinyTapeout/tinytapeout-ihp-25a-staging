module tt_um_nomuwill (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire clknet_0_clk;
 wire \izh_1.spike ;
 wire \izh_1.u[0] ;
 wire \izh_1.u[10] ;
 wire \izh_1.u[11] ;
 wire \izh_1.u[12] ;
 wire \izh_1.u[13] ;
 wire \izh_1.u[14] ;
 wire \izh_1.u[1] ;
 wire \izh_1.u[2] ;
 wire \izh_1.u[3] ;
 wire \izh_1.u[4] ;
 wire \izh_1.u[5] ;
 wire \izh_1.u[6] ;
 wire \izh_1.u[7] ;
 wire \izh_1.u[8] ;
 wire \izh_1.u[9] ;
 wire \izh_2.spike ;
 wire \izh_2.u[0] ;
 wire \izh_2.u[10] ;
 wire \izh_2.u[11] ;
 wire \izh_2.u[12] ;
 wire \izh_2.u[13] ;
 wire \izh_2.u[14] ;
 wire \izh_2.u[1] ;
 wire \izh_2.u[2] ;
 wire \izh_2.u[3] ;
 wire \izh_2.u[4] ;
 wire \izh_2.u[5] ;
 wire \izh_2.u[6] ;
 wire \izh_2.u[7] ;
 wire \izh_2.u[8] ;
 wire \izh_2.u[9] ;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;

 sg13g2_inv_1 _0971_ (.Y(_0084_),
    .A(\izh_1.u[3] ));
 sg13g2_inv_1 _0972_ (.Y(_0085_),
    .A(\izh_1.u[2] ));
 sg13g2_inv_1 _0973_ (.Y(_0086_),
    .A(\izh_2.u[3] ));
 sg13g2_inv_2 _0974_ (.Y(_0087_),
    .A(uo_out[2]));
 sg13g2_inv_1 _0975_ (.Y(_0088_),
    .A(uo_out[4]));
 sg13g2_inv_1 _0976_ (.Y(_0089_),
    .A(net208));
 sg13g2_inv_1 _0977_ (.Y(_0090_),
    .A(net200));
 sg13g2_inv_1 _0978_ (.Y(_0091_),
    .A(net248));
 sg13g2_inv_1 _0979_ (.Y(_0092_),
    .A(net230));
 sg13g2_inv_1 _0980_ (.Y(_0093_),
    .A(_0008_));
 sg13g2_inv_1 _0981_ (.Y(_0094_),
    .A(_0014_));
 sg13g2_inv_1 _0982_ (.Y(_0095_),
    .A(net95));
 sg13g2_inv_1 _0983_ (.Y(_0096_),
    .A(\izh_1.u[10] ));
 sg13g2_inv_1 _0984_ (.Y(_0097_),
    .A(net63));
 sg13g2_inv_1 _0985_ (.Y(_0098_),
    .A(\izh_1.u[12] ));
 sg13g2_inv_1 _0986_ (.Y(_0099_),
    .A(_0030_));
 sg13g2_inv_1 _0987_ (.Y(_0100_),
    .A(net93));
 sg13g2_nand2_2 _0988_ (.Y(_0101_),
    .A(net202),
    .B(net209));
 sg13g2_and2_2 _0989_ (.A(net202),
    .B(net200),
    .X(_0102_));
 sg13g2_nand2_1 _0990_ (.Y(_0103_),
    .A(net202),
    .B(net200));
 sg13g2_nand2_1 _0991_ (.Y(_0104_),
    .A(net208),
    .B(_0102_));
 sg13g2_inv_2 _0992_ (.Y(\izh_1.spike ),
    .A(net195));
 sg13g2_and2_1 _0993_ (.A(net224),
    .B(net230),
    .X(_0105_));
 sg13g2_and2_2 _0994_ (.A(net224),
    .B(net222),
    .X(_0106_));
 sg13g2_nand2_1 _0995_ (.Y(_0107_),
    .A(net225),
    .B(uio_oe[6]));
 sg13g2_nand2_1 _0996_ (.Y(_0108_),
    .A(net230),
    .B(_0106_));
 sg13g2_inv_2 _0997_ (.Y(\izh_2.spike ),
    .A(net193));
 sg13g2_and2_1 _0998_ (.A(uio_oe[7]),
    .B(net221),
    .X(_0109_));
 sg13g2_nor2_1 _0999_ (.A(uio_oe[4]),
    .B(net224),
    .Y(_0110_));
 sg13g2_and2_2 _1000_ (.A(net233),
    .B(net228),
    .X(_0111_));
 sg13g2_nand2_1 _1001_ (.Y(_0112_),
    .A(net233),
    .B(net228));
 sg13g2_xnor2_1 _1002_ (.Y(_0113_),
    .A(net232),
    .B(net228));
 sg13g2_a21oi_1 _1003_ (.A1(net240),
    .A2(uio_oe[0]),
    .Y(_0114_),
    .B1(net238));
 sg13g2_a21oi_1 _1004_ (.A1(net240),
    .A2(net235),
    .Y(_0115_),
    .B1(net232));
 sg13g2_and2_2 _1005_ (.A(net234),
    .B(net236),
    .X(_0116_));
 sg13g2_nand2_1 _1006_ (.Y(_0117_),
    .A(net233),
    .B(net238));
 sg13g2_nor2_1 _1007_ (.A(_0114_),
    .B(_0115_),
    .Y(_0118_));
 sg13g2_nand2b_1 _1008_ (.Y(_0119_),
    .B(_0118_),
    .A_N(_0113_));
 sg13g2_o21ai_1 _1009_ (.B1(net228),
    .Y(_0120_),
    .A1(net233),
    .A2(net224));
 sg13g2_o21ai_1 _1010_ (.B1(_0120_),
    .Y(_0121_),
    .A1(_0110_),
    .A2(_0119_));
 sg13g2_xor2_1 _1011_ (.B(net222),
    .A(uio_oe[5]),
    .X(_0122_));
 sg13g2_a21o_1 _1012_ (.A2(_0122_),
    .A1(_0121_),
    .B1(_0106_),
    .X(_0123_));
 sg13g2_o21ai_1 _1013_ (.B1(net230),
    .Y(_0124_),
    .A1(net222),
    .A2(_0123_));
 sg13g2_nor2_1 _1014_ (.A(_0094_),
    .B(_0124_),
    .Y(_0125_));
 sg13g2_a21o_1 _1015_ (.A2(_0123_),
    .A1(net222),
    .B1(net230),
    .X(_0126_));
 sg13g2_nand2_1 _1016_ (.Y(_0127_),
    .A(_0124_),
    .B(_0126_));
 sg13g2_or2_1 _1017_ (.X(_0128_),
    .B(_0127_),
    .A(\izh_2.u[11] ));
 sg13g2_xor2_1 _1018_ (.B(net222),
    .A(net230),
    .X(_0129_));
 sg13g2_xnor2_1 _1019_ (.Y(_0130_),
    .A(_0123_),
    .B(_0129_));
 sg13g2_nor2_1 _1020_ (.A(\izh_2.u[10] ),
    .B(_0130_),
    .Y(_0131_));
 sg13g2_xor2_1 _1021_ (.B(_0122_),
    .A(_0121_),
    .X(_0132_));
 sg13g2_nand2_1 _1022_ (.Y(_0133_),
    .A(_0011_),
    .B(_0132_));
 sg13g2_xnor2_1 _1023_ (.Y(_0134_),
    .A(net228),
    .B(net224));
 sg13g2_nand2_1 _1024_ (.Y(_0135_),
    .A(_0112_),
    .B(_0119_));
 sg13g2_xnor2_1 _1025_ (.Y(_0136_),
    .A(_0134_),
    .B(_0135_));
 sg13g2_nor2b_1 _1026_ (.A(\izh_2.u[8] ),
    .B_N(_0136_),
    .Y(_0137_));
 sg13g2_xnor2_1 _1027_ (.Y(_0138_),
    .A(_0113_),
    .B(_0118_));
 sg13g2_nand2_1 _1028_ (.Y(_0139_),
    .A(_0009_),
    .B(_0138_));
 sg13g2_o21ai_1 _1029_ (.B1(net240),
    .Y(_0140_),
    .A1(uio_oe[0]),
    .A2(net235));
 sg13g2_xor2_1 _1030_ (.B(net235),
    .A(net232),
    .X(_0141_));
 sg13g2_xnor2_1 _1031_ (.Y(_0142_),
    .A(_0140_),
    .B(_0141_));
 sg13g2_nand2b_1 _1032_ (.Y(_0143_),
    .B(_0142_),
    .A_N(\izh_2.u[6] ));
 sg13g2_nand2_1 _1033_ (.Y(_0144_),
    .A(uio_oe[0]),
    .B(net235));
 sg13g2_xnor2_1 _1034_ (.Y(_0145_),
    .A(net240),
    .B(net235));
 sg13g2_o21ai_1 _1035_ (.B1(_0144_),
    .Y(_0146_),
    .A1(uio_oe[0]),
    .A2(_0145_));
 sg13g2_nand2_1 _1036_ (.Y(_0147_),
    .A(_0005_),
    .B(_0146_));
 sg13g2_xnor2_1 _1037_ (.Y(_0148_),
    .A(net240),
    .B(uio_oe[0]));
 sg13g2_nor2_1 _1038_ (.A(\izh_2.u[4] ),
    .B(_0148_),
    .Y(_0149_));
 sg13g2_xor2_1 _1039_ (.B(_0148_),
    .A(_0006_),
    .X(_0150_));
 sg13g2_nor2_1 _1040_ (.A(\izh_2.u[1] ),
    .B(\izh_2.u[0] ),
    .Y(_0151_));
 sg13g2_a22oi_1 _1041_ (.Y(_0152_),
    .B1(_0007_),
    .B2(_0151_),
    .A2(uio_oe[0]),
    .A1(_0086_));
 sg13g2_nor2_1 _1042_ (.A(_0086_),
    .B(uio_oe[0]),
    .Y(_0153_));
 sg13g2_nor3_1 _1043_ (.A(_0150_),
    .B(_0152_),
    .C(_0153_),
    .Y(_0154_));
 sg13g2_xnor2_1 _1044_ (.Y(_0155_),
    .A(\izh_2.u[5] ),
    .B(_0146_));
 sg13g2_o21ai_1 _1045_ (.B1(_0155_),
    .Y(_0156_),
    .A1(_0149_),
    .A2(_0154_));
 sg13g2_xnor2_1 _1046_ (.Y(_0157_),
    .A(_0004_),
    .B(_0142_));
 sg13g2_a21o_1 _1047_ (.A2(_0156_),
    .A1(_0147_),
    .B1(_0157_),
    .X(_0158_));
 sg13g2_xor2_1 _1048_ (.B(_0138_),
    .A(\izh_2.u[7] ),
    .X(_0159_));
 sg13g2_a21o_1 _1049_ (.A2(_0158_),
    .A1(_0143_),
    .B1(_0159_),
    .X(_0160_));
 sg13g2_xnor2_1 _1050_ (.Y(_0161_),
    .A(_0008_),
    .B(_0136_));
 sg13g2_a21oi_1 _1051_ (.A1(_0139_),
    .A2(_0160_),
    .Y(_0162_),
    .B1(_0161_));
 sg13g2_xnor2_1 _1052_ (.Y(_0163_),
    .A(\izh_2.u[9] ),
    .B(_0132_));
 sg13g2_o21ai_1 _1053_ (.B1(_0163_),
    .Y(_0164_),
    .A1(_0137_),
    .A2(_0162_));
 sg13g2_nand2_1 _1054_ (.Y(_0165_),
    .A(_0133_),
    .B(_0164_));
 sg13g2_xnor2_1 _1055_ (.Y(_0166_),
    .A(_0010_),
    .B(_0130_));
 sg13g2_a21oi_1 _1056_ (.A1(_0165_),
    .A2(_0166_),
    .Y(_0167_),
    .B1(_0131_));
 sg13g2_xor2_1 _1057_ (.B(_0127_),
    .A(_0012_),
    .X(_0168_));
 sg13g2_o21ai_1 _1058_ (.B1(_0128_),
    .Y(_0169_),
    .A1(_0167_),
    .A2(_0168_));
 sg13g2_xor2_1 _1059_ (.B(_0124_),
    .A(\izh_2.u[12] ),
    .X(_0170_));
 sg13g2_a21o_1 _1060_ (.A2(_0170_),
    .A1(_0169_),
    .B1(_0125_),
    .X(_0171_));
 sg13g2_nor2b_1 _1061_ (.A(\izh_2.u[13] ),
    .B_N(_0171_),
    .Y(_0172_));
 sg13g2_xnor2_1 _1062_ (.Y(_0173_),
    .A(\izh_2.u[14] ),
    .B(_0172_));
 sg13g2_xor2_1 _1063_ (.B(_0171_),
    .A(_0013_),
    .X(_0174_));
 sg13g2_nand2_1 _1064_ (.Y(_0175_),
    .A(\izh_2.u[7] ),
    .B(_0174_));
 sg13g2_xnor2_1 _1065_ (.Y(_0176_),
    .A(_0169_),
    .B(_0170_));
 sg13g2_nor2_1 _1066_ (.A(_0004_),
    .B(_0176_),
    .Y(_0177_));
 sg13g2_xor2_1 _1067_ (.B(_0168_),
    .A(_0167_),
    .X(_0178_));
 sg13g2_nand2_1 _1068_ (.Y(_0179_),
    .A(\izh_2.u[5] ),
    .B(_0178_));
 sg13g2_xnor2_1 _1069_ (.Y(_0180_),
    .A(_0165_),
    .B(_0166_));
 sg13g2_nor2_1 _1070_ (.A(_0006_),
    .B(_0180_),
    .Y(_0181_));
 sg13g2_or3_1 _1071_ (.A(_0137_),
    .B(_0162_),
    .C(_0163_),
    .X(_0182_));
 sg13g2_and2_1 _1072_ (.A(_0164_),
    .B(_0182_),
    .X(_0183_));
 sg13g2_nand2_1 _1073_ (.Y(_0184_),
    .A(\izh_2.u[3] ),
    .B(_0183_));
 sg13g2_nand3_1 _1074_ (.B(_0160_),
    .C(_0161_),
    .A(_0139_),
    .Y(_0185_));
 sg13g2_nand2b_1 _1075_ (.Y(_0186_),
    .B(_0185_),
    .A_N(_0162_));
 sg13g2_nor2_1 _1076_ (.A(_0007_),
    .B(_0186_),
    .Y(_0187_));
 sg13g2_nand3_1 _1077_ (.B(_0158_),
    .C(_0159_),
    .A(_0143_),
    .Y(_0188_));
 sg13g2_nand3_1 _1078_ (.B(_0160_),
    .C(_0188_),
    .A(\izh_2.u[1] ),
    .Y(_0189_));
 sg13g2_nand3_1 _1079_ (.B(_0156_),
    .C(_0157_),
    .A(_0147_),
    .Y(_0190_));
 sg13g2_and2_1 _1080_ (.A(_0158_),
    .B(_0190_),
    .X(_0191_));
 sg13g2_nand2_1 _1081_ (.Y(_0192_),
    .A(net106),
    .B(_0191_));
 sg13g2_a21o_1 _1082_ (.A2(_0188_),
    .A1(_0160_),
    .B1(\izh_2.u[1] ),
    .X(_0193_));
 sg13g2_nand2_1 _1083_ (.Y(_0194_),
    .A(_0189_),
    .B(_0193_));
 sg13g2_o21ai_1 _1084_ (.B1(_0189_),
    .Y(_0195_),
    .A1(_0192_),
    .A2(_0194_));
 sg13g2_xnor2_1 _1085_ (.Y(_0196_),
    .A(net65),
    .B(_0186_));
 sg13g2_a21oi_1 _1086_ (.A1(_0195_),
    .A2(_0196_),
    .Y(_0197_),
    .B1(_0187_));
 sg13g2_xnor2_1 _1087_ (.Y(_0198_),
    .A(\izh_2.u[3] ),
    .B(_0183_));
 sg13g2_o21ai_1 _1088_ (.B1(_0184_),
    .Y(_0199_),
    .A1(_0197_),
    .A2(_0198_));
 sg13g2_xnor2_1 _1089_ (.Y(_0200_),
    .A(net72),
    .B(_0180_));
 sg13g2_a21oi_1 _1090_ (.A1(_0199_),
    .A2(_0200_),
    .Y(_0201_),
    .B1(_0181_));
 sg13g2_xor2_1 _1091_ (.B(_0178_),
    .A(_0005_),
    .X(_0202_));
 sg13g2_o21ai_1 _1092_ (.B1(_0179_),
    .Y(_0203_),
    .A1(_0201_),
    .A2(_0202_));
 sg13g2_xnor2_1 _1093_ (.Y(_0204_),
    .A(\izh_2.u[6] ),
    .B(_0176_));
 sg13g2_a21oi_2 _1094_ (.B1(_0177_),
    .Y(_0205_),
    .A2(_0204_),
    .A1(_0203_));
 sg13g2_xor2_1 _1095_ (.B(_0174_),
    .A(_0009_),
    .X(_0206_));
 sg13g2_o21ai_1 _1096_ (.B1(_0175_),
    .Y(_0207_),
    .A1(_0205_),
    .A2(_0206_));
 sg13g2_xor2_1 _1097_ (.B(_0173_),
    .A(net66),
    .X(_0208_));
 sg13g2_a22oi_1 _1098_ (.Y(_0209_),
    .B1(_0207_),
    .B2(_0208_),
    .A2(_0173_),
    .A1(_0093_));
 sg13g2_a21oi_1 _1099_ (.A1(net193),
    .A2(_0209_),
    .Y(_0210_),
    .B1(net61));
 sg13g2_and3_1 _1100_ (.X(_0211_),
    .A(net61),
    .B(net193),
    .C(_0209_));
 sg13g2_nor3_1 _1101_ (.A(net243),
    .B(net62),
    .C(_0211_),
    .Y(_0031_));
 sg13g2_nor2_2 _1102_ (.A(net61),
    .B(_0209_),
    .Y(_0212_));
 sg13g2_xor2_1 _1103_ (.B(_0212_),
    .A(net73),
    .X(_0213_));
 sg13g2_nand2_1 _1104_ (.Y(_0214_),
    .A(\izh_2.u[9] ),
    .B(\izh_2.u[10] ));
 sg13g2_xor2_1 _1105_ (.B(\izh_2.u[10] ),
    .A(\izh_2.u[9] ),
    .X(_0215_));
 sg13g2_o21ai_1 _1106_ (.B1(net245),
    .Y(_0216_),
    .A1(net193),
    .A2(_0215_));
 sg13g2_a21oi_1 _1107_ (.A1(net193),
    .A2(_0213_),
    .Y(_0032_),
    .B1(_0216_));
 sg13g2_a21oi_1 _1108_ (.A1(\izh_2.u[10] ),
    .A2(_0212_),
    .Y(_0217_),
    .B1(net101));
 sg13g2_and3_1 _1109_ (.X(_0218_),
    .A(\izh_2.u[10] ),
    .B(\izh_2.u[11] ),
    .C(_0212_));
 sg13g2_nor3_1 _1110_ (.A(\izh_2.spike ),
    .B(net102),
    .C(_0218_),
    .Y(_0219_));
 sg13g2_xnor2_1 _1111_ (.Y(_0220_),
    .A(_0012_),
    .B(_0214_));
 sg13g2_a21oi_1 _1112_ (.A1(\izh_2.spike ),
    .A2(_0220_),
    .Y(_0221_),
    .B1(_0219_));
 sg13g2_nor2_1 _1113_ (.A(net243),
    .B(net103),
    .Y(_0033_));
 sg13g2_nand3_1 _1114_ (.B(\izh_2.spike ),
    .C(_0214_),
    .A(_0012_),
    .Y(_0222_));
 sg13g2_o21ai_1 _1115_ (.B1(_0222_),
    .Y(_0223_),
    .A1(\izh_2.spike ),
    .A2(_0218_));
 sg13g2_o21ai_1 _1116_ (.B1(net246),
    .Y(_0224_),
    .A1(net59),
    .A2(_0223_));
 sg13g2_a21oi_1 _1117_ (.A1(net59),
    .A2(_0223_),
    .Y(_0034_),
    .B1(_0224_));
 sg13g2_and4_1 _1118_ (.A(\izh_2.u[10] ),
    .B(\izh_2.u[11] ),
    .C(\izh_2.u[12] ),
    .D(_0212_),
    .X(_0225_));
 sg13g2_a21oi_1 _1119_ (.A1(\izh_2.u[13] ),
    .A2(_0225_),
    .Y(_0226_),
    .B1(\izh_2.spike ));
 sg13g2_o21ai_1 _1120_ (.B1(_0226_),
    .Y(_0227_),
    .A1(\izh_2.u[13] ),
    .A2(_0225_));
 sg13g2_nand2b_1 _1121_ (.Y(_0228_),
    .B(_0214_),
    .A_N(\izh_2.u[11] ));
 sg13g2_nand2_1 _1122_ (.Y(_0229_),
    .A(\izh_2.u[12] ),
    .B(_0228_));
 sg13g2_inv_1 _1123_ (.Y(_0230_),
    .A(_0229_));
 sg13g2_a21oi_1 _1124_ (.A1(net88),
    .A2(_0229_),
    .Y(_0231_),
    .B1(net193));
 sg13g2_o21ai_1 _1125_ (.B1(_0231_),
    .Y(_0232_),
    .A1(net88),
    .A2(_0229_));
 sg13g2_a21oi_1 _1126_ (.A1(_0227_),
    .A2(net89),
    .Y(_0035_),
    .B1(net243));
 sg13g2_a21oi_1 _1127_ (.A1(\izh_2.u[13] ),
    .A2(_0230_),
    .Y(_0233_),
    .B1(net194));
 sg13g2_or3_1 _1128_ (.A(_0095_),
    .B(_0226_),
    .C(_0233_),
    .X(_0234_));
 sg13g2_o21ai_1 _1129_ (.B1(_0095_),
    .Y(_0235_),
    .A1(_0226_),
    .A2(_0233_));
 sg13g2_and3_1 _1130_ (.X(_0036_),
    .A(net246),
    .B(_0234_),
    .C(net96));
 sg13g2_xor2_1 _1131_ (.B(net200),
    .A(net202),
    .X(_0236_));
 sg13g2_nand2_1 _1132_ (.Y(_0237_),
    .A(net206),
    .B(net202));
 sg13g2_nor2_1 _1133_ (.A(net206),
    .B(net202),
    .Y(_0238_));
 sg13g2_xnor2_1 _1134_ (.Y(_0239_),
    .A(net211),
    .B(net206));
 sg13g2_a21oi_1 _1135_ (.A1(net216),
    .A2(net220),
    .Y(_0240_),
    .B1(net215));
 sg13g2_and2_1 _1136_ (.A(uo_out[1]),
    .B(uo_out[3]),
    .X(_0241_));
 sg13g2_nand3_1 _1137_ (.B(net220),
    .C(net211),
    .A(net216),
    .Y(_0242_));
 sg13g2_o21ai_1 _1138_ (.B1(net215),
    .Y(_0243_),
    .A1(net217),
    .A2(net211));
 sg13g2_a21oi_1 _1139_ (.A1(_0242_),
    .A2(_0243_),
    .Y(_0244_),
    .B1(_0239_));
 sg13g2_a21oi_1 _1140_ (.A1(net211),
    .A2(net206),
    .Y(_0245_),
    .B1(_0244_));
 sg13g2_a21oi_1 _1141_ (.A1(_0237_),
    .A2(_0245_),
    .Y(_0246_),
    .B1(_0238_));
 sg13g2_a21oi_1 _1142_ (.A1(_0236_),
    .A2(_0246_),
    .Y(_0247_),
    .B1(_0102_));
 sg13g2_a21oi_1 _1143_ (.A1(_0089_),
    .A2(_0090_),
    .Y(_0248_),
    .B1(_0247_));
 sg13g2_o21ai_1 _1144_ (.B1(net208),
    .Y(_0249_),
    .A1(net200),
    .A2(_0248_));
 sg13g2_nor2_1 _1145_ (.A(_0099_),
    .B(_0249_),
    .Y(_0250_));
 sg13g2_o21ai_1 _1146_ (.B1(_0249_),
    .Y(_0251_),
    .A1(net208),
    .A2(_0248_));
 sg13g2_or2_1 _1147_ (.X(_0252_),
    .B(_0251_),
    .A(\izh_1.u[11] ));
 sg13g2_xor2_1 _1148_ (.B(net200),
    .A(net208),
    .X(_0253_));
 sg13g2_xnor2_1 _1149_ (.Y(_0254_),
    .A(_0247_),
    .B(_0253_));
 sg13g2_xor2_1 _1150_ (.B(_0246_),
    .A(_0236_),
    .X(_0255_));
 sg13g2_xor2_1 _1151_ (.B(net202),
    .A(net206),
    .X(_0256_));
 sg13g2_xnor2_1 _1152_ (.Y(_0257_),
    .A(_0245_),
    .B(_0256_));
 sg13g2_nor2b_1 _1153_ (.A(\izh_1.u[8] ),
    .B_N(_0257_),
    .Y(_0258_));
 sg13g2_inv_1 _1154_ (.Y(_0259_),
    .A(_0258_));
 sg13g2_nand3_1 _1155_ (.B(_0242_),
    .C(_0243_),
    .A(_0239_),
    .Y(_0260_));
 sg13g2_nor2b_2 _1156_ (.A(_0244_),
    .B_N(_0260_),
    .Y(_0261_));
 sg13g2_nand2_1 _1157_ (.Y(_0262_),
    .A(_0025_),
    .B(_0261_));
 sg13g2_a21oi_1 _1158_ (.A1(net216),
    .A2(net215),
    .Y(_0263_),
    .B1(_0240_));
 sg13g2_xnor2_1 _1159_ (.Y(_0264_),
    .A(net211),
    .B(_0263_));
 sg13g2_or2_1 _1160_ (.X(_0265_),
    .B(_0264_),
    .A(\izh_1.u[6] ));
 sg13g2_nand2_1 _1161_ (.Y(_0266_),
    .A(net220),
    .B(net215));
 sg13g2_xnor2_1 _1162_ (.Y(_0267_),
    .A(net217),
    .B(net215));
 sg13g2_o21ai_1 _1163_ (.B1(_0266_),
    .Y(_0268_),
    .A1(net220),
    .A2(_0267_));
 sg13g2_nand2_1 _1164_ (.Y(_0269_),
    .A(_0021_),
    .B(_0268_));
 sg13g2_xor2_1 _1165_ (.B(net220),
    .A(net217),
    .X(_0270_));
 sg13g2_nor2b_1 _1166_ (.A(\izh_1.u[4] ),
    .B_N(_0270_),
    .Y(_0271_));
 sg13g2_xnor2_1 _1167_ (.Y(_0272_),
    .A(_0022_),
    .B(_0270_));
 sg13g2_nor2_1 _1168_ (.A(_0084_),
    .B(net220),
    .Y(_0273_));
 sg13g2_nor2_1 _1169_ (.A(\izh_1.u[1] ),
    .B(\izh_1.u[0] ),
    .Y(_0274_));
 sg13g2_a22oi_1 _1170_ (.Y(_0275_),
    .B1(_0023_),
    .B2(_0274_),
    .A2(net218),
    .A1(_0084_));
 sg13g2_nor3_1 _1171_ (.A(_0272_),
    .B(_0273_),
    .C(_0275_),
    .Y(_0276_));
 sg13g2_xnor2_1 _1172_ (.Y(_0277_),
    .A(\izh_1.u[5] ),
    .B(_0268_));
 sg13g2_o21ai_1 _1173_ (.B1(_0277_),
    .Y(_0278_),
    .A1(_0271_),
    .A2(_0276_));
 sg13g2_xor2_1 _1174_ (.B(_0264_),
    .A(_0020_),
    .X(_0279_));
 sg13g2_a21o_1 _1175_ (.A2(_0278_),
    .A1(_0269_),
    .B1(_0279_),
    .X(_0280_));
 sg13g2_xor2_1 _1176_ (.B(_0261_),
    .A(\izh_1.u[7] ),
    .X(_0281_));
 sg13g2_a21o_2 _1177_ (.A2(_0280_),
    .A1(_0265_),
    .B1(_0281_),
    .X(_0282_));
 sg13g2_xnor2_1 _1178_ (.Y(_0283_),
    .A(_0024_),
    .B(_0257_));
 sg13g2_a21o_2 _1179_ (.A2(_0282_),
    .A1(_0262_),
    .B1(_0283_),
    .X(_0284_));
 sg13g2_xnor2_1 _1180_ (.Y(_0285_),
    .A(\izh_1.u[9] ),
    .B(_0255_));
 sg13g2_inv_1 _1181_ (.Y(_0286_),
    .A(_0285_));
 sg13g2_a21oi_2 _1182_ (.B1(_0286_),
    .Y(_0287_),
    .A2(_0284_),
    .A1(_0259_));
 sg13g2_a21o_1 _1183_ (.A2(_0255_),
    .A1(_0027_),
    .B1(_0287_),
    .X(_0288_));
 sg13g2_xor2_1 _1184_ (.B(_0254_),
    .A(_0026_),
    .X(_0289_));
 sg13g2_a22oi_1 _1185_ (.Y(_0290_),
    .B1(_0288_),
    .B2(_0289_),
    .A2(_0254_),
    .A1(_0096_));
 sg13g2_xor2_1 _1186_ (.B(_0251_),
    .A(_0028_),
    .X(_0291_));
 sg13g2_o21ai_1 _1187_ (.B1(_0252_),
    .Y(_0292_),
    .A1(_0290_),
    .A2(_0291_));
 sg13g2_xnor2_1 _1188_ (.Y(_0293_),
    .A(_0098_),
    .B(_0249_));
 sg13g2_a21o_1 _1189_ (.A2(_0293_),
    .A1(_0292_),
    .B1(_0250_),
    .X(_0294_));
 sg13g2_nor2b_1 _1190_ (.A(\izh_1.u[13] ),
    .B_N(_0294_),
    .Y(_0295_));
 sg13g2_xnor2_1 _1191_ (.Y(_0296_),
    .A(\izh_1.u[14] ),
    .B(_0295_));
 sg13g2_nand2b_1 _1192_ (.Y(_0297_),
    .B(_0296_),
    .A_N(_0024_));
 sg13g2_xor2_1 _1193_ (.B(_0294_),
    .A(_0029_),
    .X(_0298_));
 sg13g2_xnor2_1 _1194_ (.Y(_0299_),
    .A(_0292_),
    .B(_0293_));
 sg13g2_or2_1 _1195_ (.X(_0300_),
    .B(_0299_),
    .A(_0020_));
 sg13g2_xor2_1 _1196_ (.B(_0291_),
    .A(_0290_),
    .X(_0301_));
 sg13g2_xnor2_1 _1197_ (.Y(_0302_),
    .A(_0288_),
    .B(_0289_));
 sg13g2_or2_1 _1198_ (.X(_0303_),
    .B(_0302_),
    .A(_0022_));
 sg13g2_and3_1 _1199_ (.X(_0304_),
    .A(_0259_),
    .B(_0284_),
    .C(_0286_));
 sg13g2_nor3_1 _1200_ (.A(_0084_),
    .B(_0287_),
    .C(_0304_),
    .Y(_0305_));
 sg13g2_nand3_1 _1201_ (.B(_0282_),
    .C(_0283_),
    .A(_0262_),
    .Y(_0306_));
 sg13g2_nand3b_1 _1202_ (.B(_0284_),
    .C(_0306_),
    .Y(_0307_),
    .A_N(_0023_));
 sg13g2_nand3_1 _1203_ (.B(_0280_),
    .C(_0281_),
    .A(_0265_),
    .Y(_0308_));
 sg13g2_nand3_1 _1204_ (.B(_0282_),
    .C(_0308_),
    .A(\izh_1.u[1] ),
    .Y(_0309_));
 sg13g2_nand3_1 _1205_ (.B(_0278_),
    .C(_0279_),
    .A(_0269_),
    .Y(_0310_));
 sg13g2_and2_1 _1206_ (.A(_0280_),
    .B(_0310_),
    .X(_0311_));
 sg13g2_nand2_1 _1207_ (.Y(_0312_),
    .A(\izh_1.u[0] ),
    .B(_0311_));
 sg13g2_a21oi_1 _1208_ (.A1(_0282_),
    .A2(_0308_),
    .Y(_0313_),
    .B1(\izh_1.u[1] ));
 sg13g2_a21o_1 _1209_ (.A2(_0308_),
    .A1(_0282_),
    .B1(\izh_1.u[1] ),
    .X(_0314_));
 sg13g2_nand2_1 _1210_ (.Y(_0315_),
    .A(_0309_),
    .B(_0314_));
 sg13g2_o21ai_1 _1211_ (.B1(_0309_),
    .Y(_0316_),
    .A1(_0312_),
    .A2(_0313_));
 sg13g2_a21oi_1 _1212_ (.A1(_0284_),
    .A2(_0306_),
    .Y(_0317_),
    .B1(_0085_));
 sg13g2_and3_1 _1213_ (.X(_0318_),
    .A(_0085_),
    .B(_0284_),
    .C(_0306_));
 sg13g2_or2_1 _1214_ (.X(_0319_),
    .B(_0318_),
    .A(_0317_));
 sg13g2_o21ai_1 _1215_ (.B1(_0316_),
    .Y(_0320_),
    .A1(_0317_),
    .A2(_0318_));
 sg13g2_o21ai_1 _1216_ (.B1(\izh_1.u[3] ),
    .Y(_0321_),
    .A1(_0287_),
    .A2(_0304_));
 sg13g2_or3_1 _1217_ (.A(\izh_1.u[3] ),
    .B(_0287_),
    .C(_0304_),
    .X(_0322_));
 sg13g2_a22oi_1 _1218_ (.Y(_0323_),
    .B1(_0321_),
    .B2(_0322_),
    .A2(_0320_),
    .A1(_0307_));
 sg13g2_nor2_1 _1219_ (.A(_0305_),
    .B(_0323_),
    .Y(_0324_));
 sg13g2_xor2_1 _1220_ (.B(_0302_),
    .A(net84),
    .X(_0325_));
 sg13g2_o21ai_1 _1221_ (.B1(_0303_),
    .Y(_0326_),
    .A1(_0324_),
    .A2(_0325_));
 sg13g2_xnor2_1 _1222_ (.Y(_0327_),
    .A(_0021_),
    .B(_0301_));
 sg13g2_a22oi_1 _1223_ (.Y(_0328_),
    .B1(_0326_),
    .B2(_0327_),
    .A2(_0301_),
    .A1(\izh_1.u[5] ));
 sg13g2_xor2_1 _1224_ (.B(_0299_),
    .A(net70),
    .X(_0329_));
 sg13g2_o21ai_1 _1225_ (.B1(_0300_),
    .Y(_0330_),
    .A1(_0328_),
    .A2(_0329_));
 sg13g2_xnor2_1 _1226_ (.Y(_0331_),
    .A(_0025_),
    .B(_0298_));
 sg13g2_a22oi_1 _1227_ (.Y(_0332_),
    .B1(_0330_),
    .B2(_0331_),
    .A2(_0298_),
    .A1(\izh_1.u[7] ));
 sg13g2_xnor2_1 _1228_ (.Y(_0333_),
    .A(net69),
    .B(_0296_));
 sg13g2_o21ai_1 _1229_ (.B1(_0297_),
    .Y(_0334_),
    .A1(_0332_),
    .A2(_0333_));
 sg13g2_nand2b_1 _1230_ (.Y(_0335_),
    .B(net195),
    .A_N(_0334_));
 sg13g2_o21ai_1 _1231_ (.B1(net247),
    .Y(_0336_),
    .A1(_0097_),
    .A2(_0335_));
 sg13g2_a21oi_1 _1232_ (.A1(_0097_),
    .A2(_0335_),
    .Y(_0037_),
    .B1(_0336_));
 sg13g2_and2_1 _1233_ (.A(_0097_),
    .B(_0334_),
    .X(_0337_));
 sg13g2_xor2_1 _1234_ (.B(_0337_),
    .A(net78),
    .X(_0338_));
 sg13g2_nand2_1 _1235_ (.Y(_0339_),
    .A(\izh_1.u[9] ),
    .B(\izh_1.u[10] ));
 sg13g2_xor2_1 _1236_ (.B(\izh_1.u[10] ),
    .A(\izh_1.u[9] ),
    .X(_0340_));
 sg13g2_o21ai_1 _1237_ (.B1(net248),
    .Y(_0341_),
    .A1(net195),
    .A2(_0340_));
 sg13g2_a21oi_1 _1238_ (.A1(net195),
    .A2(_0338_),
    .Y(_0038_),
    .B1(_0341_));
 sg13g2_a21oi_1 _1239_ (.A1(\izh_1.u[10] ),
    .A2(_0337_),
    .Y(_0342_),
    .B1(\izh_1.u[11] ));
 sg13g2_nand4_1 _1240_ (.B(_0097_),
    .C(\izh_1.u[11] ),
    .A(\izh_1.u[10] ),
    .Y(_0343_),
    .D(_0334_));
 sg13g2_nand2_1 _1241_ (.Y(_0344_),
    .A(net195),
    .B(_0343_));
 sg13g2_or2_1 _1242_ (.X(_0345_),
    .B(_0344_),
    .A(_0342_));
 sg13g2_xnor2_1 _1243_ (.Y(_0346_),
    .A(net99),
    .B(_0339_));
 sg13g2_nand2_1 _1244_ (.Y(_0347_),
    .A(\izh_1.spike ),
    .B(_0346_));
 sg13g2_a21oi_1 _1245_ (.A1(_0345_),
    .A2(_0347_),
    .Y(_0039_),
    .B1(net244));
 sg13g2_nand3_1 _1246_ (.B(\izh_1.spike ),
    .C(_0339_),
    .A(_0028_),
    .Y(_0348_));
 sg13g2_nand2_1 _1247_ (.Y(_0349_),
    .A(_0344_),
    .B(_0348_));
 sg13g2_o21ai_1 _1248_ (.B1(net248),
    .Y(_0350_),
    .A1(net57),
    .A2(_0349_));
 sg13g2_a21oi_1 _1249_ (.A1(net57),
    .A2(_0349_),
    .Y(_0040_),
    .B1(_0350_));
 sg13g2_nor2_1 _1250_ (.A(_0098_),
    .B(_0343_),
    .Y(_0351_));
 sg13g2_a21oi_1 _1251_ (.A1(\izh_1.u[13] ),
    .A2(_0351_),
    .Y(_0352_),
    .B1(\izh_1.spike ));
 sg13g2_o21ai_1 _1252_ (.B1(_0352_),
    .Y(_0353_),
    .A1(\izh_1.u[13] ),
    .A2(_0351_));
 sg13g2_nand2b_1 _1253_ (.Y(_0354_),
    .B(_0339_),
    .A_N(\izh_1.u[11] ));
 sg13g2_nand2_1 _1254_ (.Y(_0355_),
    .A(\izh_1.u[12] ),
    .B(_0354_));
 sg13g2_inv_1 _1255_ (.Y(_0356_),
    .A(_0355_));
 sg13g2_a21oi_1 _1256_ (.A1(net80),
    .A2(_0355_),
    .Y(_0357_),
    .B1(net195));
 sg13g2_o21ai_1 _1257_ (.B1(_0357_),
    .Y(_0358_),
    .A1(net80),
    .A2(_0355_));
 sg13g2_a21oi_1 _1258_ (.A1(_0353_),
    .A2(net81),
    .Y(_0041_),
    .B1(net244));
 sg13g2_a21oi_1 _1259_ (.A1(\izh_1.u[13] ),
    .A2(_0356_),
    .Y(_0359_),
    .B1(net195));
 sg13g2_or3_1 _1260_ (.A(_0100_),
    .B(_0352_),
    .C(_0359_),
    .X(_0360_));
 sg13g2_o21ai_1 _1261_ (.B1(_0100_),
    .Y(_0361_),
    .A1(_0352_),
    .A2(_0359_));
 sg13g2_and3_1 _1262_ (.X(_0042_),
    .A(net248),
    .B(_0360_),
    .C(net94));
 sg13g2_nand2_2 _1263_ (.Y(_0362_),
    .A(net228),
    .B(net222));
 sg13g2_inv_1 _1264_ (.Y(_0363_),
    .A(_0362_));
 sg13g2_xor2_1 _1265_ (.B(net230),
    .A(uio_oe[5]),
    .X(_0364_));
 sg13g2_xnor2_1 _1266_ (.Y(_0365_),
    .A(_0362_),
    .B(_0364_));
 sg13g2_or2_1 _1267_ (.X(_0366_),
    .B(_0144_),
    .A(_0142_));
 sg13g2_o21ai_1 _1268_ (.B1(uio_oe[1]),
    .Y(_0367_),
    .A1(net235),
    .A2(net226));
 sg13g2_a21oi_1 _1269_ (.A1(net235),
    .A2(net226),
    .Y(_0368_),
    .B1(uio_oe[5]));
 sg13g2_a21oi_2 _1270_ (.B1(net234),
    .Y(_0369_),
    .A2(net227),
    .A1(net236));
 sg13g2_nand2_1 _1271_ (.Y(_0370_),
    .A(uio_oe[3]),
    .B(net225));
 sg13g2_a21o_1 _1272_ (.A2(_0368_),
    .A1(_0367_),
    .B1(_0369_),
    .X(_0371_));
 sg13g2_o21ai_1 _1273_ (.B1(_0371_),
    .Y(_0372_),
    .A1(net226),
    .A2(_0366_));
 sg13g2_o21ai_1 _1274_ (.B1(_0362_),
    .Y(_0373_),
    .A1(net232),
    .A2(uio_oe[5]));
 sg13g2_o21ai_1 _1275_ (.B1(_0372_),
    .Y(_0374_),
    .A1(net226),
    .A2(net222));
 sg13g2_nor2_1 _1276_ (.A(_0373_),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_and2_1 _1277_ (.A(_0365_),
    .B(_0375_),
    .X(_0376_));
 sg13g2_xnor2_1 _1278_ (.Y(_0377_),
    .A(_0365_),
    .B(_0375_));
 sg13g2_nand2_1 _1279_ (.Y(_0378_),
    .A(\izh_2.u[0] ),
    .B(_0377_));
 sg13g2_xor2_1 _1280_ (.B(_0377_),
    .A(net106),
    .X(_0379_));
 sg13g2_and3_1 _1281_ (.X(_0380_),
    .A(net232),
    .B(net236),
    .C(net226));
 sg13g2_nand3_1 _1282_ (.B(net236),
    .C(net227),
    .A(uio_oe[3]),
    .Y(_0381_));
 sg13g2_and3_1 _1283_ (.X(_0382_),
    .A(uio_oe[1]),
    .B(net242),
    .C(_0380_));
 sg13g2_nand2_1 _1284_ (.Y(_0383_),
    .A(net242),
    .B(_0122_));
 sg13g2_nand2_2 _1285_ (.Y(_0384_),
    .A(uio_oe[1]),
    .B(net223));
 sg13g2_or3_1 _1286_ (.A(_0369_),
    .B(_0380_),
    .C(_0384_),
    .X(_0385_));
 sg13g2_o21ai_1 _1287_ (.B1(_0384_),
    .Y(_0386_),
    .A1(_0369_),
    .A2(_0380_));
 sg13g2_nand3_1 _1288_ (.B(_0385_),
    .C(_0386_),
    .A(_0116_),
    .Y(_0387_));
 sg13g2_a21oi_1 _1289_ (.A1(_0385_),
    .A2(_0386_),
    .Y(_0388_),
    .B1(_0116_));
 sg13g2_a21o_1 _1290_ (.A2(_0386_),
    .A1(_0385_),
    .B1(_0116_),
    .X(_0389_));
 sg13g2_and4_1 _1291_ (.A(net242),
    .B(net236),
    .C(net227),
    .D(uio_oe[6]),
    .X(_0390_));
 sg13g2_or2_1 _1292_ (.X(_0391_),
    .B(_0362_),
    .A(_0144_));
 sg13g2_a22oi_1 _1293_ (.Y(_0392_),
    .B1(uio_oe[6]),
    .B2(net242),
    .A2(net227),
    .A1(net236));
 sg13g2_nor2_1 _1294_ (.A(_0390_),
    .B(_0392_),
    .Y(_0393_));
 sg13g2_xnor2_1 _1295_ (.Y(_0394_),
    .A(_0384_),
    .B(_0393_));
 sg13g2_xor2_1 _1296_ (.B(_0393_),
    .A(_0384_),
    .X(_0395_));
 sg13g2_nand3_1 _1297_ (.B(_0389_),
    .C(_0394_),
    .A(_0387_),
    .Y(_0396_));
 sg13g2_a21o_1 _1298_ (.A2(_0389_),
    .A1(_0387_),
    .B1(_0394_),
    .X(_0397_));
 sg13g2_and4_1 _1299_ (.A(uio_oe[1]),
    .B(net226),
    .C(_0396_),
    .D(_0397_),
    .X(_0398_));
 sg13g2_nand4_1 _1300_ (.B(net226),
    .C(_0396_),
    .A(uio_oe[1]),
    .Y(_0399_),
    .D(_0397_));
 sg13g2_a22oi_1 _1301_ (.Y(_0400_),
    .B1(_0396_),
    .B2(_0397_),
    .A2(net227),
    .A1(uio_oe[1]));
 sg13g2_nor2_1 _1302_ (.A(_0398_),
    .B(_0400_),
    .Y(_0401_));
 sg13g2_xnor2_1 _1303_ (.Y(_0402_),
    .A(_0383_),
    .B(_0401_));
 sg13g2_nand2_1 _1304_ (.Y(_0403_),
    .A(net242),
    .B(net226));
 sg13g2_nor3_1 _1305_ (.A(net240),
    .B(_0366_),
    .C(_0403_),
    .Y(_0404_));
 sg13g2_o21ai_1 _1306_ (.B1(net240),
    .Y(_0405_),
    .A1(net232),
    .A2(net235));
 sg13g2_a21oi_1 _1307_ (.A1(_0117_),
    .A2(_0403_),
    .Y(_0406_),
    .B1(_0405_));
 sg13g2_nor2_1 _1308_ (.A(_0404_),
    .B(_0406_),
    .Y(_0407_));
 sg13g2_nand2_1 _1309_ (.Y(_0408_),
    .A(_0402_),
    .B(_0406_));
 sg13g2_and2_1 _1310_ (.A(_0402_),
    .B(_0404_),
    .X(_0409_));
 sg13g2_xnor2_1 _1311_ (.Y(_0410_),
    .A(_0402_),
    .B(_0407_));
 sg13g2_xnor2_1 _1312_ (.Y(_0411_),
    .A(_0382_),
    .B(_0410_));
 sg13g2_or2_1 _1313_ (.X(_0412_),
    .B(_0411_),
    .A(_0379_));
 sg13g2_nand2_2 _1314_ (.Y(_0413_),
    .A(net245),
    .B(net192));
 sg13g2_a21oi_1 _1315_ (.A1(_0379_),
    .A2(_0411_),
    .Y(_0414_),
    .B1(_0413_));
 sg13g2_and2_1 _1316_ (.A(_0412_),
    .B(_0414_),
    .X(_0043_));
 sg13g2_a21o_1 _1317_ (.A2(_0364_),
    .A1(_0363_),
    .B1(_0376_),
    .X(_0415_));
 sg13g2_xnor2_1 _1318_ (.Y(_0416_),
    .A(_0016_),
    .B(_0105_));
 sg13g2_nand2_1 _1319_ (.Y(_0417_),
    .A(_0415_),
    .B(_0416_));
 sg13g2_xor2_1 _1320_ (.B(_0416_),
    .A(_0415_),
    .X(_0418_));
 sg13g2_and2_1 _1321_ (.A(net242),
    .B(_0106_),
    .X(_0419_));
 sg13g2_o21ai_1 _1322_ (.B1(_0399_),
    .Y(_0420_),
    .A1(_0383_),
    .A2(_0400_));
 sg13g2_o21ai_1 _1323_ (.B1(_0387_),
    .Y(_0421_),
    .A1(_0388_),
    .A2(_0395_));
 sg13g2_o21ai_1 _1324_ (.B1(_0381_),
    .Y(_0422_),
    .A1(_0369_),
    .A2(_0384_));
 sg13g2_nand2_2 _1325_ (.Y(_0423_),
    .A(uio_oe[1]),
    .B(uio_oe[6]));
 sg13g2_and4_1 _1326_ (.A(uio_oe[3]),
    .B(net236),
    .C(net227),
    .D(uio_oe[5]),
    .X(_0424_));
 sg13g2_nand2_1 _1327_ (.Y(_0425_),
    .A(uio_oe[2]),
    .B(uio_oe[5]));
 sg13g2_a22oi_1 _1328_ (.Y(_0426_),
    .B1(uio_oe[5]),
    .B2(net236),
    .A2(net227),
    .A1(uio_oe[3]));
 sg13g2_or3_1 _1329_ (.A(_0423_),
    .B(_0424_),
    .C(_0426_),
    .X(_0427_));
 sg13g2_o21ai_1 _1330_ (.B1(_0423_),
    .Y(_0428_),
    .A1(_0424_),
    .A2(_0426_));
 sg13g2_nand3_1 _1331_ (.B(_0427_),
    .C(_0428_),
    .A(_0422_),
    .Y(_0429_));
 sg13g2_a21o_1 _1332_ (.A2(_0428_),
    .A1(_0427_),
    .B1(_0422_),
    .X(_0430_));
 sg13g2_nand2_1 _1333_ (.Y(_0431_),
    .A(net232),
    .B(uio_oe[7]));
 sg13g2_nand2_2 _1334_ (.Y(_0432_),
    .A(net242),
    .B(uio_oe[7]));
 sg13g2_xnor2_1 _1335_ (.Y(_0433_),
    .A(_0111_),
    .B(_0432_));
 sg13g2_nand2b_1 _1336_ (.Y(_0434_),
    .B(_0433_),
    .A_N(_0425_));
 sg13g2_xnor2_1 _1337_ (.Y(_0435_),
    .A(_0425_),
    .B(_0433_));
 sg13g2_nand3_1 _1338_ (.B(_0430_),
    .C(_0435_),
    .A(_0429_),
    .Y(_0436_));
 sg13g2_a21o_1 _1339_ (.A2(_0430_),
    .A1(_0429_),
    .B1(_0435_),
    .X(_0437_));
 sg13g2_nand3_1 _1340_ (.B(_0436_),
    .C(_0437_),
    .A(_0421_),
    .Y(_0438_));
 sg13g2_a21o_1 _1341_ (.A2(_0437_),
    .A1(_0436_),
    .B1(_0421_),
    .X(_0439_));
 sg13g2_o21ai_1 _1342_ (.B1(_0391_),
    .Y(_0440_),
    .A1(_0384_),
    .A2(_0392_));
 sg13g2_nand2b_1 _1343_ (.Y(_0441_),
    .B(_0440_),
    .A_N(_0423_));
 sg13g2_xnor2_1 _1344_ (.Y(_0442_),
    .A(_0423_),
    .B(_0440_));
 sg13g2_nand2b_1 _1345_ (.Y(_0443_),
    .B(_0442_),
    .A_N(_0432_));
 sg13g2_xnor2_1 _1346_ (.Y(_0444_),
    .A(_0432_),
    .B(_0442_));
 sg13g2_nand3_1 _1347_ (.B(_0439_),
    .C(_0444_),
    .A(_0438_),
    .Y(_0445_));
 sg13g2_a21o_1 _1348_ (.A2(_0439_),
    .A1(_0438_),
    .B1(_0444_),
    .X(_0446_));
 sg13g2_nand3_1 _1349_ (.B(_0445_),
    .C(_0446_),
    .A(_0420_),
    .Y(_0447_));
 sg13g2_a21o_1 _1350_ (.A2(_0446_),
    .A1(_0445_),
    .B1(_0420_),
    .X(_0448_));
 sg13g2_and3_1 _1351_ (.X(_0449_),
    .A(_0419_),
    .B(_0447_),
    .C(_0448_));
 sg13g2_nand3_1 _1352_ (.B(_0447_),
    .C(_0448_),
    .A(_0419_),
    .Y(_0450_));
 sg13g2_a21oi_2 _1353_ (.B1(_0419_),
    .Y(_0451_),
    .A2(_0448_),
    .A1(_0447_));
 sg13g2_o21ai_1 _1354_ (.B1(_0408_),
    .Y(_0452_),
    .A1(_0449_),
    .A2(_0451_));
 sg13g2_nor3_1 _1355_ (.A(_0408_),
    .B(_0449_),
    .C(_0451_),
    .Y(_0453_));
 sg13g2_or3_1 _1356_ (.A(_0408_),
    .B(_0449_),
    .C(_0451_),
    .X(_0454_));
 sg13g2_a21oi_1 _1357_ (.A1(_0382_),
    .A2(_0410_),
    .Y(_0455_),
    .B1(_0409_));
 sg13g2_and3_1 _1358_ (.X(_0456_),
    .A(_0452_),
    .B(_0454_),
    .C(_0455_));
 sg13g2_a21oi_1 _1359_ (.A1(_0452_),
    .A2(_0454_),
    .Y(_0457_),
    .B1(_0455_));
 sg13g2_o21ai_1 _1360_ (.B1(_0418_),
    .Y(_0458_),
    .A1(_0456_),
    .A2(_0457_));
 sg13g2_or3_1 _1361_ (.A(_0418_),
    .B(_0456_),
    .C(_0457_),
    .X(_0459_));
 sg13g2_a21o_1 _1362_ (.A2(_0459_),
    .A1(_0458_),
    .B1(_0018_),
    .X(_0460_));
 sg13g2_nand3_1 _1363_ (.B(_0458_),
    .C(_0459_),
    .A(_0018_),
    .Y(_0461_));
 sg13g2_nand3_1 _1364_ (.B(_0460_),
    .C(_0461_),
    .A(_0378_),
    .Y(_0462_));
 sg13g2_a21oi_1 _1365_ (.A1(_0460_),
    .A2(_0461_),
    .Y(_0463_),
    .B1(_0378_));
 sg13g2_a21o_1 _1366_ (.A2(_0461_),
    .A1(_0460_),
    .B1(_0378_),
    .X(_0464_));
 sg13g2_nand2_1 _1367_ (.Y(_0465_),
    .A(_0462_),
    .B(_0464_));
 sg13g2_xnor2_1 _1368_ (.Y(_0466_),
    .A(_0412_),
    .B(_0465_));
 sg13g2_nor2_1 _1369_ (.A(_0413_),
    .B(_0466_),
    .Y(_0044_));
 sg13g2_o21ai_1 _1370_ (.B1(net192),
    .Y(_0467_),
    .A1(_0092_),
    .A2(_0417_));
 sg13g2_a21oi_1 _1371_ (.A1(_0092_),
    .A2(_0417_),
    .Y(_0468_),
    .B1(_0467_));
 sg13g2_inv_1 _1372_ (.Y(_0469_),
    .A(_0468_));
 sg13g2_a221oi_1 _1373_ (.B2(_0452_),
    .C1(_0453_),
    .B1(_0409_),
    .A1(net222),
    .Y(_0470_),
    .A2(_0382_));
 sg13g2_nand2_1 _1374_ (.Y(_0471_),
    .A(_0447_),
    .B(_0450_));
 sg13g2_nand2_1 _1375_ (.Y(_0472_),
    .A(_0441_),
    .B(_0443_));
 sg13g2_nand2_1 _1376_ (.Y(_0473_),
    .A(_0438_),
    .B(_0445_));
 sg13g2_nand2_1 _1377_ (.Y(_0474_),
    .A(_0429_),
    .B(_0436_));
 sg13g2_xor2_1 _1378_ (.B(_0370_),
    .A(uio_oe[4]),
    .X(_0475_));
 sg13g2_nand2b_1 _1379_ (.Y(_0476_),
    .B(_0427_),
    .A_N(_0424_));
 sg13g2_nand2_2 _1380_ (.Y(_0477_),
    .A(net239),
    .B(uio_oe[7]));
 sg13g2_nand2_2 _1381_ (.Y(_0478_),
    .A(uio_oe[2]),
    .B(uio_oe[6]));
 sg13g2_a22oi_1 _1382_ (.Y(_0479_),
    .B1(_0370_),
    .B2(_0478_),
    .A2(_0116_),
    .A1(_0106_));
 sg13g2_nand2b_1 _1383_ (.Y(_0480_),
    .B(_0479_),
    .A_N(_0477_));
 sg13g2_xnor2_1 _1384_ (.Y(_0481_),
    .A(_0477_),
    .B(_0479_));
 sg13g2_nand2_1 _1385_ (.Y(_0482_),
    .A(_0476_),
    .B(_0481_));
 sg13g2_xnor2_1 _1386_ (.Y(_0483_),
    .A(_0476_),
    .B(_0481_));
 sg13g2_xor2_1 _1387_ (.B(_0483_),
    .A(_0475_),
    .X(_0484_));
 sg13g2_xnor2_1 _1388_ (.Y(_0485_),
    .A(_0474_),
    .B(_0484_));
 sg13g2_o21ai_1 _1389_ (.B1(_0434_),
    .Y(_0486_),
    .A1(_0112_),
    .A2(_0432_));
 sg13g2_nand2b_1 _1390_ (.Y(_0487_),
    .B(_0486_),
    .A_N(_0478_));
 sg13g2_xnor2_1 _1391_ (.Y(_0488_),
    .A(_0478_),
    .B(_0486_));
 sg13g2_nand2b_1 _1392_ (.Y(_0489_),
    .B(_0488_),
    .A_N(_0477_));
 sg13g2_xnor2_1 _1393_ (.Y(_0490_),
    .A(_0477_),
    .B(_0488_));
 sg13g2_nor2b_1 _1394_ (.A(_0485_),
    .B_N(_0490_),
    .Y(_0491_));
 sg13g2_xnor2_1 _1395_ (.Y(_0492_),
    .A(_0485_),
    .B(_0490_));
 sg13g2_xnor2_1 _1396_ (.Y(_0493_),
    .A(_0473_),
    .B(_0492_));
 sg13g2_nor2b_1 _1397_ (.A(_0493_),
    .B_N(_0472_),
    .Y(_0494_));
 sg13g2_xnor2_1 _1398_ (.Y(_0495_),
    .A(_0472_),
    .B(_0493_));
 sg13g2_nand2_1 _1399_ (.Y(_0496_),
    .A(_0471_),
    .B(_0495_));
 sg13g2_xnor2_1 _1400_ (.Y(_0497_),
    .A(_0471_),
    .B(_0495_));
 sg13g2_xnor2_1 _1401_ (.Y(_0498_),
    .A(_0470_),
    .B(_0497_));
 sg13g2_nor2_1 _1402_ (.A(_0469_),
    .B(_0498_),
    .Y(_0499_));
 sg13g2_xnor2_1 _1403_ (.Y(_0500_),
    .A(_0468_),
    .B(_0498_));
 sg13g2_xnor2_1 _1404_ (.Y(_0501_),
    .A(_0007_),
    .B(_0500_));
 sg13g2_a21oi_1 _1405_ (.A1(_0458_),
    .A2(_0461_),
    .Y(_0502_),
    .B1(_0501_));
 sg13g2_nand3_1 _1406_ (.B(_0461_),
    .C(_0501_),
    .A(_0458_),
    .Y(_0503_));
 sg13g2_nor2b_1 _1407_ (.A(_0502_),
    .B_N(_0503_),
    .Y(_0504_));
 sg13g2_o21ai_1 _1408_ (.B1(_0462_),
    .Y(_0505_),
    .A1(_0412_),
    .A2(_0463_));
 sg13g2_xnor2_1 _1409_ (.Y(_0506_),
    .A(_0504_),
    .B(_0505_));
 sg13g2_nor2_1 _1410_ (.A(_0413_),
    .B(_0506_),
    .Y(_0045_));
 sg13g2_a21oi_1 _1411_ (.A1(_0503_),
    .A2(_0505_),
    .Y(_0507_),
    .B1(_0502_));
 sg13g2_o21ai_1 _1412_ (.B1(_0496_),
    .Y(_0508_),
    .A1(_0470_),
    .A2(_0497_));
 sg13g2_a21o_1 _1413_ (.A2(_0492_),
    .A1(_0473_),
    .B1(_0494_),
    .X(_0509_));
 sg13g2_nand2_1 _1414_ (.Y(_0510_),
    .A(_0487_),
    .B(_0489_));
 sg13g2_a21o_1 _1415_ (.A2(_0484_),
    .A1(_0474_),
    .B1(_0491_),
    .X(_0511_));
 sg13g2_nand2_1 _1416_ (.Y(_0512_),
    .A(uio_oe[2]),
    .B(uio_oe[7]));
 sg13g2_a22oi_1 _1417_ (.Y(_0513_),
    .B1(_0111_),
    .B2(net224),
    .A2(uio_oe[6]),
    .A1(net232));
 sg13g2_a21o_1 _1418_ (.A2(_0111_),
    .A1(_0106_),
    .B1(_0513_),
    .X(_0514_));
 sg13g2_nor2_1 _1419_ (.A(_0512_),
    .B(_0514_),
    .Y(_0515_));
 sg13g2_xor2_1 _1420_ (.B(_0514_),
    .A(_0512_),
    .X(_0516_));
 sg13g2_inv_1 _1421_ (.Y(_0517_),
    .A(_0516_));
 sg13g2_a22oi_1 _1422_ (.Y(_0518_),
    .B1(uio_oe[6]),
    .B2(uio_oe[3]),
    .A2(uio_oe[7]),
    .A1(uio_oe[2]));
 sg13g2_a21oi_1 _1423_ (.A1(_0109_),
    .A2(_0116_),
    .Y(_0519_),
    .B1(_0518_));
 sg13g2_o21ai_1 _1424_ (.B1(_0480_),
    .Y(_0520_),
    .A1(_0107_),
    .A2(_0117_));
 sg13g2_nand2_1 _1425_ (.Y(_0521_),
    .A(_0519_),
    .B(_0520_));
 sg13g2_xnor2_1 _1426_ (.Y(_0522_),
    .A(_0519_),
    .B(_0520_));
 sg13g2_o21ai_1 _1427_ (.B1(_0482_),
    .Y(_0523_),
    .A1(_0475_),
    .A2(_0483_));
 sg13g2_nand2b_1 _1428_ (.Y(_0524_),
    .B(_0523_),
    .A_N(_0522_));
 sg13g2_xor2_1 _1429_ (.B(_0523_),
    .A(_0522_),
    .X(_0525_));
 sg13g2_xnor2_1 _1430_ (.Y(_0526_),
    .A(_0517_),
    .B(_0525_));
 sg13g2_nor2b_1 _1431_ (.A(_0526_),
    .B_N(_0511_),
    .Y(_0527_));
 sg13g2_xnor2_1 _1432_ (.Y(_0528_),
    .A(_0511_),
    .B(_0526_));
 sg13g2_xnor2_1 _1433_ (.Y(_0529_),
    .A(_0510_),
    .B(_0528_));
 sg13g2_nor2b_1 _1434_ (.A(_0529_),
    .B_N(_0509_),
    .Y(_0530_));
 sg13g2_nand2b_1 _1435_ (.Y(_0531_),
    .B(_0529_),
    .A_N(_0509_));
 sg13g2_xor2_1 _1436_ (.B(_0529_),
    .A(_0509_),
    .X(_0532_));
 sg13g2_xnor2_1 _1437_ (.Y(_0533_),
    .A(_0508_),
    .B(_0532_));
 sg13g2_and2_1 _1438_ (.A(_0467_),
    .B(_0533_),
    .X(_0534_));
 sg13g2_xor2_1 _1439_ (.B(_0533_),
    .A(_0467_),
    .X(_0535_));
 sg13g2_xnor2_1 _1440_ (.Y(_0536_),
    .A(_0017_),
    .B(_0535_));
 sg13g2_a21oi_1 _1441_ (.A1(_0007_),
    .A2(_0500_),
    .Y(_0537_),
    .B1(_0499_));
 sg13g2_or2_1 _1442_ (.X(_0538_),
    .B(_0537_),
    .A(_0536_));
 sg13g2_xnor2_1 _1443_ (.Y(_0539_),
    .A(_0536_),
    .B(_0537_));
 sg13g2_nor2_1 _1444_ (.A(_0507_),
    .B(_0539_),
    .Y(_0540_));
 sg13g2_a21oi_1 _1445_ (.A1(_0507_),
    .A2(_0539_),
    .Y(_0541_),
    .B1(_0413_));
 sg13g2_nor2b_1 _1446_ (.A(_0540_),
    .B_N(_0541_),
    .Y(_0046_));
 sg13g2_a21o_1 _1447_ (.A2(_0528_),
    .A1(_0510_),
    .B1(_0527_),
    .X(_0542_));
 sg13g2_a21oi_2 _1448_ (.B1(_0515_),
    .Y(_0543_),
    .A2(_0111_),
    .A1(_0106_));
 sg13g2_o21ai_1 _1449_ (.B1(_0524_),
    .Y(_0544_),
    .A1(_0517_),
    .A2(_0525_));
 sg13g2_nand2b_1 _1450_ (.Y(_0545_),
    .B(_0478_),
    .A_N(_0431_));
 sg13g2_inv_1 _1451_ (.Y(_0546_),
    .A(_0545_));
 sg13g2_nor2_1 _1452_ (.A(_0015_),
    .B(_0362_),
    .Y(_0547_));
 sg13g2_xor2_1 _1453_ (.B(_0362_),
    .A(_0015_),
    .X(_0548_));
 sg13g2_xnor2_1 _1454_ (.Y(_0549_),
    .A(_0545_),
    .B(_0548_));
 sg13g2_nor2b_1 _1455_ (.A(_0521_),
    .B_N(_0549_),
    .Y(_0550_));
 sg13g2_xnor2_1 _1456_ (.Y(_0551_),
    .A(_0521_),
    .B(_0549_));
 sg13g2_nand2_1 _1457_ (.Y(_0552_),
    .A(net228),
    .B(_0122_));
 sg13g2_xor2_1 _1458_ (.B(_0552_),
    .A(_0431_),
    .X(_0553_));
 sg13g2_xnor2_1 _1459_ (.Y(_0554_),
    .A(_0551_),
    .B(_0553_));
 sg13g2_nand2b_1 _1460_ (.Y(_0555_),
    .B(_0544_),
    .A_N(_0554_));
 sg13g2_xor2_1 _1461_ (.B(_0554_),
    .A(_0544_),
    .X(_0556_));
 sg13g2_xor2_1 _1462_ (.B(_0556_),
    .A(_0543_),
    .X(_0557_));
 sg13g2_nand2_1 _1463_ (.Y(_0558_),
    .A(_0542_),
    .B(_0557_));
 sg13g2_a21oi_2 _1464_ (.B1(_0530_),
    .Y(_0559_),
    .A2(_0531_),
    .A1(_0508_));
 sg13g2_xnor2_1 _1465_ (.Y(_0560_),
    .A(_0542_),
    .B(_0557_));
 sg13g2_o21ai_1 _1466_ (.B1(_0558_),
    .Y(_0561_),
    .A1(_0559_),
    .A2(_0560_));
 sg13g2_o21ai_1 _1467_ (.B1(_0555_),
    .Y(_0562_),
    .A1(_0543_),
    .A2(_0556_));
 sg13g2_nand2_1 _1468_ (.Y(_0563_),
    .A(net225),
    .B(_0363_));
 sg13g2_o21ai_1 _1469_ (.B1(_0563_),
    .Y(_0564_),
    .A1(_0431_),
    .A2(_0552_));
 sg13g2_a21oi_1 _1470_ (.A1(_0551_),
    .A2(_0553_),
    .Y(_0565_),
    .B1(_0550_));
 sg13g2_nand2_1 _1471_ (.Y(_0566_),
    .A(_0105_),
    .B(_0363_));
 sg13g2_nand2_1 _1472_ (.Y(_0567_),
    .A(net228),
    .B(net230));
 sg13g2_a22oi_1 _1473_ (.Y(_0568_),
    .B1(_0567_),
    .B2(_0107_),
    .A2(_0363_),
    .A1(_0105_));
 sg13g2_a22oi_1 _1474_ (.Y(_0569_),
    .B1(_0546_),
    .B2(_0548_),
    .A2(_0116_),
    .A1(_0109_));
 sg13g2_nor2b_1 _1475_ (.A(_0569_),
    .B_N(_0568_),
    .Y(_0570_));
 sg13g2_xnor2_1 _1476_ (.Y(_0571_),
    .A(_0568_),
    .B(_0569_));
 sg13g2_nand2_1 _1477_ (.Y(_0572_),
    .A(net224),
    .B(_0547_));
 sg13g2_o21ai_1 _1478_ (.B1(_0572_),
    .Y(_0573_),
    .A1(_0106_),
    .A2(_0547_));
 sg13g2_nor2_1 _1479_ (.A(_0567_),
    .B(_0573_),
    .Y(_0574_));
 sg13g2_xor2_1 _1480_ (.B(_0573_),
    .A(_0567_),
    .X(_0575_));
 sg13g2_xnor2_1 _1481_ (.Y(_0576_),
    .A(_0571_),
    .B(_0575_));
 sg13g2_nor2_1 _1482_ (.A(_0565_),
    .B(_0576_),
    .Y(_0577_));
 sg13g2_xor2_1 _1483_ (.B(_0576_),
    .A(_0565_),
    .X(_0578_));
 sg13g2_xnor2_1 _1484_ (.Y(_0579_),
    .A(_0564_),
    .B(_0578_));
 sg13g2_nor2b_1 _1485_ (.A(_0579_),
    .B_N(_0562_),
    .Y(_0580_));
 sg13g2_xnor2_1 _1486_ (.Y(_0581_),
    .A(_0562_),
    .B(_0579_));
 sg13g2_xnor2_1 _1487_ (.Y(_0582_),
    .A(_0561_),
    .B(_0581_));
 sg13g2_nor2_1 _1488_ (.A(_0019_),
    .B(_0582_),
    .Y(_0583_));
 sg13g2_xnor2_1 _1489_ (.Y(_0584_),
    .A(uo_out[1]),
    .B(_0582_));
 sg13g2_a21oi_1 _1490_ (.A1(_0005_),
    .A2(_0584_),
    .Y(_0585_),
    .B1(_0583_));
 sg13g2_a21oi_1 _1491_ (.A1(_0561_),
    .A2(_0581_),
    .Y(_0586_),
    .B1(_0580_));
 sg13g2_a21oi_1 _1492_ (.A1(_0564_),
    .A2(_0578_),
    .Y(_0587_),
    .B1(_0577_));
 sg13g2_a21oi_1 _1493_ (.A1(net224),
    .A2(_0547_),
    .Y(_0588_),
    .B1(_0574_));
 sg13g2_xor2_1 _1494_ (.B(_0566_),
    .A(_0016_),
    .X(_0589_));
 sg13g2_a21o_1 _1495_ (.A2(_0575_),
    .A1(_0571_),
    .B1(_0570_),
    .X(_0590_));
 sg13g2_xor2_1 _1496_ (.B(_0590_),
    .A(_0589_),
    .X(_0591_));
 sg13g2_nor2b_1 _1497_ (.A(_0588_),
    .B_N(_0591_),
    .Y(_0592_));
 sg13g2_xnor2_1 _1498_ (.Y(_0593_),
    .A(_0588_),
    .B(_0591_));
 sg13g2_nand2b_1 _1499_ (.Y(_0594_),
    .B(_0593_),
    .A_N(_0587_));
 sg13g2_xnor2_1 _1500_ (.Y(_0595_),
    .A(_0587_),
    .B(_0593_));
 sg13g2_nand2b_1 _1501_ (.Y(_0596_),
    .B(_0595_),
    .A_N(_0586_));
 sg13g2_xnor2_1 _1502_ (.Y(_0597_),
    .A(_0586_),
    .B(_0595_));
 sg13g2_and2_1 _1503_ (.A(uo_out[2]),
    .B(_0597_),
    .X(_0598_));
 sg13g2_xnor2_1 _1504_ (.Y(_0599_),
    .A(_0087_),
    .B(_0597_));
 sg13g2_xnor2_1 _1505_ (.Y(_0600_),
    .A(_0004_),
    .B(_0599_));
 sg13g2_nor2_1 _1506_ (.A(_0585_),
    .B(_0600_),
    .Y(_0601_));
 sg13g2_xor2_1 _1507_ (.B(_0600_),
    .A(_0585_),
    .X(_0602_));
 sg13g2_xnor2_1 _1508_ (.Y(_0603_),
    .A(_0005_),
    .B(_0584_));
 sg13g2_xor2_1 _1509_ (.B(_0560_),
    .A(_0559_),
    .X(_0604_));
 sg13g2_nand2_1 _1510_ (.Y(_0605_),
    .A(uo_out[0]),
    .B(_0604_));
 sg13g2_xor2_1 _1511_ (.B(_0604_),
    .A(uo_out[0]),
    .X(_0606_));
 sg13g2_nand2_1 _1512_ (.Y(_0607_),
    .A(_0006_),
    .B(_0606_));
 sg13g2_and3_1 _1513_ (.X(_0608_),
    .A(_0603_),
    .B(_0605_),
    .C(_0607_));
 sg13g2_a21o_1 _1514_ (.A2(_0607_),
    .A1(_0605_),
    .B1(_0603_),
    .X(_0609_));
 sg13g2_a21o_1 _1515_ (.A2(_0535_),
    .A1(_0017_),
    .B1(_0534_),
    .X(_0610_));
 sg13g2_xnor2_1 _1516_ (.Y(_0611_),
    .A(_0006_),
    .B(_0606_));
 sg13g2_nor2b_1 _1517_ (.A(_0611_),
    .B_N(_0610_),
    .Y(_0612_));
 sg13g2_o21ai_1 _1518_ (.B1(_0538_),
    .Y(_0613_),
    .A1(_0507_),
    .A2(_0539_));
 sg13g2_xnor2_1 _1519_ (.Y(_0614_),
    .A(_0610_),
    .B(_0611_));
 sg13g2_a21oi_2 _1520_ (.B1(_0612_),
    .Y(_0615_),
    .A2(_0614_),
    .A1(_0613_));
 sg13g2_o21ai_1 _1521_ (.B1(_0609_),
    .Y(_0616_),
    .A1(_0608_),
    .A2(_0615_));
 sg13g2_a21oi_1 _1522_ (.A1(_0602_),
    .A2(_0616_),
    .Y(_0617_),
    .B1(_0601_));
 sg13g2_a21oi_1 _1523_ (.A1(_0004_),
    .A2(_0599_),
    .Y(_0618_),
    .B1(_0598_));
 sg13g2_nand2_1 _1524_ (.Y(_0619_),
    .A(_0594_),
    .B(_0596_));
 sg13g2_a21oi_1 _1525_ (.A1(_0589_),
    .A2(_0590_),
    .Y(_0620_),
    .B1(_0592_));
 sg13g2_o21ai_1 _1526_ (.B1(_0105_),
    .Y(_0621_),
    .A1(_0016_),
    .A2(_0362_));
 sg13g2_xor2_1 _1527_ (.B(uo_out[3]),
    .A(\izh_2.u[7] ),
    .X(_0622_));
 sg13g2_xnor2_1 _1528_ (.Y(_0623_),
    .A(_0621_),
    .B(_0622_));
 sg13g2_xnor2_1 _1529_ (.Y(_0624_),
    .A(_0620_),
    .B(_0623_));
 sg13g2_xnor2_1 _1530_ (.Y(_0625_),
    .A(_0619_),
    .B(_0624_));
 sg13g2_xor2_1 _1531_ (.B(_0625_),
    .A(_0618_),
    .X(_0626_));
 sg13g2_xnor2_1 _1532_ (.Y(_0627_),
    .A(_0617_),
    .B(_0626_));
 sg13g2_nor2_1 _1533_ (.A(_0413_),
    .B(_0627_),
    .Y(_0047_));
 sg13g2_nand2_1 _1534_ (.Y(_0628_),
    .A(net191),
    .B(_0191_));
 sg13g2_xor2_1 _1535_ (.B(_0628_),
    .A(net92),
    .X(_0629_));
 sg13g2_nor2_1 _1536_ (.A(net243),
    .B(_0629_),
    .Y(_0048_));
 sg13g2_xnor2_1 _1537_ (.Y(_0630_),
    .A(_0192_),
    .B(_0194_));
 sg13g2_o21ai_1 _1538_ (.B1(net245),
    .Y(_0631_),
    .A1(net87),
    .A2(net191));
 sg13g2_a21oi_1 _1539_ (.A1(net191),
    .A2(_0630_),
    .Y(_0049_),
    .B1(_0631_));
 sg13g2_xnor2_1 _1540_ (.Y(_0632_),
    .A(_0195_),
    .B(_0196_));
 sg13g2_o21ai_1 _1541_ (.B1(net245),
    .Y(_0633_),
    .A1(net65),
    .A2(net191));
 sg13g2_a21oi_1 _1542_ (.A1(net191),
    .A2(_0632_),
    .Y(_0050_),
    .B1(_0633_));
 sg13g2_xnor2_1 _1543_ (.Y(_0634_),
    .A(_0197_),
    .B(_0198_));
 sg13g2_o21ai_1 _1544_ (.B1(net245),
    .Y(_0635_),
    .A1(net76),
    .A2(net191));
 sg13g2_a21oi_1 _1545_ (.A1(net191),
    .A2(_0634_),
    .Y(_0051_),
    .B1(_0635_));
 sg13g2_xnor2_1 _1546_ (.Y(_0636_),
    .A(_0199_),
    .B(_0200_));
 sg13g2_o21ai_1 _1547_ (.B1(net245),
    .Y(_0637_),
    .A1(net72),
    .A2(net191));
 sg13g2_a21oi_1 _1548_ (.A1(net192),
    .A2(_0636_),
    .Y(_0052_),
    .B1(_0637_));
 sg13g2_xor2_1 _1549_ (.B(_0202_),
    .A(_0201_),
    .X(_0638_));
 sg13g2_nor2_1 _1550_ (.A(\izh_2.spike ),
    .B(_0638_),
    .Y(_0639_));
 sg13g2_o21ai_1 _1551_ (.B1(net246),
    .Y(_0640_),
    .A1(net83),
    .A2(net194));
 sg13g2_nor2_1 _1552_ (.A(_0639_),
    .B(_0640_),
    .Y(_0053_));
 sg13g2_xnor2_1 _1553_ (.Y(_0641_),
    .A(_0203_),
    .B(_0204_));
 sg13g2_o21ai_1 _1554_ (.B1(net246),
    .Y(_0642_),
    .A1(net75),
    .A2(net194));
 sg13g2_a21oi_1 _1555_ (.A1(net194),
    .A2(_0641_),
    .Y(_0054_),
    .B1(_0642_));
 sg13g2_xnor2_1 _1556_ (.Y(_0643_),
    .A(_0205_),
    .B(_0206_));
 sg13g2_o21ai_1 _1557_ (.B1(net245),
    .Y(_0644_),
    .A1(net97),
    .A2(net193));
 sg13g2_a21oi_1 _1558_ (.A1(net193),
    .A2(_0643_),
    .Y(_0055_),
    .B1(_0644_));
 sg13g2_xnor2_1 _1559_ (.Y(_0645_),
    .A(_0207_),
    .B(_0208_));
 sg13g2_o21ai_1 _1560_ (.B1(net245),
    .Y(_0646_),
    .A1(net66),
    .A2(net192));
 sg13g2_a21oi_1 _1561_ (.A1(net192),
    .A2(_0645_),
    .Y(_0056_),
    .B1(_0646_));
 sg13g2_xnor2_1 _1562_ (.Y(_0647_),
    .A(_0613_),
    .B(_0614_));
 sg13g2_a21oi_1 _1563_ (.A1(net192),
    .A2(_0647_),
    .Y(_0057_),
    .B1(net243));
 sg13g2_nand2b_1 _1564_ (.Y(_0648_),
    .B(_0609_),
    .A_N(_0608_));
 sg13g2_xnor2_1 _1565_ (.Y(_0649_),
    .A(_0615_),
    .B(_0648_));
 sg13g2_a21oi_1 _1566_ (.A1(net194),
    .A2(_0649_),
    .Y(_0058_),
    .B1(net243));
 sg13g2_xnor2_1 _1567_ (.Y(_0650_),
    .A(_0602_),
    .B(_0616_));
 sg13g2_a21oi_1 _1568_ (.A1(net194),
    .A2(_0650_),
    .Y(_0059_),
    .B1(net243));
 sg13g2_xor2_1 _1569_ (.B(net209),
    .A(uo_out[5]),
    .X(_0651_));
 sg13g2_nand2b_1 _1570_ (.Y(_0652_),
    .B(_0264_),
    .A_N(_0266_));
 sg13g2_and2_1 _1571_ (.A(uo_out[2]),
    .B(net205),
    .X(_0653_));
 sg13g2_nand2_2 _1572_ (.Y(_0654_),
    .A(uo_out[2]),
    .B(uo_out[4]));
 sg13g2_a22oi_1 _1573_ (.Y(_0655_),
    .B1(uo_out[4]),
    .B2(uo_out[1]),
    .A2(uo_out[2]),
    .A1(uo_out[3]));
 sg13g2_nand4_1 _1574_ (.B(uo_out[3]),
    .C(uo_out[2]),
    .A(uo_out[1]),
    .Y(_0656_),
    .D(uo_out[4]));
 sg13g2_nor2b_1 _1575_ (.A(_0655_),
    .B_N(_0656_),
    .Y(_0657_));
 sg13g2_nand2_1 _1576_ (.Y(_0658_),
    .A(_0241_),
    .B(_0657_));
 sg13g2_nand3_1 _1577_ (.B(_0654_),
    .C(_0658_),
    .A(_0652_),
    .Y(_0659_));
 sg13g2_o21ai_1 _1578_ (.B1(_0659_),
    .Y(_0660_),
    .A1(net211),
    .A2(uo_out[5]));
 sg13g2_nand2_1 _1579_ (.Y(_0661_),
    .A(net206),
    .B(net200));
 sg13g2_a22oi_1 _1580_ (.Y(_0662_),
    .B1(uo_out[6]),
    .B2(uo_out[4]),
    .A2(uo_out[5]),
    .A1(net211));
 sg13g2_a22oi_1 _1581_ (.Y(_0663_),
    .B1(_0660_),
    .B2(_0662_),
    .A2(_0090_),
    .A1(_0088_));
 sg13g2_nand2_1 _1582_ (.Y(_0664_),
    .A(_0651_),
    .B(_0663_));
 sg13g2_xnor2_1 _1583_ (.Y(_0665_),
    .A(_0651_),
    .B(_0663_));
 sg13g2_nand2_1 _1584_ (.Y(_0666_),
    .A(\izh_1.u[0] ),
    .B(_0665_));
 sg13g2_xor2_1 _1585_ (.B(_0665_),
    .A(net107),
    .X(_0667_));
 sg13g2_nor2_1 _1586_ (.A(_0087_),
    .B(_0019_),
    .Y(_0668_));
 sg13g2_and3_1 _1587_ (.X(_0669_),
    .A(uo_out[0]),
    .B(uo_out[4]),
    .C(_0241_));
 sg13g2_a21oi_1 _1588_ (.A1(uo_out[0]),
    .A2(uo_out[4]),
    .Y(_0670_),
    .B1(_0241_));
 sg13g2_nor2_1 _1589_ (.A(_0669_),
    .B(_0670_),
    .Y(_0671_));
 sg13g2_xnor2_1 _1590_ (.Y(_0672_),
    .A(_0668_),
    .B(_0671_));
 sg13g2_nor3_1 _1591_ (.A(_0087_),
    .B(_0242_),
    .C(_0672_),
    .Y(_0673_));
 sg13g2_or3_1 _1592_ (.A(uo_out[1]),
    .B(_0652_),
    .C(_0672_),
    .X(_0674_));
 sg13g2_a21oi_1 _1593_ (.A1(_0668_),
    .A2(_0671_),
    .Y(_0675_),
    .B1(_0669_));
 sg13g2_inv_1 _1594_ (.Y(_0676_),
    .A(_0675_));
 sg13g2_nand2_1 _1595_ (.Y(_0677_),
    .A(uo_out[0]),
    .B(uo_out[5]));
 sg13g2_o21ai_1 _1596_ (.B1(_0656_),
    .Y(_0678_),
    .A1(_0655_),
    .A2(_0677_));
 sg13g2_nand2_1 _1597_ (.Y(_0679_),
    .A(uo_out[0]),
    .B(uo_out[6]));
 sg13g2_nand2b_1 _1598_ (.Y(_0680_),
    .B(_0678_),
    .A_N(_0679_));
 sg13g2_xor2_1 _1599_ (.B(_0679_),
    .A(_0678_),
    .X(_0681_));
 sg13g2_nand2_1 _1600_ (.Y(_0682_),
    .A(net217),
    .B(uo_out[5]));
 sg13g2_xnor2_1 _1601_ (.Y(_0683_),
    .A(_0000_),
    .B(_0654_));
 sg13g2_xor2_1 _1602_ (.B(_0683_),
    .A(_0682_),
    .X(_0684_));
 sg13g2_nand2_2 _1603_ (.Y(_0685_),
    .A(uo_out[1]),
    .B(uo_out[6]));
 sg13g2_and4_1 _1604_ (.A(uo_out[1]),
    .B(uo_out[0]),
    .C(uo_out[5]),
    .D(uo_out[6]),
    .X(_0686_));
 sg13g2_nand4_1 _1605_ (.B(net219),
    .C(uo_out[5]),
    .A(net217),
    .Y(_0687_),
    .D(uo_out[6]));
 sg13g2_a22oi_1 _1606_ (.Y(_0688_),
    .B1(uo_out[6]),
    .B2(net219),
    .A2(net203),
    .A1(net217));
 sg13g2_nand3b_1 _1607_ (.B(_0653_),
    .C(_0687_),
    .Y(_0689_),
    .A_N(_0688_));
 sg13g2_o21ai_1 _1608_ (.B1(_0654_),
    .Y(_0690_),
    .A1(_0686_),
    .A2(_0688_));
 sg13g2_and3_1 _1609_ (.X(_0691_),
    .A(_0678_),
    .B(_0689_),
    .C(_0690_));
 sg13g2_nand3_1 _1610_ (.B(_0689_),
    .C(_0690_),
    .A(_0678_),
    .Y(_0692_));
 sg13g2_a21o_1 _1611_ (.A2(_0690_),
    .A1(_0689_),
    .B1(_0678_),
    .X(_0693_));
 sg13g2_nand3_1 _1612_ (.B(_0692_),
    .C(_0693_),
    .A(_0684_),
    .Y(_0694_));
 sg13g2_a21o_1 _1613_ (.A2(_0693_),
    .A1(_0692_),
    .B1(_0684_),
    .X(_0695_));
 sg13g2_xnor2_1 _1614_ (.Y(_0696_),
    .A(_0657_),
    .B(_0677_));
 sg13g2_and3_1 _1615_ (.X(_0697_),
    .A(_0694_),
    .B(_0695_),
    .C(_0696_));
 sg13g2_nand3_1 _1616_ (.B(_0695_),
    .C(_0696_),
    .A(_0694_),
    .Y(_0698_));
 sg13g2_a21oi_1 _1617_ (.A1(_0694_),
    .A2(_0695_),
    .Y(_0699_),
    .B1(_0696_));
 sg13g2_o21ai_1 _1618_ (.B1(_0681_),
    .Y(_0700_),
    .A1(_0697_),
    .A2(_0699_));
 sg13g2_or3_1 _1619_ (.A(_0681_),
    .B(_0697_),
    .C(_0699_),
    .X(_0701_));
 sg13g2_and3_1 _1620_ (.X(_0702_),
    .A(_0676_),
    .B(_0700_),
    .C(_0701_));
 sg13g2_a21oi_1 _1621_ (.A1(_0700_),
    .A2(_0701_),
    .Y(_0703_),
    .B1(_0676_));
 sg13g2_nor3_1 _1622_ (.A(_0674_),
    .B(_0702_),
    .C(_0703_),
    .Y(_0704_));
 sg13g2_o21ai_1 _1623_ (.B1(_0674_),
    .Y(_0705_),
    .A1(_0702_),
    .A2(_0703_));
 sg13g2_nor2b_1 _1624_ (.A(_0704_),
    .B_N(_0705_),
    .Y(_0706_));
 sg13g2_xnor2_1 _1625_ (.Y(_0707_),
    .A(_0673_),
    .B(_0706_));
 sg13g2_or2_1 _1626_ (.X(_0708_),
    .B(_0707_),
    .A(_0667_));
 sg13g2_nand2_2 _1627_ (.Y(_0709_),
    .A(net247),
    .B(net198));
 sg13g2_a21oi_1 _1628_ (.A1(_0667_),
    .A2(_0707_),
    .Y(_0710_),
    .B1(_0709_));
 sg13g2_and2_1 _1629_ (.A(_0708_),
    .B(_0710_),
    .X(_0060_));
 sg13g2_a21oi_1 _1630_ (.A1(_0673_),
    .A2(_0705_),
    .Y(_0711_),
    .B1(_0704_));
 sg13g2_o21ai_1 _1631_ (.B1(_0698_),
    .Y(_0712_),
    .A1(_0681_),
    .A2(_0699_));
 sg13g2_a21oi_1 _1632_ (.A1(_0684_),
    .A2(_0693_),
    .Y(_0713_),
    .B1(_0691_));
 sg13g2_and2_1 _1633_ (.A(uo_out[2]),
    .B(net203),
    .X(_0714_));
 sg13g2_nand2_1 _1634_ (.Y(_0715_),
    .A(_0687_),
    .B(_0689_));
 sg13g2_and2_1 _1635_ (.A(net219),
    .B(uo_out[7]),
    .X(_0716_));
 sg13g2_nand2_1 _1636_ (.Y(_0717_),
    .A(net219),
    .B(uo_out[7]));
 sg13g2_nor2_1 _1637_ (.A(_0685_),
    .B(_0717_),
    .Y(_0718_));
 sg13g2_xnor2_1 _1638_ (.Y(_0719_),
    .A(_0685_),
    .B(_0716_));
 sg13g2_xnor2_1 _1639_ (.Y(_0720_),
    .A(_0715_),
    .B(_0719_));
 sg13g2_nor2_1 _1640_ (.A(_0713_),
    .B(_0720_),
    .Y(_0721_));
 sg13g2_xor2_1 _1641_ (.B(_0720_),
    .A(_0713_),
    .X(_0722_));
 sg13g2_nand2_1 _1642_ (.Y(_0723_),
    .A(uo_out[3]),
    .B(_0653_));
 sg13g2_o21ai_1 _1643_ (.B1(_0723_),
    .Y(_0724_),
    .A1(_0682_),
    .A2(_0683_));
 sg13g2_nor2b_1 _1644_ (.A(_0685_),
    .B_N(_0724_),
    .Y(_0725_));
 sg13g2_xnor2_1 _1645_ (.Y(_0726_),
    .A(_0685_),
    .B(_0724_));
 sg13g2_xnor2_1 _1646_ (.Y(_0727_),
    .A(_0717_),
    .B(_0726_));
 sg13g2_xnor2_1 _1647_ (.Y(_0728_),
    .A(_0722_),
    .B(_0727_));
 sg13g2_nand2b_1 _1648_ (.Y(_0729_),
    .B(_0712_),
    .A_N(_0728_));
 sg13g2_xor2_1 _1649_ (.B(_0728_),
    .A(_0712_),
    .X(_0730_));
 sg13g2_xor2_1 _1650_ (.B(_0730_),
    .A(_0680_),
    .X(_0731_));
 sg13g2_nand2_1 _1651_ (.Y(_0732_),
    .A(_0702_),
    .B(_0731_));
 sg13g2_xnor2_1 _1652_ (.Y(_0733_),
    .A(_0702_),
    .B(_0731_));
 sg13g2_xnor2_1 _1653_ (.Y(_0734_),
    .A(_0711_),
    .B(_0733_));
 sg13g2_nand2_1 _1654_ (.Y(_0735_),
    .A(_0101_),
    .B(_0664_));
 sg13g2_xor2_1 _1655_ (.B(_0735_),
    .A(_0001_),
    .X(_0736_));
 sg13g2_nor2_1 _1656_ (.A(_0734_),
    .B(_0736_),
    .Y(_0737_));
 sg13g2_xor2_1 _1657_ (.B(_0736_),
    .A(_0734_),
    .X(_0738_));
 sg13g2_xnor2_1 _1658_ (.Y(_0739_),
    .A(_0003_),
    .B(_0738_));
 sg13g2_nand2b_1 _1659_ (.Y(_0740_),
    .B(_0666_),
    .A_N(_0739_));
 sg13g2_xor2_1 _1660_ (.B(_0739_),
    .A(_0666_),
    .X(_0741_));
 sg13g2_a21oi_1 _1661_ (.A1(_0708_),
    .A2(_0741_),
    .Y(_0742_),
    .B1(_0709_));
 sg13g2_o21ai_1 _1662_ (.B1(_0742_),
    .Y(_0743_),
    .A1(_0708_),
    .A2(_0741_));
 sg13g2_inv_1 _1663_ (.Y(_0061_),
    .A(_0743_));
 sg13g2_o21ai_1 _1664_ (.B1(_0740_),
    .Y(_0744_),
    .A1(_0708_),
    .A2(_0741_));
 sg13g2_nor2_1 _1665_ (.A(_0001_),
    .B(_0664_),
    .Y(_0745_));
 sg13g2_nor2_1 _1666_ (.A(net209),
    .B(_0745_),
    .Y(_0746_));
 sg13g2_a21o_1 _1667_ (.A2(_0745_),
    .A1(net209),
    .B1(\izh_1.spike ),
    .X(_0747_));
 sg13g2_inv_1 _1668_ (.Y(_0748_),
    .A(_0747_));
 sg13g2_nor2_1 _1669_ (.A(_0746_),
    .B(_0747_),
    .Y(_0749_));
 sg13g2_o21ai_1 _1670_ (.B1(_0732_),
    .Y(_0750_),
    .A1(_0711_),
    .A2(_0733_));
 sg13g2_o21ai_1 _1671_ (.B1(_0729_),
    .Y(_0751_),
    .A1(_0680_),
    .A2(_0730_));
 sg13g2_a21oi_1 _1672_ (.A1(_0716_),
    .A2(_0726_),
    .Y(_0752_),
    .B1(_0725_));
 sg13g2_a21oi_1 _1673_ (.A1(_0722_),
    .A2(_0727_),
    .Y(_0753_),
    .B1(_0721_));
 sg13g2_nand2_1 _1674_ (.Y(_0754_),
    .A(net217),
    .B(net209));
 sg13g2_a22oi_1 _1675_ (.Y(_0755_),
    .B1(uo_out[6]),
    .B2(net215),
    .A2(net205),
    .A1(net212));
 sg13g2_nand2_1 _1676_ (.Y(_0756_),
    .A(net212),
    .B(net200));
 sg13g2_or2_1 _1677_ (.X(_0757_),
    .B(_0756_),
    .A(_0654_));
 sg13g2_nand2b_1 _1678_ (.Y(_0758_),
    .B(_0757_),
    .A_N(_0755_));
 sg13g2_xnor2_1 _1679_ (.Y(_0759_),
    .A(_0754_),
    .B(_0758_));
 sg13g2_mux2_1 _1680_ (.A0(_0714_),
    .A1(_0715_),
    .S(_0719_),
    .X(_0760_));
 sg13g2_o21ai_1 _1681_ (.B1(_0754_),
    .Y(_0761_),
    .A1(_0087_),
    .A2(_0090_));
 sg13g2_nand2_2 _1682_ (.Y(_0762_),
    .A(net215),
    .B(uo_out[7]));
 sg13g2_o21ai_1 _1683_ (.B1(_0761_),
    .Y(_0763_),
    .A1(_0685_),
    .A2(_0762_));
 sg13g2_a21o_1 _1684_ (.A2(_0719_),
    .A1(_0714_),
    .B1(_0718_),
    .X(_0764_));
 sg13g2_nor2b_1 _1685_ (.A(_0763_),
    .B_N(_0764_),
    .Y(_0765_));
 sg13g2_xnor2_1 _1686_ (.Y(_0766_),
    .A(_0763_),
    .B(_0764_));
 sg13g2_xor2_1 _1687_ (.B(_0766_),
    .A(net205),
    .X(_0767_));
 sg13g2_xnor2_1 _1688_ (.Y(_0768_),
    .A(_0760_),
    .B(_0767_));
 sg13g2_nor2_1 _1689_ (.A(_0759_),
    .B(_0768_),
    .Y(_0769_));
 sg13g2_xnor2_1 _1690_ (.Y(_0770_),
    .A(_0759_),
    .B(_0768_));
 sg13g2_xor2_1 _1691_ (.B(_0770_),
    .A(_0753_),
    .X(_0771_));
 sg13g2_nand2b_1 _1692_ (.Y(_0772_),
    .B(_0771_),
    .A_N(_0752_));
 sg13g2_xnor2_1 _1693_ (.Y(_0773_),
    .A(_0752_),
    .B(_0771_));
 sg13g2_and2_1 _1694_ (.A(_0751_),
    .B(_0773_),
    .X(_0774_));
 sg13g2_or2_1 _1695_ (.X(_0775_),
    .B(_0773_),
    .A(_0751_));
 sg13g2_xnor2_1 _1696_ (.Y(_0776_),
    .A(_0751_),
    .B(_0773_));
 sg13g2_xnor2_1 _1697_ (.Y(_0777_),
    .A(_0750_),
    .B(_0776_));
 sg13g2_and2_1 _1698_ (.A(_0749_),
    .B(_0777_),
    .X(_0778_));
 sg13g2_xor2_1 _1699_ (.B(_0777_),
    .A(_0749_),
    .X(_0779_));
 sg13g2_xnor2_1 _1700_ (.Y(_0780_),
    .A(_0023_),
    .B(_0779_));
 sg13g2_a21oi_1 _1701_ (.A1(_0003_),
    .A2(_0738_),
    .Y(_0781_),
    .B1(_0737_));
 sg13g2_nor2_1 _1702_ (.A(_0780_),
    .B(_0781_),
    .Y(_0782_));
 sg13g2_xor2_1 _1703_ (.B(_0781_),
    .A(_0780_),
    .X(_0783_));
 sg13g2_a21oi_1 _1704_ (.A1(_0744_),
    .A2(_0783_),
    .Y(_0784_),
    .B1(_0709_));
 sg13g2_o21ai_1 _1705_ (.B1(_0784_),
    .Y(_0785_),
    .A1(_0744_),
    .A2(_0783_));
 sg13g2_inv_1 _1706_ (.Y(_0062_),
    .A(_0785_));
 sg13g2_a21oi_1 _1707_ (.A1(_0744_),
    .A2(_0783_),
    .Y(_0786_),
    .B1(_0782_));
 sg13g2_a21oi_2 _1708_ (.B1(_0774_),
    .Y(_0787_),
    .A2(_0775_),
    .A1(_0750_));
 sg13g2_o21ai_1 _1709_ (.B1(_0772_),
    .Y(_0788_),
    .A1(_0753_),
    .A2(_0770_));
 sg13g2_o21ai_1 _1710_ (.B1(_0757_),
    .Y(_0789_),
    .A1(_0754_),
    .A2(_0755_));
 sg13g2_a21oi_1 _1711_ (.A1(_0760_),
    .A2(_0767_),
    .Y(_0790_),
    .B1(_0769_));
 sg13g2_nand2_1 _1712_ (.Y(_0791_),
    .A(net212),
    .B(_0236_));
 sg13g2_nor2_1 _1713_ (.A(_0762_),
    .B(_0791_),
    .Y(_0792_));
 sg13g2_xor2_1 _1714_ (.B(_0791_),
    .A(_0762_),
    .X(_0793_));
 sg13g2_a21oi_1 _1715_ (.A1(net205),
    .A2(_0766_),
    .Y(_0794_),
    .B1(_0765_));
 sg13g2_nor2b_1 _1716_ (.A(_0762_),
    .B_N(_0685_),
    .Y(_0795_));
 sg13g2_xnor2_1 _1717_ (.Y(_0796_),
    .A(_0756_),
    .B(_0795_));
 sg13g2_nor2b_1 _1718_ (.A(_0794_),
    .B_N(_0796_),
    .Y(_0797_));
 sg13g2_xnor2_1 _1719_ (.Y(_0798_),
    .A(_0794_),
    .B(_0796_));
 sg13g2_xnor2_1 _1720_ (.Y(_0799_),
    .A(_0793_),
    .B(_0798_));
 sg13g2_nor2_1 _1721_ (.A(_0790_),
    .B(_0799_),
    .Y(_0800_));
 sg13g2_xor2_1 _1722_ (.B(_0799_),
    .A(_0790_),
    .X(_0801_));
 sg13g2_xnor2_1 _1723_ (.Y(_0802_),
    .A(_0789_),
    .B(_0801_));
 sg13g2_nand2b_1 _1724_ (.Y(_0803_),
    .B(_0788_),
    .A_N(_0802_));
 sg13g2_xor2_1 _1725_ (.B(_0802_),
    .A(_0788_),
    .X(_0804_));
 sg13g2_xnor2_1 _1726_ (.Y(_0805_),
    .A(_0787_),
    .B(_0804_));
 sg13g2_nor2_1 _1727_ (.A(_0748_),
    .B(_0805_),
    .Y(_0806_));
 sg13g2_xnor2_1 _1728_ (.Y(_0807_),
    .A(_0747_),
    .B(_0805_));
 sg13g2_xnor2_1 _1729_ (.Y(_0808_),
    .A(_0002_),
    .B(_0807_));
 sg13g2_a21oi_1 _1730_ (.A1(_0023_),
    .A2(_0779_),
    .Y(_0809_),
    .B1(_0778_));
 sg13g2_or2_1 _1731_ (.X(_0810_),
    .B(_0809_),
    .A(_0808_));
 sg13g2_xnor2_1 _1732_ (.Y(_0811_),
    .A(_0808_),
    .B(_0809_));
 sg13g2_a21oi_1 _1733_ (.A1(_0786_),
    .A2(_0811_),
    .Y(_0812_),
    .B1(_0709_));
 sg13g2_o21ai_1 _1734_ (.B1(_0812_),
    .Y(_0813_),
    .A1(_0786_),
    .A2(_0811_));
 sg13g2_inv_1 _1735_ (.Y(_0063_),
    .A(_0813_));
 sg13g2_a21oi_1 _1736_ (.A1(_0789_),
    .A2(_0801_),
    .Y(_0814_),
    .B1(_0800_));
 sg13g2_a21oi_2 _1737_ (.B1(_0792_),
    .Y(_0815_),
    .A2(_0102_),
    .A1(net211));
 sg13g2_nand2_1 _1738_ (.Y(_0816_),
    .A(net212),
    .B(net208));
 sg13g2_xor2_1 _1739_ (.B(_0816_),
    .A(_0661_),
    .X(_0817_));
 sg13g2_xnor2_1 _1740_ (.Y(_0818_),
    .A(net202),
    .B(_0817_));
 sg13g2_a21oi_1 _1741_ (.A1(_0685_),
    .A2(_0756_),
    .Y(_0819_),
    .B1(_0762_));
 sg13g2_nor2b_1 _1742_ (.A(_0818_),
    .B_N(_0819_),
    .Y(_0820_));
 sg13g2_xor2_1 _1743_ (.B(_0819_),
    .A(_0818_),
    .X(_0821_));
 sg13g2_nand2_1 _1744_ (.Y(_0822_),
    .A(net207),
    .B(net208));
 sg13g2_nor2_1 _1745_ (.A(_0791_),
    .B(_0822_),
    .Y(_0823_));
 sg13g2_inv_1 _1746_ (.Y(_0824_),
    .A(_0823_));
 sg13g2_a22oi_1 _1747_ (.Y(_0825_),
    .B1(_0236_),
    .B2(net206),
    .A2(net208),
    .A1(net212));
 sg13g2_nor2_1 _1748_ (.A(_0823_),
    .B(_0825_),
    .Y(_0826_));
 sg13g2_nor2b_1 _1749_ (.A(_0821_),
    .B_N(_0826_),
    .Y(_0827_));
 sg13g2_xor2_1 _1750_ (.B(_0826_),
    .A(_0821_),
    .X(_0828_));
 sg13g2_a21oi_1 _1751_ (.A1(_0793_),
    .A2(_0798_),
    .Y(_0829_),
    .B1(_0797_));
 sg13g2_nor2_1 _1752_ (.A(_0828_),
    .B(_0829_),
    .Y(_0830_));
 sg13g2_xnor2_1 _1753_ (.Y(_0831_),
    .A(_0828_),
    .B(_0829_));
 sg13g2_nor2_1 _1754_ (.A(_0815_),
    .B(_0831_),
    .Y(_0832_));
 sg13g2_xnor2_1 _1755_ (.Y(_0833_),
    .A(_0815_),
    .B(_0831_));
 sg13g2_nor2_1 _1756_ (.A(_0814_),
    .B(_0833_),
    .Y(_0834_));
 sg13g2_o21ai_1 _1757_ (.B1(_0803_),
    .Y(_0835_),
    .A1(_0787_),
    .A2(_0804_));
 sg13g2_xor2_1 _1758_ (.B(_0833_),
    .A(_0814_),
    .X(_0836_));
 sg13g2_a21o_1 _1759_ (.A2(_0836_),
    .A1(_0835_),
    .B1(_0834_),
    .X(_0837_));
 sg13g2_nor2_1 _1760_ (.A(_0830_),
    .B(_0832_),
    .Y(_0838_));
 sg13g2_a21oi_1 _1761_ (.A1(net206),
    .A2(_0102_),
    .Y(_0839_),
    .B1(_0823_));
 sg13g2_and3_1 _1762_ (.X(_0840_),
    .A(net203),
    .B(_0817_),
    .C(_0839_));
 sg13g2_nor3_1 _1763_ (.A(_0820_),
    .B(_0827_),
    .C(_0840_),
    .Y(_0841_));
 sg13g2_nand2_1 _1764_ (.Y(_0842_),
    .A(_0827_),
    .B(_0840_));
 sg13g2_nand2b_1 _1765_ (.Y(_0843_),
    .B(_0842_),
    .A_N(_0841_));
 sg13g2_nor2_1 _1766_ (.A(_0838_),
    .B(_0843_),
    .Y(_0844_));
 sg13g2_xor2_1 _1767_ (.B(_0843_),
    .A(_0838_),
    .X(_0845_));
 sg13g2_xor2_1 _1768_ (.B(_0845_),
    .A(_0837_),
    .X(_0846_));
 sg13g2_and2_1 _1769_ (.A(net2),
    .B(_0846_),
    .X(_0847_));
 sg13g2_xor2_1 _1770_ (.B(_0846_),
    .A(net2),
    .X(_0848_));
 sg13g2_a21o_1 _1771_ (.A2(_0848_),
    .A1(_0021_),
    .B1(_0847_),
    .X(_0849_));
 sg13g2_a21oi_1 _1772_ (.A1(_0837_),
    .A2(_0845_),
    .Y(_0850_),
    .B1(_0844_));
 sg13g2_a221oi_1 _1773_ (.B2(net203),
    .C1(_0823_),
    .B1(_0817_),
    .A1(net207),
    .Y(_0851_),
    .A2(_0102_));
 sg13g2_o21ai_1 _1774_ (.B1(_0824_),
    .Y(_0852_),
    .A1(_0103_),
    .A2(_0851_));
 sg13g2_nand2_1 _1775_ (.Y(_0853_),
    .A(_0103_),
    .B(_0822_));
 sg13g2_nand2_1 _1776_ (.Y(_0854_),
    .A(_0851_),
    .B(_0853_));
 sg13g2_o21ai_1 _1777_ (.B1(_0854_),
    .Y(_0855_),
    .A1(_0101_),
    .A2(_0661_));
 sg13g2_xnor2_1 _1778_ (.Y(_0856_),
    .A(_0001_),
    .B(_0855_));
 sg13g2_xnor2_1 _1779_ (.Y(_0857_),
    .A(_0852_),
    .B(_0856_));
 sg13g2_nand2_1 _1780_ (.Y(_0858_),
    .A(_0839_),
    .B(_0842_));
 sg13g2_inv_1 _1781_ (.Y(_0859_),
    .A(_0858_));
 sg13g2_xnor2_1 _1782_ (.Y(_0860_),
    .A(_0857_),
    .B(_0858_));
 sg13g2_nand2b_1 _1783_ (.Y(_0861_),
    .B(_0860_),
    .A_N(_0850_));
 sg13g2_xnor2_1 _1784_ (.Y(_0862_),
    .A(_0850_),
    .B(_0860_));
 sg13g2_and2_1 _1785_ (.A(net3),
    .B(_0862_),
    .X(_0863_));
 sg13g2_xor2_1 _1786_ (.B(_0862_),
    .A(net3),
    .X(_0864_));
 sg13g2_xnor2_1 _1787_ (.Y(_0865_),
    .A(_0020_),
    .B(_0864_));
 sg13g2_nor2b_1 _1788_ (.A(_0865_),
    .B_N(_0849_),
    .Y(_0866_));
 sg13g2_xor2_1 _1789_ (.B(_0836_),
    .A(_0835_),
    .X(_0867_));
 sg13g2_and2_1 _1790_ (.A(net1),
    .B(_0867_),
    .X(_0868_));
 sg13g2_xor2_1 _1791_ (.B(_0867_),
    .A(net1),
    .X(_0869_));
 sg13g2_a21oi_1 _1792_ (.A1(_0022_),
    .A2(_0869_),
    .Y(_0870_),
    .B1(_0868_));
 sg13g2_xnor2_1 _1793_ (.Y(_0871_),
    .A(_0021_),
    .B(_0848_));
 sg13g2_or2_1 _1794_ (.X(_0872_),
    .B(_0871_),
    .A(_0870_));
 sg13g2_a21oi_1 _1795_ (.A1(_0002_),
    .A2(_0807_),
    .Y(_0873_),
    .B1(_0806_));
 sg13g2_xnor2_1 _1796_ (.Y(_0874_),
    .A(_0022_),
    .B(_0869_));
 sg13g2_nor2_1 _1797_ (.A(_0873_),
    .B(_0874_),
    .Y(_0875_));
 sg13g2_o21ai_1 _1798_ (.B1(_0810_),
    .Y(_0876_),
    .A1(_0786_),
    .A2(_0811_));
 sg13g2_xor2_1 _1799_ (.B(_0874_),
    .A(_0873_),
    .X(_0877_));
 sg13g2_a21oi_1 _1800_ (.A1(_0876_),
    .A2(_0877_),
    .Y(_0878_),
    .B1(_0875_));
 sg13g2_xnor2_1 _1801_ (.Y(_0879_),
    .A(_0870_),
    .B(_0871_));
 sg13g2_o21ai_1 _1802_ (.B1(_0872_),
    .Y(_0880_),
    .A1(_0878_),
    .A2(_0879_));
 sg13g2_xnor2_1 _1803_ (.Y(_0881_),
    .A(_0849_),
    .B(_0865_));
 sg13g2_a21oi_1 _1804_ (.A1(_0880_),
    .A2(_0881_),
    .Y(_0882_),
    .B1(_0866_));
 sg13g2_a21oi_1 _1805_ (.A1(_0020_),
    .A2(_0864_),
    .Y(_0883_),
    .B1(_0863_));
 sg13g2_o21ai_1 _1806_ (.B1(_0861_),
    .Y(_0884_),
    .A1(_0857_),
    .A2(_0859_));
 sg13g2_nor2_1 _1807_ (.A(_0001_),
    .B(_0854_),
    .Y(_0885_));
 sg13g2_a21oi_1 _1808_ (.A1(_0852_),
    .A2(_0856_),
    .Y(_0886_),
    .B1(_0885_));
 sg13g2_nor2_1 _1809_ (.A(_0001_),
    .B(_0661_),
    .Y(_0887_));
 sg13g2_nor2_1 _1810_ (.A(_0101_),
    .B(_0887_),
    .Y(_0888_));
 sg13g2_xor2_1 _1811_ (.B(net4),
    .A(\izh_1.u[7] ),
    .X(_0889_));
 sg13g2_xnor2_1 _1812_ (.Y(_0890_),
    .A(_0888_),
    .B(_0889_));
 sg13g2_xnor2_1 _1813_ (.Y(_0891_),
    .A(_0886_),
    .B(_0890_));
 sg13g2_xnor2_1 _1814_ (.Y(_0892_),
    .A(_0884_),
    .B(_0891_));
 sg13g2_xnor2_1 _1815_ (.Y(_0893_),
    .A(_0883_),
    .B(_0892_));
 sg13g2_xnor2_1 _1816_ (.Y(_0894_),
    .A(_0882_),
    .B(_0893_));
 sg13g2_nor2_1 _1817_ (.A(_0709_),
    .B(_0894_),
    .Y(_0064_));
 sg13g2_nand2_1 _1818_ (.Y(_0895_),
    .A(net195),
    .B(_0311_));
 sg13g2_xor2_1 _1819_ (.B(_0895_),
    .A(net91),
    .X(_0896_));
 sg13g2_nor2_1 _1820_ (.A(net244),
    .B(_0896_),
    .Y(_0065_));
 sg13g2_xnor2_1 _1821_ (.Y(_0897_),
    .A(_0312_),
    .B(_0315_));
 sg13g2_o21ai_1 _1822_ (.B1(net248),
    .Y(_0898_),
    .A1(net85),
    .A2(net196));
 sg13g2_a21oi_1 _1823_ (.A1(net196),
    .A2(_0897_),
    .Y(_0066_),
    .B1(_0898_));
 sg13g2_xnor2_1 _1824_ (.Y(_0899_),
    .A(_0316_),
    .B(_0319_));
 sg13g2_o21ai_1 _1825_ (.B1(net247),
    .Y(_0900_),
    .A1(net64),
    .A2(net198));
 sg13g2_a21oi_1 _1826_ (.A1(net198),
    .A2(_0899_),
    .Y(_0067_),
    .B1(_0900_));
 sg13g2_nand4_1 _1827_ (.B(_0320_),
    .C(_0321_),
    .A(_0307_),
    .Y(_0901_),
    .D(_0322_));
 sg13g2_nand2b_1 _1828_ (.Y(_0902_),
    .B(_0901_),
    .A_N(_0323_));
 sg13g2_o21ai_1 _1829_ (.B1(net248),
    .Y(_0903_),
    .A1(net68),
    .A2(net197));
 sg13g2_a21oi_1 _1830_ (.A1(net197),
    .A2(_0902_),
    .Y(_0068_),
    .B1(_0903_));
 sg13g2_xnor2_1 _1831_ (.Y(_0904_),
    .A(_0324_),
    .B(_0325_));
 sg13g2_o21ai_1 _1832_ (.B1(net247),
    .Y(_0905_),
    .A1(net84),
    .A2(net197));
 sg13g2_a21oi_1 _1833_ (.A1(net197),
    .A2(_0904_),
    .Y(_0069_),
    .B1(_0905_));
 sg13g2_xnor2_1 _1834_ (.Y(_0906_),
    .A(_0326_),
    .B(_0327_));
 sg13g2_o21ai_1 _1835_ (.B1(net247),
    .Y(_0907_),
    .A1(net67),
    .A2(net197));
 sg13g2_a21oi_1 _1836_ (.A1(net197),
    .A2(_0906_),
    .Y(_0070_),
    .B1(_0907_));
 sg13g2_xnor2_1 _1837_ (.Y(_0908_),
    .A(_0328_),
    .B(_0329_));
 sg13g2_o21ai_1 _1838_ (.B1(net247),
    .Y(_0909_),
    .A1(net70),
    .A2(net196));
 sg13g2_a21oi_1 _1839_ (.A1(net196),
    .A2(_0908_),
    .Y(_0071_),
    .B1(_0909_));
 sg13g2_xnor2_1 _1840_ (.Y(_0077_),
    .A(_0330_),
    .B(_0331_));
 sg13g2_o21ai_1 _1841_ (.B1(net247),
    .Y(_0078_),
    .A1(net104),
    .A2(net198));
 sg13g2_a21oi_1 _1842_ (.A1(net196),
    .A2(_0077_),
    .Y(_0072_),
    .B1(_0078_));
 sg13g2_xnor2_1 _1843_ (.Y(_0079_),
    .A(_0332_),
    .B(_0333_));
 sg13g2_o21ai_1 _1844_ (.B1(net247),
    .Y(_0080_),
    .A1(net69),
    .A2(net196));
 sg13g2_a21oi_1 _1845_ (.A1(net196),
    .A2(_0079_),
    .Y(_0073_),
    .B1(_0080_));
 sg13g2_xnor2_1 _1846_ (.Y(_0081_),
    .A(_0876_),
    .B(_0877_));
 sg13g2_a21oi_1 _1847_ (.A1(net198),
    .A2(_0081_),
    .Y(_0074_),
    .B1(net244));
 sg13g2_xnor2_1 _1848_ (.Y(_0082_),
    .A(_0878_),
    .B(_0879_));
 sg13g2_a21oi_1 _1849_ (.A1(net197),
    .A2(_0082_),
    .Y(_0075_),
    .B1(net244));
 sg13g2_xnor2_1 _1850_ (.Y(_0083_),
    .A(_0880_),
    .B(_0881_));
 sg13g2_a21oi_1 _1851_ (.A1(net197),
    .A2(_0083_),
    .Y(_0076_),
    .B1(net243));
 sg13g2_dfrbp_1 _1852_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net55),
    .D(_0031_),
    .Q_N(_0011_),
    .Q(\izh_2.u[9] ));
 sg13g2_dfrbp_1 _1853_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net36),
    .D(net74),
    .Q_N(_0010_),
    .Q(\izh_2.u[10] ));
 sg13g2_dfrbp_1 _1854_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net35),
    .D(_0033_),
    .Q_N(_0012_),
    .Q(\izh_2.u[11] ));
 sg13g2_dfrbp_1 _1855_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net34),
    .D(net60),
    .Q_N(_0014_),
    .Q(\izh_2.u[12] ));
 sg13g2_dfrbp_1 _1856_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net33),
    .D(net90),
    .Q_N(_0013_),
    .Q(\izh_2.u[13] ));
 sg13g2_dfrbp_1 _1857_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net32),
    .D(_0036_),
    .Q_N(_0924_),
    .Q(\izh_2.u[14] ));
 sg13g2_dfrbp_1 _1858_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net31),
    .D(_0037_),
    .Q_N(_0027_),
    .Q(\izh_1.u[9] ));
 sg13g2_dfrbp_1 _1859_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net30),
    .D(net79),
    .Q_N(_0026_),
    .Q(\izh_1.u[10] ));
 sg13g2_dfrbp_1 _1860_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net29),
    .D(net100),
    .Q_N(_0028_),
    .Q(\izh_1.u[11] ));
 sg13g2_dfrbp_1 _1861_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net28),
    .D(net58),
    .Q_N(_0030_),
    .Q(\izh_1.u[12] ));
 sg13g2_dfrbp_1 _1862_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net27),
    .D(net82),
    .Q_N(_0029_),
    .Q(\izh_1.u[13] ));
 sg13g2_dfrbp_1 _1863_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net26),
    .D(_0042_),
    .Q_N(_0923_),
    .Q(\izh_1.u[14] ));
 sg13g2_dfrbp_1 _1864_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net25),
    .D(_0043_),
    .Q_N(_0922_),
    .Q(net241));
 sg13g2_dfrbp_1 _1865_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net24),
    .D(_0044_),
    .Q_N(_0921_),
    .Q(net239));
 sg13g2_dfrbp_1 _1866_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net23),
    .D(_0045_),
    .Q_N(_0920_),
    .Q(net237));
 sg13g2_dfrbp_1 _1867_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net22),
    .D(_0046_),
    .Q_N(_0919_),
    .Q(net234));
 sg13g2_dfrbp_1 _1868_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net21),
    .D(_0047_),
    .Q_N(_0918_),
    .Q(net231));
 sg13g2_dfrbp_1 _1869_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net20),
    .D(_0048_),
    .Q_N(_0917_),
    .Q(\izh_2.u[0] ));
 sg13g2_dfrbp_1 _1870_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net18),
    .D(_0049_),
    .Q_N(_0018_),
    .Q(\izh_2.u[1] ));
 sg13g2_dfrbp_1 _1871_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net16),
    .D(_0050_),
    .Q_N(_0007_),
    .Q(\izh_2.u[2] ));
 sg13g2_dfrbp_1 _1872_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net14),
    .D(net77),
    .Q_N(_0017_),
    .Q(\izh_2.u[3] ));
 sg13g2_dfrbp_1 _1873_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net12),
    .D(_0052_),
    .Q_N(_0006_),
    .Q(\izh_2.u[4] ));
 sg13g2_dfrbp_1 _1874_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net56),
    .D(_0053_),
    .Q_N(_0005_),
    .Q(\izh_2.u[5] ));
 sg13g2_dfrbp_1 _1875_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net54),
    .D(_0054_),
    .Q_N(_0004_),
    .Q(\izh_2.u[6] ));
 sg13g2_dfrbp_1 _1876_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net52),
    .D(net98),
    .Q_N(_0009_),
    .Q(\izh_2.u[7] ));
 sg13g2_dfrbp_1 _1877_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net50),
    .D(_0056_),
    .Q_N(_0008_),
    .Q(\izh_2.u[8] ));
 sg13g2_dfrbp_1 _1878_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net48),
    .D(_0057_),
    .Q_N(_0916_),
    .Q(net229));
 sg13g2_dfrbp_1 _1879_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net47),
    .D(_0058_),
    .Q_N(_0015_),
    .Q(net223));
 sg13g2_dfrbp_1 _1880_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net46),
    .D(_0059_),
    .Q_N(_0016_),
    .Q(net221));
 sg13g2_dfrbp_1 _1881_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net45),
    .D(_0060_),
    .Q_N(_0915_),
    .Q(net218));
 sg13g2_dfrbp_1 _1882_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net44),
    .D(_0061_),
    .Q_N(_0019_),
    .Q(net216));
 sg13g2_dfrbp_1 _1883_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net43),
    .D(_0062_),
    .Q_N(_0914_),
    .Q(net214));
 sg13g2_dfrbp_1 _1884_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net42),
    .D(_0063_),
    .Q_N(_0000_),
    .Q(net213));
 sg13g2_dfrbp_1 _1885_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net41),
    .D(_0064_),
    .Q_N(_0913_),
    .Q(net210));
 sg13g2_dfrbp_1 _1886_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net40),
    .D(_0065_),
    .Q_N(_0912_),
    .Q(\izh_1.u[0] ));
 sg13g2_dfrbp_1 _1887_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net38),
    .D(net86),
    .Q_N(_0003_),
    .Q(\izh_1.u[1] ));
 sg13g2_dfrbp_1 _1888_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net19),
    .D(_0067_),
    .Q_N(_0023_),
    .Q(\izh_1.u[2] ));
 sg13g2_dfrbp_1 _1889_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net15),
    .D(_0068_),
    .Q_N(_0002_),
    .Q(\izh_1.u[3] ));
 sg13g2_dfrbp_1 _1890_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net11),
    .D(_0069_),
    .Q_N(_0022_),
    .Q(\izh_1.u[4] ));
 sg13g2_dfrbp_1 _1891_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net53),
    .D(_0070_),
    .Q_N(_0021_),
    .Q(\izh_1.u[5] ));
 sg13g2_dfrbp_1 _1892_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net49),
    .D(net71),
    .Q_N(_0020_),
    .Q(\izh_1.u[6] ));
 sg13g2_dfrbp_1 _1893_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net37),
    .D(net105),
    .Q_N(_0025_),
    .Q(\izh_1.u[7] ));
 sg13g2_dfrbp_1 _1894_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net13),
    .D(_0073_),
    .Q_N(_0024_),
    .Q(\izh_1.u[8] ));
 sg13g2_dfrbp_1 _1895_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net51),
    .D(_0074_),
    .Q_N(_0911_),
    .Q(net204));
 sg13g2_dfrbp_1 _1896_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net39),
    .D(_0075_),
    .Q_N(_0910_),
    .Q(net201));
 sg13g2_dfrbp_1 _1897_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net17),
    .D(_0076_),
    .Q_N(_0001_),
    .Q(net199));
 sg13g2_tiehi _1873__12 (.L_HI(net12));
 sg13g2_tiehi _1894__13 (.L_HI(net13));
 sg13g2_tiehi _1872__14 (.L_HI(net14));
 sg13g2_tiehi _1889__15 (.L_HI(net15));
 sg13g2_tiehi _1871__16 (.L_HI(net16));
 sg13g2_tiehi _1897__17 (.L_HI(net17));
 sg13g2_tiehi _1870__18 (.L_HI(net18));
 sg13g2_tiehi _1888__19 (.L_HI(net19));
 sg13g2_tiehi _1869__20 (.L_HI(net20));
 sg13g2_tiehi _1868__21 (.L_HI(net21));
 sg13g2_tiehi _1867__22 (.L_HI(net22));
 sg13g2_tiehi _1866__23 (.L_HI(net23));
 sg13g2_tiehi _1865__24 (.L_HI(net24));
 sg13g2_tiehi _1864__25 (.L_HI(net25));
 sg13g2_tiehi _1863__26 (.L_HI(net26));
 sg13g2_tiehi _1862__27 (.L_HI(net27));
 sg13g2_tiehi _1861__28 (.L_HI(net28));
 sg13g2_tiehi _1860__29 (.L_HI(net29));
 sg13g2_tiehi _1859__30 (.L_HI(net30));
 sg13g2_tiehi _1858__31 (.L_HI(net31));
 sg13g2_tiehi _1857__32 (.L_HI(net32));
 sg13g2_tiehi _1856__33 (.L_HI(net33));
 sg13g2_tiehi _1855__34 (.L_HI(net34));
 sg13g2_tiehi _1854__35 (.L_HI(net35));
 sg13g2_tiehi _1853__36 (.L_HI(net36));
 sg13g2_tiehi _1893__37 (.L_HI(net37));
 sg13g2_tiehi _1887__38 (.L_HI(net38));
 sg13g2_tiehi _1896__39 (.L_HI(net39));
 sg13g2_tiehi _1886__40 (.L_HI(net40));
 sg13g2_tiehi _1885__41 (.L_HI(net41));
 sg13g2_tiehi _1884__42 (.L_HI(net42));
 sg13g2_tiehi _1883__43 (.L_HI(net43));
 sg13g2_tiehi _1882__44 (.L_HI(net44));
 sg13g2_tiehi _1881__45 (.L_HI(net45));
 sg13g2_tiehi _1880__46 (.L_HI(net46));
 sg13g2_tiehi _1879__47 (.L_HI(net47));
 sg13g2_tiehi _1878__48 (.L_HI(net48));
 sg13g2_tiehi _1892__49 (.L_HI(net49));
 sg13g2_tiehi _1877__50 (.L_HI(net50));
 sg13g2_tiehi _1895__51 (.L_HI(net51));
 sg13g2_tiehi _1876__52 (.L_HI(net52));
 sg13g2_tiehi _1891__53 (.L_HI(net53));
 sg13g2_tiehi _1875__54 (.L_HI(net54));
 sg13g2_tiehi _1852__55 (.L_HI(net55));
 sg13g2_tiehi _1874__56 (.L_HI(net56));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_nomuwill_6 (.L_LO(net6));
 sg13g2_tielo tt_um_nomuwill_7 (.L_LO(net7));
 sg13g2_tielo tt_um_nomuwill_8 (.L_LO(net8));
 sg13g2_tielo tt_um_nomuwill_9 (.L_LO(net9));
 sg13g2_tielo tt_um_nomuwill_10 (.L_LO(net10));
 sg13g2_tiehi _1890__11 (.L_HI(net11));
 sg13g2_buf_2 _1950_ (.A(\izh_2.spike ),
    .X(uio_out[6]));
 sg13g2_buf_2 _1951_ (.A(\izh_1.spike ),
    .X(uio_out[7]));
 sg13g2_buf_2 fanout191 (.A(net192),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_0108_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(net194),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_0108_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(net196),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(net198),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(net198),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_0104_),
    .X(net198));
 sg13g2_buf_4 fanout199 (.X(uo_out[6]),
    .A(net199));
 sg13g2_buf_2 fanout200 (.A(net199),
    .X(net200));
 sg13g2_buf_4 fanout201 (.X(uo_out[5]),
    .A(net203));
 sg13g2_buf_2 fanout202 (.A(net203),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(net201),
    .X(net203));
 sg13g2_buf_4 fanout204 (.X(uo_out[4]),
    .A(net207));
 sg13g2_buf_1 fanout205 (.A(net207),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(net207),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(net204),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(net209),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(uo_out[7]),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(net210),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout211 (.X(net211),
    .A(uo_out[3]));
 sg13g2_buf_1 fanout212 (.A(uo_out[3]),
    .X(net212));
 sg13g2_buf_4 fanout213 (.X(uo_out[3]),
    .A(net213));
 sg13g2_buf_4 fanout214 (.X(uo_out[2]),
    .A(net214));
 sg13g2_buf_2 fanout215 (.A(net214),
    .X(net215));
 sg13g2_buf_4 fanout216 (.X(uo_out[1]),
    .A(net217));
 sg13g2_buf_2 fanout217 (.A(net216),
    .X(net217));
 sg13g2_buf_4 fanout218 (.X(uo_out[0]),
    .A(net220));
 sg13g2_buf_1 fanout219 (.A(net220),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(net218),
    .X(net220));
 sg13g2_buf_4 fanout221 (.X(uio_oe[6]),
    .A(net221));
 sg13g2_buf_4 fanout222 (.X(net222),
    .A(net221));
 sg13g2_buf_4 fanout223 (.X(uio_oe[5]),
    .A(net223));
 sg13g2_buf_2 fanout224 (.A(net225),
    .X(net224));
 sg13g2_buf_1 fanout225 (.A(net223),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(net229),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(net229),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(uio_oe[4]),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(net229),
    .X(uio_oe[4]));
 sg13g2_buf_2 fanout230 (.A(net231),
    .X(net230));
 sg13g2_buf_4 fanout231 (.X(uio_oe[7]),
    .A(net231));
 sg13g2_buf_4 fanout232 (.X(net232),
    .A(uio_oe[3]));
 sg13g2_buf_1 fanout233 (.A(uio_oe[3]),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(net234),
    .X(uio_oe[3]));
 sg13g2_buf_2 fanout235 (.A(net238),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(net238),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(net238),
    .X(uio_oe[2]));
 sg13g2_buf_2 fanout238 (.A(net237),
    .X(net238));
 sg13g2_buf_4 fanout239 (.X(uio_oe[1]),
    .A(net240));
 sg13g2_buf_2 fanout240 (.A(net239),
    .X(net240));
 sg13g2_buf_4 fanout241 (.X(uio_oe[0]),
    .A(net241));
 sg13g2_buf_2 fanout242 (.A(net241),
    .X(net242));
 sg13g2_buf_4 fanout243 (.X(net243),
    .A(_0091_));
 sg13g2_buf_2 fanout244 (.A(_0091_),
    .X(net244));
 sg13g2_buf_4 fanout245 (.X(net245),
    .A(rst_n));
 sg13g2_buf_1 fanout246 (.A(rst_n),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(net248),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(rst_n),
    .X(net248));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_tielo tt_um_nomuwill_5 (.L_LO(net5));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0030_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0040_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0014_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0034_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0011_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0210_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0027_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold8 (.A(\izh_1.u[2] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold9 (.A(\izh_2.u[2] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold10 (.A(\izh_2.u[8] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold11 (.A(\izh_1.u[5] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold12 (.A(\izh_1.u[3] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold13 (.A(\izh_1.u[8] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold14 (.A(\izh_1.u[6] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0071_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold16 (.A(\izh_2.u[4] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0010_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0032_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold19 (.A(\izh_2.u[6] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold20 (.A(\izh_2.u[3] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0051_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0026_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0038_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0029_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0358_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0041_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold27 (.A(\izh_2.u[5] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold28 (.A(\izh_1.u[4] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold29 (.A(\izh_1.u[1] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0066_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold31 (.A(\izh_2.u[1] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0013_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0232_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0035_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold35 (.A(\izh_1.u[0] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold36 (.A(\izh_2.u[0] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold37 (.A(\izh_1.u[14] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0361_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold39 (.A(\izh_2.u[14] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0235_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold41 (.A(\izh_2.u[7] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0055_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0028_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0039_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold45 (.A(\izh_2.u[11] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0217_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0221_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold48 (.A(\izh_1.u[7] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0072_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold50 (.A(\izh_2.u[0] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold51 (.A(\izh_1.u[0] ),
    .X(net107));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_4 FILLER_12_315 ();
 sg13g2_decap_4 FILLER_12_324 ();
 sg13g2_fill_1 FILLER_12_328 ();
 sg13g2_decap_8 FILLER_12_334 ();
 sg13g2_decap_4 FILLER_12_341 ();
 sg13g2_fill_2 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_4 FILLER_13_259 ();
 sg13g2_fill_2 FILLER_13_263 ();
 sg13g2_fill_1 FILLER_13_298 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_4 FILLER_14_126 ();
 sg13g2_fill_2 FILLER_14_130 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_fill_1 FILLER_14_151 ();
 sg13g2_decap_4 FILLER_14_175 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_decap_4 FILLER_14_185 ();
 sg13g2_fill_1 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_194 ();
 sg13g2_decap_8 FILLER_14_201 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_215 ();
 sg13g2_decap_8 FILLER_14_222 ();
 sg13g2_decap_8 FILLER_14_229 ();
 sg13g2_decap_8 FILLER_14_236 ();
 sg13g2_decap_8 FILLER_14_243 ();
 sg13g2_decap_8 FILLER_14_250 ();
 sg13g2_decap_8 FILLER_14_257 ();
 sg13g2_fill_2 FILLER_14_323 ();
 sg13g2_fill_2 FILLER_14_334 ();
 sg13g2_fill_1 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_fill_1 FILLER_15_91 ();
 sg13g2_fill_2 FILLER_15_123 ();
 sg13g2_fill_1 FILLER_15_138 ();
 sg13g2_fill_2 FILLER_15_169 ();
 sg13g2_fill_1 FILLER_15_171 ();
 sg13g2_decap_8 FILLER_15_207 ();
 sg13g2_decap_8 FILLER_15_214 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_decap_8 FILLER_15_242 ();
 sg13g2_fill_2 FILLER_15_249 ();
 sg13g2_fill_2 FILLER_15_264 ();
 sg13g2_fill_1 FILLER_15_266 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_326 ();
 sg13g2_decap_4 FILLER_15_348 ();
 sg13g2_fill_2 FILLER_15_352 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_fill_2 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_93 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_fill_2 FILLER_16_155 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_decap_4 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_215 ();
 sg13g2_decap_8 FILLER_16_222 ();
 sg13g2_decap_8 FILLER_16_229 ();
 sg13g2_decap_4 FILLER_16_236 ();
 sg13g2_fill_2 FILLER_16_286 ();
 sg13g2_fill_1 FILLER_16_288 ();
 sg13g2_decap_4 FILLER_16_300 ();
 sg13g2_decap_4 FILLER_16_312 ();
 sg13g2_fill_1 FILLER_16_316 ();
 sg13g2_decap_4 FILLER_16_322 ();
 sg13g2_fill_1 FILLER_16_339 ();
 sg13g2_fill_2 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_fill_2 FILLER_17_63 ();
 sg13g2_fill_1 FILLER_17_65 ();
 sg13g2_fill_1 FILLER_17_92 ();
 sg13g2_decap_4 FILLER_17_96 ();
 sg13g2_fill_2 FILLER_17_100 ();
 sg13g2_fill_1 FILLER_17_123 ();
 sg13g2_fill_2 FILLER_17_137 ();
 sg13g2_fill_1 FILLER_17_162 ();
 sg13g2_fill_2 FILLER_17_180 ();
 sg13g2_fill_1 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_239 ();
 sg13g2_fill_2 FILLER_17_246 ();
 sg13g2_fill_1 FILLER_17_248 ();
 sg13g2_fill_2 FILLER_17_253 ();
 sg13g2_decap_4 FILLER_17_264 ();
 sg13g2_fill_2 FILLER_17_287 ();
 sg13g2_fill_1 FILLER_17_289 ();
 sg13g2_fill_1 FILLER_17_298 ();
 sg13g2_decap_4 FILLER_17_310 ();
 sg13g2_fill_2 FILLER_17_349 ();
 sg13g2_fill_1 FILLER_17_351 ();
 sg13g2_decap_4 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_4 FILLER_18_42 ();
 sg13g2_fill_2 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_57 ();
 sg13g2_fill_1 FILLER_18_59 ();
 sg13g2_decap_8 FILLER_18_65 ();
 sg13g2_fill_2 FILLER_18_72 ();
 sg13g2_decap_4 FILLER_18_125 ();
 sg13g2_fill_2 FILLER_18_129 ();
 sg13g2_fill_2 FILLER_18_165 ();
 sg13g2_fill_1 FILLER_18_167 ();
 sg13g2_fill_2 FILLER_18_214 ();
 sg13g2_fill_2 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_294 ();
 sg13g2_decap_4 FILLER_18_311 ();
 sg13g2_fill_2 FILLER_18_315 ();
 sg13g2_fill_2 FILLER_18_322 ();
 sg13g2_fill_1 FILLER_18_324 ();
 sg13g2_fill_1 FILLER_18_329 ();
 sg13g2_fill_2 FILLER_18_338 ();
 sg13g2_fill_1 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_61 ();
 sg13g2_decap_4 FILLER_19_75 ();
 sg13g2_fill_2 FILLER_19_79 ();
 sg13g2_fill_2 FILLER_19_106 ();
 sg13g2_fill_1 FILLER_19_108 ();
 sg13g2_fill_1 FILLER_19_131 ();
 sg13g2_fill_1 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_173 ();
 sg13g2_fill_1 FILLER_19_175 ();
 sg13g2_fill_2 FILLER_19_300 ();
 sg13g2_decap_8 FILLER_19_320 ();
 sg13g2_fill_2 FILLER_19_334 ();
 sg13g2_fill_1 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_fill_2 FILLER_19_357 ();
 sg13g2_fill_2 FILLER_19_369 ();
 sg13g2_fill_1 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_fill_1 FILLER_20_45 ();
 sg13g2_decap_8 FILLER_20_50 ();
 sg13g2_fill_1 FILLER_20_57 ();
 sg13g2_fill_2 FILLER_20_75 ();
 sg13g2_fill_2 FILLER_20_80 ();
 sg13g2_fill_1 FILLER_20_82 ();
 sg13g2_fill_2 FILLER_20_103 ();
 sg13g2_fill_2 FILLER_20_110 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_decap_4 FILLER_20_157 ();
 sg13g2_fill_1 FILLER_20_161 ();
 sg13g2_fill_2 FILLER_20_178 ();
 sg13g2_fill_1 FILLER_20_184 ();
 sg13g2_fill_2 FILLER_20_211 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_238 ();
 sg13g2_fill_1 FILLER_20_243 ();
 sg13g2_fill_2 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_303 ();
 sg13g2_fill_2 FILLER_20_330 ();
 sg13g2_fill_2 FILLER_20_357 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_fill_1 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_4 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_18 ();
 sg13g2_fill_1 FILLER_21_49 ();
 sg13g2_decap_4 FILLER_21_66 ();
 sg13g2_fill_2 FILLER_21_91 ();
 sg13g2_fill_2 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_100 ();
 sg13g2_decap_8 FILLER_21_116 ();
 sg13g2_decap_4 FILLER_21_123 ();
 sg13g2_fill_2 FILLER_21_127 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_fill_2 FILLER_21_139 ();
 sg13g2_fill_1 FILLER_21_141 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_decap_4 FILLER_21_158 ();
 sg13g2_fill_1 FILLER_21_162 ();
 sg13g2_fill_2 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_216 ();
 sg13g2_decap_4 FILLER_21_223 ();
 sg13g2_fill_1 FILLER_21_227 ();
 sg13g2_fill_1 FILLER_21_254 ();
 sg13g2_fill_1 FILLER_21_285 ();
 sg13g2_decap_4 FILLER_21_304 ();
 sg13g2_decap_4 FILLER_21_317 ();
 sg13g2_decap_4 FILLER_21_334 ();
 sg13g2_fill_1 FILLER_21_346 ();
 sg13g2_fill_2 FILLER_21_360 ();
 sg13g2_fill_2 FILLER_21_369 ();
 sg13g2_decap_4 FILLER_21_389 ();
 sg13g2_fill_1 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_19 ();
 sg13g2_fill_2 FILLER_22_26 ();
 sg13g2_fill_1 FILLER_22_28 ();
 sg13g2_fill_2 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_44 ();
 sg13g2_fill_2 FILLER_22_62 ();
 sg13g2_fill_1 FILLER_22_64 ();
 sg13g2_fill_2 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_4 FILLER_22_102 ();
 sg13g2_fill_2 FILLER_22_106 ();
 sg13g2_fill_1 FILLER_22_122 ();
 sg13g2_fill_1 FILLER_22_138 ();
 sg13g2_decap_4 FILLER_22_155 ();
 sg13g2_fill_1 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_189 ();
 sg13g2_decap_4 FILLER_22_226 ();
 sg13g2_fill_1 FILLER_22_230 ();
 sg13g2_fill_2 FILLER_22_249 ();
 sg13g2_fill_1 FILLER_22_251 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_fill_2 FILLER_22_311 ();
 sg13g2_fill_1 FILLER_22_313 ();
 sg13g2_fill_1 FILLER_22_330 ();
 sg13g2_fill_2 FILLER_22_358 ();
 sg13g2_decap_4 FILLER_22_370 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_30 ();
 sg13g2_fill_2 FILLER_23_37 ();
 sg13g2_fill_1 FILLER_23_39 ();
 sg13g2_fill_2 FILLER_23_71 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_fill_2 FILLER_23_165 ();
 sg13g2_fill_1 FILLER_23_167 ();
 sg13g2_fill_1 FILLER_23_173 ();
 sg13g2_decap_4 FILLER_23_200 ();
 sg13g2_fill_1 FILLER_23_204 ();
 sg13g2_fill_1 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_215 ();
 sg13g2_decap_4 FILLER_23_222 ();
 sg13g2_fill_2 FILLER_23_226 ();
 sg13g2_fill_2 FILLER_23_245 ();
 sg13g2_fill_1 FILLER_23_247 ();
 sg13g2_fill_1 FILLER_23_274 ();
 sg13g2_fill_2 FILLER_23_286 ();
 sg13g2_fill_1 FILLER_23_288 ();
 sg13g2_fill_2 FILLER_23_298 ();
 sg13g2_fill_2 FILLER_23_313 ();
 sg13g2_fill_1 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_fill_2 FILLER_23_334 ();
 sg13g2_fill_1 FILLER_23_341 ();
 sg13g2_fill_1 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_20 ();
 sg13g2_decap_4 FILLER_24_74 ();
 sg13g2_fill_2 FILLER_24_78 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_fill_2 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_100 ();
 sg13g2_decap_4 FILLER_24_145 ();
 sg13g2_fill_1 FILLER_24_149 ();
 sg13g2_fill_2 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_172 ();
 sg13g2_fill_1 FILLER_24_179 ();
 sg13g2_decap_4 FILLER_24_196 ();
 sg13g2_fill_1 FILLER_24_200 ();
 sg13g2_fill_2 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_decap_8 FILLER_24_258 ();
 sg13g2_decap_8 FILLER_24_265 ();
 sg13g2_fill_1 FILLER_24_272 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_fill_2 FILLER_24_293 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_fill_2 FILLER_24_313 ();
 sg13g2_fill_2 FILLER_24_323 ();
 sg13g2_fill_1 FILLER_24_333 ();
 sg13g2_fill_2 FILLER_24_360 ();
 sg13g2_fill_1 FILLER_24_362 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_fill_1 FILLER_24_389 ();
 sg13g2_decap_4 FILLER_24_394 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_22 ();
 sg13g2_fill_2 FILLER_25_29 ();
 sg13g2_decap_4 FILLER_25_40 ();
 sg13g2_decap_4 FILLER_25_49 ();
 sg13g2_fill_1 FILLER_25_53 ();
 sg13g2_decap_4 FILLER_25_58 ();
 sg13g2_decap_4 FILLER_25_67 ();
 sg13g2_fill_2 FILLER_25_80 ();
 sg13g2_decap_8 FILLER_25_90 ();
 sg13g2_decap_8 FILLER_25_97 ();
 sg13g2_fill_2 FILLER_25_104 ();
 sg13g2_fill_1 FILLER_25_106 ();
 sg13g2_fill_2 FILLER_25_113 ();
 sg13g2_fill_2 FILLER_25_128 ();
 sg13g2_decap_8 FILLER_25_138 ();
 sg13g2_fill_2 FILLER_25_145 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_166 ();
 sg13g2_fill_2 FILLER_25_204 ();
 sg13g2_fill_2 FILLER_25_209 ();
 sg13g2_fill_1 FILLER_25_211 ();
 sg13g2_decap_8 FILLER_25_216 ();
 sg13g2_fill_2 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_265 ();
 sg13g2_decap_4 FILLER_25_292 ();
 sg13g2_decap_8 FILLER_25_307 ();
 sg13g2_decap_4 FILLER_25_314 ();
 sg13g2_fill_2 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_334 ();
 sg13g2_decap_4 FILLER_25_340 ();
 sg13g2_decap_4 FILLER_25_348 ();
 sg13g2_fill_1 FILLER_25_352 ();
 sg13g2_fill_2 FILLER_25_357 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_2 ();
 sg13g2_decap_4 FILLER_26_54 ();
 sg13g2_fill_1 FILLER_26_58 ();
 sg13g2_fill_1 FILLER_26_90 ();
 sg13g2_decap_4 FILLER_26_106 ();
 sg13g2_fill_1 FILLER_26_110 ();
 sg13g2_decap_4 FILLER_26_127 ();
 sg13g2_fill_1 FILLER_26_131 ();
 sg13g2_fill_2 FILLER_26_175 ();
 sg13g2_fill_1 FILLER_26_177 ();
 sg13g2_fill_1 FILLER_26_188 ();
 sg13g2_decap_4 FILLER_26_194 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_decap_4 FILLER_26_213 ();
 sg13g2_fill_2 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_fill_1 FILLER_26_249 ();
 sg13g2_fill_2 FILLER_26_255 ();
 sg13g2_fill_1 FILLER_26_257 ();
 sg13g2_decap_8 FILLER_26_268 ();
 sg13g2_decap_8 FILLER_26_285 ();
 sg13g2_fill_1 FILLER_26_292 ();
 sg13g2_fill_2 FILLER_26_314 ();
 sg13g2_fill_1 FILLER_26_316 ();
 sg13g2_decap_4 FILLER_26_342 ();
 sg13g2_fill_1 FILLER_26_346 ();
 sg13g2_fill_2 FILLER_26_368 ();
 sg13g2_fill_2 FILLER_26_375 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_23 ();
 sg13g2_decap_8 FILLER_27_50 ();
 sg13g2_decap_8 FILLER_27_57 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_105 ();
 sg13g2_decap_4 FILLER_27_138 ();
 sg13g2_fill_2 FILLER_27_142 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_fill_1 FILLER_27_161 ();
 sg13g2_decap_4 FILLER_27_167 ();
 sg13g2_fill_2 FILLER_27_171 ();
 sg13g2_decap_4 FILLER_27_218 ();
 sg13g2_fill_1 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_257 ();
 sg13g2_decap_4 FILLER_27_266 ();
 sg13g2_fill_1 FILLER_27_280 ();
 sg13g2_fill_2 FILLER_27_289 ();
 sg13g2_fill_1 FILLER_27_291 ();
 sg13g2_decap_8 FILLER_27_335 ();
 sg13g2_fill_2 FILLER_27_360 ();
 sg13g2_fill_2 FILLER_27_375 ();
 sg13g2_decap_4 FILLER_27_381 ();
 sg13g2_fill_2 FILLER_27_385 ();
 sg13g2_fill_1 FILLER_27_391 ();
 sg13g2_fill_2 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_30 ();
 sg13g2_fill_2 FILLER_28_37 ();
 sg13g2_decap_8 FILLER_28_43 ();
 sg13g2_fill_1 FILLER_28_50 ();
 sg13g2_fill_2 FILLER_28_76 ();
 sg13g2_fill_1 FILLER_28_78 ();
 sg13g2_fill_1 FILLER_28_88 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_105 ();
 sg13g2_fill_2 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_128 ();
 sg13g2_decap_8 FILLER_28_136 ();
 sg13g2_decap_8 FILLER_28_178 ();
 sg13g2_fill_2 FILLER_28_193 ();
 sg13g2_fill_1 FILLER_28_195 ();
 sg13g2_fill_1 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_223 ();
 sg13g2_decap_4 FILLER_28_230 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_fill_2 FILLER_28_245 ();
 sg13g2_fill_2 FILLER_28_251 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_decap_8 FILLER_28_257 ();
 sg13g2_decap_8 FILLER_28_264 ();
 sg13g2_decap_4 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_285 ();
 sg13g2_fill_1 FILLER_28_287 ();
 sg13g2_decap_4 FILLER_28_296 ();
 sg13g2_decap_4 FILLER_28_312 ();
 sg13g2_fill_1 FILLER_28_316 ();
 sg13g2_fill_1 FILLER_28_325 ();
 sg13g2_decap_4 FILLER_28_339 ();
 sg13g2_fill_1 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_354 ();
 sg13g2_fill_1 FILLER_28_369 ();
 sg13g2_fill_1 FILLER_28_375 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_23 ();
 sg13g2_fill_1 FILLER_29_25 ();
 sg13g2_fill_1 FILLER_29_62 ();
 sg13g2_decap_4 FILLER_29_68 ();
 sg13g2_fill_2 FILLER_29_72 ();
 sg13g2_fill_2 FILLER_29_87 ();
 sg13g2_fill_1 FILLER_29_89 ();
 sg13g2_fill_2 FILLER_29_98 ();
 sg13g2_fill_1 FILLER_29_100 ();
 sg13g2_fill_2 FILLER_29_104 ();
 sg13g2_fill_1 FILLER_29_106 ();
 sg13g2_decap_8 FILLER_29_120 ();
 sg13g2_decap_8 FILLER_29_127 ();
 sg13g2_fill_1 FILLER_29_134 ();
 sg13g2_decap_8 FILLER_29_141 ();
 sg13g2_decap_8 FILLER_29_148 ();
 sg13g2_fill_2 FILLER_29_155 ();
 sg13g2_fill_1 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_162 ();
 sg13g2_decap_4 FILLER_29_179 ();
 sg13g2_decap_4 FILLER_29_191 ();
 sg13g2_fill_1 FILLER_29_195 ();
 sg13g2_fill_2 FILLER_29_204 ();
 sg13g2_fill_1 FILLER_29_206 ();
 sg13g2_decap_4 FILLER_29_215 ();
 sg13g2_fill_2 FILLER_29_235 ();
 sg13g2_fill_1 FILLER_29_237 ();
 sg13g2_fill_1 FILLER_29_251 ();
 sg13g2_fill_1 FILLER_29_286 ();
 sg13g2_fill_2 FILLER_29_303 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_decap_8 FILLER_29_353 ();
 sg13g2_fill_2 FILLER_29_360 ();
 sg13g2_fill_1 FILLER_29_362 ();
 sg13g2_fill_1 FILLER_29_387 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_27 ();
 sg13g2_decap_8 FILLER_30_34 ();
 sg13g2_fill_1 FILLER_30_41 ();
 sg13g2_decap_4 FILLER_30_46 ();
 sg13g2_decap_8 FILLER_30_55 ();
 sg13g2_decap_4 FILLER_30_67 ();
 sg13g2_fill_2 FILLER_30_101 ();
 sg13g2_decap_4 FILLER_30_119 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_decap_4 FILLER_30_150 ();
 sg13g2_fill_2 FILLER_30_170 ();
 sg13g2_fill_1 FILLER_30_172 ();
 sg13g2_decap_8 FILLER_30_181 ();
 sg13g2_fill_2 FILLER_30_188 ();
 sg13g2_decap_8 FILLER_30_198 ();
 sg13g2_decap_8 FILLER_30_205 ();
 sg13g2_decap_8 FILLER_30_212 ();
 sg13g2_decap_4 FILLER_30_219 ();
 sg13g2_decap_4 FILLER_30_259 ();
 sg13g2_fill_1 FILLER_30_263 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_4 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_fill_2 FILLER_30_296 ();
 sg13g2_fill_1 FILLER_30_298 ();
 sg13g2_decap_8 FILLER_30_323 ();
 sg13g2_decap_4 FILLER_30_369 ();
 sg13g2_fill_2 FILLER_30_373 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_fill_1 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_39 ();
 sg13g2_decap_8 FILLER_31_78 ();
 sg13g2_fill_2 FILLER_31_85 ();
 sg13g2_fill_1 FILLER_31_87 ();
 sg13g2_decap_8 FILLER_31_103 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_4 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_130 ();
 sg13g2_fill_2 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_148 ();
 sg13g2_fill_1 FILLER_31_158 ();
 sg13g2_decap_8 FILLER_31_173 ();
 sg13g2_decap_4 FILLER_31_206 ();
 sg13g2_fill_2 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_233 ();
 sg13g2_decap_8 FILLER_31_250 ();
 sg13g2_fill_2 FILLER_31_257 ();
 sg13g2_fill_1 FILLER_31_259 ();
 sg13g2_decap_4 FILLER_31_301 ();
 sg13g2_fill_2 FILLER_31_313 ();
 sg13g2_fill_2 FILLER_31_331 ();
 sg13g2_fill_1 FILLER_31_333 ();
 sg13g2_decap_4 FILLER_31_345 ();
 sg13g2_fill_2 FILLER_31_349 ();
 sg13g2_decap_8 FILLER_31_377 ();
 sg13g2_fill_2 FILLER_31_384 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_18 ();
 sg13g2_fill_1 FILLER_32_20 ();
 sg13g2_decap_4 FILLER_32_30 ();
 sg13g2_decap_4 FILLER_32_45 ();
 sg13g2_fill_1 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_55 ();
 sg13g2_fill_2 FILLER_32_62 ();
 sg13g2_fill_1 FILLER_32_64 ();
 sg13g2_decap_8 FILLER_32_72 ();
 sg13g2_decap_4 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_102 ();
 sg13g2_decap_4 FILLER_32_127 ();
 sg13g2_fill_1 FILLER_32_131 ();
 sg13g2_decap_4 FILLER_32_149 ();
 sg13g2_fill_2 FILLER_32_153 ();
 sg13g2_fill_1 FILLER_32_177 ();
 sg13g2_fill_2 FILLER_32_199 ();
 sg13g2_decap_8 FILLER_32_206 ();
 sg13g2_decap_4 FILLER_32_213 ();
 sg13g2_fill_1 FILLER_32_217 ();
 sg13g2_fill_2 FILLER_32_230 ();
 sg13g2_decap_4 FILLER_32_256 ();
 sg13g2_fill_2 FILLER_32_260 ();
 sg13g2_decap_8 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_280 ();
 sg13g2_fill_2 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_293 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_fill_2 FILLER_32_337 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_351 ();
 sg13g2_fill_2 FILLER_32_384 ();
 sg13g2_fill_1 FILLER_32_386 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_30 ();
 sg13g2_fill_2 FILLER_33_41 ();
 sg13g2_fill_1 FILLER_33_43 ();
 sg13g2_decap_4 FILLER_33_51 ();
 sg13g2_fill_2 FILLER_33_74 ();
 sg13g2_decap_8 FILLER_33_86 ();
 sg13g2_fill_2 FILLER_33_93 ();
 sg13g2_fill_1 FILLER_33_103 ();
 sg13g2_decap_8 FILLER_33_114 ();
 sg13g2_decap_4 FILLER_33_121 ();
 sg13g2_fill_2 FILLER_33_138 ();
 sg13g2_fill_2 FILLER_33_144 ();
 sg13g2_decap_4 FILLER_33_157 ();
 sg13g2_fill_2 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_191 ();
 sg13g2_decap_4 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_241 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_fill_2 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_303 ();
 sg13g2_decap_4 FILLER_33_319 ();
 sg13g2_fill_2 FILLER_33_323 ();
 sg13g2_fill_1 FILLER_33_329 ();
 sg13g2_fill_1 FILLER_33_374 ();
 sg13g2_decap_4 FILLER_33_388 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_1 FILLER_34_36 ();
 sg13g2_fill_2 FILLER_34_60 ();
 sg13g2_decap_4 FILLER_34_92 ();
 sg13g2_fill_2 FILLER_34_96 ();
 sg13g2_decap_8 FILLER_34_107 ();
 sg13g2_decap_4 FILLER_34_114 ();
 sg13g2_decap_4 FILLER_34_144 ();
 sg13g2_fill_1 FILLER_34_148 ();
 sg13g2_fill_1 FILLER_34_162 ();
 sg13g2_fill_1 FILLER_34_176 ();
 sg13g2_decap_4 FILLER_34_182 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_decap_8 FILLER_34_205 ();
 sg13g2_decap_8 FILLER_34_212 ();
 sg13g2_decap_4 FILLER_34_219 ();
 sg13g2_fill_1 FILLER_34_228 ();
 sg13g2_fill_2 FILLER_34_246 ();
 sg13g2_fill_1 FILLER_34_248 ();
 sg13g2_decap_8 FILLER_34_268 ();
 sg13g2_decap_8 FILLER_34_275 ();
 sg13g2_decap_8 FILLER_34_297 ();
 sg13g2_fill_2 FILLER_34_304 ();
 sg13g2_fill_1 FILLER_34_306 ();
 sg13g2_decap_4 FILLER_34_326 ();
 sg13g2_decap_8 FILLER_34_339 ();
 sg13g2_decap_4 FILLER_34_346 ();
 sg13g2_fill_2 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_360 ();
 sg13g2_decap_4 FILLER_34_371 ();
 sg13g2_fill_2 FILLER_34_375 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_9 ();
 sg13g2_fill_2 FILLER_35_31 ();
 sg13g2_decap_8 FILLER_35_43 ();
 sg13g2_decap_4 FILLER_35_50 ();
 sg13g2_decap_8 FILLER_35_59 ();
 sg13g2_decap_8 FILLER_35_66 ();
 sg13g2_fill_2 FILLER_35_73 ();
 sg13g2_decap_4 FILLER_35_87 ();
 sg13g2_fill_2 FILLER_35_119 ();
 sg13g2_decap_4 FILLER_35_134 ();
 sg13g2_fill_2 FILLER_35_138 ();
 sg13g2_fill_2 FILLER_35_144 ();
 sg13g2_decap_4 FILLER_35_153 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_fill_2 FILLER_35_170 ();
 sg13g2_decap_4 FILLER_35_193 ();
 sg13g2_fill_1 FILLER_35_197 ();
 sg13g2_decap_8 FILLER_35_206 ();
 sg13g2_decap_8 FILLER_35_213 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_fill_1 FILLER_35_222 ();
 sg13g2_fill_2 FILLER_35_248 ();
 sg13g2_fill_2 FILLER_35_267 ();
 sg13g2_fill_1 FILLER_35_282 ();
 sg13g2_decap_8 FILLER_35_304 ();
 sg13g2_decap_4 FILLER_35_321 ();
 sg13g2_fill_1 FILLER_35_325 ();
 sg13g2_decap_8 FILLER_35_347 ();
 sg13g2_fill_2 FILLER_35_354 ();
 sg13g2_fill_2 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_379 ();
 sg13g2_fill_2 FILLER_35_389 ();
 sg13g2_fill_1 FILLER_35_391 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_22 ();
 sg13g2_decap_4 FILLER_36_29 ();
 sg13g2_fill_1 FILLER_36_33 ();
 sg13g2_fill_2 FILLER_36_39 ();
 sg13g2_decap_4 FILLER_36_57 ();
 sg13g2_fill_1 FILLER_36_80 ();
 sg13g2_decap_8 FILLER_36_86 ();
 sg13g2_fill_2 FILLER_36_93 ();
 sg13g2_decap_4 FILLER_36_103 ();
 sg13g2_fill_1 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_120 ();
 sg13g2_decap_8 FILLER_36_139 ();
 sg13g2_decap_8 FILLER_36_174 ();
 sg13g2_fill_2 FILLER_36_181 ();
 sg13g2_fill_1 FILLER_36_183 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_fill_2 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_228 ();
 sg13g2_decap_8 FILLER_36_242 ();
 sg13g2_decap_8 FILLER_36_249 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_263 ();
 sg13g2_decap_8 FILLER_36_283 ();
 sg13g2_decap_8 FILLER_36_297 ();
 sg13g2_fill_1 FILLER_36_325 ();
 sg13g2_fill_1 FILLER_36_331 ();
 sg13g2_fill_1 FILLER_36_358 ();
 sg13g2_decap_4 FILLER_36_366 ();
 sg13g2_fill_2 FILLER_36_378 ();
 sg13g2_fill_1 FILLER_36_380 ();
 sg13g2_fill_1 FILLER_36_385 ();
 sg13g2_fill_2 FILLER_36_391 ();
 sg13g2_fill_1 FILLER_36_393 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_fill_2 FILLER_37_25 ();
 sg13g2_fill_1 FILLER_37_27 ();
 sg13g2_fill_2 FILLER_37_47 ();
 sg13g2_decap_8 FILLER_37_68 ();
 sg13g2_decap_8 FILLER_37_92 ();
 sg13g2_fill_1 FILLER_37_99 ();
 sg13g2_fill_1 FILLER_37_113 ();
 sg13g2_decap_8 FILLER_37_208 ();
 sg13g2_decap_8 FILLER_37_215 ();
 sg13g2_decap_8 FILLER_37_222 ();
 sg13g2_fill_1 FILLER_37_229 ();
 sg13g2_fill_2 FILLER_37_238 ();
 sg13g2_fill_1 FILLER_37_240 ();
 sg13g2_fill_1 FILLER_37_282 ();
 sg13g2_fill_2 FILLER_37_301 ();
 sg13g2_fill_1 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_346 ();
 sg13g2_fill_2 FILLER_37_353 ();
 sg13g2_fill_2 FILLER_37_371 ();
 sg13g2_fill_1 FILLER_37_373 ();
 sg13g2_fill_1 FILLER_37_390 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_29 ();
 sg13g2_decap_4 FILLER_38_40 ();
 sg13g2_fill_2 FILLER_38_44 ();
 sg13g2_fill_2 FILLER_38_69 ();
 sg13g2_decap_8 FILLER_38_97 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_126 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_fill_2 FILLER_38_184 ();
 sg13g2_decap_8 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_decap_4 FILLER_38_227 ();
 sg13g2_fill_2 FILLER_38_231 ();
 sg13g2_fill_2 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_245 ();
 sg13g2_fill_2 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_fill_2 FILLER_38_299 ();
 sg13g2_fill_1 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_319 ();
 sg13g2_decap_8 FILLER_38_326 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_373 ();
 sg13g2_fill_1 FILLER_38_380 ();
 sg13g2_decap_4 FILLER_38_389 ();
 sg13g2_fill_1 FILLER_38_393 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_out[0] = net5;
 assign uio_out[1] = net6;
 assign uio_out[2] = net7;
 assign uio_out[3] = net8;
 assign uio_out[4] = net9;
 assign uio_out[5] = net10;
endmodule

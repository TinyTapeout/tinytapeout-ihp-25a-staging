module tt_um_a1k0n_nyancat (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire audio_pwm;
 wire \audio_pwm_accum[0] ;
 wire \audio_pwm_accum[1] ;
 wire \audio_pwm_accum[2] ;
 wire \audio_pwm_accum[3] ;
 wire \audio_pwm_accum[4] ;
 wire \audio_pwm_accum[5] ;
 wire \audio_pwm_accum[6] ;
 wire \audio_pwm_accum[7] ;
 wire \audio_pwm_accum[8] ;
 wire \audio_pwm_accum[9] ;
 wire \audio_pwm_accum_next[0] ;
 wire \audio_pwm_accum_next[1] ;
 wire \audio_pwm_accum_next[2] ;
 wire \audio_pwm_accum_next[3] ;
 wire \audio_pwm_accum_next[4] ;
 wire \audio_pwm_accum_next[5] ;
 wire \audio_pwm_accum_next[6] ;
 wire \audio_pwm_accum_next[7] ;
 wire \audio_pwm_accum_next[8] ;
 wire \audio_pwm_accum_next[9] ;
 wire \audio_sample_lpf[0] ;
 wire \audio_sample_lpf[1] ;
 wire \audio_sample_lpf[2] ;
 wire \audio_sample_lpf[3] ;
 wire \audio_sample_lpf[4] ;
 wire \audio_sample_lpf[5] ;
 wire \audio_sample_lpf[6] ;
 wire \audio_sample_lpf[7] ;
 wire \audio_sample_lpf[8] ;
 wire \audio_sample_lpf[9] ;
 wire \bass_pha[0] ;
 wire \bass_pha[10] ;
 wire \bass_pha[11] ;
 wire \bass_pha[12] ;
 wire \bass_pha[13] ;
 wire \bass_pha[14] ;
 wire \bass_pha[15] ;
 wire \bass_pha[1] ;
 wire \bass_pha[2] ;
 wire \bass_pha[3] ;
 wire \bass_pha[4] ;
 wire \bass_pha[5] ;
 wire \bass_pha[6] ;
 wire \bass_pha[7] ;
 wire \bass_pha[8] ;
 wire \bass_pha[9] ;
 wire \bass_vol[0] ;
 wire \bass_vol[1] ;
 wire \bass_vol[2] ;
 wire \bass_vol[3] ;
 wire \bass_vol[4] ;
 wire \bass_vol[5] ;
 wire \cos[0] ;
 wire \cos[1] ;
 wire \cos[2] ;
 wire \cos[3] ;
 wire \cos[4] ;
 wire \cos[5] ;
 wire \cos[6] ;
 wire \frame_count[0] ;
 wire \frame_count[1] ;
 wire \frame_count[2] ;
 wire \frame_count[3] ;
 wire \frame_count[4] ;
 wire \frame_count[5] ;
 wire \frame_count[6] ;
 wire \frame_count[7] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \kick_ctr[0] ;
 wire \kick_ctr[1] ;
 wire \kick_osci[0] ;
 wire \kick_osci[1] ;
 wire \kick_osci[2] ;
 wire \kick_osci[3] ;
 wire \kick_osci[4] ;
 wire \kick_osci[5] ;
 wire \kick_osci[6] ;
 wire \kick_osci[7] ;
 wire \kick_osci[8] ;
 wire \line_lfsr[0] ;
 wire \line_lfsr[1] ;
 wire \line_lfsr[2] ;
 wire \line_lfsr[3] ;
 wire \line_lfsr[4] ;
 wire \line_lfsr[5] ;
 wire \line_lfsr[6] ;
 wire \nyan_x_offset[0] ;
 wire \nyan_x_offset[1] ;
 wire \nyan_x_offset[2] ;
 wire \nyan_x_offset[3] ;
 wire \nyan_x_offset[4] ;
 wire \nyanframe[0] ;
 wire \nyanframe[1] ;
 wire \nyanframe[2] ;
 wire \sample_beat_ctr[0] ;
 wire \sample_beat_ctr[1] ;
 wire \sample_beat_ctr[2] ;
 wire \sin[0] ;
 wire \sin[6] ;
 wire song_loops;
 wire \songpos[0] ;
 wire \songpos[1] ;
 wire \songpos[2] ;
 wire \songpos[3] ;
 wire \songpos[4] ;
 wire \songpos[5] ;
 wire \songpos[6] ;
 wire \songpos[7] ;
 wire \songpos[8] ;
 wire \sqr_pha[0] ;
 wire \sqr_pha[10] ;
 wire \sqr_pha[11] ;
 wire \sqr_pha[12] ;
 wire \sqr_pha[1] ;
 wire \sqr_pha[2] ;
 wire \sqr_pha[3] ;
 wire \sqr_pha[4] ;
 wire \sqr_pha[5] ;
 wire \sqr_pha[6] ;
 wire \sqr_pha[7] ;
 wire \sqr_pha[8] ;
 wire \sqr_pha[9] ;
 wire \sqr_vol[0] ;
 wire \sqr_vol[1] ;
 wire \sqr_vol[2] ;
 wire \sqr_vol[3] ;
 wire \sqr_vol[4] ;
 wire \sqr_vol[5] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;

 sg13g2_inv_1 _2329_ (.Y(_1522_),
    .A(net76));
 sg13g2_inv_1 _2330_ (.Y(_1523_),
    .A(net116));
 sg13g2_inv_1 _2331_ (.Y(_1524_),
    .A(\kick_ctr[0] ));
 sg13g2_inv_1 _2332_ (.Y(_1525_),
    .A(\kick_osci[3] ));
 sg13g2_inv_1 _2333_ (.Y(_1526_),
    .A(net967));
 sg13g2_inv_1 _2334_ (.Y(_1527_),
    .A(net951));
 sg13g2_inv_4 _2335_ (.A(net946),
    .Y(_1528_));
 sg13g2_inv_4 _2336_ (.A(net948),
    .Y(_1529_));
 sg13g2_inv_2 _2337_ (.Y(_1530_),
    .A(net943));
 sg13g2_inv_2 _2338_ (.Y(_1531_),
    .A(net945));
 sg13g2_inv_1 _2339_ (.Y(_1532_),
    .A(net272));
 sg13g2_inv_1 _2340_ (.Y(_1533_),
    .A(net942));
 sg13g2_inv_4 _2341_ (.A(net988),
    .Y(_1534_));
 sg13g2_inv_2 _2342_ (.Y(_1535_),
    .A(net979));
 sg13g2_inv_1 _2343_ (.Y(_1536_),
    .A(net984));
 sg13g2_inv_1 _2344_ (.Y(_1537_),
    .A(\songpos[8] ));
 sg13g2_inv_1 _2345_ (.Y(_1538_),
    .A(net962));
 sg13g2_inv_1 _2346_ (.Y(_1539_),
    .A(\nyanframe[2] ));
 sg13g2_inv_1 _2347_ (.Y(_1540_),
    .A(net966));
 sg13g2_inv_1 _2348_ (.Y(_1541_),
    .A(\nyanframe[1] ));
 sg13g2_inv_1 _2349_ (.Y(_1542_),
    .A(_0032_));
 sg13g2_inv_1 _2350_ (.Y(_1543_),
    .A(_0034_));
 sg13g2_inv_1 _2351_ (.Y(_1544_),
    .A(net255));
 sg13g2_inv_1 _2352_ (.Y(_1545_),
    .A(net236));
 sg13g2_inv_1 _2353_ (.Y(_1546_),
    .A(net238));
 sg13g2_inv_1 _2354_ (.Y(_1547_),
    .A(net250));
 sg13g2_inv_1 _2355_ (.Y(_1548_),
    .A(net197));
 sg13g2_inv_1 _2356_ (.Y(_1549_),
    .A(\bass_vol[4] ));
 sg13g2_inv_1 _2357_ (.Y(_1550_),
    .A(net187));
 sg13g2_inv_1 _2358_ (.Y(_1551_),
    .A(net149));
 sg13g2_inv_1 _2359_ (.Y(_1552_),
    .A(net122));
 sg13g2_inv_1 _2360_ (.Y(_1553_),
    .A(net161));
 sg13g2_inv_1 _2361_ (.Y(_1554_),
    .A(net94));
 sg13g2_inv_1 _2362_ (.Y(_1555_),
    .A(\sqr_pha[12] ));
 sg13g2_inv_1 _2363_ (.Y(_1556_),
    .A(net145));
 sg13g2_inv_1 _2364_ (.Y(_1557_),
    .A(_0014_));
 sg13g2_inv_1 _2365_ (.Y(_1558_),
    .A(_0015_));
 sg13g2_inv_1 _2366_ (.Y(_1559_),
    .A(net210));
 sg13g2_inv_1 _2367_ (.Y(_1560_),
    .A(_0016_));
 sg13g2_inv_1 _2368_ (.Y(_1561_),
    .A(net159));
 sg13g2_inv_1 _2369_ (.Y(_1562_),
    .A(\kick_osci[6] ));
 sg13g2_inv_1 _2370_ (.Y(_1563_),
    .A(net226));
 sg13g2_inv_1 _2371_ (.Y(_1564_),
    .A(_0021_));
 sg13g2_inv_1 _2372_ (.Y(_1565_),
    .A(_0022_));
 sg13g2_inv_1 _2373_ (.Y(_1566_),
    .A(\bass_pha[15] ));
 sg13g2_inv_1 _2374_ (.Y(_1567_),
    .A(\cos[5] ));
 sg13g2_inv_1 _2375_ (.Y(_1568_),
    .A(_0024_));
 sg13g2_inv_1 _2376_ (.Y(_1569_),
    .A(_0025_));
 sg13g2_nor2_1 _2377_ (.A(net941),
    .B(_1529_),
    .Y(_1570_));
 sg13g2_nand2_1 _2378_ (.Y(_1571_),
    .A(net951),
    .B(net948));
 sg13g2_nor3_2 _2379_ (.A(net946),
    .B(net945),
    .C(net919),
    .Y(_1572_));
 sg13g2_nand2b_1 _2380_ (.Y(_1573_),
    .B(\hvsync_gen.vpos[7] ),
    .A_N(_1572_));
 sg13g2_xnor2_1 _2381_ (.Y(_1574_),
    .A(net943),
    .B(_1572_));
 sg13g2_xnor2_1 _2382_ (.Y(_1575_),
    .A(_1530_),
    .B(_1572_));
 sg13g2_nand2_1 _2383_ (.Y(_1576_),
    .A(\hvsync_gen.vpos[5] ),
    .B(net933));
 sg13g2_xnor2_1 _2384_ (.Y(_1577_),
    .A(_1528_),
    .B(net933));
 sg13g2_xnor2_1 _2385_ (.Y(_1578_),
    .A(\hvsync_gen.vpos[5] ),
    .B(net933));
 sg13g2_nor2_1 _2386_ (.A(net966),
    .B(net916),
    .Y(_1579_));
 sg13g2_nand2_2 _2387_ (.Y(_1580_),
    .A(net935),
    .B(net914));
 sg13g2_and2_1 _2388_ (.A(\hvsync_gen.hpos[2] ),
    .B(\nyan_x_offset[2] ),
    .X(_1581_));
 sg13g2_nand2_1 _2389_ (.Y(_1582_),
    .A(\nyan_x_offset[3] ),
    .B(\hvsync_gen.hpos[3] ));
 sg13g2_xor2_1 _2390_ (.B(\hvsync_gen.hpos[3] ),
    .A(\nyan_x_offset[3] ),
    .X(_1583_));
 sg13g2_and2_1 _2391_ (.A(_1581_),
    .B(_1583_),
    .X(_1584_));
 sg13g2_xor2_1 _2392_ (.B(_1583_),
    .A(_1581_),
    .X(_1585_));
 sg13g2_xor2_1 _2393_ (.B(\nyan_x_offset[2] ),
    .A(\hvsync_gen.hpos[2] ),
    .X(_1586_));
 sg13g2_nor2_1 _2394_ (.A(\hvsync_gen.hpos[1] ),
    .B(\nyan_x_offset[1] ),
    .Y(_1587_));
 sg13g2_nor2b_1 _2395_ (.A(_1587_),
    .B_N(_1586_),
    .Y(_1588_));
 sg13g2_xnor2_1 _2396_ (.Y(_1589_),
    .A(_1586_),
    .B(_1587_));
 sg13g2_xnor2_1 _2397_ (.Y(_1590_),
    .A(\hvsync_gen.hpos[1] ),
    .B(\nyan_x_offset[1] ));
 sg13g2_and3_1 _2398_ (.X(_1591_),
    .A(\hvsync_gen.hpos[0] ),
    .B(\nyan_x_offset[0] ),
    .C(_1590_));
 sg13g2_a21oi_1 _2399_ (.A1(_1589_),
    .A2(_1591_),
    .Y(_1592_),
    .B1(_1588_));
 sg13g2_xnor2_1 _2400_ (.Y(_1593_),
    .A(_1585_),
    .B(_1592_));
 sg13g2_xor2_1 _2401_ (.B(_1592_),
    .A(_1585_),
    .X(_1594_));
 sg13g2_nand2b_1 _2402_ (.Y(_1595_),
    .B(net963),
    .A_N(net971));
 sg13g2_and2_1 _2403_ (.A(net970),
    .B(_1595_),
    .X(_1596_));
 sg13g2_xor2_1 _2404_ (.B(_1595_),
    .A(net970),
    .X(_1597_));
 sg13g2_nand2_1 _2405_ (.Y(_1598_),
    .A(net972),
    .B(\nyan_x_offset[4] ));
 sg13g2_xor2_1 _2406_ (.B(\nyan_x_offset[4] ),
    .A(net972),
    .X(_1599_));
 sg13g2_nand2b_2 _2407_ (.Y(_1600_),
    .B(_1599_),
    .A_N(_1582_));
 sg13g2_xor2_1 _2408_ (.B(_1599_),
    .A(_1582_),
    .X(_1601_));
 sg13g2_inv_1 _2409_ (.Y(_1602_),
    .A(_1601_));
 sg13g2_and3_1 _2410_ (.X(_1603_),
    .A(_1585_),
    .B(_1589_),
    .C(_1591_));
 sg13g2_nand3_1 _2411_ (.B(_1589_),
    .C(_1591_),
    .A(_1585_),
    .Y(_1604_));
 sg13g2_a21o_1 _2412_ (.A2(_1588_),
    .A1(_1583_),
    .B1(_1584_),
    .X(_1605_));
 sg13g2_o21ai_1 _2413_ (.B1(_1583_),
    .Y(_1606_),
    .A1(_1581_),
    .A2(_1588_));
 sg13g2_a21oi_2 _2414_ (.B1(_1601_),
    .Y(_1607_),
    .A2(_1606_),
    .A1(_1604_));
 sg13g2_o21ai_1 _2415_ (.B1(_1602_),
    .Y(_1608_),
    .A1(_1603_),
    .A2(_1605_));
 sg13g2_xnor2_1 _2416_ (.Y(_1609_),
    .A(net971),
    .B(net963));
 sg13g2_xnor2_1 _2417_ (.Y(_1610_),
    .A(_1598_),
    .B(_1609_));
 sg13g2_inv_1 _2418_ (.Y(_1611_),
    .A(_1610_));
 sg13g2_nor2_2 _2419_ (.A(_1600_),
    .B(_1609_),
    .Y(_1612_));
 sg13g2_a21oi_1 _2420_ (.A1(_1598_),
    .A2(_1600_),
    .Y(_1613_),
    .B1(_1609_));
 sg13g2_a21oi_1 _2421_ (.A1(_1607_),
    .A2(_1611_),
    .Y(_1614_),
    .B1(_1613_));
 sg13g2_a21o_1 _2422_ (.A2(_1611_),
    .A1(_1607_),
    .B1(_1613_),
    .X(_1615_));
 sg13g2_a21oi_2 _2423_ (.B1(_1596_),
    .Y(_1616_),
    .A2(_1615_),
    .A1(_1597_));
 sg13g2_a21o_1 _2424_ (.A2(_1615_),
    .A1(_1597_),
    .B1(_1596_),
    .X(_1617_));
 sg13g2_nand3_1 _2425_ (.B(_1543_),
    .C(_1617_),
    .A(_1526_),
    .Y(_1618_));
 sg13g2_o21ai_1 _2426_ (.B1(net967),
    .Y(_1619_),
    .A1(_0034_),
    .A2(_1616_));
 sg13g2_nand3_1 _2427_ (.B(_1543_),
    .C(_1617_),
    .A(net967),
    .Y(_1620_));
 sg13g2_o21ai_1 _2428_ (.B1(_1526_),
    .Y(_1621_),
    .A1(_0034_),
    .A2(_1616_));
 sg13g2_nand2_1 _2429_ (.Y(_1622_),
    .A(_1620_),
    .B(_1621_));
 sg13g2_nand2_1 _2430_ (.Y(_1623_),
    .A(net827),
    .B(net824));
 sg13g2_xnor2_1 _2431_ (.Y(_1624_),
    .A(_1543_),
    .B(_1616_));
 sg13g2_xnor2_1 _2432_ (.Y(_1625_),
    .A(_0034_),
    .B(_1616_));
 sg13g2_nand3_1 _2433_ (.B(_1604_),
    .C(_1606_),
    .A(_1601_),
    .Y(_1626_));
 sg13g2_o21ai_1 _2434_ (.B1(_1601_),
    .Y(_1627_),
    .A1(_1603_),
    .A2(_1605_));
 sg13g2_nand3_1 _2435_ (.B(_1604_),
    .C(_1606_),
    .A(_1602_),
    .Y(_1628_));
 sg13g2_nand2_1 _2436_ (.Y(_1629_),
    .A(_1627_),
    .B(_1628_));
 sg13g2_nand2_2 _2437_ (.Y(_1630_),
    .A(_1608_),
    .B(_1626_));
 sg13g2_xnor2_1 _2438_ (.Y(_1631_),
    .A(_1597_),
    .B(_1614_));
 sg13g2_xnor2_1 _2439_ (.Y(_1632_),
    .A(_1597_),
    .B(_1615_));
 sg13g2_xnor2_1 _2440_ (.Y(_1633_),
    .A(_1607_),
    .B(_1611_));
 sg13g2_a21oi_1 _2441_ (.A1(_1600_),
    .A2(_1633_),
    .Y(_1634_),
    .B1(_1612_));
 sg13g2_a21o_2 _2442_ (.A2(_1633_),
    .A1(_1600_),
    .B1(_1612_),
    .X(_1635_));
 sg13g2_nor2_1 _2443_ (.A(net855),
    .B(net839),
    .Y(_1636_));
 sg13g2_nand2_2 _2444_ (.Y(_1637_),
    .A(net845),
    .B(net835));
 sg13g2_nand2_2 _2445_ (.Y(_1638_),
    .A(_1630_),
    .B(net836));
 sg13g2_nor3_2 _2446_ (.A(net872),
    .B(net854),
    .C(net841),
    .Y(_1639_));
 sg13g2_nor2_2 _2447_ (.A(net879),
    .B(net871),
    .Y(_1640_));
 sg13g2_nand3_1 _2448_ (.B(_1627_),
    .C(_1628_),
    .A(net878),
    .Y(_1641_));
 sg13g2_nor3_2 _2449_ (.A(net860),
    .B(net843),
    .C(net869),
    .Y(_1642_));
 sg13g2_nand3_1 _2450_ (.B(net838),
    .C(_1640_),
    .A(net851),
    .Y(_1643_));
 sg13g2_and4_2 _2451_ (.A(net828),
    .B(net825),
    .C(net822),
    .D(_1642_),
    .X(_1644_));
 sg13g2_nand4_1 _2452_ (.B(net825),
    .C(net822),
    .A(net828),
    .Y(_1645_),
    .D(_1642_));
 sg13g2_xnor2_1 _2453_ (.Y(_1646_),
    .A(net969),
    .B(_1616_));
 sg13g2_xnor2_1 _2454_ (.Y(_1647_),
    .A(net969),
    .B(_1617_));
 sg13g2_nor2_1 _2455_ (.A(net845),
    .B(net809),
    .Y(_1648_));
 sg13g2_nand2_2 _2456_ (.Y(_1649_),
    .A(net859),
    .B(net806));
 sg13g2_a21oi_2 _2457_ (.B1(net805),
    .Y(_1650_),
    .A2(net825),
    .A1(net828));
 sg13g2_a221oi_1 _2458_ (.B2(_1600_),
    .C1(_1612_),
    .B1(_1633_),
    .A1(_1627_),
    .Y(_1651_),
    .A2(_1628_));
 sg13g2_nand2_2 _2459_ (.Y(_1652_),
    .A(net871),
    .B(net839));
 sg13g2_nor2_2 _2460_ (.A(net878),
    .B(net870),
    .Y(_1653_));
 sg13g2_nand3_1 _2461_ (.B(_1608_),
    .C(_1626_),
    .A(net880),
    .Y(_1654_));
 sg13g2_nor2_1 _2462_ (.A(net837),
    .B(net867),
    .Y(_1655_));
 sg13g2_nand2_1 _2463_ (.Y(_1656_),
    .A(net843),
    .B(net831));
 sg13g2_a22oi_1 _2464_ (.Y(_1657_),
    .B1(net806),
    .B2(_1656_),
    .A2(net826),
    .A1(net829));
 sg13g2_nand2_1 _2465_ (.Y(_1658_),
    .A(_1649_),
    .B(_1657_));
 sg13g2_nand2_2 _2466_ (.Y(_1659_),
    .A(net837),
    .B(net867));
 sg13g2_nor3_2 _2467_ (.A(net859),
    .B(net844),
    .C(net831),
    .Y(_1660_));
 sg13g2_nand3_1 _2468_ (.B(net836),
    .C(net866),
    .A(net846),
    .Y(_1661_));
 sg13g2_nand2_1 _2469_ (.Y(_1662_),
    .A(net819),
    .B(_1660_));
 sg13g2_nand3_1 _2470_ (.B(_1657_),
    .C(_1662_),
    .A(_1649_),
    .Y(_1663_));
 sg13g2_nand2_1 _2471_ (.Y(_1664_),
    .A(_1645_),
    .B(_1663_));
 sg13g2_nor2_1 _2472_ (.A(\hvsync_gen.vpos[5] ),
    .B(_1664_),
    .Y(_1665_));
 sg13g2_nor2_2 _2473_ (.A(net951),
    .B(net948),
    .Y(_1666_));
 sg13g2_nand2_1 _2474_ (.Y(_1667_),
    .A(net939),
    .B(_1529_));
 sg13g2_nand2_1 _2475_ (.Y(_1668_),
    .A(net871),
    .B(net854));
 sg13g2_nor2_2 _2476_ (.A(_1594_),
    .B(net851),
    .Y(_1669_));
 sg13g2_nand2_2 _2477_ (.Y(_1670_),
    .A(net879),
    .B(net855));
 sg13g2_nand2_1 _2478_ (.Y(_1671_),
    .A(net855),
    .B(net839));
 sg13g2_a21oi_1 _2479_ (.A1(net878),
    .A2(net834),
    .Y(_1672_),
    .B1(net847));
 sg13g2_o21ai_1 _2480_ (.B1(net856),
    .Y(_1673_),
    .A1(net879),
    .A2(net840));
 sg13g2_nor2_2 _2481_ (.A(net811),
    .B(_1672_),
    .Y(_1674_));
 sg13g2_a21oi_2 _2482_ (.B1(net848),
    .Y(_1675_),
    .A2(net835),
    .A1(net870));
 sg13g2_nand2_2 _2483_ (.Y(_1676_),
    .A(net856),
    .B(net869));
 sg13g2_nor2_1 _2484_ (.A(net845),
    .B(_1640_),
    .Y(_1677_));
 sg13g2_nand2_1 _2485_ (.Y(_1678_),
    .A(net803),
    .B(_1676_));
 sg13g2_nor3_2 _2486_ (.A(net816),
    .B(_1669_),
    .C(_1675_),
    .Y(_1679_));
 sg13g2_nand3_1 _2487_ (.B(_1671_),
    .C(_1676_),
    .A(net800),
    .Y(_1680_));
 sg13g2_or2_1 _2488_ (.X(_1681_),
    .B(net832),
    .A(net857));
 sg13g2_nor2_2 _2489_ (.A(net854),
    .B(net832),
    .Y(_1682_));
 sg13g2_o21ai_1 _2490_ (.B1(net850),
    .Y(_1683_),
    .A1(net837),
    .A2(net867));
 sg13g2_a21oi_2 _2491_ (.B1(net859),
    .Y(_1684_),
    .A2(net831),
    .A1(net843));
 sg13g2_a21oi_1 _2492_ (.A1(net829),
    .A2(net824),
    .Y(_1685_),
    .B1(_1684_));
 sg13g2_nand2_1 _2493_ (.Y(_1686_),
    .A(_1679_),
    .B(_1685_));
 sg13g2_a21oi_1 _2494_ (.A1(_1679_),
    .A2(_1685_),
    .Y(_1687_),
    .B1(net911));
 sg13g2_nand2_1 _2495_ (.Y(_1688_),
    .A(_1637_),
    .B(_1650_));
 sg13g2_nor2_1 _2496_ (.A(net919),
    .B(_1666_),
    .Y(_1689_));
 sg13g2_nand2_1 _2497_ (.Y(_1690_),
    .A(net933),
    .B(net912));
 sg13g2_nand2_1 _2498_ (.Y(_1691_),
    .A(net841),
    .B(net866));
 sg13g2_nor2_2 _2499_ (.A(net879),
    .B(net870),
    .Y(_1692_));
 sg13g2_nand2_2 _2500_ (.Y(_1693_),
    .A(net878),
    .B(net871));
 sg13g2_nor2_1 _2501_ (.A(net839),
    .B(_1692_),
    .Y(_1694_));
 sg13g2_a21oi_2 _2502_ (.B1(net847),
    .Y(_1695_),
    .A2(_1693_),
    .A1(net834));
 sg13g2_a21oi_2 _2503_ (.B1(_1682_),
    .Y(_1696_),
    .A2(_1695_),
    .A1(net798));
 sg13g2_nor2_2 _2504_ (.A(net953),
    .B(net800),
    .Y(_1697_));
 sg13g2_nand2b_1 _2505_ (.Y(_1698_),
    .B(_1697_),
    .A_N(_1696_));
 sg13g2_nor2_2 _2506_ (.A(net846),
    .B(net799),
    .Y(_1699_));
 sg13g2_nand2_1 _2507_ (.Y(_1700_),
    .A(net859),
    .B(net817));
 sg13g2_nor3_2 _2508_ (.A(net849),
    .B(net836),
    .C(net866),
    .Y(_1701_));
 sg13g2_nand2_2 _2509_ (.Y(_1702_),
    .A(net833),
    .B(_1669_));
 sg13g2_a22oi_1 _2510_ (.Y(_1703_),
    .B1(net810),
    .B2(_1701_),
    .A2(net824),
    .A1(net827));
 sg13g2_nand2_2 _2511_ (.Y(_1704_),
    .A(net872),
    .B(net834));
 sg13g2_nor2_2 _2512_ (.A(net840),
    .B(net866),
    .Y(_1705_));
 sg13g2_nand2_2 _2513_ (.Y(_1706_),
    .A(net834),
    .B(net831));
 sg13g2_nor2_2 _2514_ (.A(net955),
    .B(net820),
    .Y(_1707_));
 sg13g2_nor2_1 _2515_ (.A(net858),
    .B(net809),
    .Y(_1708_));
 sg13g2_a22oi_1 _2516_ (.Y(_1709_),
    .B1(_1705_),
    .B2(_1707_),
    .A2(_1684_),
    .A1(net800));
 sg13g2_nand3_1 _2517_ (.B(_1703_),
    .C(_1709_),
    .A(_1698_),
    .Y(_1710_));
 sg13g2_a221oi_1 _2518_ (.B2(_1710_),
    .C1(_1665_),
    .B1(net889),
    .A1(_1687_),
    .Y(_1711_),
    .A2(_1688_));
 sg13g2_nor2_1 _2519_ (.A(net953),
    .B(_1529_),
    .Y(_1712_));
 sg13g2_nand2_1 _2520_ (.Y(_1713_),
    .A(net939),
    .B(net950));
 sg13g2_a221oi_1 _2521_ (.B2(_1600_),
    .C1(_1612_),
    .B1(_1633_),
    .A1(net878),
    .Y(_1714_),
    .A2(net870));
 sg13g2_nand2_1 _2522_ (.Y(_1715_),
    .A(net843),
    .B(net869));
 sg13g2_nor2_1 _2523_ (.A(net854),
    .B(_1714_),
    .Y(_1716_));
 sg13g2_a221oi_1 _2524_ (.B2(_1715_),
    .C1(net800),
    .B1(net846),
    .A1(net829),
    .Y(_1717_),
    .A2(net826));
 sg13g2_a221oi_1 _2525_ (.B2(_1600_),
    .C1(_1612_),
    .B1(_1633_),
    .A1(_1608_),
    .Y(_1718_),
    .A2(_1626_));
 sg13g2_nand2_2 _2526_ (.Y(_1719_),
    .A(net870),
    .B(net841));
 sg13g2_nand3_1 _2527_ (.B(_1704_),
    .C(_1719_),
    .A(_1677_),
    .Y(_1720_));
 sg13g2_a21oi_2 _2528_ (.B1(net810),
    .Y(_1721_),
    .A2(net824),
    .A1(net827));
 sg13g2_a22oi_1 _2529_ (.Y(_1722_),
    .B1(net787),
    .B2(_1696_),
    .A2(_1720_),
    .A1(_1717_));
 sg13g2_nor2_1 _2530_ (.A(net941),
    .B(net948),
    .Y(_1723_));
 sg13g2_nand2_1 _2531_ (.Y(_1724_),
    .A(net953),
    .B(_1529_));
 sg13g2_nand2_2 _2532_ (.Y(_1725_),
    .A(net799),
    .B(_1682_));
 sg13g2_a21oi_1 _2533_ (.A1(_1703_),
    .A2(_1725_),
    .Y(_1726_),
    .B1(net900));
 sg13g2_a22oi_1 _2534_ (.Y(_1727_),
    .B1(net822),
    .B2(_1639_),
    .A2(_1621_),
    .A1(_1620_));
 sg13g2_a21o_1 _2535_ (.A2(_1639_),
    .A1(net822),
    .B1(net790),
    .X(_1728_));
 sg13g2_a22oi_1 _2536_ (.Y(_1729_),
    .B1(net822),
    .B2(_1642_),
    .A2(_1621_),
    .A1(_1620_));
 sg13g2_a21oi_2 _2537_ (.B1(net831),
    .Y(_1730_),
    .A2(net835),
    .A1(net872));
 sg13g2_or3_1 _2538_ (.A(net857),
    .B(net813),
    .C(_1730_),
    .X(_1731_));
 sg13g2_a22oi_1 _2539_ (.Y(_1732_),
    .B1(net809),
    .B2(_1661_),
    .A2(net824),
    .A1(net827));
 sg13g2_a21o_1 _2540_ (.A2(_1732_),
    .A1(_1731_),
    .B1(_1729_),
    .X(_1733_));
 sg13g2_a21oi_1 _2541_ (.A1(_1687_),
    .A2(_1688_),
    .Y(_1734_),
    .B1(net916));
 sg13g2_a221oi_1 _2542_ (.B2(net917),
    .C1(_1726_),
    .B1(_1733_),
    .A1(net907),
    .Y(_1735_),
    .A2(_1722_));
 sg13g2_nand2_1 _2543_ (.Y(_1736_),
    .A(net836),
    .B(_1640_));
 sg13g2_and2_1 _2544_ (.A(net868),
    .B(net866),
    .X(_1737_));
 sg13g2_or2_2 _2545_ (.X(_1738_),
    .B(_1737_),
    .A(net841));
 sg13g2_nand4_1 _2546_ (.B(net810),
    .C(_1719_),
    .A(net854),
    .Y(_1739_),
    .D(_1738_));
 sg13g2_nand3_1 _2547_ (.B(_1677_),
    .C(net798),
    .A(net799),
    .Y(_1740_));
 sg13g2_nand4_1 _2548_ (.B(_1681_),
    .C(_1739_),
    .A(net788),
    .Y(_1741_),
    .D(_1740_));
 sg13g2_nor2_2 _2549_ (.A(_0039_),
    .B(net889),
    .Y(_1742_));
 sg13g2_nand2_1 _2550_ (.Y(_1743_),
    .A(net916),
    .B(_1742_));
 sg13g2_o21ai_1 _2551_ (.B1(net966),
    .Y(_1744_),
    .A1(_1741_),
    .A2(_1743_));
 sg13g2_a21oi_1 _2552_ (.A1(_1734_),
    .A2(_1735_),
    .Y(_1745_),
    .B1(_1744_));
 sg13g2_nor2_2 _2553_ (.A(net965),
    .B(net914),
    .Y(_1746_));
 sg13g2_nand2_2 _2554_ (.Y(_1747_),
    .A(net936),
    .B(net915));
 sg13g2_a21o_2 _2555_ (.A2(net835),
    .A1(net870),
    .B1(_1714_),
    .X(_1748_));
 sg13g2_o21ai_1 _2556_ (.B1(_1683_),
    .Y(_1749_),
    .A1(_1700_),
    .A2(_1730_));
 sg13g2_nor4_1 _2557_ (.A(_0039_),
    .B(net795),
    .C(net889),
    .D(_1749_),
    .Y(_1750_));
 sg13g2_o21ai_1 _2558_ (.B1(_1750_),
    .Y(_1751_),
    .A1(_1649_),
    .A2(_1748_));
 sg13g2_a21oi_1 _2559_ (.A1(_1746_),
    .A2(_1751_),
    .Y(_1752_),
    .B1(_1745_));
 sg13g2_o21ai_1 _2560_ (.B1(_1752_),
    .Y(_1753_),
    .A1(_1580_),
    .A2(_1711_));
 sg13g2_nand2_1 _2561_ (.Y(_1754_),
    .A(_0035_),
    .B(net933));
 sg13g2_xnor2_1 _2562_ (.Y(_1755_),
    .A(_1531_),
    .B(_1754_));
 sg13g2_xnor2_1 _2563_ (.Y(_1756_),
    .A(net944),
    .B(_1754_));
 sg13g2_nor4_2 _2564_ (.A(net878),
    .B(net871),
    .C(net857),
    .Y(_1757_),
    .D(net840));
 sg13g2_nand2_1 _2565_ (.Y(_1758_),
    .A(net879),
    .B(_1639_));
 sg13g2_a21oi_2 _2566_ (.B1(net790),
    .Y(_1759_),
    .A2(_1757_),
    .A1(net823));
 sg13g2_a221oi_1 _2567_ (.B2(_1669_),
    .C1(net807),
    .B1(net833),
    .A1(_1630_),
    .Y(_1760_),
    .A2(net851));
 sg13g2_nand2_2 _2568_ (.Y(_1761_),
    .A(net839),
    .B(_1693_));
 sg13g2_nor2_2 _2569_ (.A(net856),
    .B(net834),
    .Y(_1762_));
 sg13g2_nand2_1 _2570_ (.Y(_1763_),
    .A(net847),
    .B(net839));
 sg13g2_a21oi_2 _2571_ (.B1(net856),
    .Y(_1764_),
    .A2(net834),
    .A1(net871));
 sg13g2_a221oi_1 _2572_ (.B2(net797),
    .C1(net818),
    .B1(_1761_),
    .A1(net859),
    .Y(_1765_),
    .A2(_1706_));
 sg13g2_nor3_1 _2573_ (.A(net794),
    .B(_1760_),
    .C(_1765_),
    .Y(_1766_));
 sg13g2_o21ai_1 _2574_ (.B1(net908),
    .Y(_1767_),
    .A1(_1759_),
    .A2(_1766_));
 sg13g2_a21oi_2 _2575_ (.B1(net845),
    .Y(_1768_),
    .A2(net835),
    .A1(net871));
 sg13g2_or3_2 _2576_ (.A(_1660_),
    .B(_1669_),
    .C(_1768_),
    .X(_1769_));
 sg13g2_nand2_1 _2577_ (.Y(_1770_),
    .A(net807),
    .B(_1769_));
 sg13g2_nand2_1 _2578_ (.Y(_1771_),
    .A(net786),
    .B(_1769_));
 sg13g2_a22oi_1 _2579_ (.Y(_1772_),
    .B1(_1639_),
    .B2(net813),
    .A2(net824),
    .A1(net827));
 sg13g2_a21oi_2 _2580_ (.B1(_1727_),
    .Y(_1773_),
    .A2(_1650_),
    .A1(_1639_));
 sg13g2_o21ai_1 _2581_ (.B1(net850),
    .Y(_1774_),
    .A1(net843),
    .A2(net869));
 sg13g2_nand2_1 _2582_ (.Y(_1775_),
    .A(net940),
    .B(net787));
 sg13g2_nand3_1 _2583_ (.B(net786),
    .C(_1774_),
    .A(net939),
    .Y(_1776_));
 sg13g2_nand3_1 _2584_ (.B(net786),
    .C(_1769_),
    .A(net957),
    .Y(_1777_));
 sg13g2_nand3_1 _2585_ (.B(_1776_),
    .C(_1777_),
    .A(_1773_),
    .Y(_1778_));
 sg13g2_nand2_1 _2586_ (.Y(_1779_),
    .A(net888),
    .B(_1778_));
 sg13g2_a21oi_1 _2587_ (.A1(_1767_),
    .A2(_1779_),
    .Y(_1780_),
    .B1(_1747_));
 sg13g2_nor2_1 _2588_ (.A(net946),
    .B(net950),
    .Y(_1781_));
 sg13g2_nor2_2 _2589_ (.A(net947),
    .B(net901),
    .Y(_1782_));
 sg13g2_nor2_2 _2590_ (.A(net850),
    .B(net833),
    .Y(_1783_));
 sg13g2_nor4_1 _2591_ (.A(_1642_),
    .B(net818),
    .C(_1669_),
    .D(_1783_),
    .Y(_1784_));
 sg13g2_nor3_1 _2592_ (.A(net795),
    .B(_1760_),
    .C(_1784_),
    .Y(_1785_));
 sg13g2_o21ai_1 _2593_ (.B1(_1782_),
    .Y(_1786_),
    .A1(_1759_),
    .A2(_1785_));
 sg13g2_nand2_1 _2594_ (.Y(_1787_),
    .A(_1575_),
    .B(_1786_));
 sg13g2_nand3_1 _2595_ (.B(_1663_),
    .C(net931),
    .A(_1645_),
    .Y(_1788_));
 sg13g2_nor2_1 _2596_ (.A(net939),
    .B(_1644_),
    .Y(_1789_));
 sg13g2_nor2_2 _2597_ (.A(_1644_),
    .B(net900),
    .Y(_1790_));
 sg13g2_o21ai_1 _2598_ (.B1(net857),
    .Y(_1791_),
    .A1(net836),
    .A2(_1641_));
 sg13g2_a21oi_1 _2599_ (.A1(net841),
    .A2(_1640_),
    .Y(_1792_),
    .B1(net845));
 sg13g2_nand2_2 _2600_ (.Y(_1793_),
    .A(_1683_),
    .B(_1791_));
 sg13g2_nand2_1 _2601_ (.Y(_1794_),
    .A(net806),
    .B(_1793_));
 sg13g2_nand3_1 _2602_ (.B(_1662_),
    .C(_1794_),
    .A(net790),
    .Y(_1795_));
 sg13g2_a21oi_1 _2603_ (.A1(net828),
    .A2(net825),
    .Y(_1796_),
    .B1(_1624_));
 sg13g2_nor3_1 _2604_ (.A(_1594_),
    .B(net860),
    .C(net838),
    .Y(_1797_));
 sg13g2_and2_2 _2605_ (.A(net847),
    .B(_1714_),
    .X(_1798_));
 sg13g2_a22oi_1 _2606_ (.Y(_1799_),
    .B1(_1797_),
    .B2(net964),
    .A2(net833),
    .A1(net851));
 sg13g2_nor2_2 _2607_ (.A(_1526_),
    .B(net822),
    .Y(_1800_));
 sg13g2_nand2_1 _2608_ (.Y(_1801_),
    .A(_1624_),
    .B(_1757_));
 sg13g2_a22oi_1 _2609_ (.Y(_1802_),
    .B1(_1800_),
    .B2(_1757_),
    .A2(_1799_),
    .A1(net784));
 sg13g2_a21oi_1 _2610_ (.A1(_1728_),
    .A2(_1802_),
    .Y(_1803_),
    .B1(net905));
 sg13g2_nand2_1 _2611_ (.Y(_1804_),
    .A(_1657_),
    .B(_1659_));
 sg13g2_nor2_1 _2612_ (.A(net934),
    .B(_1644_),
    .Y(_1805_));
 sg13g2_a221oi_1 _2613_ (.B2(_1805_),
    .C1(_1803_),
    .B1(_1804_),
    .A1(_1790_),
    .Y(_1806_),
    .A2(_1795_));
 sg13g2_a21oi_1 _2614_ (.A1(_1788_),
    .A2(_1806_),
    .Y(_1807_),
    .B1(net915));
 sg13g2_nor2_2 _2615_ (.A(net936),
    .B(net913),
    .Y(_1808_));
 sg13g2_nand2_2 _2616_ (.Y(_1809_),
    .A(net965),
    .B(net915));
 sg13g2_nor2_1 _2617_ (.A(net842),
    .B(_1640_),
    .Y(_1810_));
 sg13g2_nand2_2 _2618_ (.Y(_1811_),
    .A(net835),
    .B(net868));
 sg13g2_nand2b_2 _2619_ (.Y(_1812_),
    .B(net842),
    .A_N(_1737_));
 sg13g2_a21oi_1 _2620_ (.A1(_1811_),
    .A2(_1812_),
    .Y(_1813_),
    .B1(net818));
 sg13g2_a221oi_1 _2621_ (.B2(_1812_),
    .C1(net818),
    .B1(_1811_),
    .A1(net860),
    .Y(_1814_),
    .A2(_1706_));
 sg13g2_nor3_1 _2622_ (.A(net795),
    .B(_1760_),
    .C(_1814_),
    .Y(_1815_));
 sg13g2_o21ai_1 _2623_ (.B1(net910),
    .Y(_1816_),
    .A1(_1759_),
    .A2(_1815_));
 sg13g2_a21oi_1 _2624_ (.A1(_1771_),
    .A2(_1773_),
    .Y(_1817_),
    .B1(net934));
 sg13g2_nand2_1 _2625_ (.Y(_1818_),
    .A(net850),
    .B(_1638_));
 sg13g2_nand3_1 _2626_ (.B(_1700_),
    .C(_1818_),
    .A(net790),
    .Y(_1819_));
 sg13g2_a21oi_1 _2627_ (.A1(_1728_),
    .A2(_1819_),
    .Y(_1820_),
    .B1(net912));
 sg13g2_nor2_1 _2628_ (.A(_1817_),
    .B(_1820_),
    .Y(_1821_));
 sg13g2_a21oi_1 _2629_ (.A1(_1816_),
    .A2(_1821_),
    .Y(_1822_),
    .B1(_1809_));
 sg13g2_or4_1 _2630_ (.A(_1780_),
    .B(_1787_),
    .C(_1807_),
    .D(_1822_),
    .X(_1823_));
 sg13g2_nand2_1 _2631_ (.Y(_1824_),
    .A(_1575_),
    .B(_1755_));
 sg13g2_nor2_1 _2632_ (.A(net793),
    .B(_1679_),
    .Y(_1825_));
 sg13g2_nand2_1 _2633_ (.Y(_1826_),
    .A(net816),
    .B(_1675_));
 sg13g2_nand3_1 _2634_ (.B(_1680_),
    .C(_1826_),
    .A(net790),
    .Y(_1827_));
 sg13g2_nor2_2 _2635_ (.A(net850),
    .B(net869),
    .Y(_1828_));
 sg13g2_nor3_2 _2636_ (.A(net847),
    .B(net840),
    .C(net868),
    .Y(_1829_));
 sg13g2_nand3_1 _2637_ (.B(net838),
    .C(_1640_),
    .A(net861),
    .Y(_1830_));
 sg13g2_a22oi_1 _2638_ (.Y(_1831_),
    .B1(net805),
    .B2(_1830_),
    .A2(net825),
    .A1(net828));
 sg13g2_nand3_1 _2639_ (.B(net860),
    .C(net838),
    .A(_1594_),
    .Y(_1832_));
 sg13g2_nor2_1 _2640_ (.A(net870),
    .B(_1832_),
    .Y(_1833_));
 sg13g2_o21ai_1 _2641_ (.B1(net818),
    .Y(_1834_),
    .A1(_1630_),
    .A2(_1832_));
 sg13g2_nand2_1 _2642_ (.Y(_1835_),
    .A(_1831_),
    .B(_1834_));
 sg13g2_a221oi_1 _2643_ (.B2(net902),
    .C1(net919),
    .B1(_1835_),
    .A1(net930),
    .Y(_1836_),
    .A2(_1827_));
 sg13g2_nand2_1 _2644_ (.Y(_1837_),
    .A(net809),
    .B(_1706_));
 sg13g2_a21oi_2 _2645_ (.B1(net806),
    .Y(_1838_),
    .A2(_1705_),
    .A1(net860));
 sg13g2_o21ai_1 _2646_ (.B1(net908),
    .Y(_1839_),
    .A1(net782),
    .A2(_1838_));
 sg13g2_nand2_1 _2647_ (.Y(_1840_),
    .A(_1836_),
    .B(_1839_));
 sg13g2_nand2_1 _2648_ (.Y(_1841_),
    .A(net913),
    .B(_1840_));
 sg13g2_nand2_2 _2649_ (.Y(_1842_),
    .A(_1643_),
    .B(net818));
 sg13g2_nand3_1 _2650_ (.B(net818),
    .C(_1706_),
    .A(_1643_),
    .Y(_1843_));
 sg13g2_and3_1 _2651_ (.X(_1844_),
    .A(_1649_),
    .B(_1657_),
    .C(_1843_));
 sg13g2_nand2b_1 _2652_ (.Y(_1845_),
    .B(net919),
    .A_N(_1844_));
 sg13g2_o21ai_1 _2653_ (.B1(_1683_),
    .Y(_1846_),
    .A1(net850),
    .A2(_1705_));
 sg13g2_a21oi_2 _2654_ (.B1(net794),
    .Y(_1847_),
    .A2(_1846_),
    .A1(net807));
 sg13g2_a221oi_1 _2655_ (.B2(_1846_),
    .C1(_1838_),
    .B1(net806),
    .A1(net828),
    .Y(_1848_),
    .A2(net825));
 sg13g2_nand2b_1 _2656_ (.Y(_1849_),
    .B(net930),
    .A_N(_1848_));
 sg13g2_nand2_1 _2657_ (.Y(_1850_),
    .A(_1845_),
    .B(_1849_));
 sg13g2_a22oi_1 _2658_ (.Y(_1851_),
    .B1(_1763_),
    .B2(_1668_),
    .A2(_1692_),
    .A1(_1671_));
 sg13g2_nand3_1 _2659_ (.B(_1657_),
    .C(_1851_),
    .A(_1649_),
    .Y(_1852_));
 sg13g2_nand2_1 _2660_ (.Y(_1853_),
    .A(net902),
    .B(_1852_));
 sg13g2_nand2_2 _2661_ (.Y(_1854_),
    .A(_1645_),
    .B(net908));
 sg13g2_a21oi_2 _2662_ (.B1(net806),
    .Y(_1855_),
    .A2(_1793_),
    .A1(_1659_));
 sg13g2_nor2_1 _2663_ (.A(net782),
    .B(_1855_),
    .Y(_1856_));
 sg13g2_o21ai_1 _2664_ (.B1(_1853_),
    .Y(_1857_),
    .A1(_1854_),
    .A2(_1856_));
 sg13g2_o21ai_1 _2665_ (.B1(net915),
    .Y(_1858_),
    .A1(_1850_),
    .A2(_1857_));
 sg13g2_a21oi_1 _2666_ (.A1(_1841_),
    .A2(_1858_),
    .Y(_1859_),
    .B1(_1824_));
 sg13g2_a21oi_1 _2667_ (.A1(_1756_),
    .A2(_1823_),
    .Y(_1860_),
    .B1(_1541_));
 sg13g2_a21oi_1 _2668_ (.A1(net881),
    .A2(_1753_),
    .Y(_1861_),
    .B1(_1859_));
 sg13g2_nor2_1 _2669_ (.A(net915),
    .B(_1756_),
    .Y(_1862_));
 sg13g2_nand2_1 _2670_ (.Y(_1863_),
    .A(net914),
    .B(_1755_));
 sg13g2_nand3_1 _2671_ (.B(_1686_),
    .C(_1688_),
    .A(net917),
    .Y(_1864_));
 sg13g2_a21oi_1 _2672_ (.A1(_1703_),
    .A2(_1725_),
    .Y(_1865_),
    .B1(net911));
 sg13g2_a221oi_1 _2673_ (.B2(net907),
    .C1(_1865_),
    .B1(_1741_),
    .A1(_1722_),
    .Y(_1866_),
    .A2(net904));
 sg13g2_nand3_1 _2674_ (.B(_1864_),
    .C(_1866_),
    .A(net966),
    .Y(_1867_));
 sg13g2_nand2_1 _2675_ (.Y(_1868_),
    .A(net854),
    .B(net832));
 sg13g2_a221oi_1 _2676_ (.B2(net799),
    .C1(net917),
    .B1(_1716_),
    .A1(net832),
    .Y(_1869_),
    .A2(_1699_));
 sg13g2_nor4_1 _2677_ (.A(net941),
    .B(net845),
    .C(net842),
    .D(net868),
    .Y(_1870_));
 sg13g2_o21ai_1 _2678_ (.B1(net804),
    .Y(_1871_),
    .A1(net857),
    .A2(_1652_));
 sg13g2_and4_1 _2679_ (.A(net953),
    .B(_1661_),
    .C(_1702_),
    .D(_1871_),
    .X(_1872_));
 sg13g2_or4_1 _2680_ (.A(net889),
    .B(_1869_),
    .C(_1870_),
    .D(_1872_),
    .X(_1873_));
 sg13g2_nor2_2 _2681_ (.A(net966),
    .B(net792),
    .Y(_1874_));
 sg13g2_nand2_1 _2682_ (.Y(_1875_),
    .A(net935),
    .B(net788));
 sg13g2_o21ai_1 _2683_ (.B1(net940),
    .Y(_1876_),
    .A1(_1716_),
    .A2(_1768_));
 sg13g2_nor2_1 _2684_ (.A(net846),
    .B(_1810_),
    .Y(_1877_));
 sg13g2_nand2_1 _2685_ (.Y(_1878_),
    .A(_1792_),
    .B(_1811_));
 sg13g2_nand4_1 _2686_ (.B(net810),
    .C(_1876_),
    .A(_1637_),
    .Y(_1879_),
    .D(_1878_));
 sg13g2_a21oi_1 _2687_ (.A1(net798),
    .A2(_1695_),
    .Y(_1880_),
    .B1(_1716_));
 sg13g2_nand4_1 _2688_ (.B(net854),
    .C(_1719_),
    .A(net949),
    .Y(_1881_),
    .D(_1738_));
 sg13g2_nand3_1 _2689_ (.B(_1880_),
    .C(_1881_),
    .A(net799),
    .Y(_1882_));
 sg13g2_nand3_1 _2690_ (.B(_1879_),
    .C(_1882_),
    .A(net889),
    .Y(_1883_));
 sg13g2_nand3_1 _2691_ (.B(_1874_),
    .C(_1883_),
    .A(_1873_),
    .Y(_1884_));
 sg13g2_a21oi_1 _2692_ (.A1(_1867_),
    .A2(_1884_),
    .Y(_1885_),
    .B1(_1863_));
 sg13g2_o21ai_1 _2693_ (.B1(_1541_),
    .Y(_1886_),
    .A1(_1575_),
    .A2(_1885_));
 sg13g2_nand2_1 _2694_ (.Y(_1887_),
    .A(_1659_),
    .B(_1812_));
 sg13g2_a21oi_2 _2695_ (.B1(net849),
    .Y(_1888_),
    .A2(net866),
    .A1(net836));
 sg13g2_o21ai_1 _2696_ (.B1(net859),
    .Y(_1889_),
    .A1(net843),
    .A2(net831));
 sg13g2_nor2_1 _2697_ (.A(net859),
    .B(net867),
    .Y(_1890_));
 sg13g2_nand2_1 _2698_ (.Y(_1891_),
    .A(net850),
    .B(_1659_));
 sg13g2_o21ai_1 _2699_ (.B1(net867),
    .Y(_1892_),
    .A1(net837),
    .A2(net869));
 sg13g2_a22oi_1 _2700_ (.Y(_1893_),
    .B1(_1892_),
    .B2(net851),
    .A2(_1888_),
    .A1(_1812_));
 sg13g2_o21ai_1 _2701_ (.B1(net931),
    .Y(_1894_),
    .A1(net782),
    .A2(_1893_));
 sg13g2_nor3_2 _2702_ (.A(net852),
    .B(net844),
    .C(net831),
    .Y(_1895_));
 sg13g2_o21ai_1 _2703_ (.B1(net847),
    .Y(_1896_),
    .A1(net834),
    .A2(net831));
 sg13g2_a21oi_2 _2704_ (.B1(_1895_),
    .Y(_1897_),
    .A2(net797),
    .A1(net798));
 sg13g2_inv_1 _2705_ (.Y(_1898_),
    .A(_1897_));
 sg13g2_a21oi_2 _2706_ (.B1(net845),
    .Y(_1899_),
    .A2(net832),
    .A1(net879));
 sg13g2_o21ai_1 _2707_ (.B1(net860),
    .Y(_1900_),
    .A1(net837),
    .A2(net867));
 sg13g2_a21oi_1 _2708_ (.A1(_1650_),
    .A2(_1897_),
    .Y(_1901_),
    .B1(net905));
 sg13g2_nand3_1 _2709_ (.B(_1813_),
    .C(_1900_),
    .A(net791),
    .Y(_1902_));
 sg13g2_a21oi_2 _2710_ (.B1(net964),
    .Y(_1903_),
    .A2(_1902_),
    .A1(_1901_));
 sg13g2_nand2_1 _2711_ (.Y(_1904_),
    .A(_1673_),
    .B(_1681_));
 sg13g2_a21oi_2 _2712_ (.B1(net803),
    .Y(_1905_),
    .A2(_1904_),
    .A1(_1638_));
 sg13g2_o21ai_1 _2713_ (.B1(net902),
    .Y(_1906_),
    .A1(net782),
    .A2(_1905_));
 sg13g2_nand3_1 _2714_ (.B(_1903_),
    .C(_1906_),
    .A(_1894_),
    .Y(_1907_));
 sg13g2_nand2_1 _2715_ (.Y(_1908_),
    .A(net930),
    .B(_1852_));
 sg13g2_nand2b_1 _2716_ (.Y(_1909_),
    .B(_1804_),
    .A_N(_1854_));
 sg13g2_o21ai_1 _2717_ (.B1(_1790_),
    .Y(_1910_),
    .A1(net782),
    .A2(_1855_));
 sg13g2_nand4_1 _2718_ (.B(_1908_),
    .C(_1909_),
    .A(net964),
    .Y(_1911_),
    .D(_1910_));
 sg13g2_nand2b_1 _2719_ (.Y(_1912_),
    .B(net920),
    .A_N(_1848_));
 sg13g2_a21oi_1 _2720_ (.A1(_1907_),
    .A2(_1911_),
    .Y(_1913_),
    .B1(net913));
 sg13g2_a21oi_1 _2721_ (.A1(_1831_),
    .A2(_1834_),
    .Y(_1914_),
    .B1(net957));
 sg13g2_nand2_1 _2722_ (.Y(_1915_),
    .A(net957),
    .B(_1827_));
 sg13g2_a21oi_1 _2723_ (.A1(net957),
    .A2(_1827_),
    .Y(_1916_),
    .B1(_1914_));
 sg13g2_a21o_1 _2724_ (.A2(_1844_),
    .A1(net890),
    .B1(_1916_),
    .X(_1917_));
 sg13g2_a21oi_1 _2725_ (.A1(net890),
    .A2(_1916_),
    .Y(_1918_),
    .B1(net915));
 sg13g2_a221oi_1 _2726_ (.B2(_1918_),
    .C1(_1824_),
    .B1(_1917_),
    .A1(_1912_),
    .Y(_1919_),
    .A2(_1913_));
 sg13g2_nand2_2 _2727_ (.Y(_1920_),
    .A(net964),
    .B(net913));
 sg13g2_a21oi_1 _2728_ (.A1(_1639_),
    .A2(net814),
    .Y(_1921_),
    .B1(net955));
 sg13g2_and2_1 _2729_ (.A(_1638_),
    .B(_1673_),
    .X(_1922_));
 sg13g2_o21ai_1 _2730_ (.B1(_1921_),
    .Y(_1923_),
    .A1(net817),
    .A2(_1922_));
 sg13g2_nand2_1 _2731_ (.Y(_1924_),
    .A(net823),
    .B(_1774_));
 sg13g2_nand3_1 _2732_ (.B(_1801_),
    .C(_1924_),
    .A(net955),
    .Y(_1925_));
 sg13g2_nand3_1 _2733_ (.B(_1923_),
    .C(_1925_),
    .A(net789),
    .Y(_1926_));
 sg13g2_a21o_1 _2734_ (.A2(_1926_),
    .A1(_1728_),
    .B1(net887),
    .X(_1927_));
 sg13g2_a221oi_1 _2735_ (.B2(_1812_),
    .C1(net809),
    .B1(_1811_),
    .A1(net953),
    .Y(_1928_),
    .A2(_1731_));
 sg13g2_a221oi_1 _2736_ (.B2(_1928_),
    .C1(net792),
    .B1(_1791_),
    .A1(net814),
    .Y(_1929_),
    .A2(_1661_));
 sg13g2_o21ai_1 _2737_ (.B1(net888),
    .Y(_1930_),
    .A1(_1729_),
    .A2(_1929_));
 sg13g2_nand4_1 _2738_ (.B(net914),
    .C(_1927_),
    .A(net966),
    .Y(_1931_),
    .D(_1930_));
 sg13g2_a21oi_1 _2739_ (.A1(net786),
    .A2(_1891_),
    .Y(_1932_),
    .B1(net933));
 sg13g2_a21oi_1 _2740_ (.A1(net957),
    .A2(_1846_),
    .Y(_1933_),
    .B1(net819));
 sg13g2_nor3_1 _2741_ (.A(net794),
    .B(_1760_),
    .C(_1933_),
    .Y(_1934_));
 sg13g2_a21oi_2 _2742_ (.B1(_1775_),
    .Y(_1935_),
    .A2(_1714_),
    .A1(_1670_));
 sg13g2_nor4_1 _2743_ (.A(net949),
    .B(_1759_),
    .C(_1934_),
    .D(_1935_),
    .Y(_1936_));
 sg13g2_a221oi_1 _2744_ (.B2(_1932_),
    .C1(_1936_),
    .B1(_1773_),
    .A1(_1664_),
    .Y(_1937_),
    .A2(net909));
 sg13g2_nand2b_1 _2745_ (.Y(_1938_),
    .B(_1808_),
    .A_N(_1937_));
 sg13g2_o21ai_1 _2746_ (.B1(_1868_),
    .Y(_1939_),
    .A1(_1681_),
    .A2(_1737_));
 sg13g2_nand2_1 _2747_ (.Y(_1940_),
    .A(net817),
    .B(_1939_));
 sg13g2_nand2_1 _2748_ (.Y(_1941_),
    .A(_1847_),
    .B(_1940_));
 sg13g2_nor2_1 _2749_ (.A(_1644_),
    .B(net890),
    .Y(_1942_));
 sg13g2_nand2_1 _2750_ (.Y(_1943_),
    .A(_1645_),
    .B(net887));
 sg13g2_nor2_2 _2751_ (.A(net940),
    .B(_1762_),
    .Y(_1944_));
 sg13g2_nand2_1 _2752_ (.Y(_1945_),
    .A(net832),
    .B(_1670_));
 sg13g2_a221oi_1 _2753_ (.B2(_1707_),
    .C1(net794),
    .B1(_1945_),
    .A1(_1842_),
    .Y(_1946_),
    .A2(_1944_));
 sg13g2_o21ai_1 _2754_ (.B1(_1946_),
    .Y(_1947_),
    .A1(net958),
    .A2(_1940_));
 sg13g2_a22oi_1 _2755_ (.Y(_1948_),
    .B1(_1942_),
    .B2(_1947_),
    .A2(_1941_),
    .A1(_1790_));
 sg13g2_a21o_1 _2756_ (.A2(net819),
    .A1(_1639_),
    .B1(net782),
    .X(_1949_));
 sg13g2_a21oi_1 _2757_ (.A1(net908),
    .A2(_1949_),
    .Y(_1950_),
    .B1(_1747_));
 sg13g2_nor2_2 _2758_ (.A(net881),
    .B(_1755_),
    .Y(_1951_));
 sg13g2_a21oi_1 _2759_ (.A1(net787),
    .A2(_1818_),
    .Y(_1952_),
    .B1(_1729_));
 sg13g2_o21ai_1 _2760_ (.B1(_1579_),
    .Y(_1953_),
    .A1(net900),
    .A2(_1952_));
 sg13g2_nor2_2 _2761_ (.A(net794),
    .B(_1642_),
    .Y(_1954_));
 sg13g2_a21oi_2 _2762_ (.B1(_1644_),
    .Y(_1955_),
    .A2(_1954_),
    .A1(_1770_));
 sg13g2_a21oi_1 _2763_ (.A1(_1676_),
    .A2(_1736_),
    .Y(_1956_),
    .B1(net814));
 sg13g2_nor2_2 _2764_ (.A(net939),
    .B(net819),
    .Y(_1957_));
 sg13g2_mux2_2 _2765_ (.A0(net868),
    .A1(_1693_),
    .S(net839),
    .X(_1958_));
 sg13g2_nand2_2 _2766_ (.Y(_1959_),
    .A(net848),
    .B(_1958_));
 sg13g2_a21oi_1 _2767_ (.A1(_1957_),
    .A2(_1959_),
    .Y(_1960_),
    .B1(_1956_));
 sg13g2_nand2_1 _2768_ (.Y(_1961_),
    .A(_1772_),
    .B(_1960_));
 sg13g2_a221oi_1 _2769_ (.B2(net887),
    .C1(_1953_),
    .B1(_1961_),
    .A1(net909),
    .Y(_1962_),
    .A2(_1955_));
 sg13g2_a21oi_1 _2770_ (.A1(_1948_),
    .A2(_1950_),
    .Y(_1963_),
    .B1(_1962_));
 sg13g2_nand4_1 _2771_ (.B(_1938_),
    .C(_1951_),
    .A(_1931_),
    .Y(_1964_),
    .D(_1963_));
 sg13g2_nor2_1 _2772_ (.A(_1886_),
    .B(_1919_),
    .Y(_1965_));
 sg13g2_a221oi_1 _2773_ (.B2(_1965_),
    .C1(\nyanframe[2] ),
    .B1(_1964_),
    .A1(_1860_),
    .Y(_1966_),
    .A2(_1861_));
 sg13g2_nor2_1 _2774_ (.A(net967),
    .B(\hvsync_gen.hpos[9] ),
    .Y(_1967_));
 sg13g2_nand2_1 _2775_ (.Y(_1968_),
    .A(net967),
    .B(\hvsync_gen.hpos[9] ));
 sg13g2_nor2b_1 _2776_ (.A(_1967_),
    .B_N(_1968_),
    .Y(_1969_));
 sg13g2_nand3_1 _2777_ (.B(_0033_),
    .C(_1617_),
    .A(_1543_),
    .Y(_1970_));
 sg13g2_xnor2_1 _2778_ (.Y(_1971_),
    .A(_1969_),
    .B(_1970_));
 sg13g2_o21ai_1 _2779_ (.B1(_1755_),
    .Y(_1972_),
    .A1(net947),
    .A2(net919));
 sg13g2_nand2_1 _2780_ (.Y(_1973_),
    .A(\hvsync_gen.vpos[8] ),
    .B(_1533_));
 sg13g2_a21oi_1 _2781_ (.A1(_0037_),
    .A2(_1973_),
    .Y(_1974_),
    .B1(_1573_));
 sg13g2_or2_1 _2782_ (.X(_1975_),
    .B(net189),
    .A(net942));
 sg13g2_a221oi_1 _2783_ (.B2(_1975_),
    .C1(_1974_),
    .B1(_1573_),
    .A1(_1532_),
    .Y(_1976_),
    .A2(net942));
 sg13g2_a21oi_1 _2784_ (.A1(net881),
    .A2(_1972_),
    .Y(_1977_),
    .B1(_1727_));
 sg13g2_nand3_1 _2785_ (.B(_1976_),
    .C(_1977_),
    .A(_1971_),
    .Y(_1978_));
 sg13g2_a221oi_1 _2786_ (.B2(_1897_),
    .C1(net941),
    .B1(_1800_),
    .A1(_1655_),
    .Y(_1979_),
    .A2(net785));
 sg13g2_nand2_2 _2787_ (.Y(_1980_),
    .A(net866),
    .B(_1714_));
 sg13g2_nand2b_1 _2788_ (.Y(_1981_),
    .B(_1980_),
    .A_N(_1774_));
 sg13g2_nand2_1 _2789_ (.Y(_1982_),
    .A(_1707_),
    .B(_1981_));
 sg13g2_o21ai_1 _2790_ (.B1(_1982_),
    .Y(_1983_),
    .A1(net949),
    .A2(_1772_));
 sg13g2_o21ai_1 _2791_ (.B1(net887),
    .Y(_1984_),
    .A1(_1979_),
    .A2(_1983_));
 sg13g2_o21ai_1 _2792_ (.B1(_1772_),
    .Y(_1985_),
    .A1(net817),
    .A2(_1791_));
 sg13g2_a21o_1 _2793_ (.A2(net859),
    .A1(net823),
    .B1(_1729_),
    .X(_1986_));
 sg13g2_a22oi_1 _2794_ (.Y(_1987_),
    .B1(_1986_),
    .B2(net910),
    .A2(_1985_),
    .A1(net904));
 sg13g2_a21oi_1 _2795_ (.A1(_1984_),
    .A2(_1987_),
    .Y(_1988_),
    .B1(_1580_));
 sg13g2_nand2b_1 _2796_ (.Y(_1989_),
    .B(_1954_),
    .A_N(_1956_));
 sg13g2_nand2_1 _2797_ (.Y(_1990_),
    .A(net909),
    .B(_1952_));
 sg13g2_a22oi_1 _2798_ (.Y(_1991_),
    .B1(_1990_),
    .B2(net900),
    .A2(_1989_),
    .A1(_1789_));
 sg13g2_o21ai_1 _2799_ (.B1(_1957_),
    .Y(_1992_),
    .A1(_1730_),
    .A2(_1899_));
 sg13g2_and4_1 _2800_ (.A(net887),
    .B(_1772_),
    .C(_1982_),
    .D(_1992_),
    .X(_1993_));
 sg13g2_nor3_1 _2801_ (.A(_1920_),
    .B(_1991_),
    .C(_1993_),
    .Y(_1994_));
 sg13g2_a21oi_1 _2802_ (.A1(_1650_),
    .A2(_1939_),
    .Y(_1995_),
    .B1(_1729_));
 sg13g2_xnor2_1 _2803_ (.Y(_1996_),
    .A(net879),
    .B(net855));
 sg13g2_or2_2 _2804_ (.X(_1997_),
    .B(_1996_),
    .A(_1652_));
 sg13g2_a221oi_1 _2805_ (.B2(net787),
    .C1(_1729_),
    .B1(_1997_),
    .A1(_1650_),
    .Y(_1998_),
    .A2(_1939_));
 sg13g2_nor2b_1 _2806_ (.A(_1998_),
    .B_N(_1782_),
    .Y(_1999_));
 sg13g2_or2_1 _2807_ (.X(_2000_),
    .B(_1798_),
    .A(net818));
 sg13g2_o21ai_1 _2808_ (.B1(_1995_),
    .Y(_2001_),
    .A1(net794),
    .A2(_2000_));
 sg13g2_nor2_1 _2809_ (.A(net822),
    .B(_1639_),
    .Y(_2002_));
 sg13g2_o21ai_1 _2810_ (.B1(net909),
    .Y(_2003_),
    .A1(_1624_),
    .A2(_1846_));
 sg13g2_nand2_1 _2811_ (.Y(_2004_),
    .A(net794),
    .B(net909));
 sg13g2_o21ai_1 _2812_ (.B1(_2004_),
    .Y(_2005_),
    .A1(_2002_),
    .A2(_2003_));
 sg13g2_a221oi_1 _2813_ (.B2(net931),
    .C1(_2005_),
    .B1(_2001_),
    .A1(net919),
    .Y(_2006_),
    .A2(_1955_));
 sg13g2_nor2_1 _2814_ (.A(_1809_),
    .B(_2006_),
    .Y(_2007_));
 sg13g2_nand2b_1 _2815_ (.Y(_2008_),
    .B(_1941_),
    .A_N(_1854_));
 sg13g2_a21oi_1 _2816_ (.A1(_1643_),
    .A2(_2000_),
    .Y(_2009_),
    .B1(net958));
 sg13g2_nand3b_1 _2817_ (.B(net955),
    .C(net822),
    .Y(_2010_),
    .A_N(_1922_));
 sg13g2_o21ai_1 _2818_ (.B1(_2010_),
    .Y(_2011_),
    .A1(net785),
    .A2(_1954_));
 sg13g2_o21ai_1 _2819_ (.B1(_1942_),
    .Y(_2012_),
    .A1(_2009_),
    .A2(_2011_));
 sg13g2_a21oi_1 _2820_ (.A1(_2008_),
    .A2(_2012_),
    .Y(_2013_),
    .B1(_1747_));
 sg13g2_or4_1 _2821_ (.A(_1988_),
    .B(_1994_),
    .C(_1999_),
    .D(_2013_),
    .X(_2014_));
 sg13g2_o21ai_1 _2822_ (.B1(_1756_),
    .Y(_2015_),
    .A1(_2007_),
    .A2(_2014_));
 sg13g2_nor4_1 _2823_ (.A(net953),
    .B(net809),
    .C(_1791_),
    .D(_1810_),
    .Y(_2016_));
 sg13g2_o21ai_1 _2824_ (.B1(_1671_),
    .Y(_2017_),
    .A1(_1705_),
    .A2(_1896_));
 sg13g2_a221oi_1 _2825_ (.B2(_2017_),
    .C1(_2016_),
    .B1(_1697_),
    .A1(_1636_),
    .Y(_2018_),
    .A2(net799));
 sg13g2_nand2_2 _2826_ (.Y(_2019_),
    .A(net947),
    .B(net891));
 sg13g2_a21oi_1 _2827_ (.A1(net843),
    .A2(_1699_),
    .Y(_2020_),
    .B1(_2019_));
 sg13g2_nand2_1 _2828_ (.Y(_2021_),
    .A(_2018_),
    .B(_2020_));
 sg13g2_nor3_1 _2829_ (.A(net809),
    .B(_1798_),
    .C(_1829_),
    .Y(_2022_));
 sg13g2_a21oi_1 _2830_ (.A1(_1637_),
    .A2(_1868_),
    .Y(_2023_),
    .B1(net799));
 sg13g2_nor3_1 _2831_ (.A(net953),
    .B(_2022_),
    .C(_2023_),
    .Y(_2024_));
 sg13g2_nor2_1 _2832_ (.A(net916),
    .B(net889),
    .Y(_2025_));
 sg13g2_o21ai_1 _2833_ (.B1(_2025_),
    .Y(_2026_),
    .A1(_1872_),
    .A2(_2024_));
 sg13g2_or2_2 _2834_ (.X(_2027_),
    .B(_1718_),
    .A(net858));
 sg13g2_a221oi_1 _2835_ (.B2(net858),
    .C1(_1743_),
    .B1(_1811_),
    .A1(net798),
    .Y(_2028_),
    .A2(_1708_));
 sg13g2_o21ai_1 _2836_ (.B1(_2028_),
    .Y(_2029_),
    .A1(_1837_),
    .A2(_2027_));
 sg13g2_nand3_1 _2837_ (.B(_2026_),
    .C(_2029_),
    .A(_2021_),
    .Y(_2030_));
 sg13g2_a21oi_1 _2838_ (.A1(net788),
    .A2(_2030_),
    .Y(_2031_),
    .B1(net935));
 sg13g2_a21oi_1 _2839_ (.A1(net832),
    .A2(_1699_),
    .Y(_2032_),
    .B1(net792));
 sg13g2_a21oi_1 _2840_ (.A1(_2018_),
    .A2(_2032_),
    .Y(_2033_),
    .B1(net887));
 sg13g2_nor4_1 _2841_ (.A(net792),
    .B(_1660_),
    .C(_1701_),
    .D(_2022_),
    .Y(_2034_));
 sg13g2_nor2_1 _2842_ (.A(net911),
    .B(_2034_),
    .Y(_2035_));
 sg13g2_a21oi_1 _2843_ (.A1(_1772_),
    .A2(_1871_),
    .Y(_2036_),
    .B1(net934));
 sg13g2_nor4_1 _2844_ (.A(net916),
    .B(_2033_),
    .C(_2035_),
    .D(_2036_),
    .Y(_2037_));
 sg13g2_nand2_1 _2845_ (.Y(_2038_),
    .A(_1648_),
    .B(_1748_));
 sg13g2_a221oi_1 _2846_ (.B2(net809),
    .C1(net914),
    .B1(_1877_),
    .A1(net845),
    .Y(_2039_),
    .A2(_1691_));
 sg13g2_nand4_1 _2847_ (.B(_1742_),
    .C(_2038_),
    .A(net788),
    .Y(_2040_),
    .D(_2039_));
 sg13g2_nand2_1 _2848_ (.Y(_2041_),
    .A(net935),
    .B(_2040_));
 sg13g2_o21ai_1 _2849_ (.B1(_1755_),
    .Y(_2042_),
    .A1(_2037_),
    .A2(_2041_));
 sg13g2_o21ai_1 _2850_ (.B1(net881),
    .Y(_2043_),
    .A1(_2031_),
    .A2(_2042_));
 sg13g2_or2_1 _2851_ (.X(_2044_),
    .B(_1798_),
    .A(_1660_));
 sg13g2_a221oi_1 _2852_ (.B2(net817),
    .C1(net958),
    .B1(_2044_),
    .A1(_1699_),
    .Y(_2045_),
    .A2(_1887_));
 sg13g2_a22oi_1 _2853_ (.Y(_2046_),
    .B1(_1847_),
    .B2(_2045_),
    .A2(_1845_),
    .A1(net912));
 sg13g2_a21o_1 _2854_ (.A2(_1764_),
    .A1(_1761_),
    .B1(_1895_),
    .X(_2047_));
 sg13g2_a221oi_1 _2855_ (.B2(net958),
    .C1(net782),
    .B1(_2047_),
    .A1(_1697_),
    .Y(_2048_),
    .A2(_1898_));
 sg13g2_nor2_1 _2856_ (.A(net888),
    .B(_2048_),
    .Y(_2049_));
 sg13g2_o21ai_1 _2857_ (.B1(_1808_),
    .Y(_2050_),
    .A1(_2046_),
    .A2(_2049_));
 sg13g2_o21ai_1 _2858_ (.B1(net908),
    .Y(_2051_),
    .A1(net782),
    .A2(_1905_));
 sg13g2_o21ai_1 _2859_ (.B1(net902),
    .Y(_2052_),
    .A1(_1658_),
    .A2(_1893_));
 sg13g2_nand4_1 _2860_ (.B(_1849_),
    .C(_2051_),
    .A(_1845_),
    .Y(_2053_),
    .D(_2052_));
 sg13g2_a22oi_1 _2861_ (.Y(_2054_),
    .B1(_2053_),
    .B2(_1746_),
    .A2(_1840_),
    .A1(net913));
 sg13g2_a21o_1 _2862_ (.A2(_2054_),
    .A1(_2050_),
    .B1(_1824_),
    .X(_2055_));
 sg13g2_and2_1 _2863_ (.A(_2043_),
    .B(_2055_),
    .X(_2056_));
 sg13g2_a21oi_1 _2864_ (.A1(_2015_),
    .A2(_2056_),
    .Y(_2057_),
    .B1(_1539_));
 sg13g2_nor3_1 _2865_ (.A(_1966_),
    .B(_1978_),
    .C(_2057_),
    .Y(_2058_));
 sg13g2_nor3_1 _2866_ (.A(_1669_),
    .B(_1684_),
    .C(_1768_),
    .Y(_2059_));
 sg13g2_o21ai_1 _2867_ (.B1(_1831_),
    .Y(_2060_),
    .A1(net805),
    .A2(_2059_));
 sg13g2_o21ai_1 _2868_ (.B1(net891),
    .Y(_2061_),
    .A1(_1914_),
    .A2(_2060_));
 sg13g2_a22oi_1 _2869_ (.Y(_2062_),
    .B1(net851),
    .B2(net805),
    .A2(net825),
    .A1(net828));
 sg13g2_nand2_1 _2870_ (.Y(_2063_),
    .A(net805),
    .B(_1738_));
 sg13g2_nand3_1 _2871_ (.B(_2062_),
    .C(_2063_),
    .A(_1834_),
    .Y(_2064_));
 sg13g2_a21oi_1 _2872_ (.A1(net930),
    .A2(_2064_),
    .Y(_2065_),
    .B1(net913));
 sg13g2_nand4_1 _2873_ (.B(net861),
    .C(net837),
    .A(net870),
    .Y(_2066_),
    .D(net786));
 sg13g2_nand2_1 _2874_ (.Y(_2067_),
    .A(net852),
    .B(_1738_));
 sg13g2_nor2_1 _2875_ (.A(_1828_),
    .B(_1888_),
    .Y(_2068_));
 sg13g2_nand3_1 _2876_ (.B(_2067_),
    .C(_2068_),
    .A(_1650_),
    .Y(_2069_));
 sg13g2_nand3_1 _2877_ (.B(_2066_),
    .C(_2069_),
    .A(net947),
    .Y(_2070_));
 sg13g2_nand3_1 _2878_ (.B(_2065_),
    .C(_2070_),
    .A(_2061_),
    .Y(_2071_));
 sg13g2_nand2_1 _2879_ (.Y(_2072_),
    .A(net790),
    .B(_1895_));
 sg13g2_a21oi_1 _2880_ (.A1(net939),
    .A2(_2072_),
    .Y(_2073_),
    .B1(_2019_));
 sg13g2_a21oi_1 _2881_ (.A1(_1915_),
    .A2(_2073_),
    .Y(_2074_),
    .B1(_1756_));
 sg13g2_a21oi_1 _2882_ (.A1(_2071_),
    .A2(_2074_),
    .Y(_2075_),
    .B1(_1574_));
 sg13g2_nor2_1 _2883_ (.A(net794),
    .B(_1832_),
    .Y(_2076_));
 sg13g2_a22oi_1 _2884_ (.Y(_2077_),
    .B1(net806),
    .B2(_1832_),
    .A2(net825),
    .A1(net828));
 sg13g2_nor3_2 _2885_ (.A(net855),
    .B(net834),
    .C(_1693_),
    .Y(_2078_));
 sg13g2_nor2_1 _2886_ (.A(_1670_),
    .B(_1719_),
    .Y(_2079_));
 sg13g2_o21ai_1 _2887_ (.B1(net814),
    .Y(_2080_),
    .A1(_1670_),
    .A2(_1719_));
 sg13g2_o21ai_1 _2888_ (.B1(_2077_),
    .Y(_2081_),
    .A1(_2078_),
    .A2(_2080_));
 sg13g2_nand2_2 _2889_ (.Y(_2082_),
    .A(net784),
    .B(_1829_));
 sg13g2_a21oi_1 _2890_ (.A1(net784),
    .A2(_1829_),
    .Y(_2083_),
    .B1(net949));
 sg13g2_a21oi_2 _2891_ (.B1(net912),
    .Y(_2084_),
    .A2(_1829_),
    .A1(net784));
 sg13g2_a21oi_1 _2892_ (.A1(net920),
    .A2(_2081_),
    .Y(_2085_),
    .B1(_2084_));
 sg13g2_a221oi_1 _2893_ (.B2(_2027_),
    .C1(net808),
    .B1(_1900_),
    .A1(net829),
    .Y(_2086_),
    .A2(net826));
 sg13g2_nor3_2 _2894_ (.A(net847),
    .B(net839),
    .C(_1692_),
    .Y(_2087_));
 sg13g2_a221oi_1 _2895_ (.B2(_1694_),
    .C1(net811),
    .B1(net855),
    .A1(net827),
    .Y(_2088_),
    .A2(net824));
 sg13g2_or3_2 _2896_ (.A(_1729_),
    .B(_2086_),
    .C(_2088_),
    .X(_2089_));
 sg13g2_and2_1 _2897_ (.A(net908),
    .B(_2089_),
    .X(_2090_));
 sg13g2_nand2_2 _2898_ (.Y(_2091_),
    .A(net801),
    .B(_1958_));
 sg13g2_nand2_1 _2899_ (.Y(_2092_),
    .A(_2062_),
    .B(_2091_));
 sg13g2_a21oi_1 _2900_ (.A1(_2062_),
    .A2(_2091_),
    .Y(_2093_),
    .B1(_1644_));
 sg13g2_o21ai_1 _2901_ (.B1(net903),
    .Y(_2094_),
    .A1(_2086_),
    .A2(_2093_));
 sg13g2_nand3_1 _2902_ (.B(_2085_),
    .C(_2094_),
    .A(_1577_),
    .Y(_2095_));
 sg13g2_nand2_1 _2903_ (.Y(_2096_),
    .A(_1702_),
    .B(_1830_));
 sg13g2_a22oi_1 _2904_ (.Y(_2097_),
    .B1(_2096_),
    .B2(net784),
    .A2(_1833_),
    .A1(_1800_));
 sg13g2_o21ai_1 _2905_ (.B1(net888),
    .Y(_2098_),
    .A1(_2083_),
    .A2(_2097_));
 sg13g2_a21oi_1 _2906_ (.A1(_1831_),
    .A2(_1842_),
    .Y(_2099_),
    .B1(net905));
 sg13g2_a21oi_1 _2907_ (.A1(_1721_),
    .A2(_1828_),
    .Y(_2100_),
    .B1(net901));
 sg13g2_nor3_1 _2908_ (.A(net916),
    .B(_2099_),
    .C(_2100_),
    .Y(_2101_));
 sg13g2_and2_1 _2909_ (.A(_2098_),
    .B(_2101_),
    .X(_2102_));
 sg13g2_o21ai_1 _2910_ (.B1(_1756_),
    .Y(_2103_),
    .A1(_2090_),
    .A2(_2095_));
 sg13g2_o21ai_1 _2911_ (.B1(_2075_),
    .Y(_2104_),
    .A1(_2102_),
    .A2(_2103_));
 sg13g2_nor2_1 _2912_ (.A(_1575_),
    .B(_1863_),
    .Y(_2105_));
 sg13g2_nand2_2 _2913_ (.Y(_2106_),
    .A(net881),
    .B(_1862_));
 sg13g2_a21oi_1 _2914_ (.A1(net784),
    .A2(_1895_),
    .Y(_2107_),
    .B1(net939));
 sg13g2_nor3_1 _2915_ (.A(net891),
    .B(_2106_),
    .C(_2107_),
    .Y(_2108_));
 sg13g2_a221oi_1 _2916_ (.B2(_1674_),
    .C1(net792),
    .B1(_1668_),
    .A1(_1637_),
    .Y(_2109_),
    .A2(net810));
 sg13g2_o21ai_1 _2917_ (.B1(_2108_),
    .Y(_2110_),
    .A1(net957),
    .A2(_2109_));
 sg13g2_nand2_1 _2918_ (.Y(_2111_),
    .A(_2104_),
    .B(_2110_));
 sg13g2_nand2_2 _2919_ (.Y(_2112_),
    .A(_1539_),
    .B(\nyanframe[1] ));
 sg13g2_a21oi_1 _2920_ (.A1(net784),
    .A2(_1895_),
    .Y(_2113_),
    .B1(net906));
 sg13g2_nor3_2 _2921_ (.A(_1660_),
    .B(_1783_),
    .C(_1798_),
    .Y(_2114_));
 sg13g2_nor2_1 _2922_ (.A(net806),
    .B(_2114_),
    .Y(_2115_));
 sg13g2_o21ai_1 _2923_ (.B1(net930),
    .Y(_2116_),
    .A1(_2092_),
    .A2(_2115_));
 sg13g2_a22oi_1 _2924_ (.Y(_2117_),
    .B1(_2114_),
    .B2(_1800_),
    .A2(_2087_),
    .A1(net785));
 sg13g2_a21oi_1 _2925_ (.A1(net902),
    .A2(_2117_),
    .Y(_2118_),
    .B1(_1747_));
 sg13g2_o21ai_1 _2926_ (.B1(net930),
    .Y(_2119_),
    .A1(_2086_),
    .A2(_2093_));
 sg13g2_a21oi_1 _2927_ (.A1(net902),
    .A2(_2089_),
    .Y(_2120_),
    .B1(_1809_));
 sg13g2_a22oi_1 _2928_ (.Y(_2121_),
    .B1(_2119_),
    .B2(_2120_),
    .A2(_2118_),
    .A1(_2116_));
 sg13g2_o21ai_1 _2929_ (.B1(net811),
    .Y(_2122_),
    .A1(_1719_),
    .A2(_1996_));
 sg13g2_a21oi_1 _2930_ (.A1(_2077_),
    .A2(_2122_),
    .Y(_2123_),
    .B1(net965));
 sg13g2_a21oi_1 _2931_ (.A1(net965),
    .A2(_2081_),
    .Y(_2124_),
    .B1(_2123_));
 sg13g2_a21oi_1 _2932_ (.A1(_1721_),
    .A2(_1828_),
    .Y(_2125_),
    .B1(net911));
 sg13g2_a21oi_1 _2933_ (.A1(_1831_),
    .A2(_1842_),
    .Y(_2126_),
    .B1(net901));
 sg13g2_nor3_1 _2934_ (.A(net915),
    .B(_2125_),
    .C(_2126_),
    .Y(_2127_));
 sg13g2_o21ai_1 _2935_ (.B1(_2127_),
    .Y(_2128_),
    .A1(net905),
    .A2(_2124_));
 sg13g2_o21ai_1 _2936_ (.B1(_2128_),
    .Y(_2129_),
    .A1(_2113_),
    .A2(_2121_));
 sg13g2_nand3_1 _2937_ (.B(net950),
    .C(_2082_),
    .A(net957),
    .Y(_2130_));
 sg13g2_nand3_1 _2938_ (.B(_2129_),
    .C(_2130_),
    .A(_1951_),
    .Y(_2131_));
 sg13g2_nand3_1 _2939_ (.B(_2066_),
    .C(_2069_),
    .A(net908),
    .Y(_2132_));
 sg13g2_a221oi_1 _2940_ (.B2(net902),
    .C1(_1576_),
    .B1(_2072_),
    .A1(net930),
    .Y(_2133_),
    .A2(_1827_));
 sg13g2_a221oi_1 _2941_ (.B2(net930),
    .C1(net913),
    .B1(_2060_),
    .A1(net902),
    .Y(_2134_),
    .A2(_1835_));
 sg13g2_a22oi_1 _2942_ (.Y(_2135_),
    .B1(_2097_),
    .B2(net908),
    .A2(_2064_),
    .A1(net919));
 sg13g2_a22oi_1 _2943_ (.Y(_2136_),
    .B1(_2134_),
    .B2(_2135_),
    .A2(_2133_),
    .A1(_2132_));
 sg13g2_or2_1 _2944_ (.X(_2137_),
    .B(_2136_),
    .A(_1824_));
 sg13g2_nand3_1 _2945_ (.B(net821),
    .C(_1653_),
    .A(net936),
    .Y(_2138_));
 sg13g2_nand4_1 _2946_ (.B(_2105_),
    .C(_2109_),
    .A(_1742_),
    .Y(_2139_),
    .D(_2138_));
 sg13g2_nand4_1 _2947_ (.B(_2131_),
    .C(_2137_),
    .A(_1539_),
    .Y(_2140_),
    .D(_2139_));
 sg13g2_a22oi_1 _2948_ (.Y(_2141_),
    .B1(_2112_),
    .B2(_2140_),
    .A2(_2111_),
    .A1(\nyanframe[1] ));
 sg13g2_a21oi_1 _2949_ (.A1(_2077_),
    .A2(_2122_),
    .Y(_2142_),
    .B1(net933));
 sg13g2_a221oi_1 _2950_ (.B2(_1800_),
    .C1(net905),
    .B1(_2114_),
    .A1(net785),
    .Y(_2143_),
    .A2(_2087_));
 sg13g2_nor4_1 _2951_ (.A(net913),
    .B(_2084_),
    .C(_2142_),
    .D(_2143_),
    .Y(_2144_));
 sg13g2_nor3_1 _2952_ (.A(net964),
    .B(_2102_),
    .C(_2144_),
    .Y(_2145_));
 sg13g2_o21ai_1 _2953_ (.B1(_1831_),
    .Y(_2146_),
    .A1(_1642_),
    .A2(_2122_));
 sg13g2_nand2_1 _2954_ (.Y(_2147_),
    .A(net910),
    .B(_2146_));
 sg13g2_a21oi_1 _2955_ (.A1(net786),
    .A2(_2096_),
    .Y(_2148_),
    .B1(net933));
 sg13g2_nor3_1 _2956_ (.A(_2084_),
    .B(_2100_),
    .C(_2148_),
    .Y(_2149_));
 sg13g2_a21o_1 _2957_ (.A2(_2149_),
    .A1(_2147_),
    .B1(_1920_),
    .X(_2150_));
 sg13g2_o21ai_1 _2958_ (.B1(_1782_),
    .Y(_2151_),
    .A1(_2092_),
    .A2(_2115_));
 sg13g2_a21oi_1 _2959_ (.A1(net786),
    .A2(_2087_),
    .Y(_2152_),
    .B1(net905));
 sg13g2_nor2b_1 _2960_ (.A(_2115_),
    .B_N(_1831_),
    .Y(_2153_));
 sg13g2_a221oi_1 _2961_ (.B2(net939),
    .C1(net891),
    .B1(_2153_),
    .A1(_1957_),
    .Y(_2154_),
    .A2(_2076_));
 sg13g2_o21ai_1 _2962_ (.B1(_1808_),
    .Y(_2155_),
    .A1(_2152_),
    .A2(_2154_));
 sg13g2_nand3_1 _2963_ (.B(_2151_),
    .C(_2155_),
    .A(_2150_),
    .Y(_2156_));
 sg13g2_o21ai_1 _2964_ (.B1(_1756_),
    .Y(_2157_),
    .A1(_2145_),
    .A2(_2156_));
 sg13g2_a21o_1 _2965_ (.A2(_2138_),
    .A1(_2109_),
    .B1(net957),
    .X(_2158_));
 sg13g2_a221oi_1 _2966_ (.B2(_2108_),
    .C1(_1539_),
    .B1(_2158_),
    .A1(_2075_),
    .Y(_2159_),
    .A2(_2157_));
 sg13g2_nor3_1 _2967_ (.A(_1978_),
    .B(_2141_),
    .C(_2159_),
    .Y(_2160_));
 sg13g2_or2_1 _2968_ (.X(_2161_),
    .B(_1695_),
    .A(net811));
 sg13g2_or2_1 _2969_ (.X(_2162_),
    .B(_2078_),
    .A(_1757_));
 sg13g2_o21ai_1 _2970_ (.B1(net868),
    .Y(_2163_),
    .A1(net871),
    .A2(net840));
 sg13g2_a221oi_1 _2971_ (.B2(_1672_),
    .C1(_1757_),
    .B1(_2163_),
    .A1(_1692_),
    .Y(_2164_),
    .A2(_1762_));
 sg13g2_nand2b_1 _2972_ (.Y(_2165_),
    .B(net812),
    .A_N(_2164_));
 sg13g2_o21ai_1 _2973_ (.B1(_2161_),
    .Y(_2166_),
    .A1(net802),
    .A2(_2164_));
 sg13g2_nor2_1 _2974_ (.A(net793),
    .B(_2166_),
    .Y(_2167_));
 sg13g2_nor2_1 _2975_ (.A(net900),
    .B(_2167_),
    .Y(_2168_));
 sg13g2_a22oi_1 _2976_ (.Y(_2169_),
    .B1(net800),
    .B2(_1889_),
    .A2(net826),
    .A1(net827));
 sg13g2_nor3_2 _2977_ (.A(net855),
    .B(net840),
    .C(_1693_),
    .Y(_2170_));
 sg13g2_nand2_1 _2978_ (.Y(_2171_),
    .A(_1636_),
    .B(_1692_));
 sg13g2_a221oi_1 _2979_ (.B2(net856),
    .C1(_2170_),
    .B1(_1980_),
    .A1(net872),
    .Y(_2172_),
    .A2(_1762_));
 sg13g2_o21ai_1 _2980_ (.B1(_2169_),
    .Y(_2173_),
    .A1(net800),
    .A2(_2172_));
 sg13g2_nand2_1 _2981_ (.Y(_2174_),
    .A(net907),
    .B(_2173_));
 sg13g2_a22oi_1 _2982_ (.Y(_2175_),
    .B1(_1737_),
    .B2(net797),
    .A2(_1695_),
    .A1(_1652_));
 sg13g2_nand2b_1 _2983_ (.Y(_2176_),
    .B(net812),
    .A_N(_2175_));
 sg13g2_o21ai_1 _2984_ (.B1(_1680_),
    .Y(_2177_),
    .A1(net801),
    .A2(_2175_));
 sg13g2_a21oi_2 _2985_ (.B1(net812),
    .Y(_2178_),
    .A2(_1958_),
    .A1(net856));
 sg13g2_nand2b_1 _2986_ (.Y(_2179_),
    .B(_1758_),
    .A_N(_2178_));
 sg13g2_a221oi_1 _2987_ (.B2(_1529_),
    .C1(net793),
    .B1(_2179_),
    .A1(net954),
    .Y(_2180_),
    .A2(_2177_));
 sg13g2_o21ai_1 _2988_ (.B1(_2174_),
    .Y(_2181_),
    .A1(net890),
    .A2(_2180_));
 sg13g2_o21ai_1 _2989_ (.B1(_1746_),
    .Y(_2182_),
    .A1(_2168_),
    .A2(_2181_));
 sg13g2_nand3_1 _2990_ (.B(_1673_),
    .C(_1980_),
    .A(net802),
    .Y(_2183_));
 sg13g2_inv_1 _2991_ (.Y(_2184_),
    .A(_2183_));
 sg13g2_o21ai_1 _2992_ (.B1(net812),
    .Y(_0186_),
    .A1(_2079_),
    .A2(_2162_));
 sg13g2_a21oi_1 _2993_ (.A1(_2183_),
    .A2(_0186_),
    .Y(_0187_),
    .B1(net906));
 sg13g2_nand3_1 _2994_ (.B(_1676_),
    .C(_1719_),
    .A(net803),
    .Y(_0188_));
 sg13g2_a22oi_1 _2995_ (.Y(_0189_),
    .B1(_1772_),
    .B2(_0188_),
    .A2(net900),
    .A1(net789));
 sg13g2_nor3_1 _2996_ (.A(_1660_),
    .B(_1798_),
    .C(_1828_),
    .Y(_0190_));
 sg13g2_o21ai_1 _2997_ (.B1(net813),
    .Y(_0191_),
    .A1(_1701_),
    .A2(_2170_));
 sg13g2_o21ai_1 _2998_ (.B1(_0191_),
    .Y(_0192_),
    .A1(net814),
    .A2(_0190_));
 sg13g2_nand3_1 _2999_ (.B(_1673_),
    .C(_1704_),
    .A(net802),
    .Y(_0193_));
 sg13g2_or3_2 _3000_ (.A(net801),
    .B(_1694_),
    .C(_1896_),
    .X(_0194_));
 sg13g2_nand4_1 _3001_ (.B(net811),
    .C(net798),
    .A(net856),
    .Y(_0195_),
    .D(_1706_));
 sg13g2_nand2_1 _3002_ (.Y(_0196_),
    .A(_0194_),
    .B(_0195_));
 sg13g2_nand3_1 _3003_ (.B(_0194_),
    .C(_0195_),
    .A(_0193_),
    .Y(_0197_));
 sg13g2_a221oi_1 _3004_ (.B2(net918),
    .C1(_0189_),
    .B1(_0197_),
    .A1(net932),
    .Y(_0198_),
    .A2(_0192_));
 sg13g2_nand2b_1 _3005_ (.Y(_0199_),
    .B(_0198_),
    .A_N(_0187_));
 sg13g2_a21oi_1 _3006_ (.A1(_1579_),
    .A2(_0199_),
    .Y(_0200_),
    .B1(_1755_));
 sg13g2_a21oi_2 _3007_ (.B1(net801),
    .Y(_0201_),
    .A2(_2171_),
    .A1(_1997_));
 sg13g2_nand3_1 _3008_ (.B(net798),
    .C(_1706_),
    .A(_1670_),
    .Y(_0202_));
 sg13g2_o21ai_1 _3009_ (.B1(net940),
    .Y(_0203_),
    .A1(net812),
    .A2(_0202_));
 sg13g2_a21oi_1 _3010_ (.A1(net812),
    .A2(_2170_),
    .Y(_0204_),
    .B1(net954));
 sg13g2_nand3_1 _3011_ (.B(_1636_),
    .C(net811),
    .A(net878),
    .Y(_0205_));
 sg13g2_nand3_1 _3012_ (.B(_0193_),
    .C(_0205_),
    .A(net954),
    .Y(_0206_));
 sg13g2_o21ai_1 _3013_ (.B1(_0206_),
    .Y(_0207_),
    .A1(_0201_),
    .A2(_0203_));
 sg13g2_nand2_1 _3014_ (.Y(_0208_),
    .A(_1645_),
    .B(net889));
 sg13g2_a21o_1 _3015_ (.A2(_0207_),
    .A1(net788),
    .B1(_0208_),
    .X(_0209_));
 sg13g2_nand3_1 _3016_ (.B(net813),
    .C(_1705_),
    .A(net849),
    .Y(_0210_));
 sg13g2_o21ai_1 _3017_ (.B1(net803),
    .Y(_0211_),
    .A1(_1640_),
    .A2(net797));
 sg13g2_nand3_1 _3018_ (.B(_0210_),
    .C(_0211_),
    .A(net789),
    .Y(_0212_));
 sg13g2_nand2_1 _3019_ (.Y(_0213_),
    .A(net836),
    .B(_1699_));
 sg13g2_nand3_1 _3020_ (.B(_0210_),
    .C(_0213_),
    .A(_1825_),
    .Y(_0214_));
 sg13g2_a22oi_1 _3021_ (.Y(_0215_),
    .B1(_0214_),
    .B2(net917),
    .A2(_0212_),
    .A1(net932));
 sg13g2_a21o_1 _3022_ (.A2(_0215_),
    .A1(_0209_),
    .B1(_1920_),
    .X(_0216_));
 sg13g2_a221oi_1 _3023_ (.B2(_1888_),
    .C1(_2170_),
    .B1(_1812_),
    .A1(net849),
    .Y(_0217_),
    .A2(net832));
 sg13g2_nor2_1 _3024_ (.A(net802),
    .B(_0217_),
    .Y(_0218_));
 sg13g2_nand2_1 _3025_ (.Y(_0219_),
    .A(net848),
    .B(_1980_));
 sg13g2_nor2_1 _3026_ (.A(net940),
    .B(_1829_),
    .Y(_0220_));
 sg13g2_a22oi_1 _3027_ (.Y(_0221_),
    .B1(_0219_),
    .B2(_0220_),
    .A2(net812),
    .A1(net954));
 sg13g2_nand2b_1 _3028_ (.Y(_0222_),
    .B(_0204_),
    .A_N(_2178_));
 sg13g2_o21ai_1 _3029_ (.B1(_0222_),
    .Y(_0223_),
    .A1(_0218_),
    .A2(_0221_));
 sg13g2_a21oi_1 _3030_ (.A1(net788),
    .A2(_0223_),
    .Y(_0224_),
    .B1(_1943_));
 sg13g2_a21o_1 _3031_ (.A2(net835),
    .A1(net878),
    .B1(_1718_),
    .X(_0225_));
 sg13g2_nand4_1 _3032_ (.B(net868),
    .C(net811),
    .A(net855),
    .Y(_0226_),
    .D(_0225_));
 sg13g2_nand3_1 _3033_ (.B(_0194_),
    .C(_0226_),
    .A(_2161_),
    .Y(_0227_));
 sg13g2_o21ai_1 _3034_ (.B1(_1790_),
    .Y(_0228_),
    .A1(net792),
    .A2(_0227_));
 sg13g2_o21ai_1 _3035_ (.B1(net817),
    .Y(_0229_),
    .A1(_1783_),
    .A2(_1890_));
 sg13g2_nand2_1 _3036_ (.Y(_0230_),
    .A(_2169_),
    .B(_0229_));
 sg13g2_nand2_1 _3037_ (.Y(_0231_),
    .A(net907),
    .B(_0230_));
 sg13g2_nand2_1 _3038_ (.Y(_0232_),
    .A(_0228_),
    .B(_0231_));
 sg13g2_o21ai_1 _3039_ (.B1(_1808_),
    .Y(_0233_),
    .A1(_0224_),
    .A2(_0232_));
 sg13g2_nand4_1 _3040_ (.B(_0200_),
    .C(_0216_),
    .A(_2182_),
    .Y(_0234_),
    .D(_0233_));
 sg13g2_nand2_1 _3041_ (.Y(_0235_),
    .A(_1830_),
    .B(_2067_));
 sg13g2_a22oi_1 _3042_ (.Y(_0236_),
    .B1(_0235_),
    .B2(_1650_),
    .A2(net786),
    .A1(_1675_));
 sg13g2_and2_1 _3043_ (.A(_1700_),
    .B(_2169_),
    .X(_0237_));
 sg13g2_nand2_1 _3044_ (.Y(_0238_),
    .A(net903),
    .B(_0237_));
 sg13g2_o21ai_1 _3045_ (.B1(_0238_),
    .Y(_0239_),
    .A1(net905),
    .A2(_0236_));
 sg13g2_a21oi_1 _3046_ (.A1(net816),
    .A2(_1892_),
    .Y(_0240_),
    .B1(_1827_));
 sg13g2_a21o_1 _3047_ (.A2(_0225_),
    .A1(net868),
    .B1(net854),
    .X(_0241_));
 sg13g2_a21oi_1 _3048_ (.A1(_1748_),
    .A2(_1899_),
    .Y(_0242_),
    .B1(net799));
 sg13g2_a221oi_1 _3049_ (.B2(_0242_),
    .C1(net792),
    .B1(_0241_),
    .A1(_1668_),
    .Y(_0243_),
    .A2(_1674_));
 sg13g2_nand2b_1 _3050_ (.Y(_0244_),
    .B(net903),
    .A_N(_0243_));
 sg13g2_o21ai_1 _3051_ (.B1(_0244_),
    .Y(_0245_),
    .A1(net911),
    .A2(_0240_));
 sg13g2_and2_1 _3052_ (.A(_1736_),
    .B(_1899_),
    .X(_0246_));
 sg13g2_a21oi_1 _3053_ (.A1(_1736_),
    .A2(_1899_),
    .Y(_0247_),
    .B1(net813));
 sg13g2_a22oi_1 _3054_ (.Y(_0248_),
    .B1(_1768_),
    .B2(net866),
    .A2(_1693_),
    .A1(net847));
 sg13g2_a21oi_2 _3055_ (.B1(_0247_),
    .Y(_0249_),
    .A2(_0248_),
    .A1(net813));
 sg13g2_a22oi_1 _3056_ (.Y(_0250_),
    .B1(_1874_),
    .B2(_0249_),
    .A2(net906),
    .A1(net936));
 sg13g2_nand3_1 _3057_ (.B(_1652_),
    .C(_1675_),
    .A(net813),
    .Y(_0251_));
 sg13g2_nand4_1 _3058_ (.B(net817),
    .C(_1659_),
    .A(net850),
    .Y(_0252_),
    .D(_1761_));
 sg13g2_nand4_1 _3059_ (.B(_1680_),
    .C(_0251_),
    .A(net789),
    .Y(_0253_),
    .D(_0252_));
 sg13g2_nand2_1 _3060_ (.Y(_0254_),
    .A(net904),
    .B(_0253_));
 sg13g2_nor2_1 _3061_ (.A(net805),
    .B(_1761_),
    .Y(_0255_));
 sg13g2_o21ai_1 _3062_ (.B1(net931),
    .Y(_0256_),
    .A1(_1827_),
    .A2(_0255_));
 sg13g2_a21oi_1 _3063_ (.A1(_1675_),
    .A2(_1715_),
    .Y(_0257_),
    .B1(_1890_));
 sg13g2_a22oi_1 _3064_ (.Y(_0258_),
    .B1(_0257_),
    .B2(_1650_),
    .A2(_0246_),
    .A1(net787));
 sg13g2_a21oi_2 _3065_ (.B1(net935),
    .Y(_0259_),
    .A2(_0258_),
    .A1(net910));
 sg13g2_nand3_1 _3066_ (.B(_0256_),
    .C(_0259_),
    .A(_0254_),
    .Y(_0260_));
 sg13g2_o21ai_1 _3067_ (.B1(_0260_),
    .Y(_0261_),
    .A1(_0245_),
    .A2(_0250_));
 sg13g2_or2_1 _3068_ (.X(_0262_),
    .B(_1738_),
    .A(net821));
 sg13g2_nand3_1 _3069_ (.B(_2062_),
    .C(_0262_),
    .A(_1826_),
    .Y(_0263_));
 sg13g2_nand2_1 _3070_ (.Y(_0264_),
    .A(net915),
    .B(_1755_));
 sg13g2_a21oi_1 _3071_ (.A1(net947),
    .A2(_0263_),
    .Y(_0265_),
    .B1(_0264_));
 sg13g2_a22oi_1 _3072_ (.Y(_0266_),
    .B1(_0261_),
    .B2(_0265_),
    .A2(_0239_),
    .A1(_1862_));
 sg13g2_a21oi_1 _3073_ (.A1(_0234_),
    .A2(_0266_),
    .Y(_0267_),
    .B1(net881));
 sg13g2_a221oi_1 _3074_ (.B2(_1792_),
    .C1(_1682_),
    .B1(_1706_),
    .A1(net827),
    .Y(_0268_),
    .A2(net824));
 sg13g2_nor2_1 _3075_ (.A(net787),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_o21ai_1 _3076_ (.B1(_1683_),
    .Y(_0270_),
    .A1(_1676_),
    .A2(_1718_));
 sg13g2_a21oi_1 _3077_ (.A1(net804),
    .A2(_0270_),
    .Y(_0271_),
    .B1(_0269_));
 sg13g2_nor2b_1 _3078_ (.A(_0039_),
    .B_N(_0271_),
    .Y(_0272_));
 sg13g2_nand2_1 _3079_ (.Y(_0273_),
    .A(_1702_),
    .B(_1717_));
 sg13g2_a221oi_1 _3080_ (.B2(net917),
    .C1(net935),
    .B1(_0273_),
    .A1(net932),
    .Y(_0274_),
    .A2(_1686_));
 sg13g2_o21ai_1 _3081_ (.B1(_0274_),
    .Y(_0275_),
    .A1(net887),
    .A2(_0272_));
 sg13g2_a21oi_1 _3082_ (.A1(net846),
    .A2(_1980_),
    .Y(_0276_),
    .B1(_1768_));
 sg13g2_nor2_1 _3083_ (.A(net800),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_a21o_1 _3084_ (.A2(_1719_),
    .A1(_1648_),
    .B1(_0039_),
    .X(_0278_));
 sg13g2_o21ai_1 _3085_ (.B1(net889),
    .Y(_0279_),
    .A1(_0277_),
    .A2(_0278_));
 sg13g2_nor2_1 _3086_ (.A(net911),
    .B(_1679_),
    .Y(_0280_));
 sg13g2_nand3_1 _3087_ (.B(net810),
    .C(_1868_),
    .A(_1637_),
    .Y(_0281_));
 sg13g2_a21oi_1 _3088_ (.A1(net917),
    .A2(_0281_),
    .Y(_0282_),
    .B1(_0280_));
 sg13g2_nand4_1 _3089_ (.B(_1874_),
    .C(_0279_),
    .A(_1725_),
    .Y(_0283_),
    .D(_0282_));
 sg13g2_a21oi_1 _3090_ (.A1(_0275_),
    .A2(_0283_),
    .Y(_0284_),
    .B1(_2106_));
 sg13g2_or2_1 _3091_ (.X(_0285_),
    .B(_0284_),
    .A(\nyanframe[2] ));
 sg13g2_o21ai_1 _3092_ (.B1(_2112_),
    .Y(_0286_),
    .A1(_0267_),
    .A2(_0285_));
 sg13g2_and4_1 _3093_ (.A(net801),
    .B(_1676_),
    .C(net798),
    .D(_1706_),
    .X(_0287_));
 sg13g2_o21ai_1 _3094_ (.B1(net932),
    .Y(_0288_),
    .A1(_0218_),
    .A2(_0287_));
 sg13g2_nand3_1 _3095_ (.B(_1670_),
    .C(_1748_),
    .A(net801),
    .Y(_0289_));
 sg13g2_o21ai_1 _3096_ (.B1(_0289_),
    .Y(_0290_),
    .A1(net801),
    .A2(_2171_));
 sg13g2_o21ai_1 _3097_ (.B1(net918),
    .Y(_0291_),
    .A1(_1674_),
    .A2(_0201_));
 sg13g2_a22oi_1 _3098_ (.Y(_0292_),
    .B1(_0290_),
    .B2(net904),
    .A2(_0227_),
    .A1(net907));
 sg13g2_nand3_1 _3099_ (.B(_0291_),
    .C(_0292_),
    .A(_0288_),
    .Y(_0293_));
 sg13g2_a21oi_1 _3100_ (.A1(net812),
    .A2(_2171_),
    .Y(_0294_),
    .B1(net900));
 sg13g2_o21ai_1 _3101_ (.B1(_0294_),
    .Y(_0295_),
    .A1(net797),
    .A2(_2091_));
 sg13g2_o21ai_1 _3102_ (.B1(net801),
    .Y(_0296_),
    .A1(net797),
    .A2(_2087_));
 sg13g2_nand3_1 _3103_ (.B(_0226_),
    .C(_0296_),
    .A(_0194_),
    .Y(_0297_));
 sg13g2_nand2_1 _3104_ (.Y(_0298_),
    .A(net907),
    .B(_0297_));
 sg13g2_o21ai_1 _3105_ (.B1(net918),
    .Y(_0299_),
    .A1(_2184_),
    .A2(_0201_));
 sg13g2_nand4_1 _3106_ (.B(_0295_),
    .C(_0298_),
    .A(_0288_),
    .Y(_0300_),
    .D(_0299_));
 sg13g2_nor2_1 _3107_ (.A(net935),
    .B(net793),
    .Y(_0301_));
 sg13g2_a22oi_1 _3108_ (.Y(_0302_),
    .B1(_0300_),
    .B2(_0301_),
    .A2(_0293_),
    .A1(_1874_));
 sg13g2_nor2_1 _3109_ (.A(net914),
    .B(_1729_),
    .Y(_0303_));
 sg13g2_a21oi_1 _3110_ (.A1(_1825_),
    .A2(_0205_),
    .Y(_0304_),
    .B1(_1854_));
 sg13g2_nand3_1 _3111_ (.B(_1678_),
    .C(_0210_),
    .A(net789),
    .Y(_0305_));
 sg13g2_a221oi_1 _3112_ (.B2(net904),
    .C1(_0304_),
    .B1(_0305_),
    .A1(net932),
    .Y(_0306_),
    .A2(_0214_));
 sg13g2_a21oi_1 _3113_ (.A1(net918),
    .A2(_0258_),
    .Y(_0307_),
    .B1(net916));
 sg13g2_a22oi_1 _3114_ (.Y(_0308_),
    .B1(_0306_),
    .B2(_0307_),
    .A2(_0303_),
    .A1(_0302_));
 sg13g2_nor2b_1 _3115_ (.A(_0308_),
    .B_N(_1951_),
    .Y(_0309_));
 sg13g2_or2_1 _3116_ (.X(_0310_),
    .B(_0271_),
    .A(net951));
 sg13g2_a21oi_1 _3117_ (.A1(net956),
    .A2(_1686_),
    .Y(_0311_),
    .B1(net935));
 sg13g2_a21o_1 _3118_ (.A2(_1899_),
    .A1(_1748_),
    .B1(net816),
    .X(_0312_));
 sg13g2_a221oi_1 _3119_ (.B2(net816),
    .C1(_1875_),
    .B1(_0270_),
    .A1(net956),
    .Y(_0313_),
    .A2(_2082_));
 sg13g2_a221oi_1 _3120_ (.B2(_0313_),
    .C1(net887),
    .B1(_0312_),
    .A1(_0310_),
    .Y(_0314_),
    .A2(_0311_));
 sg13g2_a221oi_1 _3121_ (.B2(net932),
    .C1(_2106_),
    .B1(_0273_),
    .A1(net917),
    .Y(_0315_),
    .A2(_0230_));
 sg13g2_nand2b_1 _3122_ (.Y(_0316_),
    .B(_0315_),
    .A_N(_0314_));
 sg13g2_a22oi_1 _3123_ (.Y(_0317_),
    .B1(_0263_),
    .B2(net931),
    .A2(_0236_),
    .A1(net919));
 sg13g2_o21ai_1 _3124_ (.B1(net903),
    .Y(_0318_),
    .A1(_1827_),
    .A2(_0255_));
 sg13g2_nand2_1 _3125_ (.Y(_0319_),
    .A(net909),
    .B(_0253_));
 sg13g2_and3_1 _3126_ (.X(_0320_),
    .A(_0317_),
    .B(_0318_),
    .C(_0319_));
 sg13g2_nand3_1 _3127_ (.B(_1755_),
    .C(_0237_),
    .A(net909),
    .Y(_0321_));
 sg13g2_a21oi_1 _3128_ (.A1(_0264_),
    .A2(_0321_),
    .Y(_0322_),
    .B1(net881));
 sg13g2_o21ai_1 _3129_ (.B1(_0322_),
    .Y(_0323_),
    .A1(net914),
    .A2(_0320_));
 sg13g2_nand2_1 _3130_ (.Y(_0324_),
    .A(_0316_),
    .B(_0323_));
 sg13g2_o21ai_1 _3131_ (.B1(\nyanframe[1] ),
    .Y(_0325_),
    .A1(_0309_),
    .A2(_0324_));
 sg13g2_o21ai_1 _3132_ (.B1(net823),
    .Y(_0326_),
    .A1(_1640_),
    .A2(net797));
 sg13g2_nand3_1 _3133_ (.B(_1801_),
    .C(_0326_),
    .A(net954),
    .Y(_0327_));
 sg13g2_a21oi_1 _3134_ (.A1(_1761_),
    .A2(net797),
    .Y(_0328_),
    .B1(_2079_));
 sg13g2_nor2_1 _3135_ (.A(net954),
    .B(_0287_),
    .Y(_0329_));
 sg13g2_o21ai_1 _3136_ (.B1(_0329_),
    .Y(_0330_),
    .A1(net802),
    .A2(_0328_));
 sg13g2_nand3_1 _3137_ (.B(_0327_),
    .C(_0330_),
    .A(net890),
    .Y(_0331_));
 sg13g2_o21ai_1 _3138_ (.B1(net918),
    .Y(_0332_),
    .A1(_0196_),
    .A2(_0247_));
 sg13g2_nor3_1 _3139_ (.A(net823),
    .B(_1701_),
    .C(_2170_),
    .Y(_0333_));
 sg13g2_a21oi_1 _3140_ (.A1(_1673_),
    .A2(_1704_),
    .Y(_0334_),
    .B1(_1624_));
 sg13g2_nor3_1 _3141_ (.A(net911),
    .B(_0333_),
    .C(_0334_),
    .Y(_0335_));
 sg13g2_nor3_1 _3142_ (.A(net793),
    .B(_1920_),
    .C(_0335_),
    .Y(_0336_));
 sg13g2_nand3_1 _3143_ (.B(_0332_),
    .C(_0336_),
    .A(_0331_),
    .Y(_0337_));
 sg13g2_nor2_1 _3144_ (.A(net949),
    .B(_2178_),
    .Y(_0338_));
 sg13g2_and2_1 _3145_ (.A(net949),
    .B(_2183_),
    .X(_0339_));
 sg13g2_a22oi_1 _3146_ (.Y(_0340_),
    .B1(_0339_),
    .B2(_2176_),
    .A2(_0338_),
    .A1(_2165_));
 sg13g2_mux2_1 _3147_ (.A0(_1695_),
    .A1(_2172_),
    .S(_1624_),
    .X(_0341_));
 sg13g2_a22oi_1 _3148_ (.Y(_0342_),
    .B1(_0341_),
    .B2(net907),
    .A2(_0280_),
    .A1(_1758_));
 sg13g2_o21ai_1 _3149_ (.B1(_0342_),
    .Y(_0343_),
    .A1(net940),
    .A2(_0340_));
 sg13g2_nand4_1 _3150_ (.B(_1680_),
    .C(_0194_),
    .A(net940),
    .Y(_0344_),
    .D(_0195_));
 sg13g2_o21ai_1 _3151_ (.B1(net911),
    .Y(_0345_),
    .A1(net934),
    .A2(_0249_));
 sg13g2_nand2b_1 _3152_ (.Y(_0346_),
    .B(_1704_),
    .A_N(_0188_));
 sg13g2_nand3_1 _3153_ (.B(_1676_),
    .C(_1811_),
    .A(net803),
    .Y(_0347_));
 sg13g2_nand3_1 _3154_ (.B(_0191_),
    .C(_0347_),
    .A(net954),
    .Y(_0348_));
 sg13g2_a21oi_1 _3155_ (.A1(_1921_),
    .A2(_0346_),
    .Y(_0349_),
    .B1(net888));
 sg13g2_a221oi_1 _3156_ (.B2(_0349_),
    .C1(_1580_),
    .B1(_0348_),
    .A1(_0344_),
    .Y(_0350_),
    .A2(_0345_));
 sg13g2_o21ai_1 _3157_ (.B1(_1674_),
    .Y(_0351_),
    .A1(net880),
    .A2(_1652_));
 sg13g2_a21o_1 _3158_ (.A2(_0351_),
    .A1(_0186_),
    .B1(_1528_),
    .X(_0352_));
 sg13g2_nand2_1 _3159_ (.Y(_0353_),
    .A(net907),
    .B(_2166_));
 sg13g2_a221oi_1 _3160_ (.B2(net904),
    .C1(_1747_),
    .B1(_2179_),
    .A1(net932),
    .Y(_0354_),
    .A2(_2177_));
 sg13g2_and2_1 _3161_ (.A(_0353_),
    .B(_0354_),
    .X(_0355_));
 sg13g2_a221oi_1 _3162_ (.B2(_0355_),
    .C1(_0350_),
    .B1(_0352_),
    .A1(_1808_),
    .Y(_0356_),
    .A2(_0343_));
 sg13g2_o21ai_1 _3163_ (.B1(_0337_),
    .Y(_0357_),
    .A1(net792),
    .A2(_0356_));
 sg13g2_nand3_1 _3164_ (.B(_2027_),
    .C(_2068_),
    .A(net816),
    .Y(_0358_));
 sg13g2_a21oi_1 _3165_ (.A1(net805),
    .A2(_0276_),
    .Y(_0359_),
    .B1(net906));
 sg13g2_a21oi_1 _3166_ (.A1(_0358_),
    .A2(_0359_),
    .Y(_0360_),
    .B1(_2106_));
 sg13g2_nand2b_1 _3167_ (.Y(_0361_),
    .B(net788),
    .A_N(_0281_));
 sg13g2_a21oi_1 _3168_ (.A1(net949),
    .A2(net788),
    .Y(_0362_),
    .B1(net953));
 sg13g2_a21oi_1 _3169_ (.A1(net787),
    .A2(_1798_),
    .Y(_0363_),
    .B1(net900));
 sg13g2_a22oi_1 _3170_ (.Y(_0364_),
    .B1(_1889_),
    .B2(net805),
    .A2(_1699_),
    .A1(net833));
 sg13g2_a21oi_1 _3171_ (.A1(_0210_),
    .A2(_0364_),
    .Y(_0365_),
    .B1(net934));
 sg13g2_a21oi_1 _3172_ (.A1(_1834_),
    .A2(_2000_),
    .Y(_0366_),
    .B1(net901));
 sg13g2_a22oi_1 _3173_ (.Y(_0367_),
    .B1(net784),
    .B2(_2078_),
    .A2(net912),
    .A1(net790));
 sg13g2_nor3_1 _3174_ (.A(_0365_),
    .B(_0366_),
    .C(_0367_),
    .Y(_0368_));
 sg13g2_nor2_1 _3175_ (.A(net936),
    .B(_0368_),
    .Y(_0369_));
 sg13g2_a221oi_1 _3176_ (.B2(_0362_),
    .C1(_0363_),
    .B1(_0361_),
    .A1(net917),
    .Y(_0370_),
    .A2(_2173_));
 sg13g2_o21ai_1 _3177_ (.B1(_0360_),
    .Y(_0371_),
    .A1(net966),
    .A2(_0370_));
 sg13g2_o21ai_1 _3178_ (.B1(\nyanframe[2] ),
    .Y(_0372_),
    .A1(_0369_),
    .A2(_0371_));
 sg13g2_nor2_1 _3179_ (.A(net901),
    .B(_0240_),
    .Y(_0373_));
 sg13g2_o21ai_1 _3180_ (.B1(_0317_),
    .Y(_0374_),
    .A1(net905),
    .A2(_0243_));
 sg13g2_o21ai_1 _3181_ (.B1(_1746_),
    .Y(_0375_),
    .A1(_0373_),
    .A2(_0374_));
 sg13g2_nand3_1 _3182_ (.B(net813),
    .C(_0248_),
    .A(net949),
    .Y(_0376_));
 sg13g2_a221oi_1 _3183_ (.B2(_1675_),
    .C1(_2170_),
    .B1(_1980_),
    .A1(net879),
    .Y(_0377_),
    .A2(_1762_));
 sg13g2_nand3b_1 _3184_ (.B(net811),
    .C(net954),
    .Y(_0378_),
    .A_N(_0377_));
 sg13g2_nand3_1 _3185_ (.B(_0376_),
    .C(_0378_),
    .A(_1825_),
    .Y(_0379_));
 sg13g2_and4_1 _3186_ (.A(net817),
    .B(_1659_),
    .C(net932),
    .D(_1715_),
    .X(_0380_));
 sg13g2_a21oi_2 _3187_ (.B1(_0380_),
    .Y(_0381_),
    .A2(_0379_),
    .A1(net890));
 sg13g2_a21oi_1 _3188_ (.A1(_0317_),
    .A2(_0381_),
    .Y(_0382_),
    .B1(_1809_));
 sg13g2_nor2b_1 _3189_ (.A(_0382_),
    .B_N(_0322_),
    .Y(_0383_));
 sg13g2_a221oi_1 _3190_ (.B2(_0383_),
    .C1(_0372_),
    .B1(_0375_),
    .A1(_1951_),
    .Y(_0384_),
    .A2(_0357_));
 sg13g2_or2_1 _3191_ (.X(_0385_),
    .B(_0384_),
    .A(_1978_));
 sg13g2_a21oi_2 _3192_ (.B1(_0385_),
    .Y(_0386_),
    .A2(_0325_),
    .A1(_0286_));
 sg13g2_a21o_1 _3193_ (.A2(_0325_),
    .A1(_0286_),
    .B1(_0385_),
    .X(_0387_));
 sg13g2_nor2_1 _3194_ (.A(net776),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_and2_1 _3195_ (.A(net777),
    .B(_0386_),
    .X(_0389_));
 sg13g2_nor2_1 _3196_ (.A(net776),
    .B(_0386_),
    .Y(_0390_));
 sg13g2_o21ai_1 _3197_ (.B1(net881),
    .Y(_0391_),
    .A1(net890),
    .A2(_1863_));
 sg13g2_nand3_1 _3198_ (.B(\hvsync_gen.hpos[2] ),
    .C(net971),
    .A(\hvsync_gen.hpos[3] ),
    .Y(_0392_));
 sg13g2_nor2_1 _3199_ (.A(net970),
    .B(net969),
    .Y(_0393_));
 sg13g2_nand2_1 _3200_ (.Y(_0394_),
    .A(net972),
    .B(net971));
 sg13g2_nand3_1 _3201_ (.B(_0393_),
    .C(_0394_),
    .A(_0392_),
    .Y(_0395_));
 sg13g2_a21oi_2 _3202_ (.B1(\hvsync_gen.hpos[9] ),
    .Y(_0396_),
    .A2(_0395_),
    .A1(net968));
 sg13g2_nand3_1 _3203_ (.B(_0391_),
    .C(_0396_),
    .A(_1976_),
    .Y(_0397_));
 sg13g2_nor4_1 _3204_ (.A(net777),
    .B(net776),
    .C(_0386_),
    .D(_0397_),
    .Y(_0398_));
 sg13g2_nand2_1 _3205_ (.Y(_0399_),
    .A(\hvsync_gen.hpos[5] ),
    .B(\frame_count[3] ));
 sg13g2_xnor2_1 _3206_ (.Y(_0400_),
    .A(\hvsync_gen.hpos[5] ),
    .B(\frame_count[3] ));
 sg13g2_and2_1 _3207_ (.A(net973),
    .B(\frame_count[2] ),
    .X(_0401_));
 sg13g2_nand2_1 _3208_ (.Y(_0402_),
    .A(\hvsync_gen.hpos[3] ),
    .B(\frame_count[1] ));
 sg13g2_xnor2_1 _3209_ (.Y(_0403_),
    .A(\hvsync_gen.hpos[3] ),
    .B(\frame_count[1] ));
 sg13g2_nand2_1 _3210_ (.Y(_0404_),
    .A(\frame_count[0] ),
    .B(\hvsync_gen.hpos[2] ));
 sg13g2_o21ai_1 _3211_ (.B1(_0402_),
    .Y(_0405_),
    .A1(_0403_),
    .A2(_0404_));
 sg13g2_xor2_1 _3212_ (.B(\frame_count[2] ),
    .A(net973),
    .X(_0406_));
 sg13g2_a21oi_1 _3213_ (.A1(_0405_),
    .A2(_0406_),
    .Y(_0407_),
    .B1(_0401_));
 sg13g2_o21ai_1 _3214_ (.B1(_0399_),
    .Y(_0408_),
    .A1(_0400_),
    .A2(_0407_));
 sg13g2_and2_1 _3215_ (.A(\hvsync_gen.hpos[6] ),
    .B(\frame_count[4] ),
    .X(_0409_));
 sg13g2_xor2_1 _3216_ (.B(\frame_count[4] ),
    .A(net970),
    .X(_0410_));
 sg13g2_xnor2_1 _3217_ (.Y(_0411_),
    .A(_0408_),
    .B(_0410_));
 sg13g2_and2_1 _3218_ (.A(net941),
    .B(_0411_),
    .X(_0412_));
 sg13g2_a21o_1 _3219_ (.A2(_0411_),
    .A1(_1666_),
    .B1(_1528_),
    .X(_0413_));
 sg13g2_nand2_1 _3220_ (.Y(_0414_),
    .A(_1781_),
    .B(_0412_));
 sg13g2_and2_1 _3221_ (.A(_0413_),
    .B(_0414_),
    .X(_0415_));
 sg13g2_xnor2_1 _3222_ (.Y(_0416_),
    .A(net944),
    .B(_0413_));
 sg13g2_xnor2_1 _3223_ (.Y(_0417_),
    .A(_0036_),
    .B(_0412_));
 sg13g2_inv_1 _3224_ (.Y(_0418_),
    .A(_0417_));
 sg13g2_nand2b_1 _3225_ (.Y(_0419_),
    .B(_0418_),
    .A_N(_0415_));
 sg13g2_or2_1 _3226_ (.X(_0420_),
    .B(_0419_),
    .A(_0416_));
 sg13g2_xor2_1 _3227_ (.B(\hvsync_gen.hpos[0] ),
    .A(\frame_count[0] ),
    .X(_0421_));
 sg13g2_inv_1 _3228_ (.Y(_0422_),
    .A(_0421_));
 sg13g2_xor2_1 _3229_ (.B(\frame_count[0] ),
    .A(\hvsync_gen.vpos[0] ),
    .X(_0423_));
 sg13g2_nor2_1 _3230_ (.A(_0421_),
    .B(_0423_),
    .Y(_0424_));
 sg13g2_xnor2_1 _3231_ (.Y(_0425_),
    .A(\hvsync_gen.vpos[0] ),
    .B(\hvsync_gen.hpos[0] ));
 sg13g2_nor2_1 _3232_ (.A(_0420_),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_a22oi_1 _3233_ (.Y(_0427_),
    .B1(net773),
    .B2(_0426_),
    .A2(_0388_),
    .A1(net777));
 sg13g2_nand2b_1 _3234_ (.Y(_0428_),
    .B(net948),
    .A_N(net995));
 sg13g2_xor2_1 _3235_ (.B(net995),
    .A(net948),
    .X(_0429_));
 sg13g2_nand2_1 _3236_ (.Y(_0430_),
    .A(net951),
    .B(net1000));
 sg13g2_xor2_1 _3237_ (.B(net1000),
    .A(net951),
    .X(_0431_));
 sg13g2_nand3_1 _3238_ (.B(net1005),
    .C(_0431_),
    .A(net960),
    .Y(_0432_));
 sg13g2_nand3_1 _3239_ (.B(_0430_),
    .C(_0432_),
    .A(_0429_),
    .Y(_0433_));
 sg13g2_a21o_1 _3240_ (.A2(_0432_),
    .A1(_0430_),
    .B1(_0429_),
    .X(_0434_));
 sg13g2_nand2_1 _3241_ (.Y(_0435_),
    .A(net976),
    .B(\songpos[6] ));
 sg13g2_o21ai_1 _3242_ (.B1(_1537_),
    .Y(_0436_),
    .A1(_1535_),
    .A2(_0435_));
 sg13g2_inv_1 _3243_ (.Y(_0437_),
    .A(_0436_));
 sg13g2_and2_1 _3244_ (.A(net961),
    .B(_0436_),
    .X(_0438_));
 sg13g2_nand2_2 _3245_ (.Y(_0439_),
    .A(net961),
    .B(_0436_));
 sg13g2_nor2b_2 _3246_ (.A(\nyanframe[1] ),
    .B_N(net261),
    .Y(_0440_));
 sg13g2_nand2_2 _3247_ (.Y(_0441_),
    .A(net952),
    .B(_0440_));
 sg13g2_inv_1 _3248_ (.Y(_0442_),
    .A(_0441_));
 sg13g2_xnor2_1 _3249_ (.Y(_0443_),
    .A(_1529_),
    .B(_0441_));
 sg13g2_nor2b_1 _3250_ (.A(net951),
    .B_N(net1000),
    .Y(_0444_));
 sg13g2_nor2_1 _3251_ (.A(_0429_),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_nand2_1 _3252_ (.Y(_0446_),
    .A(_0429_),
    .B(_0444_));
 sg13g2_nand2b_1 _3253_ (.Y(_0447_),
    .B(_0446_),
    .A_N(_0445_));
 sg13g2_nand2b_1 _3254_ (.Y(_0448_),
    .B(net1005),
    .A_N(net960));
 sg13g2_nor2_1 _3255_ (.A(_0431_),
    .B(_0448_),
    .Y(_0449_));
 sg13g2_xnor2_1 _3256_ (.Y(_0450_),
    .A(net960),
    .B(net1004));
 sg13g2_xor2_1 _3257_ (.B(_0450_),
    .A(\hvsync_gen.vpos[1] ),
    .X(_0451_));
 sg13g2_or2_1 _3258_ (.X(_0452_),
    .B(_0451_),
    .A(_1542_));
 sg13g2_nor2_1 _3259_ (.A(_0032_),
    .B(_0450_),
    .Y(_0453_));
 sg13g2_a21oi_1 _3260_ (.A1(_0431_),
    .A2(_0448_),
    .Y(_0454_),
    .B1(_0453_));
 sg13g2_a21oi_2 _3261_ (.B1(_0449_),
    .Y(_0455_),
    .A2(_0454_),
    .A1(_0452_));
 sg13g2_xnor2_1 _3262_ (.Y(_0456_),
    .A(_0447_),
    .B(_0455_));
 sg13g2_a22oi_1 _3263_ (.Y(_0457_),
    .B1(_0456_),
    .B2(_0436_),
    .A2(_0443_),
    .A1(net961));
 sg13g2_a21oi_1 _3264_ (.A1(_0433_),
    .A2(_0434_),
    .Y(_0458_),
    .B1(_0439_));
 sg13g2_a21o_1 _3265_ (.A2(_0457_),
    .A1(_0439_),
    .B1(_0458_),
    .X(_0459_));
 sg13g2_a21o_1 _3266_ (.A2(net1004),
    .A1(net960),
    .B1(_0431_),
    .X(_0460_));
 sg13g2_nand3_1 _3267_ (.B(_0436_),
    .C(_0460_),
    .A(_0432_),
    .Y(_0461_));
 sg13g2_nor2_1 _3268_ (.A(net951),
    .B(_0440_),
    .Y(_0462_));
 sg13g2_o21ai_1 _3269_ (.B1(net961),
    .Y(_0463_),
    .A1(_0442_),
    .A2(_0462_));
 sg13g2_nand2_1 _3270_ (.Y(_0464_),
    .A(_0439_),
    .B(_0463_));
 sg13g2_nor2b_1 _3271_ (.A(net1004),
    .B_N(net960),
    .Y(_0465_));
 sg13g2_xnor2_1 _3272_ (.Y(_0466_),
    .A(_0431_),
    .B(_0465_));
 sg13g2_a21oi_1 _3273_ (.A1(_0436_),
    .A2(_0466_),
    .Y(_0467_),
    .B1(net961));
 sg13g2_a21oi_2 _3274_ (.B1(_0467_),
    .Y(_0468_),
    .A2(_0464_),
    .A1(_0461_));
 sg13g2_inv_1 _3275_ (.Y(_0469_),
    .A(_0468_));
 sg13g2_xor2_1 _3276_ (.B(_1591_),
    .A(_1589_),
    .X(_0470_));
 sg13g2_nor2_1 _3277_ (.A(net880),
    .B(net886),
    .Y(_0471_));
 sg13g2_nor2_1 _3278_ (.A(net869),
    .B(net885),
    .Y(_0472_));
 sg13g2_nand2b_1 _3279_ (.Y(_0473_),
    .B(net843),
    .A_N(_0472_));
 sg13g2_xnor2_1 _3280_ (.Y(_0474_),
    .A(net880),
    .B(net886));
 sg13g2_nand2_1 _3281_ (.Y(_0475_),
    .A(net964),
    .B(_0440_));
 sg13g2_nand3_1 _3282_ (.B(_2112_),
    .C(_0475_),
    .A(song_loops),
    .Y(_0476_));
 sg13g2_nor2b_2 _3283_ (.A(_0476_),
    .B_N(_0474_),
    .Y(_0477_));
 sg13g2_xnor2_1 _3284_ (.Y(_0478_),
    .A(net872),
    .B(_0471_));
 sg13g2_nand2b_2 _3285_ (.Y(_0479_),
    .B(_0477_),
    .A_N(_0478_));
 sg13g2_xnor2_1 _3286_ (.Y(_0480_),
    .A(net837),
    .B(_0472_));
 sg13g2_nor2_1 _3287_ (.A(_0479_),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_o21ai_1 _3288_ (.B1(_0473_),
    .Y(_0482_),
    .A1(_0479_),
    .A2(_0480_));
 sg13g2_xnor2_1 _3289_ (.Y(_0483_),
    .A(net861),
    .B(_0482_));
 sg13g2_xnor2_1 _3290_ (.Y(_0484_),
    .A(net852),
    .B(_0482_));
 sg13g2_xor2_1 _3291_ (.B(_0480_),
    .A(_0479_),
    .X(_0485_));
 sg13g2_xnor2_1 _3292_ (.Y(_0486_),
    .A(_0479_),
    .B(_0480_));
 sg13g2_xnor2_1 _3293_ (.Y(_0487_),
    .A(_0477_),
    .B(_0478_));
 sg13g2_xor2_1 _3294_ (.B(_0476_),
    .A(_0474_),
    .X(_0488_));
 sg13g2_nor2_1 _3295_ (.A(_0485_),
    .B(net796),
    .Y(_0489_));
 sg13g2_and2_1 _3296_ (.A(_0488_),
    .B(_0489_),
    .X(_0490_));
 sg13g2_nand2_1 _3297_ (.Y(_0491_),
    .A(net885),
    .B(net796));
 sg13g2_nor2_1 _3298_ (.A(net837),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_xor2_1 _3299_ (.B(_0488_),
    .A(net796),
    .X(_0493_));
 sg13g2_o21ai_1 _3300_ (.B1(_0484_),
    .Y(_0494_),
    .A1(_0486_),
    .A2(_0493_));
 sg13g2_nor3_1 _3301_ (.A(_0490_),
    .B(_0492_),
    .C(_0494_),
    .Y(_0495_));
 sg13g2_nor2_1 _3302_ (.A(net885),
    .B(_0487_),
    .Y(_0496_));
 sg13g2_a21oi_1 _3303_ (.A1(_0487_),
    .A2(_0488_),
    .Y(_0497_),
    .B1(_0496_));
 sg13g2_a21oi_1 _3304_ (.A1(_1542_),
    .A2(_0451_),
    .Y(_0498_),
    .B1(_0437_));
 sg13g2_nand2_1 _3305_ (.Y(_0499_),
    .A(_0030_),
    .B(_0437_));
 sg13g2_a22oi_1 _3306_ (.Y(_0500_),
    .B1(_0499_),
    .B2(net961),
    .A2(_0498_),
    .A1(_0452_));
 sg13g2_a21o_2 _3307_ (.A2(_0450_),
    .A1(_0438_),
    .B1(_0500_),
    .X(_0501_));
 sg13g2_inv_1 _3308_ (.Y(_0502_),
    .A(_0501_));
 sg13g2_nor3_1 _3309_ (.A(_0486_),
    .B(_0488_),
    .C(_0491_),
    .Y(_0503_));
 sg13g2_nand2_1 _3310_ (.Y(_0504_),
    .A(net886),
    .B(_0486_));
 sg13g2_nor2_1 _3311_ (.A(_0493_),
    .B(_0504_),
    .Y(_0505_));
 sg13g2_o21ai_1 _3312_ (.B1(_0484_),
    .Y(_0506_),
    .A1(_0503_),
    .A2(_0505_));
 sg13g2_nand2_1 _3313_ (.Y(_0507_),
    .A(net885),
    .B(_0488_));
 sg13g2_or2_1 _3314_ (.X(_0508_),
    .B(_0507_),
    .A(net796));
 sg13g2_o21ai_1 _3315_ (.B1(_0506_),
    .Y(_0509_),
    .A1(_0484_),
    .A2(_0508_));
 sg13g2_o21ai_1 _3316_ (.B1(_0468_),
    .Y(_0510_),
    .A1(_0484_),
    .A2(_0497_));
 sg13g2_nor2_1 _3317_ (.A(_0495_),
    .B(_0510_),
    .Y(_0511_));
 sg13g2_a21oi_1 _3318_ (.A1(_0469_),
    .A2(_0509_),
    .Y(_0512_),
    .B1(_0511_));
 sg13g2_nand2_1 _3319_ (.Y(_0513_),
    .A(_0468_),
    .B(_0501_));
 sg13g2_nor2_1 _3320_ (.A(net885),
    .B(_0484_),
    .Y(_0514_));
 sg13g2_nand2_1 _3321_ (.Y(_0515_),
    .A(_0493_),
    .B(_0514_));
 sg13g2_nor2_1 _3322_ (.A(net885),
    .B(_0488_),
    .Y(_0516_));
 sg13g2_nor3_1 _3323_ (.A(_0485_),
    .B(net796),
    .C(_0516_),
    .Y(_0517_));
 sg13g2_nand2_1 _3324_ (.Y(_0518_),
    .A(_0507_),
    .B(_0517_));
 sg13g2_nand3_1 _3325_ (.B(net796),
    .C(_0488_),
    .A(net885),
    .Y(_0519_));
 sg13g2_nand3b_1 _3326_ (.B(_0519_),
    .C(_0485_),
    .Y(_0520_),
    .A_N(_0516_));
 sg13g2_o21ai_1 _3327_ (.B1(_0491_),
    .Y(_0521_),
    .A1(_0478_),
    .A2(_0488_));
 sg13g2_a21oi_1 _3328_ (.A1(_0486_),
    .A2(_0521_),
    .Y(_0522_),
    .B1(_0483_));
 sg13g2_nand3_1 _3329_ (.B(_0520_),
    .C(_0522_),
    .A(_0518_),
    .Y(_0523_));
 sg13g2_a21o_1 _3330_ (.A2(_0523_),
    .A1(_0515_),
    .B1(_0513_),
    .X(_0524_));
 sg13g2_o21ai_1 _3331_ (.B1(_0524_),
    .Y(_0525_),
    .A1(_0501_),
    .A2(_0512_));
 sg13g2_nand2_1 _3332_ (.Y(_0526_),
    .A(_0483_),
    .B(_0485_));
 sg13g2_nor2_1 _3333_ (.A(\hvsync_gen.vpos[8] ),
    .B(net977),
    .Y(_0527_));
 sg13g2_xnor2_1 _3334_ (.Y(_0528_),
    .A(\hvsync_gen.vpos[8] ),
    .B(net977));
 sg13g2_nand2_1 _3335_ (.Y(_0529_),
    .A(_1530_),
    .B(_1535_));
 sg13g2_and2_1 _3336_ (.A(_0528_),
    .B(_0529_),
    .X(_0530_));
 sg13g2_nand2_1 _3337_ (.Y(_0531_),
    .A(net945),
    .B(net985));
 sg13g2_xnor2_1 _3338_ (.Y(_0532_),
    .A(net943),
    .B(net979));
 sg13g2_nand2b_1 _3339_ (.Y(_0533_),
    .B(_0532_),
    .A_N(_0531_));
 sg13g2_xnor2_1 _3340_ (.Y(_0534_),
    .A(_0531_),
    .B(_0532_));
 sg13g2_nand2_1 _3341_ (.Y(_0535_),
    .A(net946),
    .B(net990));
 sg13g2_xnor2_1 _3342_ (.Y(_0536_),
    .A(net945),
    .B(net985));
 sg13g2_nor2_1 _3343_ (.A(_0535_),
    .B(_0536_),
    .Y(_0537_));
 sg13g2_xor2_1 _3344_ (.B(net990),
    .A(net946),
    .X(_0538_));
 sg13g2_or2_1 _3345_ (.X(_0539_),
    .B(net995),
    .A(net948));
 sg13g2_xnor2_1 _3346_ (.Y(_0540_),
    .A(_0538_),
    .B(_0539_));
 sg13g2_nor2_1 _3347_ (.A(_0434_),
    .B(_0540_),
    .Y(_0541_));
 sg13g2_a21oi_1 _3348_ (.A1(_0538_),
    .A2(_0539_),
    .Y(_0542_),
    .B1(_0541_));
 sg13g2_xnor2_1 _3349_ (.Y(_0543_),
    .A(_0535_),
    .B(_0536_));
 sg13g2_nor2_1 _3350_ (.A(_0542_),
    .B(_0543_),
    .Y(_0544_));
 sg13g2_o21ai_1 _3351_ (.B1(_0534_),
    .Y(_0545_),
    .A1(_0537_),
    .A2(_0544_));
 sg13g2_nand2_1 _3352_ (.Y(_0546_),
    .A(_0533_),
    .B(_0545_));
 sg13g2_nor2_1 _3353_ (.A(_0530_),
    .B(_0546_),
    .Y(_0547_));
 sg13g2_nor2_1 _3354_ (.A(_0528_),
    .B(_0529_),
    .Y(_0548_));
 sg13g2_o21ai_1 _3355_ (.B1(_0546_),
    .Y(_0549_),
    .A1(_0530_),
    .A2(_0548_));
 sg13g2_xor2_1 _3356_ (.B(net976),
    .A(net942),
    .X(_0550_));
 sg13g2_xor2_1 _3357_ (.B(_0550_),
    .A(_0527_),
    .X(_0551_));
 sg13g2_a21oi_1 _3358_ (.A1(_0549_),
    .A2(_0551_),
    .Y(_0552_),
    .B1(_0547_));
 sg13g2_or3_1 _3359_ (.A(_0534_),
    .B(_0537_),
    .C(_0544_),
    .X(_0553_));
 sg13g2_nand2_1 _3360_ (.Y(_0554_),
    .A(_0545_),
    .B(_0553_));
 sg13g2_xnor2_1 _3361_ (.Y(_0555_),
    .A(_0542_),
    .B(_0543_));
 sg13g2_nand2_1 _3362_ (.Y(_0556_),
    .A(_0434_),
    .B(_0540_));
 sg13g2_nand3b_1 _3363_ (.B(_0556_),
    .C(song_loops),
    .Y(_0557_),
    .A_N(_0541_));
 sg13g2_a21o_1 _3364_ (.A2(_0441_),
    .A1(_0036_),
    .B1(_0035_),
    .X(_0558_));
 sg13g2_nand3_1 _3365_ (.B(_0035_),
    .C(_0441_),
    .A(_0036_),
    .Y(_0559_));
 sg13g2_nand3_1 _3366_ (.B(_0558_),
    .C(_0559_),
    .A(song_loops),
    .Y(_0560_));
 sg13g2_o21ai_1 _3367_ (.B1(net946),
    .Y(_0561_),
    .A1(net950),
    .A2(_0442_));
 sg13g2_nor2_1 _3368_ (.A(net943),
    .B(net944),
    .Y(_0562_));
 sg13g2_nand2b_1 _3369_ (.Y(_0563_),
    .B(_0562_),
    .A_N(_1973_));
 sg13g2_nand2_1 _3370_ (.Y(_0564_),
    .A(net943),
    .B(net944));
 sg13g2_nor3_1 _3371_ (.A(\hvsync_gen.vpos[8] ),
    .B(\hvsync_gen.vpos[9] ),
    .C(_0564_),
    .Y(_0565_));
 sg13g2_o21ai_1 _3372_ (.B1(_0439_),
    .Y(_0566_),
    .A1(_0561_),
    .A2(_0565_));
 sg13g2_a21oi_1 _3373_ (.A1(_0561_),
    .A2(_0563_),
    .Y(_0567_),
    .B1(_0566_));
 sg13g2_a22oi_1 _3374_ (.Y(_0568_),
    .B1(_0560_),
    .B2(_0567_),
    .A2(_0557_),
    .A1(_0436_));
 sg13g2_nand2_1 _3375_ (.Y(_0569_),
    .A(_0469_),
    .B(_0501_));
 sg13g2_a21oi_1 _3376_ (.A1(_0469_),
    .A2(_0501_),
    .Y(_0570_),
    .B1(_0459_));
 sg13g2_nor2_1 _3377_ (.A(net943),
    .B(_1535_),
    .Y(_0571_));
 sg13g2_xnor2_1 _3378_ (.Y(_0572_),
    .A(_0528_),
    .B(_0571_));
 sg13g2_nor2_1 _3379_ (.A(_0428_),
    .B(_0538_),
    .Y(_0573_));
 sg13g2_xnor2_1 _3380_ (.Y(_0574_),
    .A(_0428_),
    .B(_0538_));
 sg13g2_a21oi_2 _3381_ (.B1(_0445_),
    .Y(_0575_),
    .A2(_0455_),
    .A1(_0446_));
 sg13g2_nor2_1 _3382_ (.A(_0574_),
    .B(_0575_),
    .Y(_0576_));
 sg13g2_nor2_1 _3383_ (.A(_0573_),
    .B(_0576_),
    .Y(_0577_));
 sg13g2_nor2_1 _3384_ (.A(_1528_),
    .B(net990),
    .Y(_0578_));
 sg13g2_nor2_1 _3385_ (.A(_0536_),
    .B(_0578_),
    .Y(_0579_));
 sg13g2_o21ai_1 _3386_ (.B1(_0532_),
    .Y(_0580_),
    .A1(_1531_),
    .A2(net985));
 sg13g2_inv_1 _3387_ (.Y(_0581_),
    .A(_0580_));
 sg13g2_nand2_1 _3388_ (.Y(_0582_),
    .A(_0536_),
    .B(_0578_));
 sg13g2_or3_1 _3389_ (.A(_1531_),
    .B(net985),
    .C(_0532_),
    .X(_0583_));
 sg13g2_nand2_1 _3390_ (.Y(_0584_),
    .A(_0582_),
    .B(_0583_));
 sg13g2_nor4_1 _3391_ (.A(_0577_),
    .B(_0579_),
    .C(_0581_),
    .D(_0584_),
    .Y(_0585_));
 sg13g2_o21ai_1 _3392_ (.B1(_0583_),
    .Y(_0586_),
    .A1(_0581_),
    .A2(_0582_));
 sg13g2_o21ai_1 _3393_ (.B1(_0572_),
    .Y(_0587_),
    .A1(_0585_),
    .A2(_0586_));
 sg13g2_mux2_1 _3394_ (.A0(_0572_),
    .A1(_0584_),
    .S(_0580_),
    .X(_0588_));
 sg13g2_a21oi_1 _3395_ (.A1(_0577_),
    .A2(_0588_),
    .Y(_0589_),
    .B1(_0585_));
 sg13g2_xnor2_1 _3396_ (.Y(_0590_),
    .A(_0574_),
    .B(_0575_));
 sg13g2_a21o_1 _3397_ (.A2(_0583_),
    .A1(_0580_),
    .B1(_0579_),
    .X(_0591_));
 sg13g2_nor2b_1 _3398_ (.A(\hvsync_gen.vpos[8] ),
    .B_N(net977),
    .Y(_0592_));
 sg13g2_xnor2_1 _3399_ (.Y(_0593_),
    .A(_0550_),
    .B(_0592_));
 sg13g2_nand4_1 _3400_ (.B(_0590_),
    .C(_0591_),
    .A(_0436_),
    .Y(_0594_),
    .D(_0593_));
 sg13g2_nor2_1 _3401_ (.A(_0589_),
    .B(_0594_),
    .Y(_0595_));
 sg13g2_a21oi_1 _3402_ (.A1(_0587_),
    .A2(_0595_),
    .Y(_0596_),
    .B1(net961));
 sg13g2_nand2_1 _3403_ (.Y(_0597_),
    .A(net852),
    .B(_0473_));
 sg13g2_nor2_1 _3404_ (.A(net821),
    .B(_0597_),
    .Y(_0598_));
 sg13g2_a21oi_1 _3405_ (.A1(_0481_),
    .A2(_0598_),
    .Y(_0599_),
    .B1(_0596_));
 sg13g2_a22oi_1 _3406_ (.Y(_0600_),
    .B1(_0597_),
    .B2(net816),
    .A2(_0481_),
    .A1(net852));
 sg13g2_nand2_1 _3407_ (.Y(_0601_),
    .A(net790),
    .B(_0600_));
 sg13g2_o21ai_1 _3408_ (.B1(net795),
    .Y(_0602_),
    .A1(net816),
    .A2(_0597_));
 sg13g2_a21oi_1 _3409_ (.A1(_0554_),
    .A2(_0555_),
    .Y(_0603_),
    .B1(_0439_));
 sg13g2_nor3_1 _3410_ (.A(_0568_),
    .B(_0570_),
    .C(_0603_),
    .Y(_0604_));
 sg13g2_mux2_1 _3411_ (.A0(_0547_),
    .A1(_0550_),
    .S(_0548_),
    .X(_0605_));
 sg13g2_o21ai_1 _3412_ (.B1(_0438_),
    .Y(_0606_),
    .A1(_0552_),
    .A2(_0605_));
 sg13g2_and4_1 _3413_ (.A(_1971_),
    .B(_0602_),
    .C(_0604_),
    .D(_0606_),
    .X(_0607_));
 sg13g2_and4_1 _3414_ (.A(_0526_),
    .B(_0599_),
    .C(_0601_),
    .D(_0607_),
    .X(_0608_));
 sg13g2_a21oi_1 _3415_ (.A1(net796),
    .A2(_0516_),
    .Y(_0609_),
    .B1(_0486_));
 sg13g2_nand2b_1 _3416_ (.Y(_0610_),
    .B(_0484_),
    .A_N(_0517_));
 sg13g2_a21oi_1 _3417_ (.A1(_0508_),
    .A2(_0609_),
    .Y(_0611_),
    .B1(_0610_));
 sg13g2_a21oi_1 _3418_ (.A1(net796),
    .A2(_0507_),
    .Y(_0612_),
    .B1(_0484_));
 sg13g2_nor3_1 _3419_ (.A(_0459_),
    .B(_0611_),
    .C(_0612_),
    .Y(_0613_));
 sg13g2_nand2b_1 _3420_ (.Y(_0614_),
    .B(_0608_),
    .A_N(_0613_));
 sg13g2_a21oi_2 _3421_ (.B1(_0614_),
    .Y(_0615_),
    .A2(_0525_),
    .A1(_0459_));
 sg13g2_nand2_1 _3422_ (.Y(_0616_),
    .A(_0484_),
    .B(_0492_));
 sg13g2_nand3_1 _3423_ (.B(_0483_),
    .C(_0489_),
    .A(net885),
    .Y(_0617_));
 sg13g2_nand4_1 _3424_ (.B(_0502_),
    .C(_0616_),
    .A(_0468_),
    .Y(_0618_),
    .D(_0617_));
 sg13g2_nand3_1 _3425_ (.B(_0569_),
    .C(_0618_),
    .A(_0459_),
    .Y(_0619_));
 sg13g2_or3_1 _3426_ (.A(_0503_),
    .B(_0505_),
    .C(_0617_),
    .X(_0620_));
 sg13g2_nand3_1 _3427_ (.B(_0506_),
    .C(_0620_),
    .A(_0469_),
    .Y(_0621_));
 sg13g2_nor2_1 _3428_ (.A(_0517_),
    .B(_0609_),
    .Y(_0622_));
 sg13g2_a221oi_1 _3429_ (.B2(_0622_),
    .C1(_0513_),
    .B1(_0522_),
    .A1(_0490_),
    .Y(_0623_),
    .A2(_0514_));
 sg13g2_nand2_1 _3430_ (.Y(_0624_),
    .A(_0608_),
    .B(_0621_));
 sg13g2_nor3_2 _3431_ (.A(_0619_),
    .B(_0623_),
    .C(_0624_),
    .Y(_0625_));
 sg13g2_or2_1 _3432_ (.X(_0626_),
    .B(_0625_),
    .A(_0615_));
 sg13g2_nor3_1 _3433_ (.A(_0424_),
    .B(_0427_),
    .C(_0626_),
    .Y(_0627_));
 sg13g2_nand2_1 _3434_ (.Y(_0628_),
    .A(net968),
    .B(\frame_count[6] ));
 sg13g2_xnor2_1 _3435_ (.Y(_0629_),
    .A(\hvsync_gen.hpos[7] ),
    .B(\frame_count[5] ));
 sg13g2_a21oi_1 _3436_ (.A1(_0408_),
    .A2(_0410_),
    .Y(_0630_),
    .B1(_0409_));
 sg13g2_nor2_1 _3437_ (.A(_0629_),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_a21oi_1 _3438_ (.A1(\hvsync_gen.hpos[7] ),
    .A2(\frame_count[5] ),
    .Y(_0632_),
    .B1(_0631_));
 sg13g2_xnor2_1 _3439_ (.Y(_0633_),
    .A(net968),
    .B(\frame_count[6] ));
 sg13g2_o21ai_1 _3440_ (.B1(_0628_),
    .Y(_0634_),
    .A1(_0632_),
    .A2(_0633_));
 sg13g2_xor2_1 _3441_ (.B(\frame_count[7] ),
    .A(\hvsync_gen.hpos[9] ),
    .X(_0635_));
 sg13g2_xnor2_1 _3442_ (.Y(_0636_),
    .A(_0634_),
    .B(_0635_));
 sg13g2_xnor2_1 _3443_ (.Y(_0637_),
    .A(_0632_),
    .B(_0633_));
 sg13g2_xnor2_1 _3444_ (.Y(_0638_),
    .A(_0629_),
    .B(_0630_));
 sg13g2_and2_1 _3445_ (.A(\line_lfsr[3] ),
    .B(_0411_),
    .X(_0639_));
 sg13g2_xnor2_1 _3446_ (.Y(_0640_),
    .A(_0400_),
    .B(_0407_));
 sg13g2_xnor2_1 _3447_ (.Y(_0641_),
    .A(_0403_),
    .B(_0404_));
 sg13g2_xnor2_1 _3448_ (.Y(_0642_),
    .A(\line_lfsr[0] ),
    .B(_0641_));
 sg13g2_xnor2_1 _3449_ (.Y(_0643_),
    .A(_0405_),
    .B(_0406_));
 sg13g2_xnor2_1 _3450_ (.Y(_0644_),
    .A(\line_lfsr[1] ),
    .B(_0643_));
 sg13g2_nor2_1 _3451_ (.A(_0642_),
    .B(_0644_),
    .Y(_0645_));
 sg13g2_nand2_1 _3452_ (.Y(_0646_),
    .A(\line_lfsr[2] ),
    .B(_0640_));
 sg13g2_o21ai_1 _3453_ (.B1(_0645_),
    .Y(_0647_),
    .A1(\line_lfsr[2] ),
    .A2(_0640_));
 sg13g2_o21ai_1 _3454_ (.B1(_0646_),
    .Y(_0648_),
    .A1(\line_lfsr[3] ),
    .A2(_0411_));
 sg13g2_xnor2_1 _3455_ (.Y(_0649_),
    .A(\line_lfsr[4] ),
    .B(_0638_));
 sg13g2_nor4_1 _3456_ (.A(_0639_),
    .B(_0647_),
    .C(_0648_),
    .D(_0649_),
    .Y(_0650_));
 sg13g2_o21ai_1 _3457_ (.B1(_0650_),
    .Y(_0651_),
    .A1(\line_lfsr[5] ),
    .A2(_0637_));
 sg13g2_a221oi_1 _3458_ (.B2(\line_lfsr[5] ),
    .C1(_0651_),
    .B1(_0637_),
    .A1(\line_lfsr[6] ),
    .Y(_0652_),
    .A2(_0636_));
 sg13g2_o21ai_1 _3459_ (.B1(_0652_),
    .Y(_0653_),
    .A1(\line_lfsr[6] ),
    .A2(_0636_));
 sg13g2_nor4_2 _3460_ (.A(_2058_),
    .B(net775),
    .C(_0386_),
    .Y(_0654_),
    .D(_0653_));
 sg13g2_nor2_1 _3461_ (.A(net774),
    .B(_0654_),
    .Y(_0655_));
 sg13g2_or2_1 _3462_ (.X(_0656_),
    .B(_0654_),
    .A(net773));
 sg13g2_nand2_1 _3463_ (.Y(_0657_),
    .A(_0416_),
    .B(_0417_));
 sg13g2_o21ai_1 _3464_ (.B1(_0419_),
    .Y(_0658_),
    .A1(_0416_),
    .A2(_0418_));
 sg13g2_a221oi_1 _3465_ (.B2(net773),
    .C1(_0615_),
    .B1(_0658_),
    .A1(_0390_),
    .Y(_0659_),
    .A2(_0655_));
 sg13g2_or2_1 _3466_ (.X(_0660_),
    .B(_0659_),
    .A(_0625_));
 sg13g2_nand2_1 _3467_ (.Y(_0661_),
    .A(_0627_),
    .B(_0660_));
 sg13g2_nor2_1 _3468_ (.A(net969),
    .B(net968),
    .Y(_0662_));
 sg13g2_nor3_2 _3469_ (.A(_1528_),
    .B(_1532_),
    .C(_0564_),
    .Y(_0663_));
 sg13g2_nor2_1 _3470_ (.A(net942),
    .B(_0663_),
    .Y(_0664_));
 sg13g2_o21ai_1 _3471_ (.B1(_0664_),
    .Y(_0665_),
    .A1(_0008_),
    .A2(_0662_));
 sg13g2_inv_1 _3472_ (.Y(_0666_),
    .A(_0665_));
 sg13g2_o21ai_1 _3473_ (.B1(_0666_),
    .Y(_0667_),
    .A1(_0627_),
    .A2(_0660_));
 sg13g2_nor2b_1 _3474_ (.A(_0667_),
    .B_N(_0661_),
    .Y(_0004_));
 sg13g2_nand2b_1 _3475_ (.Y(_0668_),
    .B(_0386_),
    .A_N(net777));
 sg13g2_nand3b_1 _3476_ (.B(_0655_),
    .C(_0668_),
    .Y(_0669_),
    .A_N(net775));
 sg13g2_nand2_1 _3477_ (.Y(_0670_),
    .A(_0416_),
    .B(_0419_));
 sg13g2_nand2_1 _3478_ (.Y(_0671_),
    .A(net773),
    .B(_0670_));
 sg13g2_a21oi_1 _3479_ (.A1(net774),
    .A2(_0670_),
    .Y(_0672_),
    .B1(_0615_));
 sg13g2_a21oi_1 _3480_ (.A1(_0669_),
    .A2(_0672_),
    .Y(_0673_),
    .B1(_0625_));
 sg13g2_a21oi_1 _3481_ (.A1(_0661_),
    .A2(_0673_),
    .Y(_0005_),
    .B1(_0665_));
 sg13g2_xnor2_1 _3482_ (.Y(_0674_),
    .A(_1531_),
    .B(_0414_));
 sg13g2_a221oi_1 _3483_ (.B2(net773),
    .C1(_0615_),
    .B1(_0674_),
    .A1(_0387_),
    .Y(_0675_),
    .A2(_0655_));
 sg13g2_or2_1 _3484_ (.X(_0676_),
    .B(_0675_),
    .A(_0625_));
 sg13g2_o21ai_1 _3485_ (.B1(net777),
    .Y(_0677_),
    .A1(net776),
    .A2(_0387_));
 sg13g2_nor2b_1 _3486_ (.A(_0654_),
    .B_N(_0677_),
    .Y(_0678_));
 sg13g2_xnor2_1 _3487_ (.Y(_0679_),
    .A(_0416_),
    .B(_0417_));
 sg13g2_or2_1 _3488_ (.X(_0680_),
    .B(_0626_),
    .A(_0422_));
 sg13g2_a21oi_1 _3489_ (.A1(net773),
    .A2(_0679_),
    .Y(_0681_),
    .B1(_0680_));
 sg13g2_o21ai_1 _3490_ (.B1(_0681_),
    .Y(_0682_),
    .A1(net773),
    .A2(_0678_));
 sg13g2_nand2_1 _3491_ (.Y(_0683_),
    .A(_0425_),
    .B(_0682_));
 sg13g2_xnor2_1 _3492_ (.Y(_0684_),
    .A(net777),
    .B(_0386_));
 sg13g2_a21oi_1 _3493_ (.A1(net775),
    .A2(_0684_),
    .Y(_0685_),
    .B1(_0654_));
 sg13g2_a221oi_1 _3494_ (.B2(net775),
    .C1(_0654_),
    .B1(_0684_),
    .A1(net777),
    .Y(_0686_),
    .A2(_0390_));
 sg13g2_nand2_1 _3495_ (.Y(_0687_),
    .A(_0420_),
    .B(_0657_));
 sg13g2_a21oi_1 _3496_ (.A1(net773),
    .A2(_0687_),
    .Y(_0688_),
    .B1(_0626_));
 sg13g2_o21ai_1 _3497_ (.B1(_0688_),
    .Y(_0689_),
    .A1(net774),
    .A2(_0686_));
 sg13g2_o21ai_1 _3498_ (.B1(_0689_),
    .Y(_0690_),
    .A1(_0425_),
    .A2(_0682_));
 sg13g2_a21o_1 _3499_ (.A2(_0690_),
    .A1(_0683_),
    .B1(_0676_),
    .X(_0691_));
 sg13g2_nand3_1 _3500_ (.B(_0683_),
    .C(_0690_),
    .A(_0676_),
    .Y(_0692_));
 sg13g2_and3_1 _3501_ (.X(_0002_),
    .A(_0666_),
    .B(_0691_),
    .C(_0692_));
 sg13g2_nand2b_1 _3502_ (.Y(_0693_),
    .B(_0685_),
    .A_N(net774));
 sg13g2_nand3_1 _3503_ (.B(_0416_),
    .C(_0417_),
    .A(_0415_),
    .Y(_0694_));
 sg13g2_and2_1 _3504_ (.A(_0420_),
    .B(_0694_),
    .X(_0695_));
 sg13g2_a21oi_1 _3505_ (.A1(net774),
    .A2(_0695_),
    .Y(_0696_),
    .B1(_0615_));
 sg13g2_a21oi_1 _3506_ (.A1(_0693_),
    .A2(_0696_),
    .Y(_0697_),
    .B1(_0625_));
 sg13g2_a21oi_1 _3507_ (.A1(_0692_),
    .A2(_0697_),
    .Y(_0003_),
    .B1(_0665_));
 sg13g2_a21oi_1 _3508_ (.A1(net775),
    .A2(_0389_),
    .Y(_0698_),
    .B1(_0656_));
 sg13g2_o21ai_1 _3509_ (.B1(_0421_),
    .Y(_0699_),
    .A1(net775),
    .A2(_0389_));
 sg13g2_nor2_1 _3510_ (.A(net775),
    .B(_0684_),
    .Y(_0700_));
 sg13g2_o21ai_1 _3511_ (.B1(_0699_),
    .Y(_0701_),
    .A1(_0425_),
    .A2(_0700_));
 sg13g2_a21oi_1 _3512_ (.A1(_0415_),
    .A2(_0417_),
    .Y(_0702_),
    .B1(_0416_));
 sg13g2_nor3_1 _3513_ (.A(_0425_),
    .B(_0671_),
    .C(_0702_),
    .Y(_0703_));
 sg13g2_a21oi_1 _3514_ (.A1(_0698_),
    .A2(_0701_),
    .Y(_0704_),
    .B1(_0703_));
 sg13g2_or2_1 _3515_ (.X(_0705_),
    .B(_0704_),
    .A(_0626_));
 sg13g2_nor2b_1 _3516_ (.A(_0671_),
    .B_N(_0420_),
    .Y(_0706_));
 sg13g2_a21oi_1 _3517_ (.A1(net777),
    .A2(_0390_),
    .Y(_0707_),
    .B1(net774));
 sg13g2_nor3_1 _3518_ (.A(_0625_),
    .B(_0706_),
    .C(_0707_),
    .Y(_0708_));
 sg13g2_nor3_1 _3519_ (.A(_0615_),
    .B(_0665_),
    .C(_0708_),
    .Y(_0709_));
 sg13g2_and2_1 _3520_ (.A(_0705_),
    .B(_0709_),
    .X(_0000_));
 sg13g2_o21ai_1 _3521_ (.B1(_0698_),
    .Y(_0710_),
    .A1(net775),
    .A2(_0668_));
 sg13g2_nand2_1 _3522_ (.Y(_0711_),
    .A(_0419_),
    .B(_0702_));
 sg13g2_a21oi_1 _3523_ (.A1(net774),
    .A2(_0711_),
    .Y(_0712_),
    .B1(_0615_));
 sg13g2_a21oi_1 _3524_ (.A1(_0710_),
    .A2(_0712_),
    .Y(_0713_),
    .B1(_0625_));
 sg13g2_a21oi_1 _3525_ (.A1(_0705_),
    .A2(_0713_),
    .Y(_0001_),
    .B1(_0665_));
 sg13g2_nor2_1 _3526_ (.A(net960),
    .B(net942),
    .Y(_0714_));
 sg13g2_nand4_1 _3527_ (.B(net904),
    .C(_0663_),
    .A(net252),
    .Y(_0007_),
    .D(_0714_));
 sg13g2_nor3_1 _3528_ (.A(net972),
    .B(net971),
    .C(net970),
    .Y(_0715_));
 sg13g2_nor2b_1 _3529_ (.A(net967),
    .B_N(\hvsync_gen.hpos[9] ),
    .Y(_0716_));
 sg13g2_nand3b_1 _3530_ (.B(_0716_),
    .C(net969),
    .Y(_0717_),
    .A_N(_0715_));
 sg13g2_nand4_1 _3531_ (.B(net971),
    .C(net970),
    .A(net973),
    .Y(_0718_),
    .D(net969));
 sg13g2_a21oi_1 _3532_ (.A1(_0716_),
    .A2(_0718_),
    .Y(_0719_),
    .B1(net264));
 sg13g2_a21o_2 _3533_ (.A2(_0717_),
    .A1(_1968_),
    .B1(_0719_),
    .X(_0006_));
 sg13g2_nand2_1 _3534_ (.Y(_0720_),
    .A(net84),
    .B(net190));
 sg13g2_xor2_1 _3535_ (.B(\audio_sample_lpf[0] ),
    .A(net84),
    .X(\audio_pwm_accum_next[0] ));
 sg13g2_nand2_1 _3536_ (.Y(_0721_),
    .A(net206),
    .B(\audio_sample_lpf[1] ));
 sg13g2_nor2_1 _3537_ (.A(\audio_pwm_accum[1] ),
    .B(\audio_sample_lpf[1] ),
    .Y(_0722_));
 sg13g2_xor2_1 _3538_ (.B(\audio_sample_lpf[1] ),
    .A(net206),
    .X(_0723_));
 sg13g2_xnor2_1 _3539_ (.Y(\audio_pwm_accum_next[1] ),
    .A(_0720_),
    .B(net207));
 sg13g2_o21ai_1 _3540_ (.B1(_0721_),
    .Y(_0724_),
    .A1(_0720_),
    .A2(_0722_));
 sg13g2_xnor2_1 _3541_ (.Y(_0725_),
    .A(net242),
    .B(net200));
 sg13g2_nor2b_1 _3542_ (.A(_0725_),
    .B_N(_0724_),
    .Y(_0726_));
 sg13g2_xnor2_1 _3543_ (.Y(\audio_pwm_accum_next[2] ),
    .A(_0724_),
    .B(_0725_));
 sg13g2_a21o_1 _3544_ (.A2(net200),
    .A1(net242),
    .B1(_0726_),
    .X(_0727_));
 sg13g2_xnor2_1 _3545_ (.Y(_0728_),
    .A(net246),
    .B(\audio_sample_lpf[3] ));
 sg13g2_nor2b_1 _3546_ (.A(_0728_),
    .B_N(_0727_),
    .Y(_0729_));
 sg13g2_xnor2_1 _3547_ (.Y(\audio_pwm_accum_next[3] ),
    .A(_0727_),
    .B(net247));
 sg13g2_a21o_1 _3548_ (.A2(\audio_sample_lpf[3] ),
    .A1(net246),
    .B1(_0729_),
    .X(_0730_));
 sg13g2_xnor2_1 _3549_ (.Y(_0731_),
    .A(net254),
    .B(net205));
 sg13g2_nor2b_1 _3550_ (.A(_0731_),
    .B_N(_0730_),
    .Y(_0732_));
 sg13g2_xnor2_1 _3551_ (.Y(\audio_pwm_accum_next[4] ),
    .A(_0730_),
    .B(_0731_));
 sg13g2_a21o_1 _3552_ (.A2(\audio_sample_lpf[4] ),
    .A1(\audio_pwm_accum[4] ),
    .B1(_0732_),
    .X(_0733_));
 sg13g2_nand2_1 _3553_ (.Y(_0734_),
    .A(net232),
    .B(net228));
 sg13g2_xnor2_1 _3554_ (.Y(_0735_),
    .A(net232),
    .B(net228));
 sg13g2_xnor2_1 _3555_ (.Y(\audio_pwm_accum_next[5] ),
    .A(_0733_),
    .B(_0735_));
 sg13g2_xnor2_1 _3556_ (.Y(_0736_),
    .A(net265),
    .B(\audio_sample_lpf[6] ));
 sg13g2_o21ai_1 _3557_ (.B1(_0733_),
    .Y(_0737_),
    .A1(\audio_pwm_accum[5] ),
    .A2(\audio_sample_lpf[5] ));
 sg13g2_a21oi_1 _3558_ (.A1(_0734_),
    .A2(_0737_),
    .Y(_0738_),
    .B1(net266));
 sg13g2_nand3_1 _3559_ (.B(_0736_),
    .C(_0737_),
    .A(_0734_),
    .Y(_0739_));
 sg13g2_nor2b_1 _3560_ (.A(net267),
    .B_N(_0739_),
    .Y(\audio_pwm_accum_next[6] ));
 sg13g2_a21oi_1 _3561_ (.A1(\audio_pwm_accum[6] ),
    .A2(net221),
    .Y(_0740_),
    .B1(_0738_));
 sg13g2_nand2_1 _3562_ (.Y(_0741_),
    .A(net244),
    .B(\audio_sample_lpf[7] ));
 sg13g2_nor2_1 _3563_ (.A(\audio_pwm_accum[7] ),
    .B(\audio_sample_lpf[7] ),
    .Y(_0742_));
 sg13g2_xor2_1 _3564_ (.B(net239),
    .A(net244),
    .X(_0743_));
 sg13g2_xnor2_1 _3565_ (.Y(\audio_pwm_accum_next[7] ),
    .A(_0740_),
    .B(_0743_));
 sg13g2_o21ai_1 _3566_ (.B1(_0741_),
    .Y(_0744_),
    .A1(_0740_),
    .A2(_0742_));
 sg13g2_xnor2_1 _3567_ (.Y(_0745_),
    .A(net248),
    .B(net175));
 sg13g2_nor2b_1 _3568_ (.A(_0745_),
    .B_N(_0744_),
    .Y(_0746_));
 sg13g2_xnor2_1 _3569_ (.Y(\audio_pwm_accum_next[8] ),
    .A(_0744_),
    .B(_0745_));
 sg13g2_nand2_1 _3570_ (.Y(_0747_),
    .A(\audio_pwm_accum[9] ),
    .B(\audio_sample_lpf[9] ));
 sg13g2_nor2_1 _3571_ (.A(\audio_pwm_accum[9] ),
    .B(\audio_sample_lpf[9] ),
    .Y(_0748_));
 sg13g2_xor2_1 _3572_ (.B(net217),
    .A(net259),
    .X(_0749_));
 sg13g2_a21oi_1 _3573_ (.A1(net248),
    .A2(net175),
    .Y(_0750_),
    .B1(_0746_));
 sg13g2_xnor2_1 _3574_ (.Y(\audio_pwm_accum_next[9] ),
    .A(_0749_),
    .B(_0750_));
 sg13g2_o21ai_1 _3575_ (.B1(_0747_),
    .Y(audio_pwm),
    .A1(_0748_),
    .A2(_0750_));
 sg13g2_nor3_1 _3576_ (.A(\hvsync_gen.hpos[3] ),
    .B(\hvsync_gen.hpos[2] ),
    .C(net969),
    .Y(_0751_));
 sg13g2_nor2_1 _3577_ (.A(net253),
    .B(\hvsync_gen.hpos[0] ),
    .Y(_0752_));
 sg13g2_and4_1 _3578_ (.A(_1967_),
    .B(_0715_),
    .C(_0751_),
    .D(_0752_),
    .X(_0753_));
 sg13g2_nand4_1 _3579_ (.B(_0715_),
    .C(_0751_),
    .A(_1967_),
    .Y(_0754_),
    .D(_0752_));
 sg13g2_nor2_2 _3580_ (.A(\hvsync_gen.vpos[0] ),
    .B(\hvsync_gen.vpos[1] ),
    .Y(_0755_));
 sg13g2_nand3_1 _3581_ (.B(_0562_),
    .C(_0755_),
    .A(_1781_),
    .Y(_0756_));
 sg13g2_nor4_1 _3582_ (.A(\hvsync_gen.vpos[2] ),
    .B(net952),
    .C(\hvsync_gen.vpos[8] ),
    .D(net942),
    .Y(_0757_));
 sg13g2_nor2b_2 _3583_ (.A(_0756_),
    .B_N(_0757_),
    .Y(_0758_));
 sg13g2_and2_1 _3584_ (.A(net899),
    .B(net884),
    .X(_0759_));
 sg13g2_nand2_1 _3585_ (.Y(_0760_),
    .A(net899),
    .B(net884));
 sg13g2_nand3_1 _3586_ (.B(net198),
    .C(net877),
    .A(\sample_beat_ctr[0] ),
    .Y(_0761_));
 sg13g2_nand2_1 _3587_ (.Y(_0762_),
    .A(\sample_beat_ctr[0] ),
    .B(net198));
 sg13g2_nor2_2 _3588_ (.A(net194),
    .B(_0762_),
    .Y(_0763_));
 sg13g2_or2_2 _3589_ (.X(_0764_),
    .B(_0762_),
    .A(\sample_beat_ctr[1] ));
 sg13g2_nor2_1 _3590_ (.A(net874),
    .B(_0764_),
    .Y(_0765_));
 sg13g2_mux2_1 _3591_ (.A0(net97),
    .A1(net1005),
    .S(net864),
    .X(_0059_));
 sg13g2_nor2_1 _3592_ (.A(net90),
    .B(net865),
    .Y(_0766_));
 sg13g2_nand2_2 _3593_ (.Y(_0767_),
    .A(net1003),
    .B(net998));
 sg13g2_xor2_1 _3594_ (.B(net999),
    .A(net1001),
    .X(_0768_));
 sg13g2_a21oi_1 _3595_ (.A1(net865),
    .A2(net928),
    .Y(_0060_),
    .B1(_0766_));
 sg13g2_nor2_1 _3596_ (.A(net103),
    .B(net865),
    .Y(_0769_));
 sg13g2_and2_1 _3597_ (.A(net1002),
    .B(net996),
    .X(_0770_));
 sg13g2_nand2_2 _3598_ (.Y(_0771_),
    .A(net1001),
    .B(net995));
 sg13g2_nand2_1 _3599_ (.Y(_0772_),
    .A(net998),
    .B(net927));
 sg13g2_nor2_2 _3600_ (.A(net1003),
    .B(net993),
    .Y(_0773_));
 sg13g2_or2_2 _3601_ (.X(_0774_),
    .B(net996),
    .A(net1004));
 sg13g2_nor2_2 _3602_ (.A(net1000),
    .B(net995),
    .Y(_0775_));
 sg13g2_a21oi_2 _3603_ (.B1(net992),
    .Y(_0776_),
    .A2(net997),
    .A1(net1003));
 sg13g2_a21oi_1 _3604_ (.A1(net997),
    .A2(net926),
    .Y(_0777_),
    .B1(_0776_));
 sg13g2_a21oi_1 _3605_ (.A1(net865),
    .A2(_0777_),
    .Y(_0061_),
    .B1(_0769_));
 sg13g2_nor2_1 _3606_ (.A(net93),
    .B(net865),
    .Y(_0778_));
 sg13g2_and2_2 _3607_ (.A(net998),
    .B(net991),
    .X(_0779_));
 sg13g2_nand2_1 _3608_ (.Y(_0780_),
    .A(net926),
    .B(_0779_));
 sg13g2_nand2_2 _3609_ (.Y(_0781_),
    .A(net998),
    .B(net995));
 sg13g2_nor2_1 _3610_ (.A(net1001),
    .B(net987),
    .Y(_0782_));
 sg13g2_or2_1 _3611_ (.X(_0783_),
    .B(net988),
    .A(net1003));
 sg13g2_a21oi_2 _3612_ (.B1(net988),
    .Y(_0784_),
    .A2(net926),
    .A1(net997));
 sg13g2_a21oi_2 _3613_ (.B1(_0784_),
    .Y(_0785_),
    .A2(_0779_),
    .A1(net927));
 sg13g2_a21oi_1 _3614_ (.A1(net865),
    .A2(_0785_),
    .Y(_0062_),
    .B1(_0778_));
 sg13g2_nor2_1 _3615_ (.A(net88),
    .B(net865),
    .Y(_0786_));
 sg13g2_and2_1 _3616_ (.A(net986),
    .B(net980),
    .X(_0787_));
 sg13g2_nand2_2 _3617_ (.Y(_0788_),
    .A(net989),
    .B(net983));
 sg13g2_nor2_2 _3618_ (.A(_0772_),
    .B(_0788_),
    .Y(_0789_));
 sg13g2_xnor2_1 _3619_ (.Y(_0790_),
    .A(\songpos[4] ),
    .B(_0780_));
 sg13g2_xnor2_1 _3620_ (.Y(_0791_),
    .A(net938),
    .B(_0780_));
 sg13g2_a21oi_1 _3621_ (.A1(net865),
    .A2(_0790_),
    .Y(_0063_),
    .B1(_0786_));
 sg13g2_nand2_1 _3622_ (.Y(_0792_),
    .A(net979),
    .B(_0789_));
 sg13g2_inv_1 _3623_ (.Y(_0793_),
    .A(_0792_));
 sg13g2_xnor2_1 _3624_ (.Y(_0794_),
    .A(net979),
    .B(_0789_));
 sg13g2_mux2_1 _3625_ (.A0(net91),
    .A1(_0794_),
    .S(net864),
    .X(_0064_));
 sg13g2_nor2_1 _3626_ (.A(net109),
    .B(net864),
    .Y(_0795_));
 sg13g2_xnor2_1 _3627_ (.Y(_0796_),
    .A(\songpos[6] ),
    .B(_0792_));
 sg13g2_a21oi_1 _3628_ (.A1(net864),
    .A2(_0796_),
    .Y(_0065_),
    .B1(_0795_));
 sg13g2_nor2_1 _3629_ (.A(net124),
    .B(_0765_),
    .Y(_0797_));
 sg13g2_nor2_2 _3630_ (.A(_0435_),
    .B(_0792_),
    .Y(_0798_));
 sg13g2_a21oi_1 _3631_ (.A1(\songpos[6] ),
    .A2(_0793_),
    .Y(_0799_),
    .B1(net976));
 sg13g2_nor2_2 _3632_ (.A(_0798_),
    .B(_0799_),
    .Y(_0800_));
 sg13g2_or2_1 _3633_ (.X(_0801_),
    .B(_0799_),
    .A(_0798_));
 sg13g2_a21oi_1 _3634_ (.A1(net864),
    .A2(_0800_),
    .Y(_0066_),
    .B1(_0797_));
 sg13g2_nor2_1 _3635_ (.A(net92),
    .B(net864),
    .Y(_0802_));
 sg13g2_nor2_2 _3636_ (.A(net978),
    .B(net977),
    .Y(_0803_));
 sg13g2_or2_2 _3637_ (.X(_0804_),
    .B(net977),
    .A(net978));
 sg13g2_nor2_2 _3638_ (.A(net974),
    .B(_0804_),
    .Y(_0805_));
 sg13g2_nand3_1 _3639_ (.B(_0789_),
    .C(_0805_),
    .A(\songpos[8] ),
    .Y(_0806_));
 sg13g2_xnor2_1 _3640_ (.Y(_0807_),
    .A(net937),
    .B(_0798_));
 sg13g2_and2_1 _3641_ (.A(_0806_),
    .B(_0807_),
    .X(_0808_));
 sg13g2_nand2_1 _3642_ (.Y(_0809_),
    .A(_0806_),
    .B(_0807_));
 sg13g2_a21oi_1 _3643_ (.A1(net864),
    .A2(_0808_),
    .Y(_0067_),
    .B1(_0802_));
 sg13g2_nand2_1 _3644_ (.Y(_0810_),
    .A(net1017),
    .B(net899));
 sg13g2_inv_2 _3645_ (.Y(_0811_),
    .A(net882));
 sg13g2_nor2_2 _3646_ (.A(\kick_ctr[0] ),
    .B(\kick_ctr[1] ),
    .Y(_0812_));
 sg13g2_or2_1 _3647_ (.X(_0813_),
    .B(\kick_ctr[1] ),
    .A(\kick_ctr[0] ));
 sg13g2_o21ai_1 _3648_ (.B1(net1009),
    .Y(_0814_),
    .A1(_0763_),
    .A2(net924));
 sg13g2_nor2_2 _3649_ (.A(net874),
    .B(_0763_),
    .Y(_0815_));
 sg13g2_nand2b_2 _3650_ (.Y(_0816_),
    .B(net863),
    .A_N(_0814_));
 sg13g2_nor2_1 _3651_ (.A(net74),
    .B(_0816_),
    .Y(_0817_));
 sg13g2_nand2_2 _3652_ (.Y(_0818_),
    .A(net998),
    .B(_0774_));
 sg13g2_nor2_1 _3653_ (.A(_0794_),
    .B(_0818_),
    .Y(_0819_));
 sg13g2_nand2_1 _3654_ (.Y(_0820_),
    .A(net985),
    .B(_0785_));
 sg13g2_o21ai_1 _3655_ (.B1(_0781_),
    .Y(_0821_),
    .A1(_0771_),
    .A2(_0820_));
 sg13g2_o21ai_1 _3656_ (.B1(_0767_),
    .Y(_0822_),
    .A1(_0771_),
    .A2(_0820_));
 sg13g2_nor2b_1 _3657_ (.A(net1002),
    .B_N(net999),
    .Y(_0823_));
 sg13g2_nand2b_1 _3658_ (.Y(_0824_),
    .B(net1004),
    .A_N(net1000));
 sg13g2_nor2b_1 _3659_ (.A(net997),
    .B_N(net992),
    .Y(_0825_));
 sg13g2_nand2b_2 _3660_ (.Y(_0826_),
    .B(net992),
    .A_N(net997));
 sg13g2_nor2_1 _3661_ (.A(net998),
    .B(_0773_),
    .Y(_0827_));
 sg13g2_nor2b_2 _3662_ (.A(net1003),
    .B_N(net993),
    .Y(_0828_));
 sg13g2_or2_1 _3663_ (.X(_0829_),
    .B(_0828_),
    .A(net928));
 sg13g2_nand3_1 _3664_ (.B(_0790_),
    .C(_0829_),
    .A(net989),
    .Y(_0830_));
 sg13g2_nand3_1 _3665_ (.B(_0785_),
    .C(_0818_),
    .A(\songpos[4] ),
    .Y(_0831_));
 sg13g2_nand2_1 _3666_ (.Y(_0832_),
    .A(_0772_),
    .B(_0788_));
 sg13g2_nor2b_2 _3667_ (.A(net994),
    .B_N(net999),
    .Y(_0833_));
 sg13g2_xnor2_1 _3668_ (.Y(_0834_),
    .A(net999),
    .B(net994));
 sg13g2_nor2b_2 _3669_ (.A(net989),
    .B_N(net996),
    .Y(_0835_));
 sg13g2_nand2b_1 _3670_ (.Y(_0836_),
    .B(net1004),
    .A_N(_0835_));
 sg13g2_nand4_1 _3671_ (.B(net983),
    .C(net928),
    .A(net995),
    .Y(_0837_),
    .D(_0785_));
 sg13g2_a22oi_1 _3672_ (.Y(_0838_),
    .B1(_0794_),
    .B2(_0837_),
    .A2(_0767_),
    .A1(net979));
 sg13g2_xor2_1 _3673_ (.B(_0821_),
    .A(_0819_),
    .X(_0839_));
 sg13g2_a22oi_1 _3674_ (.Y(_0840_),
    .B1(_0830_),
    .B2(_0819_),
    .A2(_0822_),
    .A1(_0794_));
 sg13g2_o21ai_1 _3675_ (.B1(_0796_),
    .Y(_0841_),
    .A1(_0800_),
    .A2(_0840_));
 sg13g2_a21oi_1 _3676_ (.A1(_0800_),
    .A2(_0839_),
    .Y(_0842_),
    .B1(_0841_));
 sg13g2_o21ai_1 _3677_ (.B1(_0794_),
    .Y(_0843_),
    .A1(_0834_),
    .A2(_0836_));
 sg13g2_a21oi_1 _3678_ (.A1(_0831_),
    .A2(_0832_),
    .Y(_0844_),
    .B1(_0794_));
 sg13g2_nor2_1 _3679_ (.A(_0801_),
    .B(_0844_),
    .Y(_0845_));
 sg13g2_a221oi_1 _3680_ (.B2(_0845_),
    .C1(_0796_),
    .B1(_0843_),
    .A1(_0801_),
    .Y(_0846_),
    .A2(_0838_));
 sg13g2_nor3_1 _3681_ (.A(_0808_),
    .B(_0842_),
    .C(_0846_),
    .Y(_0847_));
 sg13g2_nor3_1 _3682_ (.A(_0773_),
    .B(_0809_),
    .C(_0820_),
    .Y(_0848_));
 sg13g2_nor3_1 _3683_ (.A(_0764_),
    .B(_0847_),
    .C(_0848_),
    .Y(_0849_));
 sg13g2_or3_1 _3684_ (.A(net874),
    .B(_0814_),
    .C(_0849_),
    .X(_0850_));
 sg13g2_a21oi_1 _3685_ (.A1(_1524_),
    .A2(net779),
    .Y(_0068_),
    .B1(_0817_));
 sg13g2_nor2_1 _3686_ (.A(_1524_),
    .B(net779),
    .Y(_0851_));
 sg13g2_nor2_2 _3687_ (.A(_0764_),
    .B(net779),
    .Y(_0852_));
 sg13g2_xnor2_1 _3688_ (.Y(_0853_),
    .A(net173),
    .B(_0851_));
 sg13g2_nor2_1 _3689_ (.A(_0852_),
    .B(net174),
    .Y(_0069_));
 sg13g2_and2_1 _3690_ (.A(net253),
    .B(\hvsync_gen.hpos[0] ),
    .X(_0854_));
 sg13g2_and2_1 _3691_ (.A(\hvsync_gen.hpos[2] ),
    .B(_0854_),
    .X(_0855_));
 sg13g2_and2_2 _3692_ (.A(\hvsync_gen.hpos[3] ),
    .B(_0855_),
    .X(_0856_));
 sg13g2_nand3_1 _3693_ (.B(_0393_),
    .C(_0856_),
    .A(net972),
    .Y(_0857_));
 sg13g2_nor3_2 _3694_ (.A(net971),
    .B(_1968_),
    .C(_0857_),
    .Y(_0858_));
 sg13g2_nor2b_2 _3695_ (.A(_0858_),
    .B_N(net1014),
    .Y(_0859_));
 sg13g2_nand2b_2 _3696_ (.Y(_0860_),
    .B(net1014),
    .A_N(_0858_));
 sg13g2_and2_1 _3697_ (.A(net66),
    .B(net830),
    .X(_0070_));
 sg13g2_nor3_1 _3698_ (.A(_0752_),
    .B(_0854_),
    .C(_0860_),
    .Y(_0071_));
 sg13g2_nor2_1 _3699_ (.A(net263),
    .B(_0854_),
    .Y(_0861_));
 sg13g2_nor3_1 _3700_ (.A(_0855_),
    .B(_0860_),
    .C(_0861_),
    .Y(_0072_));
 sg13g2_o21ai_1 _3701_ (.B1(net1014),
    .Y(_0862_),
    .A1(net277),
    .A2(_0855_));
 sg13g2_nor2_1 _3702_ (.A(_0856_),
    .B(_0862_),
    .Y(_0073_));
 sg13g2_o21ai_1 _3703_ (.B1(net1014),
    .Y(_0863_),
    .A1(net972),
    .A2(_0856_));
 sg13g2_a21oi_1 _3704_ (.A1(net972),
    .A2(_0856_),
    .Y(_0074_),
    .B1(_0863_));
 sg13g2_nor2b_1 _3705_ (.A(_0394_),
    .B_N(_0856_),
    .Y(_0864_));
 sg13g2_a21oi_1 _3706_ (.A1(net972),
    .A2(_0856_),
    .Y(_0865_),
    .B1(net971));
 sg13g2_nor3_1 _3707_ (.A(_0860_),
    .B(_0864_),
    .C(_0865_),
    .Y(_0075_));
 sg13g2_and2_1 _3708_ (.A(net970),
    .B(_0864_),
    .X(_0866_));
 sg13g2_nor2_1 _3709_ (.A(net970),
    .B(_0864_),
    .Y(_0867_));
 sg13g2_nor3_1 _3710_ (.A(_0860_),
    .B(_0866_),
    .C(_0867_),
    .Y(_0076_));
 sg13g2_nor2_1 _3711_ (.A(net969),
    .B(_0866_),
    .Y(_0868_));
 sg13g2_nor2b_2 _3712_ (.A(_0718_),
    .B_N(_0856_),
    .Y(_0869_));
 sg13g2_nor3_1 _3713_ (.A(_0860_),
    .B(_0868_),
    .C(_0869_),
    .Y(_0077_));
 sg13g2_o21ai_1 _3714_ (.B1(net830),
    .Y(_0870_),
    .A1(net967),
    .A2(_0869_));
 sg13g2_a21oi_1 _3715_ (.A1(net967),
    .A2(_0869_),
    .Y(_0078_),
    .B1(_0870_));
 sg13g2_nor2b_1 _3716_ (.A(net183),
    .B_N(_0869_),
    .Y(_0871_));
 sg13g2_o21ai_1 _3717_ (.B1(net830),
    .Y(_0872_),
    .A1(\hvsync_gen.hpos[9] ),
    .A2(_0871_));
 sg13g2_a21oi_1 _3718_ (.A1(\hvsync_gen.hpos[9] ),
    .A2(_0871_),
    .Y(_0079_),
    .B1(_0872_));
 sg13g2_mux2_1 _3719_ (.A0(\frame_count[0] ),
    .A1(net70),
    .S(_0759_),
    .X(_0080_));
 sg13g2_nand2_1 _3720_ (.Y(_0873_),
    .A(\frame_count[0] ),
    .B(net877));
 sg13g2_or3_2 _3721_ (.A(\frame_count[0] ),
    .B(\frame_count[1] ),
    .C(net874),
    .X(_0874_));
 sg13g2_and3_1 _3722_ (.X(_0875_),
    .A(\frame_count[0] ),
    .B(\frame_count[1] ),
    .C(net877));
 sg13g2_xnor2_1 _3723_ (.Y(_0081_),
    .A(net192),
    .B(_0873_));
 sg13g2_xor2_1 _3724_ (.B(_0875_),
    .A(net179),
    .X(_0082_));
 sg13g2_a21oi_1 _3725_ (.A1(\frame_count[2] ),
    .A2(_0875_),
    .Y(_0876_),
    .B1(net142));
 sg13g2_and3_2 _3726_ (.X(_0877_),
    .A(net179),
    .B(net142),
    .C(_0875_));
 sg13g2_nor2_1 _3727_ (.A(net143),
    .B(_0877_),
    .Y(_0083_));
 sg13g2_xor2_1 _3728_ (.B(_0877_),
    .A(net229),
    .X(_0084_));
 sg13g2_a21oi_1 _3729_ (.A1(\frame_count[4] ),
    .A2(_0877_),
    .Y(_0878_),
    .B1(net203));
 sg13g2_nand3_1 _3730_ (.B(net203),
    .C(_0877_),
    .A(net278),
    .Y(_0879_));
 sg13g2_nor2b_1 _3731_ (.A(net204),
    .B_N(_0879_),
    .Y(_0085_));
 sg13g2_xnor2_1 _3732_ (.Y(_0086_),
    .A(net177),
    .B(_0879_));
 sg13g2_nand4_1 _3733_ (.B(\frame_count[5] ),
    .C(\frame_count[6] ),
    .A(\frame_count[4] ),
    .Y(_0880_),
    .D(_0877_));
 sg13g2_xnor2_1 _3734_ (.Y(_0087_),
    .A(net131),
    .B(_0880_));
 sg13g2_a21oi_2 _3735_ (.B1(net884),
    .Y(_0881_),
    .A2(_0755_),
    .A1(_0030_));
 sg13g2_nor2_2 _3736_ (.A(net883),
    .B(_0881_),
    .Y(_0882_));
 sg13g2_nor2b_1 _3737_ (.A(_0758_),
    .B_N(net154),
    .Y(_0883_));
 sg13g2_mux2_1 _3738_ (.A0(net225),
    .A1(_0883_),
    .S(net862),
    .X(_0088_));
 sg13g2_nor2_1 _3739_ (.A(\line_lfsr[2] ),
    .B(_0758_),
    .Y(_0884_));
 sg13g2_nor2_1 _3740_ (.A(net154),
    .B(net862),
    .Y(_0885_));
 sg13g2_a21oi_1 _3741_ (.A1(net862),
    .A2(_0884_),
    .Y(_0089_),
    .B1(_0885_));
 sg13g2_nor2b_1 _3742_ (.A(net884),
    .B_N(net162),
    .Y(_0886_));
 sg13g2_mux2_1 _3743_ (.A0(net170),
    .A1(_0886_),
    .S(net862),
    .X(_0090_));
 sg13g2_nor2_1 _3744_ (.A(\line_lfsr[4] ),
    .B(net884),
    .Y(_0887_));
 sg13g2_nor2_1 _3745_ (.A(net162),
    .B(net862),
    .Y(_0888_));
 sg13g2_a21oi_1 _3746_ (.A1(_0882_),
    .A2(_0887_),
    .Y(_0091_),
    .B1(_0888_));
 sg13g2_nor2_1 _3747_ (.A(net168),
    .B(net884),
    .Y(_0889_));
 sg13g2_nor2_1 _3748_ (.A(net181),
    .B(_0882_),
    .Y(_0890_));
 sg13g2_a21oi_1 _3749_ (.A1(net862),
    .A2(_0889_),
    .Y(_0092_),
    .B1(net182));
 sg13g2_xnor2_1 _3750_ (.Y(_0891_),
    .A(\line_lfsr[0] ),
    .B(\line_lfsr[6] ));
 sg13g2_nor2_1 _3751_ (.A(net884),
    .B(_0891_),
    .Y(_0892_));
 sg13g2_mux2_1 _3752_ (.A0(net168),
    .A1(_0892_),
    .S(net862),
    .X(_0093_));
 sg13g2_nor2_1 _3753_ (.A(\line_lfsr[0] ),
    .B(net884),
    .Y(_0893_));
 sg13g2_nor2_1 _3754_ (.A(net185),
    .B(net862),
    .Y(_0894_));
 sg13g2_a21oi_1 _3755_ (.A1(_0882_),
    .A2(_0893_),
    .Y(_0094_),
    .B1(_0894_));
 sg13g2_nand2_1 _3756_ (.Y(_0895_),
    .A(net964),
    .B(_1541_));
 sg13g2_o21ai_1 _3757_ (.B1(net67),
    .Y(_0896_),
    .A1(_0031_),
    .A2(_0895_));
 sg13g2_nand2_1 _3758_ (.Y(_0897_),
    .A(net964),
    .B(_0874_));
 sg13g2_o21ai_1 _3759_ (.B1(_0897_),
    .Y(_0095_),
    .A1(_0874_),
    .A2(net68));
 sg13g2_or2_1 _3760_ (.X(_0898_),
    .B(_0874_),
    .A(net936));
 sg13g2_nor2_1 _3761_ (.A(_0440_),
    .B(_0898_),
    .Y(_0899_));
 sg13g2_a21oi_1 _3762_ (.A1(_1541_),
    .A2(_0898_),
    .Y(_0096_),
    .B1(_0899_));
 sg13g2_o21ai_1 _3763_ (.B1(net222),
    .Y(_0900_),
    .A1(_0440_),
    .A2(_0898_));
 sg13g2_o21ai_1 _3764_ (.B1(net223),
    .Y(_0097_),
    .A1(_2112_),
    .A2(_0898_));
 sg13g2_nor2_1 _3765_ (.A(net101),
    .B(net875),
    .Y(_0901_));
 sg13g2_nand2b_1 _3766_ (.Y(_0902_),
    .B(\nyan_x_offset[3] ),
    .A_N(\cos[0] ));
 sg13g2_xor2_1 _3767_ (.B(\nyan_x_offset[3] ),
    .A(\cos[0] ),
    .X(_0903_));
 sg13g2_a21oi_1 _3768_ (.A1(net875),
    .A2(_0903_),
    .Y(_0098_),
    .B1(_0901_));
 sg13g2_nor2b_1 _3769_ (.A(\nyan_x_offset[4] ),
    .B_N(\cos[1] ),
    .Y(_0904_));
 sg13g2_xnor2_1 _3770_ (.Y(_0905_),
    .A(\nyan_x_offset[4] ),
    .B(\cos[1] ));
 sg13g2_xor2_1 _3771_ (.B(_0905_),
    .A(_0902_),
    .X(_0906_));
 sg13g2_nor2_1 _3772_ (.A(net127),
    .B(net875),
    .Y(_0907_));
 sg13g2_a21oi_1 _3773_ (.A1(net875),
    .A2(_0906_),
    .Y(_0099_),
    .B1(_0907_));
 sg13g2_xor2_1 _3774_ (.B(\cos[2] ),
    .A(net962),
    .X(_0908_));
 sg13g2_a21oi_1 _3775_ (.A1(_0902_),
    .A2(_0905_),
    .Y(_0909_),
    .B1(_0904_));
 sg13g2_nand2_1 _3776_ (.Y(_0910_),
    .A(_0908_),
    .B(_0909_));
 sg13g2_nor2_1 _3777_ (.A(_0908_),
    .B(_0909_),
    .Y(_0911_));
 sg13g2_nor2_1 _3778_ (.A(net873),
    .B(_0911_),
    .Y(_0912_));
 sg13g2_a22oi_1 _3779_ (.Y(_0100_),
    .B1(_0910_),
    .B2(_0912_),
    .A2(net873),
    .A1(_1523_));
 sg13g2_nor2_1 _3780_ (.A(net106),
    .B(net875),
    .Y(_0913_));
 sg13g2_a21oi_1 _3781_ (.A1(_1538_),
    .A2(\cos[2] ),
    .Y(_0914_),
    .B1(_0911_));
 sg13g2_nand2_1 _3782_ (.Y(_0915_),
    .A(_1538_),
    .B(\cos[3] ));
 sg13g2_nor2_1 _3783_ (.A(_1538_),
    .B(\cos[3] ),
    .Y(_0916_));
 sg13g2_xnor2_1 _3784_ (.Y(_0917_),
    .A(net962),
    .B(\cos[3] ));
 sg13g2_xnor2_1 _3785_ (.Y(_0918_),
    .A(_0914_),
    .B(_0917_));
 sg13g2_a21oi_1 _3786_ (.A1(net875),
    .A2(_0918_),
    .Y(_0101_),
    .B1(_0913_));
 sg13g2_nor2b_1 _3787_ (.A(net962),
    .B_N(\cos[4] ),
    .Y(_0919_));
 sg13g2_nand2b_1 _3788_ (.Y(_0920_),
    .B(net962),
    .A_N(\cos[4] ));
 sg13g2_nand2b_1 _3789_ (.Y(_0921_),
    .B(_0920_),
    .A_N(_0919_));
 sg13g2_a21oi_1 _3790_ (.A1(_0914_),
    .A2(_0915_),
    .Y(_0922_),
    .B1(_0916_));
 sg13g2_xnor2_1 _3791_ (.Y(_0923_),
    .A(_0921_),
    .B(_0922_));
 sg13g2_nand2_1 _3792_ (.Y(_0924_),
    .A(net875),
    .B(_0923_));
 sg13g2_o21ai_1 _3793_ (.B1(_0924_),
    .Y(_0925_),
    .A1(net165),
    .A2(net875));
 sg13g2_inv_1 _3794_ (.Y(_0102_),
    .A(_0925_));
 sg13g2_nand2_1 _3795_ (.Y(_0926_),
    .A(net80),
    .B(net873));
 sg13g2_a21oi_1 _3796_ (.A1(_0920_),
    .A2(_0922_),
    .Y(_0927_),
    .B1(_0919_));
 sg13g2_xnor2_1 _3797_ (.Y(_0928_),
    .A(net962),
    .B(\cos[5] ));
 sg13g2_xnor2_1 _3798_ (.Y(_0929_),
    .A(_0927_),
    .B(_0928_));
 sg13g2_o21ai_1 _3799_ (.B1(_0926_),
    .Y(_0103_),
    .A1(net873),
    .A2(_0929_));
 sg13g2_a21oi_1 _3800_ (.A1(net962),
    .A2(_1567_),
    .Y(_0930_),
    .B1(_0927_));
 sg13g2_a21oi_1 _3801_ (.A1(_1538_),
    .A2(\cos[5] ),
    .Y(_0931_),
    .B1(_0930_));
 sg13g2_xnor2_1 _3802_ (.Y(_0932_),
    .A(net962),
    .B(\cos[6] ));
 sg13g2_xnor2_1 _3803_ (.Y(_0933_),
    .A(_0931_),
    .B(_0932_));
 sg13g2_mux2_1 _3804_ (.A0(net133),
    .A1(net781),
    .S(net876),
    .X(_0104_));
 sg13g2_nand2_1 _3805_ (.Y(_0934_),
    .A(net118),
    .B(_0923_));
 sg13g2_xnor2_1 _3806_ (.Y(_0105_),
    .A(net118),
    .B(_0924_));
 sg13g2_nor2_1 _3807_ (.A(net214),
    .B(net876),
    .Y(_0935_));
 sg13g2_nand2_1 _3808_ (.Y(_0936_),
    .A(net279),
    .B(_0929_));
 sg13g2_xor2_1 _3809_ (.B(_0929_),
    .A(\nyan_x_offset[0] ),
    .X(_0937_));
 sg13g2_nand2b_1 _3810_ (.Y(_0938_),
    .B(_0937_),
    .A_N(_0934_));
 sg13g2_xor2_1 _3811_ (.B(_0937_),
    .A(_0934_),
    .X(_0939_));
 sg13g2_a21oi_1 _3812_ (.A1(net876),
    .A2(_0939_),
    .Y(_0106_),
    .B1(_0935_));
 sg13g2_xnor2_1 _3813_ (.Y(_0940_),
    .A(\nyan_x_offset[1] ),
    .B(net780));
 sg13g2_a21oi_1 _3814_ (.A1(_0936_),
    .A2(_0938_),
    .Y(_0941_),
    .B1(_0940_));
 sg13g2_nand3_1 _3815_ (.B(_0938_),
    .C(_0940_),
    .A(_0936_),
    .Y(_0942_));
 sg13g2_nand2_1 _3816_ (.Y(_0943_),
    .A(net202),
    .B(net873));
 sg13g2_nand2_1 _3817_ (.Y(_0944_),
    .A(net876),
    .B(_0942_));
 sg13g2_o21ai_1 _3818_ (.B1(_0943_),
    .Y(_0107_),
    .A1(_0941_),
    .A2(_0944_));
 sg13g2_nand2_1 _3819_ (.Y(_0945_),
    .A(\nyan_x_offset[2] ),
    .B(net780));
 sg13g2_xnor2_1 _3820_ (.Y(_0946_),
    .A(\nyan_x_offset[2] ),
    .B(net780));
 sg13g2_a21oi_1 _3821_ (.A1(\nyan_x_offset[1] ),
    .A2(net780),
    .Y(_0947_),
    .B1(_0941_));
 sg13g2_inv_1 _3822_ (.Y(_0948_),
    .A(_0947_));
 sg13g2_xnor2_1 _3823_ (.Y(_0949_),
    .A(_0946_),
    .B(_0947_));
 sg13g2_nand2_1 _3824_ (.Y(_0950_),
    .A(net208),
    .B(net873));
 sg13g2_o21ai_1 _3825_ (.B1(_0950_),
    .Y(_0108_),
    .A1(net874),
    .A2(_0949_));
 sg13g2_xnor2_1 _3826_ (.Y(_0951_),
    .A(\nyan_x_offset[3] ),
    .B(net781));
 sg13g2_o21ai_1 _3827_ (.B1(_0948_),
    .Y(_0952_),
    .A1(\nyan_x_offset[2] ),
    .A2(net780));
 sg13g2_and3_1 _3828_ (.X(_0953_),
    .A(_0945_),
    .B(_0951_),
    .C(_0952_));
 sg13g2_a21oi_2 _3829_ (.B1(_0951_),
    .Y(_0954_),
    .A2(_0952_),
    .A1(_0945_));
 sg13g2_nor3_1 _3830_ (.A(net873),
    .B(_0953_),
    .C(_0954_),
    .Y(_0955_));
 sg13g2_a21o_1 _3831_ (.A2(net873),
    .A1(net270),
    .B1(_0955_),
    .X(_0109_));
 sg13g2_a21oi_1 _3832_ (.A1(\nyan_x_offset[3] ),
    .A2(net781),
    .Y(_0956_),
    .B1(_0954_));
 sg13g2_o21ai_1 _3833_ (.B1(net780),
    .Y(_0957_),
    .A1(\nyan_x_offset[3] ),
    .A2(_0954_));
 sg13g2_o21ai_1 _3834_ (.B1(net876),
    .Y(_0958_),
    .A1(net780),
    .A2(_0954_));
 sg13g2_nand2b_1 _3835_ (.Y(_0959_),
    .B(_0957_),
    .A_N(_0958_));
 sg13g2_xnor2_1 _3836_ (.Y(_0110_),
    .A(net260),
    .B(_0959_));
 sg13g2_a21oi_1 _3837_ (.A1(\nyan_x_offset[4] ),
    .A2(net780),
    .Y(_0960_),
    .B1(_0958_));
 sg13g2_o21ai_1 _3838_ (.B1(_0960_),
    .Y(_0961_),
    .A1(\nyan_x_offset[4] ),
    .A2(_0956_));
 sg13g2_xnor2_1 _3839_ (.Y(_0111_),
    .A(net963),
    .B(_0961_));
 sg13g2_o21ai_1 _3840_ (.B1(net974),
    .Y(_0962_),
    .A1(net978),
    .A2(net977));
 sg13g2_and2_2 _3841_ (.A(net937),
    .B(_0962_),
    .X(_0963_));
 sg13g2_nand2_2 _3842_ (.Y(_0964_),
    .A(net937),
    .B(_0962_));
 sg13g2_nor2b_2 _3843_ (.A(net986),
    .B_N(net980),
    .Y(_0965_));
 sg13g2_nand2b_2 _3844_ (.Y(_0966_),
    .B(net992),
    .A_N(net980));
 sg13g2_nor2b_2 _3845_ (.A(net981),
    .B_N(net986),
    .Y(_0967_));
 sg13g2_nand2b_1 _3846_ (.Y(_0968_),
    .B(net986),
    .A_N(net980));
 sg13g2_nand2_1 _3847_ (.Y(_0969_),
    .A(_0966_),
    .B(_0968_));
 sg13g2_a22oi_1 _3848_ (.Y(_0970_),
    .B1(_0966_),
    .B2(_0968_),
    .A2(net992),
    .A1(net986));
 sg13g2_nor3_1 _3849_ (.A(_0964_),
    .B(_0965_),
    .C(_0970_),
    .Y(_0971_));
 sg13g2_nand2_2 _3850_ (.Y(_0972_),
    .A(net937),
    .B(_0805_));
 sg13g2_nor2_2 _3851_ (.A(_1534_),
    .B(net993),
    .Y(_0973_));
 sg13g2_nand2_1 _3852_ (.Y(_0974_),
    .A(net987),
    .B(_0826_));
 sg13g2_nand2_2 _3853_ (.Y(_0975_),
    .A(net986),
    .B(_0834_));
 sg13g2_inv_1 _3854_ (.Y(_0976_),
    .A(_0975_));
 sg13g2_nand2_2 _3855_ (.Y(_0977_),
    .A(net998),
    .B(_1534_));
 sg13g2_nor2_1 _3856_ (.A(net989),
    .B(_0775_),
    .Y(_0978_));
 sg13g2_o21ai_1 _3857_ (.B1(net983),
    .Y(_0979_),
    .A1(net988),
    .A2(_0775_));
 sg13g2_nand2b_1 _3858_ (.Y(_0980_),
    .B(_0975_),
    .A_N(_0979_));
 sg13g2_a21oi_1 _3859_ (.A1(_0826_),
    .A2(_0967_),
    .Y(_0981_),
    .B1(_0963_));
 sg13g2_a221oi_1 _3860_ (.B2(_0981_),
    .C1(_0971_),
    .B1(_0980_),
    .A1(net937),
    .Y(_0982_),
    .A2(_0805_));
 sg13g2_nand3b_1 _3861_ (.B(_0966_),
    .C(_0963_),
    .Y(_0983_),
    .A_N(_0965_));
 sg13g2_nor2_1 _3862_ (.A(net980),
    .B(_0833_),
    .Y(_0984_));
 sg13g2_nor2_1 _3863_ (.A(net999),
    .B(net988),
    .Y(_0985_));
 sg13g2_or2_1 _3864_ (.X(_0986_),
    .B(net989),
    .A(net1000));
 sg13g2_o21ai_1 _3865_ (.B1(net981),
    .Y(_0987_),
    .A1(net997),
    .A2(net986));
 sg13g2_inv_1 _3866_ (.Y(_0988_),
    .A(_0987_));
 sg13g2_nor2_1 _3867_ (.A(_0825_),
    .B(_0987_),
    .Y(_0989_));
 sg13g2_o21ai_1 _3868_ (.B1(_0964_),
    .Y(_0990_),
    .A1(_0984_),
    .A2(_0989_));
 sg13g2_nand3_1 _3869_ (.B(_0983_),
    .C(_0990_),
    .A(_0972_),
    .Y(_0991_));
 sg13g2_nor2_1 _3870_ (.A(net921),
    .B(_0991_),
    .Y(_0992_));
 sg13g2_a22oi_1 _3871_ (.Y(_0993_),
    .B1(_0834_),
    .B2(_0987_),
    .A2(_0833_),
    .A1(net980));
 sg13g2_o21ai_1 _3872_ (.B1(_0963_),
    .Y(_0994_),
    .A1(net992),
    .A2(net925));
 sg13g2_nand2_1 _3873_ (.Y(_0995_),
    .A(_0964_),
    .B(_0993_));
 sg13g2_nand3_1 _3874_ (.B(_0994_),
    .C(_0995_),
    .A(_0972_),
    .Y(_0996_));
 sg13g2_nor2_1 _3875_ (.A(net921),
    .B(_0996_),
    .Y(_0997_));
 sg13g2_a21oi_2 _3876_ (.B1(net921),
    .Y(_0998_),
    .A2(_0996_),
    .A1(_0991_));
 sg13g2_nand2b_1 _3877_ (.Y(_0999_),
    .B(_0812_),
    .A_N(_0982_));
 sg13g2_nor2b_1 _3878_ (.A(_0982_),
    .B_N(_0998_),
    .Y(_1000_));
 sg13g2_a21oi_1 _3879_ (.A1(_0012_),
    .A2(net921),
    .Y(_1001_),
    .B1(_0992_));
 sg13g2_nor2b_1 _3880_ (.A(_1000_),
    .B_N(_1001_),
    .Y(_1002_));
 sg13g2_nand2_1 _3881_ (.Y(_1003_),
    .A(net897),
    .B(_1002_));
 sg13g2_xnor2_1 _3882_ (.Y(_0112_),
    .A(net129),
    .B(_1003_));
 sg13g2_nand2b_1 _3883_ (.Y(_1004_),
    .B(net922),
    .A_N(_0013_));
 sg13g2_a221oi_1 _3884_ (.B2(_1004_),
    .C1(_0992_),
    .B1(_0999_),
    .A1(_0812_),
    .Y(_1005_),
    .A2(_0996_));
 sg13g2_nand2_1 _3885_ (.Y(_1006_),
    .A(\bass_pha[1] ),
    .B(_1005_));
 sg13g2_xnor2_1 _3886_ (.Y(_1007_),
    .A(_1556_),
    .B(_1005_));
 sg13g2_nand3_1 _3887_ (.B(_1002_),
    .C(_1007_),
    .A(net129),
    .Y(_1008_));
 sg13g2_a21o_1 _3888_ (.A2(_1002_),
    .A1(net129),
    .B1(_1007_),
    .X(_1009_));
 sg13g2_a21oi_1 _3889_ (.A1(_1008_),
    .A2(_1009_),
    .Y(_1010_),
    .B1(net892));
 sg13g2_a21oi_1 _3890_ (.A1(_1556_),
    .A2(net892),
    .Y(_0113_),
    .B1(_1010_));
 sg13g2_a21oi_2 _3891_ (.B1(_1000_),
    .Y(_1011_),
    .A2(net921),
    .A1(_1557_));
 sg13g2_nor2b_1 _3892_ (.A(_1011_),
    .B_N(\bass_pha[2] ),
    .Y(_1012_));
 sg13g2_xor2_1 _3893_ (.B(_1011_),
    .A(net125),
    .X(_1013_));
 sg13g2_a21oi_1 _3894_ (.A1(_1006_),
    .A2(_1008_),
    .Y(_1014_),
    .B1(_1013_));
 sg13g2_nand3_1 _3895_ (.B(_1008_),
    .C(_1013_),
    .A(_1006_),
    .Y(_1015_));
 sg13g2_nand2_1 _3896_ (.Y(_1016_),
    .A(net897),
    .B(_1015_));
 sg13g2_nand2_1 _3897_ (.Y(_1017_),
    .A(net125),
    .B(net892));
 sg13g2_o21ai_1 _3898_ (.B1(_1017_),
    .Y(_0114_),
    .A1(_1014_),
    .A2(_1016_));
 sg13g2_nand2_1 _3899_ (.Y(_1018_),
    .A(net141),
    .B(net892));
 sg13g2_nand2_1 _3900_ (.Y(_1019_),
    .A(_0982_),
    .B(_0996_));
 sg13g2_a22oi_1 _3901_ (.Y(_1020_),
    .B1(_0992_),
    .B2(_1019_),
    .A2(net921),
    .A1(_1558_));
 sg13g2_nand2b_1 _3902_ (.Y(_1021_),
    .B(net141),
    .A_N(_1020_));
 sg13g2_xnor2_1 _3903_ (.Y(_1022_),
    .A(net141),
    .B(_1020_));
 sg13g2_nor3_1 _3904_ (.A(_1012_),
    .B(_1014_),
    .C(_1022_),
    .Y(_1023_));
 sg13g2_o21ai_1 _3905_ (.B1(_1022_),
    .Y(_1024_),
    .A1(_1012_),
    .A2(_1014_));
 sg13g2_nand2_1 _3906_ (.Y(_1025_),
    .A(net897),
    .B(_1024_));
 sg13g2_o21ai_1 _3907_ (.B1(_1018_),
    .Y(_0115_),
    .A1(_1023_),
    .A2(_1025_));
 sg13g2_a22oi_1 _3908_ (.Y(_1026_),
    .B1(_0991_),
    .B2(_0997_),
    .A2(net921),
    .A1(_1560_));
 sg13g2_nor2_1 _3909_ (.A(_1561_),
    .B(_1026_),
    .Y(_1027_));
 sg13g2_xnor2_1 _3910_ (.Y(_1028_),
    .A(_1561_),
    .B(_1026_));
 sg13g2_a21o_1 _3911_ (.A2(_1024_),
    .A1(_1021_),
    .B1(_1028_),
    .X(_1029_));
 sg13g2_nand3_1 _3912_ (.B(_1024_),
    .C(_1028_),
    .A(_1021_),
    .Y(_1030_));
 sg13g2_a21oi_1 _3913_ (.A1(_1029_),
    .A2(_1030_),
    .Y(_1031_),
    .B1(net892));
 sg13g2_a21oi_1 _3914_ (.A1(_1561_),
    .A2(net892),
    .Y(_0116_),
    .B1(_1031_));
 sg13g2_nor2b_1 _3915_ (.A(_1027_),
    .B_N(_1029_),
    .Y(_1032_));
 sg13g2_and2_1 _3916_ (.A(_0992_),
    .B(_0996_),
    .X(_1033_));
 sg13g2_nor2_2 _3917_ (.A(_0017_),
    .B(_0812_),
    .Y(_1034_));
 sg13g2_nor3_1 _3918_ (.A(\bass_pha[5] ),
    .B(_1033_),
    .C(_1034_),
    .Y(_1035_));
 sg13g2_o21ai_1 _3919_ (.B1(\bass_pha[5] ),
    .Y(_1036_),
    .A1(_1033_),
    .A2(_1034_));
 sg13g2_nor2b_1 _3920_ (.A(_1035_),
    .B_N(_1036_),
    .Y(_1037_));
 sg13g2_xnor2_1 _3921_ (.Y(_1038_),
    .A(_1032_),
    .B(_1037_));
 sg13g2_mux2_1 _3922_ (.A0(net146),
    .A1(_1038_),
    .S(net897),
    .X(_0117_));
 sg13g2_nand2_1 _3923_ (.Y(_1039_),
    .A(net134),
    .B(net892));
 sg13g2_nor2_1 _3924_ (.A(_0018_),
    .B(_0812_),
    .Y(_1040_));
 sg13g2_nor3_1 _3925_ (.A(\bass_pha[6] ),
    .B(_0998_),
    .C(_1040_),
    .Y(_1041_));
 sg13g2_o21ai_1 _3926_ (.B1(\bass_pha[6] ),
    .Y(_1042_),
    .A1(_0998_),
    .A2(_1040_));
 sg13g2_nor2b_1 _3927_ (.A(_1041_),
    .B_N(_1042_),
    .Y(_1043_));
 sg13g2_o21ai_1 _3928_ (.B1(_1036_),
    .Y(_1044_),
    .A1(_1032_),
    .A2(_1035_));
 sg13g2_nand2_1 _3929_ (.Y(_1045_),
    .A(_1043_),
    .B(_1044_));
 sg13g2_xnor2_1 _3930_ (.Y(_1046_),
    .A(_1043_),
    .B(_1044_));
 sg13g2_o21ai_1 _3931_ (.B1(_1039_),
    .Y(_0118_),
    .A1(net892),
    .A2(_1046_));
 sg13g2_a21oi_1 _3932_ (.A1(_0019_),
    .A2(net921),
    .Y(_1047_),
    .B1(_0998_));
 sg13g2_and2_1 _3933_ (.A(\bass_pha[7] ),
    .B(_1047_),
    .X(_1048_));
 sg13g2_xnor2_1 _3934_ (.Y(_1049_),
    .A(\bass_pha[7] ),
    .B(_1047_));
 sg13g2_and3_1 _3935_ (.X(_1050_),
    .A(_1042_),
    .B(_1045_),
    .C(_1049_));
 sg13g2_a21oi_2 _3936_ (.B1(_1049_),
    .Y(_1051_),
    .A2(_1045_),
    .A1(_1042_));
 sg13g2_nor3_1 _3937_ (.A(net895),
    .B(_1050_),
    .C(_1051_),
    .Y(_1052_));
 sg13g2_a21o_1 _3938_ (.A2(net895),
    .A1(net160),
    .B1(_1052_),
    .X(_0119_));
 sg13g2_nand3_1 _3939_ (.B(\bass_pha[8] ),
    .C(net922),
    .A(\kick_osci[8] ),
    .Y(_1053_));
 sg13g2_a21o_1 _3940_ (.A2(net922),
    .A1(\kick_osci[8] ),
    .B1(\bass_pha[8] ),
    .X(_1054_));
 sg13g2_and2_1 _3941_ (.A(_1053_),
    .B(_1054_),
    .X(_1055_));
 sg13g2_o21ai_1 _3942_ (.B1(_1055_),
    .Y(_1056_),
    .A1(_1048_),
    .A2(_1051_));
 sg13g2_or3_1 _3943_ (.A(_1048_),
    .B(_1051_),
    .C(_1055_),
    .X(_1057_));
 sg13g2_and3_1 _3944_ (.X(_1058_),
    .A(net898),
    .B(_1056_),
    .C(_1057_));
 sg13g2_a21o_1 _3945_ (.A2(net896),
    .A1(net153),
    .B1(_1058_),
    .X(_0120_));
 sg13g2_a21oi_2 _3946_ (.B1(_0020_),
    .Y(_1059_),
    .A2(_1056_),
    .A1(_1053_));
 sg13g2_nand3_1 _3947_ (.B(_1053_),
    .C(_1056_),
    .A(_0020_),
    .Y(_1060_));
 sg13g2_nor2b_1 _3948_ (.A(_1059_),
    .B_N(_1060_),
    .Y(_1061_));
 sg13g2_mux2_1 _3949_ (.A0(net95),
    .A1(_1061_),
    .S(net898),
    .X(_0121_));
 sg13g2_and2_1 _3950_ (.A(net898),
    .B(_1059_),
    .X(_1062_));
 sg13g2_nand2_1 _3951_ (.Y(_1063_),
    .A(\bass_pha[10] ),
    .B(_1062_));
 sg13g2_xor2_1 _3952_ (.B(_1062_),
    .A(net147),
    .X(_0122_));
 sg13g2_nand3_1 _3953_ (.B(\bass_pha[11] ),
    .C(_1059_),
    .A(\bass_pha[10] ),
    .Y(_1064_));
 sg13g2_xnor2_1 _3954_ (.Y(_0123_),
    .A(net135),
    .B(_1063_));
 sg13g2_nand2_1 _3955_ (.Y(_1065_),
    .A(net99),
    .B(net896));
 sg13g2_xnor2_1 _3956_ (.Y(_1066_),
    .A(_0021_),
    .B(_1064_));
 sg13g2_o21ai_1 _3957_ (.B1(_1065_),
    .Y(_0124_),
    .A1(net896),
    .A2(_1066_));
 sg13g2_and4_1 _3958_ (.A(\bass_pha[10] ),
    .B(\bass_pha[11] ),
    .C(\bass_pha[12] ),
    .D(_1062_),
    .X(_1067_));
 sg13g2_nand2_1 _3959_ (.Y(_1068_),
    .A(net86),
    .B(_1067_));
 sg13g2_xor2_1 _3960_ (.B(_1067_),
    .A(net86),
    .X(_0125_));
 sg13g2_xnor2_1 _3961_ (.Y(_0126_),
    .A(net78),
    .B(_1068_));
 sg13g2_nor2_1 _3962_ (.A(net113),
    .B(_1068_),
    .Y(_1069_));
 sg13g2_xnor2_1 _3963_ (.Y(_0127_),
    .A(_1566_),
    .B(_1069_));
 sg13g2_nor3_1 _3964_ (.A(net1000),
    .B(net974),
    .C(_0804_),
    .Y(_1070_));
 sg13g2_a21oi_1 _3965_ (.A1(_0809_),
    .A2(_1070_),
    .Y(_1071_),
    .B1(net874));
 sg13g2_a21oi_2 _3966_ (.B1(net863),
    .Y(_1072_),
    .A2(_1071_),
    .A1(net1005));
 sg13g2_inv_1 _3967_ (.Y(_1073_),
    .A(_1072_));
 sg13g2_nand2b_1 _3968_ (.Y(_1074_),
    .B(net280),
    .A_N(net156));
 sg13g2_a21oi_1 _3969_ (.A1(_0764_),
    .A2(_1074_),
    .Y(_1075_),
    .B1(_1072_));
 sg13g2_o21ai_1 _3970_ (.B1(net156),
    .Y(_1076_),
    .A1(_1546_),
    .A2(_1072_));
 sg13g2_nand2b_1 _3971_ (.Y(_0128_),
    .B(net157),
    .A_N(_1075_));
 sg13g2_nand2_1 _3972_ (.Y(_1077_),
    .A(_1547_),
    .B(\bass_vol[1] ));
 sg13g2_xnor2_1 _3973_ (.Y(_1078_),
    .A(\bass_vol[3] ),
    .B(net197));
 sg13g2_nand2_1 _3974_ (.Y(_1079_),
    .A(_1074_),
    .B(_1078_));
 sg13g2_xnor2_1 _3975_ (.Y(_1080_),
    .A(_1074_),
    .B(_1078_));
 sg13g2_a22oi_1 _3976_ (.Y(_0129_),
    .B1(_1080_),
    .B2(net863),
    .A2(_1072_),
    .A1(_1548_));
 sg13g2_xor2_1 _3977_ (.B(\bass_vol[4] ),
    .A(\bass_vol[2] ),
    .X(_1081_));
 sg13g2_and3_1 _3978_ (.X(_1082_),
    .A(_1077_),
    .B(_1079_),
    .C(_1081_));
 sg13g2_a21oi_1 _3979_ (.A1(_1077_),
    .A2(_1079_),
    .Y(_1083_),
    .B1(_1081_));
 sg13g2_or2_1 _3980_ (.X(_1084_),
    .B(_1083_),
    .A(_1082_));
 sg13g2_a22oi_1 _3981_ (.Y(_0130_),
    .B1(_1084_),
    .B2(net863),
    .A2(_1072_),
    .A1(_1546_));
 sg13g2_nand2_1 _3982_ (.Y(_1085_),
    .A(\bass_vol[3] ),
    .B(_1550_));
 sg13g2_xor2_1 _3983_ (.B(\bass_vol[5] ),
    .A(\bass_vol[3] ),
    .X(_1086_));
 sg13g2_a21oi_1 _3984_ (.A1(\bass_vol[2] ),
    .A2(_1549_),
    .Y(_1087_),
    .B1(_1083_));
 sg13g2_xnor2_1 _3985_ (.Y(_1088_),
    .A(_1086_),
    .B(_1087_));
 sg13g2_a22oi_1 _3986_ (.Y(_0131_),
    .B1(_1088_),
    .B2(_0815_),
    .A2(_1072_),
    .A1(_1547_));
 sg13g2_o21ai_1 _3987_ (.B1(_1085_),
    .Y(_1089_),
    .A1(_1086_),
    .A2(_1087_));
 sg13g2_nor2_1 _3988_ (.A(\bass_vol[4] ),
    .B(_1089_),
    .Y(_1090_));
 sg13g2_o21ai_1 _3989_ (.B1(_1073_),
    .Y(_1091_),
    .A1(_0763_),
    .A2(_1090_));
 sg13g2_o21ai_1 _3990_ (.B1(net213),
    .Y(_1092_),
    .A1(_1072_),
    .A2(_1089_));
 sg13g2_nand2_1 _3991_ (.Y(_0132_),
    .A(_1091_),
    .B(_1092_));
 sg13g2_a22oi_1 _3992_ (.Y(_0133_),
    .B1(_1091_),
    .B2(_1550_),
    .A2(_1090_),
    .A1(net863));
 sg13g2_a221oi_1 _3993_ (.B2(net928),
    .C1(_1536_),
    .B1(_0835_),
    .A1(_0774_),
    .Y(_1093_),
    .A2(_0779_));
 sg13g2_o21ai_1 _3994_ (.B1(_0986_),
    .Y(_1094_),
    .A1(_1534_),
    .A2(net927));
 sg13g2_nor2_1 _3995_ (.A(net983),
    .B(_0823_),
    .Y(_1095_));
 sg13g2_nand2_1 _3996_ (.Y(_1096_),
    .A(net938),
    .B(_0977_));
 sg13g2_and2_1 _3997_ (.A(_1094_),
    .B(_1095_),
    .X(_1097_));
 sg13g2_or3_1 _3998_ (.A(net937),
    .B(_1093_),
    .C(_1097_),
    .X(_1098_));
 sg13g2_a21oi_1 _3999_ (.A1(net1001),
    .A2(_0976_),
    .Y(_1099_),
    .B1(_1096_));
 sg13g2_nand2_1 _4000_ (.Y(_1100_),
    .A(_0782_),
    .B(_0833_));
 sg13g2_nor2_1 _4001_ (.A(net994),
    .B(_0823_),
    .Y(_1101_));
 sg13g2_a21oi_1 _4002_ (.A1(net994),
    .A2(net929),
    .Y(_1102_),
    .B1(_1101_));
 sg13g2_nor2b_1 _4003_ (.A(net987),
    .B_N(net1001),
    .Y(_1103_));
 sg13g2_a221oi_1 _4004_ (.B2(_1102_),
    .C1(net938),
    .B1(_1100_),
    .A1(net926),
    .Y(_1104_),
    .A2(_0985_));
 sg13g2_o21ai_1 _4005_ (.B1(net978),
    .Y(_1105_),
    .A1(_1099_),
    .A2(_1104_));
 sg13g2_nand3b_1 _4006_ (.B(net988),
    .C(_0774_),
    .Y(_1106_),
    .A_N(net999));
 sg13g2_nand2_1 _4007_ (.Y(_1107_),
    .A(net985),
    .B(_1106_));
 sg13g2_a21oi_1 _4008_ (.A1(_1534_),
    .A2(_1102_),
    .Y(_1108_),
    .B1(_1107_));
 sg13g2_o21ai_1 _4009_ (.B1(_1094_),
    .Y(_1109_),
    .A1(net1002),
    .A2(_0834_));
 sg13g2_a21oi_1 _4010_ (.A1(net938),
    .A2(_1109_),
    .Y(_1110_),
    .B1(_1108_));
 sg13g2_nor2b_2 _4011_ (.A(net978),
    .B_N(net977),
    .Y(_1111_));
 sg13g2_nand2_1 _4012_ (.Y(_1112_),
    .A(net987),
    .B(_0833_));
 sg13g2_inv_1 _4013_ (.Y(_1113_),
    .A(_1112_));
 sg13g2_a22oi_1 _4014_ (.Y(_1114_),
    .B1(_1113_),
    .B2(net1001),
    .A2(_0835_),
    .A1(net929));
 sg13g2_a21o_1 _4015_ (.A2(_1114_),
    .A1(net982),
    .B1(_1097_),
    .X(_1115_));
 sg13g2_a22oi_1 _4016_ (.Y(_1116_),
    .B1(_1111_),
    .B2(_1115_),
    .A2(_1110_),
    .A1(_0803_));
 sg13g2_nand2_1 _4017_ (.Y(_1117_),
    .A(_1105_),
    .B(_1116_));
 sg13g2_nand2_1 _4018_ (.Y(_1118_),
    .A(net975),
    .B(_1117_));
 sg13g2_nand2b_1 _4019_ (.Y(_1119_),
    .B(_1111_),
    .A_N(_1110_));
 sg13g2_nor2_1 _4020_ (.A(net926),
    .B(_0827_),
    .Y(_1120_));
 sg13g2_a221oi_1 _4021_ (.B2(_0975_),
    .C1(_1535_),
    .B1(_0969_),
    .A1(_0828_),
    .Y(_1121_),
    .A2(_0965_));
 sg13g2_o21ai_1 _4022_ (.B1(_1121_),
    .Y(_1122_),
    .A1(_0788_),
    .A2(_1120_));
 sg13g2_nand2_1 _4023_ (.Y(_1123_),
    .A(_0966_),
    .B(_1096_));
 sg13g2_nand2_2 _4024_ (.Y(_1124_),
    .A(net988),
    .B(_0781_));
 sg13g2_o21ai_1 _4025_ (.B1(_1123_),
    .Y(_1125_),
    .A1(net1001),
    .A2(_1124_));
 sg13g2_o21ai_1 _4026_ (.B1(_0988_),
    .Y(_1126_),
    .A1(net929),
    .A2(_0974_));
 sg13g2_nand3_1 _4027_ (.B(_1125_),
    .C(_1126_),
    .A(_0803_),
    .Y(_1127_));
 sg13g2_nand3_1 _4028_ (.B(_1122_),
    .C(_1127_),
    .A(_1119_),
    .Y(_1128_));
 sg13g2_o21ai_1 _4029_ (.B1(_1118_),
    .Y(_1129_),
    .A1(net975),
    .A2(_1128_));
 sg13g2_o21ai_1 _4030_ (.B1(_1098_),
    .Y(_1130_),
    .A1(\songpos[8] ),
    .A2(_1129_));
 sg13g2_a21oi_1 _4031_ (.A1(_0771_),
    .A2(_0977_),
    .Y(_1131_),
    .B1(_1103_));
 sg13g2_nor2_1 _4032_ (.A(net982),
    .B(_1131_),
    .Y(_1132_));
 sg13g2_nand2_1 _4033_ (.Y(_1133_),
    .A(_1112_),
    .B(_1132_));
 sg13g2_nor2_1 _4034_ (.A(_0773_),
    .B(_0974_),
    .Y(_1134_));
 sg13g2_nand2b_1 _4035_ (.Y(_1135_),
    .B(_1103_),
    .A_N(_0834_));
 sg13g2_nand2_1 _4036_ (.Y(_1136_),
    .A(net982),
    .B(_1135_));
 sg13g2_o21ai_1 _4037_ (.B1(_1133_),
    .Y(_1137_),
    .A1(_1134_),
    .A2(_1136_));
 sg13g2_o21ai_1 _4038_ (.B1(net938),
    .Y(_1138_),
    .A1(net997),
    .A2(_0773_));
 sg13g2_a21oi_1 _4039_ (.A1(net993),
    .A2(_0783_),
    .Y(_1139_),
    .B1(_1138_));
 sg13g2_o21ai_1 _4040_ (.B1(net925),
    .Y(_1140_),
    .A1(net1003),
    .A2(_0775_));
 sg13g2_a221oi_1 _4041_ (.B2(_0825_),
    .C1(_1139_),
    .B1(_0967_),
    .A1(_0818_),
    .Y(_1141_),
    .A2(_0965_));
 sg13g2_a21oi_1 _4042_ (.A1(_1140_),
    .A2(_1141_),
    .Y(_1142_),
    .B1(_0804_));
 sg13g2_o21ai_1 _4043_ (.B1(_0984_),
    .Y(_1143_),
    .A1(_0784_),
    .A2(_1134_));
 sg13g2_o21ai_1 _4044_ (.B1(_0771_),
    .Y(_1144_),
    .A1(_0773_),
    .A2(_0985_));
 sg13g2_nor2_1 _4045_ (.A(_0779_),
    .B(_1144_),
    .Y(_1145_));
 sg13g2_o21ai_1 _4046_ (.B1(net984),
    .Y(_1146_),
    .A1(_1534_),
    .A2(_0771_));
 sg13g2_o21ai_1 _4047_ (.B1(_1143_),
    .Y(_1147_),
    .A1(_1145_),
    .A2(_1146_));
 sg13g2_nor2_1 _4048_ (.A(net993),
    .B(net929),
    .Y(_1148_));
 sg13g2_nor4_1 _4049_ (.A(net926),
    .B(_1096_),
    .C(_1103_),
    .D(_1148_),
    .Y(_1149_));
 sg13g2_a221oi_1 _4050_ (.B2(_0776_),
    .C1(_1149_),
    .B1(_0965_),
    .A1(net925),
    .Y(_1150_),
    .A2(_0827_));
 sg13g2_inv_1 _4051_ (.Y(_1151_),
    .A(_1150_));
 sg13g2_a221oi_1 _4052_ (.B2(_1111_),
    .C1(_1142_),
    .B1(_1150_),
    .A1(net978),
    .Y(_1152_),
    .A2(_1147_));
 sg13g2_nor2_1 _4053_ (.A(net975),
    .B(_1152_),
    .Y(_1153_));
 sg13g2_a21o_1 _4054_ (.A2(_1124_),
    .A1(net929),
    .B1(_1148_),
    .X(_1154_));
 sg13g2_o21ai_1 _4055_ (.B1(net988),
    .Y(_1155_),
    .A1(net1002),
    .A2(net999));
 sg13g2_nand2_1 _4056_ (.Y(_1156_),
    .A(net928),
    .B(_0973_));
 sg13g2_a22oi_1 _4057_ (.Y(_1157_),
    .B1(_1156_),
    .B2(_1132_),
    .A2(_1154_),
    .A1(net982));
 sg13g2_o21ai_1 _4058_ (.B1(net975),
    .Y(_1158_),
    .A1(_1535_),
    .A2(_1157_));
 sg13g2_a221oi_1 _4059_ (.B2(_0803_),
    .C1(_1158_),
    .B1(_1151_),
    .A1(_1111_),
    .Y(_1159_),
    .A2(_1137_));
 sg13g2_nor3_1 _4060_ (.A(\songpos[8] ),
    .B(_1153_),
    .C(_1159_),
    .Y(_1160_));
 sg13g2_a21o_2 _4061_ (.A2(_1137_),
    .A1(\songpos[8] ),
    .B1(_1160_),
    .X(_1161_));
 sg13g2_o21ai_1 _4062_ (.B1(_1536_),
    .Y(_1162_),
    .A1(_1534_),
    .A2(_0834_));
 sg13g2_nor3_1 _4063_ (.A(_1534_),
    .B(net926),
    .C(_0834_),
    .Y(_1163_));
 sg13g2_nor2b_1 _4064_ (.A(net992),
    .B_N(net980),
    .Y(_1164_));
 sg13g2_a21oi_1 _4065_ (.A1(net928),
    .A2(_1164_),
    .Y(_1165_),
    .B1(_0965_));
 sg13g2_o21ai_1 _4066_ (.B1(_1165_),
    .Y(_1166_),
    .A1(net980),
    .A2(_1163_));
 sg13g2_nor3_1 _4067_ (.A(net981),
    .B(_0834_),
    .C(_1163_),
    .Y(_1167_));
 sg13g2_nor2_1 _4068_ (.A(_0833_),
    .B(_1165_),
    .Y(_1168_));
 sg13g2_or2_1 _4069_ (.X(_1169_),
    .B(_1168_),
    .A(_1167_));
 sg13g2_a21oi_1 _4070_ (.A1(net986),
    .A2(_1166_),
    .Y(_1170_),
    .B1(_1169_));
 sg13g2_nand2_1 _4071_ (.Y(_1171_),
    .A(_0767_),
    .B(_0835_));
 sg13g2_a21oi_1 _4072_ (.A1(_0975_),
    .A2(_1171_),
    .Y(_1172_),
    .B1(net983));
 sg13g2_a22oi_1 _4073_ (.Y(_1173_),
    .B1(_0781_),
    .B2(_1534_),
    .A2(_0774_),
    .A1(_0771_));
 sg13g2_o21ai_1 _4074_ (.B1(net983),
    .Y(_1174_),
    .A1(_0783_),
    .A2(_0826_));
 sg13g2_nor2_1 _4075_ (.A(_1173_),
    .B(_1174_),
    .Y(_1175_));
 sg13g2_nor2_1 _4076_ (.A(_1172_),
    .B(_1175_),
    .Y(_1176_));
 sg13g2_nor3_1 _4077_ (.A(net927),
    .B(_0833_),
    .C(_1155_),
    .Y(_1177_));
 sg13g2_or2_1 _4078_ (.X(_1178_),
    .B(_1177_),
    .A(net984));
 sg13g2_a21oi_1 _4079_ (.A1(_0771_),
    .A2(_0978_),
    .Y(_1179_),
    .B1(_1178_));
 sg13g2_nand3_1 _4080_ (.B(_1100_),
    .C(_1106_),
    .A(net983),
    .Y(_1180_));
 sg13g2_a21oi_1 _4081_ (.A1(net927),
    .A2(_0985_),
    .Y(_1181_),
    .B1(_1180_));
 sg13g2_nor2_2 _4082_ (.A(_1179_),
    .B(_1181_),
    .Y(_1182_));
 sg13g2_a221oi_1 _4083_ (.B2(_1111_),
    .C1(net974),
    .B1(_1182_),
    .A1(net978),
    .Y(_1183_),
    .A2(_1176_));
 sg13g2_o21ai_1 _4084_ (.B1(_1183_),
    .Y(_1184_),
    .A1(_0804_),
    .A2(_1170_));
 sg13g2_nand2_1 _4085_ (.Y(_1185_),
    .A(_0803_),
    .B(_1182_));
 sg13g2_o21ai_1 _4086_ (.B1(net925),
    .Y(_1186_),
    .A1(net928),
    .A2(_0773_));
 sg13g2_a21oi_1 _4087_ (.A1(_0829_),
    .A2(_0967_),
    .Y(_1187_),
    .B1(_1535_));
 sg13g2_nand2_1 _4088_ (.Y(_1188_),
    .A(_1186_),
    .B(_1187_));
 sg13g2_nand2_1 _4089_ (.Y(_1189_),
    .A(_0776_),
    .B(net925));
 sg13g2_nand2_1 _4090_ (.Y(_1190_),
    .A(net997),
    .B(net938));
 sg13g2_nand2_1 _4091_ (.Y(_1191_),
    .A(net938),
    .B(_1113_));
 sg13g2_nand3_1 _4092_ (.B(_1189_),
    .C(_1191_),
    .A(_1111_),
    .Y(_1192_));
 sg13g2_nand4_1 _4093_ (.B(_1185_),
    .C(_1188_),
    .A(net975),
    .Y(_1193_),
    .D(_1192_));
 sg13g2_nand3_1 _4094_ (.B(_1184_),
    .C(_1193_),
    .A(net937),
    .Y(_1194_));
 sg13g2_nand2_1 _4095_ (.Y(_1195_),
    .A(net925),
    .B(_0826_));
 sg13g2_a21o_1 _4096_ (.A2(_0833_),
    .A1(net1001),
    .B1(_1195_),
    .X(_1196_));
 sg13g2_nand3_1 _4097_ (.B(_1191_),
    .C(_1196_),
    .A(\songpos[8] ),
    .Y(_1197_));
 sg13g2_nand2_2 _4098_ (.Y(_1198_),
    .A(_1194_),
    .B(_1197_));
 sg13g2_nor2b_1 _4099_ (.A(_1198_),
    .B_N(_1161_),
    .Y(_1199_));
 sg13g2_nor3_1 _4100_ (.A(net894),
    .B(_1130_),
    .C(_1199_),
    .Y(_1200_));
 sg13g2_xor2_1 _4101_ (.B(_1200_),
    .A(net108),
    .X(_0134_));
 sg13g2_nand2_1 _4102_ (.Y(_1201_),
    .A(net82),
    .B(net894));
 sg13g2_nor2_1 _4103_ (.A(\sqr_pha[0] ),
    .B(_1199_),
    .Y(_1202_));
 sg13g2_nor3_2 _4104_ (.A(_0010_),
    .B(_1130_),
    .C(_1202_),
    .Y(_1203_));
 sg13g2_o21ai_1 _4105_ (.B1(_0010_),
    .Y(_1204_),
    .A1(_1130_),
    .A2(_1202_));
 sg13g2_nand2_1 _4106_ (.Y(_1205_),
    .A(net898),
    .B(_1204_));
 sg13g2_o21ai_1 _4107_ (.B1(_1201_),
    .Y(_0135_),
    .A1(_1203_),
    .A2(_1205_));
 sg13g2_a21oi_1 _4108_ (.A1(_1130_),
    .A2(_1161_),
    .Y(_1206_),
    .B1(_1199_));
 sg13g2_nor2b_1 _4109_ (.A(_1206_),
    .B_N(\sqr_pha[2] ),
    .Y(_1207_));
 sg13g2_xnor2_1 _4110_ (.Y(_1208_),
    .A(net120),
    .B(_1206_));
 sg13g2_and2_1 _4111_ (.A(_1203_),
    .B(_1208_),
    .X(_1209_));
 sg13g2_o21ai_1 _4112_ (.B1(net897),
    .Y(_1210_),
    .A1(_1203_),
    .A2(_1208_));
 sg13g2_nand2_1 _4113_ (.Y(_1211_),
    .A(net120),
    .B(net894));
 sg13g2_o21ai_1 _4114_ (.B1(_1211_),
    .Y(_0136_),
    .A1(_1209_),
    .A2(_1210_));
 sg13g2_nand2b_1 _4115_ (.Y(_1212_),
    .B(_1198_),
    .A_N(_1161_));
 sg13g2_xnor2_1 _4116_ (.Y(_1213_),
    .A(_1130_),
    .B(_1212_));
 sg13g2_nand2_1 _4117_ (.Y(_1214_),
    .A(\sqr_pha[3] ),
    .B(_1213_));
 sg13g2_xor2_1 _4118_ (.B(_1213_),
    .A(\sqr_pha[3] ),
    .X(_1215_));
 sg13g2_o21ai_1 _4119_ (.B1(_1215_),
    .Y(_1216_),
    .A1(_1207_),
    .A2(_1209_));
 sg13g2_nor3_1 _4120_ (.A(_1207_),
    .B(_1209_),
    .C(_1215_),
    .Y(_1217_));
 sg13g2_and2_1 _4121_ (.A(net237),
    .B(net893),
    .X(_1218_));
 sg13g2_nor2_1 _4122_ (.A(net893),
    .B(_1217_),
    .Y(_1219_));
 sg13g2_a21o_1 _4123_ (.A2(_1219_),
    .A1(_1216_),
    .B1(_1218_),
    .X(_0137_));
 sg13g2_a21o_1 _4124_ (.A2(_1198_),
    .A1(_1161_),
    .B1(_1130_),
    .X(_1220_));
 sg13g2_or2_1 _4125_ (.X(_1221_),
    .B(_1220_),
    .A(_1551_));
 sg13g2_xnor2_1 _4126_ (.Y(_1222_),
    .A(_1551_),
    .B(_1220_));
 sg13g2_a21o_1 _4127_ (.A2(_1216_),
    .A1(_1214_),
    .B1(_1222_),
    .X(_1223_));
 sg13g2_nand3_1 _4128_ (.B(_1216_),
    .C(_1222_),
    .A(_1214_),
    .Y(_1224_));
 sg13g2_a21oi_1 _4129_ (.A1(_1223_),
    .A2(_1224_),
    .Y(_1225_),
    .B1(net893));
 sg13g2_a21oi_1 _4130_ (.A1(_1551_),
    .A2(net893),
    .Y(_0138_),
    .B1(_1225_));
 sg13g2_nand2b_1 _4131_ (.Y(_1226_),
    .B(_1161_),
    .A_N(_1130_));
 sg13g2_nand2_1 _4132_ (.Y(_1227_),
    .A(_1198_),
    .B(_1226_));
 sg13g2_nor2_1 _4133_ (.A(_0011_),
    .B(_1227_),
    .Y(_1228_));
 sg13g2_xnor2_1 _4134_ (.Y(_1229_),
    .A(_0011_),
    .B(_1227_));
 sg13g2_nand3_1 _4135_ (.B(_1223_),
    .C(_1229_),
    .A(_1221_),
    .Y(_1230_));
 sg13g2_a21oi_1 _4136_ (.A1(_1221_),
    .A2(_1223_),
    .Y(_1231_),
    .B1(_1229_));
 sg13g2_nand3b_1 _4137_ (.B(net897),
    .C(_1230_),
    .Y(_1232_),
    .A_N(_1231_));
 sg13g2_o21ai_1 _4138_ (.B1(_1232_),
    .Y(_0139_),
    .A1(_1552_),
    .A2(net897));
 sg13g2_nor2b_2 _4139_ (.A(_1226_),
    .B_N(_1198_),
    .Y(_1233_));
 sg13g2_nand2b_1 _4140_ (.Y(_1234_),
    .B(\sqr_pha[6] ),
    .A_N(_1233_));
 sg13g2_xnor2_1 _4141_ (.Y(_1235_),
    .A(\sqr_pha[6] ),
    .B(_1233_));
 sg13g2_o21ai_1 _4142_ (.B1(_1235_),
    .Y(_1236_),
    .A1(_1228_),
    .A2(_1231_));
 sg13g2_or3_1 _4143_ (.A(_1228_),
    .B(_1231_),
    .C(_1235_),
    .X(_1237_));
 sg13g2_a21oi_1 _4144_ (.A1(_1236_),
    .A2(_1237_),
    .Y(_1238_),
    .B1(net893));
 sg13g2_a21oi_1 _4145_ (.A1(_1553_),
    .A2(net893),
    .Y(_0140_),
    .B1(_1238_));
 sg13g2_and2_1 _4146_ (.A(\sqr_pha[7] ),
    .B(_1233_),
    .X(_1239_));
 sg13g2_xnor2_1 _4147_ (.Y(_1240_),
    .A(\sqr_pha[7] ),
    .B(_1233_));
 sg13g2_and3_1 _4148_ (.X(_1241_),
    .A(_1234_),
    .B(_1236_),
    .C(_1240_));
 sg13g2_a21oi_1 _4149_ (.A1(_1234_),
    .A2(_1236_),
    .Y(_1242_),
    .B1(_1240_));
 sg13g2_nor3_1 _4150_ (.A(net893),
    .B(_1241_),
    .C(_1242_),
    .Y(_1243_));
 sg13g2_a21o_1 _4151_ (.A2(net893),
    .A1(net172),
    .B1(_1243_),
    .X(_0141_));
 sg13g2_o21ai_1 _4152_ (.B1(net897),
    .Y(_1244_),
    .A1(_1239_),
    .A2(_1242_));
 sg13g2_nor2_2 _4153_ (.A(_1554_),
    .B(_1244_),
    .Y(_1245_));
 sg13g2_xnor2_1 _4154_ (.Y(_0142_),
    .A(net94),
    .B(_1244_));
 sg13g2_xor2_1 _4155_ (.B(_1245_),
    .A(net115),
    .X(_0143_));
 sg13g2_a21oi_1 _4156_ (.A1(net115),
    .A2(_1245_),
    .Y(_1246_),
    .B1(net119));
 sg13g2_and2_1 _4157_ (.A(net115),
    .B(net119),
    .X(_1247_));
 sg13g2_a21oi_1 _4158_ (.A1(_1245_),
    .A2(_1247_),
    .Y(_0144_),
    .B1(_1246_));
 sg13g2_a21oi_1 _4159_ (.A1(_1245_),
    .A2(_1247_),
    .Y(_1248_),
    .B1(net111));
 sg13g2_nand3_1 _4160_ (.B(_1245_),
    .C(_1247_),
    .A(net111),
    .Y(_1249_));
 sg13g2_nor2b_1 _4161_ (.A(net112),
    .B_N(_1249_),
    .Y(_0145_));
 sg13g2_xnor2_1 _4162_ (.Y(_0146_),
    .A(net104),
    .B(_1249_));
 sg13g2_and2_1 _4163_ (.A(net989),
    .B(_0775_),
    .X(_1250_));
 sg13g2_nor3_1 _4164_ (.A(net1004),
    .B(_0978_),
    .C(_1250_),
    .Y(_1251_));
 sg13g2_nor3_1 _4165_ (.A(net990),
    .B(net985),
    .C(_0774_),
    .Y(_1252_));
 sg13g2_a21oi_1 _4166_ (.A1(_0790_),
    .A2(_1251_),
    .Y(_1253_),
    .B1(_1252_));
 sg13g2_o21ai_1 _4167_ (.B1(_1124_),
    .Y(_1254_),
    .A1(_0823_),
    .A2(_0828_));
 sg13g2_nor2_1 _4168_ (.A(net989),
    .B(_0781_),
    .Y(_1255_));
 sg13g2_nor3_1 _4169_ (.A(_0790_),
    .B(_1254_),
    .C(_1255_),
    .Y(_1256_));
 sg13g2_nor3_1 _4170_ (.A(_0783_),
    .B(_0791_),
    .C(_0833_),
    .Y(_1257_));
 sg13g2_o21ai_1 _4171_ (.B1(_0791_),
    .Y(_1258_),
    .A1(net1004),
    .A2(_0986_));
 sg13g2_nor3_1 _4172_ (.A(net1002),
    .B(_0973_),
    .C(_0978_),
    .Y(_1259_));
 sg13g2_o21ai_1 _4173_ (.B1(_1258_),
    .Y(_1260_),
    .A1(_0791_),
    .A2(_1259_));
 sg13g2_nor3_1 _4174_ (.A(_0796_),
    .B(_1256_),
    .C(_1257_),
    .Y(_1261_));
 sg13g2_a21oi_1 _4175_ (.A1(_0796_),
    .A2(_1253_),
    .Y(_1262_),
    .B1(_1261_));
 sg13g2_nand2_1 _4176_ (.Y(_1263_),
    .A(_0801_),
    .B(_1262_));
 sg13g2_nand2b_1 _4177_ (.Y(_1264_),
    .B(_1253_),
    .A_N(_0796_));
 sg13g2_nand2_1 _4178_ (.Y(_1265_),
    .A(_0796_),
    .B(_1260_));
 sg13g2_nand3_1 _4179_ (.B(_1264_),
    .C(_1265_),
    .A(_0800_),
    .Y(_1266_));
 sg13g2_nand3_1 _4180_ (.B(_1263_),
    .C(_1266_),
    .A(_0794_),
    .Y(_1267_));
 sg13g2_o21ai_1 _4181_ (.B1(_0790_),
    .Y(_1268_),
    .A1(net989),
    .A2(_0774_));
 sg13g2_o21ai_1 _4182_ (.B1(_0824_),
    .Y(_1269_),
    .A1(_0835_),
    .A2(_1250_));
 sg13g2_o21ai_1 _4183_ (.B1(_0836_),
    .Y(_1270_),
    .A1(_0775_),
    .A2(_0791_));
 sg13g2_nand2b_1 _4184_ (.Y(_1271_),
    .B(_1269_),
    .A_N(_1270_));
 sg13g2_nand3_1 _4185_ (.B(_1258_),
    .C(_1268_),
    .A(_0800_),
    .Y(_1272_));
 sg13g2_o21ai_1 _4186_ (.B1(_1272_),
    .Y(_1273_),
    .A1(_0800_),
    .A2(_1271_));
 sg13g2_nor2_1 _4187_ (.A(_0794_),
    .B(_1273_),
    .Y(_1274_));
 sg13g2_nor2_1 _4188_ (.A(_0808_),
    .B(_1274_),
    .Y(_1275_));
 sg13g2_o21ai_1 _4189_ (.B1(net877),
    .Y(_1276_),
    .A1(_0809_),
    .A2(_1260_));
 sg13g2_a21oi_2 _4190_ (.B1(_1276_),
    .Y(_1277_),
    .A2(_1275_),
    .A1(_1267_));
 sg13g2_nor2_2 _4191_ (.A(_0815_),
    .B(_1277_),
    .Y(_1278_));
 sg13g2_o21ai_1 _4192_ (.B1(\sqr_vol[3] ),
    .Y(_1279_),
    .A1(net863),
    .A2(_1277_));
 sg13g2_nand2b_1 _4193_ (.Y(_1280_),
    .B(net230),
    .A_N(\sqr_vol[0] ));
 sg13g2_a21oi_1 _4194_ (.A1(_0764_),
    .A2(_1280_),
    .Y(_1281_),
    .B1(_1278_));
 sg13g2_nand2_1 _4195_ (.Y(_1282_),
    .A(_0763_),
    .B(_1277_));
 sg13g2_a21o_1 _4196_ (.A2(_1279_),
    .A1(net151),
    .B1(_1281_),
    .X(_0147_));
 sg13g2_nand2b_1 _4197_ (.Y(_1283_),
    .B(\sqr_vol[1] ),
    .A_N(\sqr_vol[4] ));
 sg13g2_xnor2_1 _4198_ (.Y(_1284_),
    .A(\sqr_vol[1] ),
    .B(\sqr_vol[4] ));
 sg13g2_nand2_1 _4199_ (.Y(_1285_),
    .A(_1280_),
    .B(_1284_));
 sg13g2_xnor2_1 _4200_ (.Y(_1286_),
    .A(_1280_),
    .B(_1284_));
 sg13g2_a22oi_1 _4201_ (.Y(_0148_),
    .B1(_1286_),
    .B2(net863),
    .A2(_1278_),
    .A1(_1544_));
 sg13g2_nor2_1 _4202_ (.A(\sqr_vol[5] ),
    .B(_1545_),
    .Y(_1287_));
 sg13g2_xor2_1 _4203_ (.B(\sqr_vol[2] ),
    .A(\sqr_vol[5] ),
    .X(_1288_));
 sg13g2_and3_1 _4204_ (.X(_1289_),
    .A(_1283_),
    .B(_1285_),
    .C(_1288_));
 sg13g2_a21oi_1 _4205_ (.A1(_1283_),
    .A2(_1285_),
    .Y(_1290_),
    .B1(_1288_));
 sg13g2_or2_1 _4206_ (.X(_1291_),
    .B(_1290_),
    .A(_1289_));
 sg13g2_a22oi_1 _4207_ (.Y(_0149_),
    .B1(_1291_),
    .B2(net863),
    .A2(_1278_),
    .A1(_1545_));
 sg13g2_nor3_1 _4208_ (.A(_1278_),
    .B(_1287_),
    .C(_1290_),
    .Y(_1292_));
 sg13g2_xnor2_1 _4209_ (.Y(_1293_),
    .A(net230),
    .B(_1292_));
 sg13g2_nand2_1 _4210_ (.Y(_0150_),
    .A(_1282_),
    .B(_1293_));
 sg13g2_nand2_1 _4211_ (.Y(_1294_),
    .A(net219),
    .B(_1292_));
 sg13g2_nor2_1 _4212_ (.A(\sqr_vol[4] ),
    .B(_1294_),
    .Y(_1295_));
 sg13g2_xor2_1 _4213_ (.B(_1294_),
    .A(\sqr_vol[4] ),
    .X(_1296_));
 sg13g2_nand2_1 _4214_ (.Y(_0151_),
    .A(_1282_),
    .B(net220));
 sg13g2_xnor2_1 _4215_ (.Y(_1297_),
    .A(net240),
    .B(_1295_));
 sg13g2_nand2_1 _4216_ (.Y(_0152_),
    .A(_1282_),
    .B(net241));
 sg13g2_nor2_1 _4217_ (.A(_1525_),
    .B(net778),
    .Y(_1298_));
 sg13g2_xnor2_1 _4218_ (.Y(_1299_),
    .A(net166),
    .B(_1298_));
 sg13g2_nor2_1 _4219_ (.A(_0852_),
    .B(net167),
    .Y(_0153_));
 sg13g2_nand2_1 _4220_ (.Y(_1300_),
    .A(net138),
    .B(net778));
 sg13g2_nor2_2 _4221_ (.A(_1525_),
    .B(\kick_osci[0] ),
    .Y(_1301_));
 sg13g2_nand2_1 _4222_ (.Y(_1302_),
    .A(\kick_osci[1] ),
    .B(_1559_));
 sg13g2_xor2_1 _4223_ (.B(\kick_osci[4] ),
    .A(net138),
    .X(_1303_));
 sg13g2_xnor2_1 _4224_ (.Y(_1304_),
    .A(_1301_),
    .B(_1303_));
 sg13g2_o21ai_1 _4225_ (.B1(_1300_),
    .Y(_0154_),
    .A1(_0816_),
    .A2(_1304_));
 sg13g2_nand2_1 _4226_ (.Y(_1305_),
    .A(net140),
    .B(net778));
 sg13g2_o21ai_1 _4227_ (.B1(_1302_),
    .Y(_1306_),
    .A1(_1301_),
    .A2(_1303_));
 sg13g2_nor2b_1 _4228_ (.A(\kick_osci[5] ),
    .B_N(\kick_osci[2] ),
    .Y(_1307_));
 sg13g2_xnor2_1 _4229_ (.Y(_1308_),
    .A(net140),
    .B(\kick_osci[5] ));
 sg13g2_xnor2_1 _4230_ (.Y(_1309_),
    .A(_1306_),
    .B(_1308_));
 sg13g2_o21ai_1 _4231_ (.B1(_1305_),
    .Y(_0155_),
    .A1(_0816_),
    .A2(_1309_));
 sg13g2_nand2_1 _4232_ (.Y(_1310_),
    .A(net171),
    .B(net778));
 sg13g2_a21oi_1 _4233_ (.A1(_1306_),
    .A2(_1308_),
    .Y(_1311_),
    .B1(_1307_));
 sg13g2_xor2_1 _4234_ (.B(\kick_osci[6] ),
    .A(\kick_osci[3] ),
    .X(_1312_));
 sg13g2_nor2_1 _4235_ (.A(_1311_),
    .B(_1312_),
    .Y(_1313_));
 sg13g2_a21o_1 _4236_ (.A2(_1312_),
    .A1(_1311_),
    .B1(_0816_),
    .X(_1314_));
 sg13g2_o21ai_1 _4237_ (.B1(_1310_),
    .Y(_0156_),
    .A1(_1313_),
    .A2(_1314_));
 sg13g2_xnor2_1 _4238_ (.Y(_1315_),
    .A(\kick_osci[4] ),
    .B(\kick_osci[7] ));
 sg13g2_a21oi_2 _4239_ (.B1(_1313_),
    .Y(_1316_),
    .A2(_1562_),
    .A1(\kick_osci[3] ));
 sg13g2_nor2b_1 _4240_ (.A(_1316_),
    .B_N(_1315_),
    .Y(_1317_));
 sg13g2_xnor2_1 _4241_ (.Y(_1318_),
    .A(_1315_),
    .B(_1316_));
 sg13g2_a21oi_1 _4242_ (.A1(_0764_),
    .A2(_1318_),
    .Y(_1319_),
    .B1(net778));
 sg13g2_a21oi_1 _4243_ (.A1(_1559_),
    .A2(net779),
    .Y(_0157_),
    .B1(_1319_));
 sg13g2_nand2_1 _4244_ (.Y(_1320_),
    .A(net164),
    .B(net778));
 sg13g2_nor2b_1 _4245_ (.A(\kick_osci[5] ),
    .B_N(\kick_osci[8] ),
    .Y(_1321_));
 sg13g2_nand2b_1 _4246_ (.Y(_1322_),
    .B(\kick_osci[5] ),
    .A_N(\kick_osci[8] ));
 sg13g2_nand2b_1 _4247_ (.Y(_1323_),
    .B(_1322_),
    .A_N(_1321_));
 sg13g2_a21oi_1 _4248_ (.A1(\kick_osci[4] ),
    .A2(_1563_),
    .Y(_1324_),
    .B1(_1317_));
 sg13g2_xnor2_1 _4249_ (.Y(_1325_),
    .A(_1323_),
    .B(_1324_));
 sg13g2_o21ai_1 _4250_ (.B1(_1320_),
    .Y(_0158_),
    .A1(_0816_),
    .A2(_1325_));
 sg13g2_o21ai_1 _4251_ (.B1(_1322_),
    .Y(_1326_),
    .A1(_1321_),
    .A2(_1324_));
 sg13g2_nor3_2 _4252_ (.A(net271),
    .B(net778),
    .C(_1326_),
    .Y(_1327_));
 sg13g2_o21ai_1 _4253_ (.B1(net271),
    .Y(_1328_),
    .A1(net778),
    .A2(_1326_));
 sg13g2_nor2b_1 _4254_ (.A(_1327_),
    .B_N(_1328_),
    .Y(_1329_));
 sg13g2_nor2_1 _4255_ (.A(_0852_),
    .B(_1329_),
    .Y(_0159_));
 sg13g2_nand2_1 _4256_ (.Y(_1330_),
    .A(_1563_),
    .B(_1327_));
 sg13g2_a21oi_1 _4257_ (.A1(_1563_),
    .A2(_1327_),
    .Y(_1331_),
    .B1(_0852_));
 sg13g2_o21ai_1 _4258_ (.B1(_1331_),
    .Y(_0160_),
    .A1(_1563_),
    .A2(_1327_));
 sg13g2_a21o_1 _4259_ (.A2(_1330_),
    .A1(net215),
    .B1(_0852_),
    .X(_0161_));
 sg13g2_xnor2_1 _4260_ (.Y(_1332_),
    .A(net974),
    .B(net977));
 sg13g2_a21o_1 _4261_ (.A2(_1180_),
    .A1(_1178_),
    .B1(_1332_),
    .X(_1333_));
 sg13g2_nor2_1 _4262_ (.A(net995),
    .B(_0435_),
    .Y(_1334_));
 sg13g2_o21ai_1 _4263_ (.B1(_1334_),
    .Y(_1335_),
    .A1(_0779_),
    .A2(net925));
 sg13g2_a21oi_2 _4264_ (.B1(net978),
    .Y(_1336_),
    .A2(_1335_),
    .A1(_1333_));
 sg13g2_nand2b_1 _4265_ (.Y(_1337_),
    .B(_0835_),
    .A_N(_0767_));
 sg13g2_nand2b_1 _4266_ (.Y(_1338_),
    .B(_1337_),
    .A_N(_1162_));
 sg13g2_a221oi_1 _4267_ (.B2(_0825_),
    .C1(net938),
    .B1(_0782_),
    .A1(net987),
    .Y(_1339_),
    .A2(net926));
 sg13g2_nor2_1 _4268_ (.A(net974),
    .B(_1339_),
    .Y(_1340_));
 sg13g2_o21ai_1 _4269_ (.B1(_0967_),
    .Y(_1341_),
    .A1(net992),
    .A2(net928));
 sg13g2_and2_1 _4270_ (.A(_1189_),
    .B(_1341_),
    .X(_1342_));
 sg13g2_a221oi_1 _4271_ (.B2(net974),
    .C1(_1535_),
    .B1(_1342_),
    .A1(_1338_),
    .Y(_1343_),
    .A2(_1340_));
 sg13g2_a21oi_1 _4272_ (.A1(_0805_),
    .A2(_1166_),
    .Y(_1344_),
    .B1(\songpos[8] ));
 sg13g2_nand2b_1 _4273_ (.Y(_1345_),
    .B(_1344_),
    .A_N(_1343_));
 sg13g2_and3_1 _4274_ (.X(_1346_),
    .A(\songpos[8] ),
    .B(_1112_),
    .C(_1195_));
 sg13g2_inv_1 _4275_ (.Y(_1347_),
    .A(_1346_));
 sg13g2_o21ai_1 _4276_ (.B1(_1347_),
    .Y(_1348_),
    .A1(_1336_),
    .A2(_1345_));
 sg13g2_or2_1 _4277_ (.X(_1349_),
    .B(_1348_),
    .A(\sqr_pha[10] ));
 sg13g2_nor2_1 _4278_ (.A(_0972_),
    .B(_1166_),
    .Y(_1350_));
 sg13g2_o21ai_1 _4279_ (.B1(\sqr_pha[11] ),
    .Y(_1351_),
    .A1(_0972_),
    .A2(_1166_));
 sg13g2_a21oi_1 _4280_ (.A1(_1555_),
    .A2(_1348_),
    .Y(_1352_),
    .B1(_1351_));
 sg13g2_a22oi_1 _4281_ (.Y(_1353_),
    .B1(_1352_),
    .B2(_1349_),
    .A2(_1350_),
    .A1(_1247_));
 sg13g2_nand2b_1 _4282_ (.Y(_1354_),
    .B(\sqr_vol[0] ),
    .A_N(net783));
 sg13g2_nand2_1 _4283_ (.Y(_1355_),
    .A(_0775_),
    .B(_0787_));
 sg13g2_a21oi_1 _4284_ (.A1(_0977_),
    .A2(_1190_),
    .Y(_1356_),
    .B1(_0964_));
 sg13g2_a221oi_1 _4285_ (.B2(_1355_),
    .C1(_1356_),
    .B1(_0964_),
    .A1(net937),
    .Y(_1357_),
    .A2(_0805_));
 sg13g2_nor2_1 _4286_ (.A(net983),
    .B(_0781_),
    .Y(_1358_));
 sg13g2_a21oi_1 _4287_ (.A1(_0775_),
    .A2(net925),
    .Y(_1359_),
    .B1(_1358_));
 sg13g2_a21oi_1 _4288_ (.A1(_0804_),
    .A2(_1359_),
    .Y(_1360_),
    .B1(net974));
 sg13g2_or2_1 _4289_ (.X(_1361_),
    .B(_0987_),
    .A(_0779_));
 sg13g2_nand3_1 _4290_ (.B(_1190_),
    .C(_1361_),
    .A(_0963_),
    .Y(_1362_));
 sg13g2_or2_1 _4291_ (.X(_1363_),
    .B(_1359_),
    .A(_0963_));
 sg13g2_o21ai_1 _4292_ (.B1(_1363_),
    .Y(_1364_),
    .A1(_1360_),
    .A2(_1362_));
 sg13g2_mux4_1 _4293_ (.S0(_1364_),
    .A0(_1569_),
    .A1(_1564_),
    .A2(_1568_),
    .A3(_1565_),
    .S1(_1357_),
    .X(_1365_));
 sg13g2_nand3_1 _4294_ (.B(_0812_),
    .C(_1365_),
    .A(\bass_vol[0] ),
    .Y(_1366_));
 sg13g2_o21ai_1 _4295_ (.B1(_1366_),
    .Y(_1367_),
    .A1(_1566_),
    .A2(_0812_));
 sg13g2_nor2_1 _4296_ (.A(\audio_sample_lpf[0] ),
    .B(_1367_),
    .Y(_1368_));
 sg13g2_xor2_1 _4297_ (.B(_1367_),
    .A(\audio_sample_lpf[0] ),
    .X(_1369_));
 sg13g2_nor2_1 _4298_ (.A(_1354_),
    .B(_1369_),
    .Y(_1370_));
 sg13g2_xnor2_1 _4299_ (.Y(_1371_),
    .A(_1354_),
    .B(_1369_));
 sg13g2_nor2_1 _4300_ (.A(\audio_sample_lpf[3] ),
    .B(_1371_),
    .Y(_1372_));
 sg13g2_xnor2_1 _4301_ (.Y(_1373_),
    .A(\audio_sample_lpf[3] ),
    .B(_1371_));
 sg13g2_nand2_1 _4302_ (.Y(_1374_),
    .A(net190),
    .B(net882));
 sg13g2_o21ai_1 _4303_ (.B1(_1374_),
    .Y(_0162_),
    .A1(net882),
    .A2(_1373_));
 sg13g2_nor2_1 _4304_ (.A(_1370_),
    .B(_1372_),
    .Y(_1375_));
 sg13g2_nand2_1 _4305_ (.Y(_1376_),
    .A(_0024_),
    .B(net923));
 sg13g2_and2_1 _4306_ (.A(\bass_vol[1] ),
    .B(_1365_),
    .X(_1377_));
 sg13g2_o21ai_1 _4307_ (.B1(_1376_),
    .Y(_1378_),
    .A1(net923),
    .A2(_1377_));
 sg13g2_nor3_1 _4308_ (.A(_1544_),
    .B(net783),
    .C(_1378_),
    .Y(_1379_));
 sg13g2_or3_1 _4309_ (.A(_1544_),
    .B(net783),
    .C(_1378_),
    .X(_1380_));
 sg13g2_o21ai_1 _4310_ (.B1(_1378_),
    .Y(_1381_),
    .A1(_1544_),
    .A2(net783));
 sg13g2_and3_1 _4311_ (.X(_1382_),
    .A(\audio_sample_lpf[1] ),
    .B(_1380_),
    .C(_1381_));
 sg13g2_a21oi_1 _4312_ (.A1(_1380_),
    .A2(_1381_),
    .Y(_1383_),
    .B1(\audio_sample_lpf[1] ));
 sg13g2_nor3_1 _4313_ (.A(_1368_),
    .B(_1382_),
    .C(_1383_),
    .Y(_1384_));
 sg13g2_or3_1 _4314_ (.A(_1368_),
    .B(_1382_),
    .C(_1383_),
    .X(_1385_));
 sg13g2_o21ai_1 _4315_ (.B1(_1368_),
    .Y(_1386_),
    .A1(_1382_),
    .A2(_1383_));
 sg13g2_and3_1 _4316_ (.X(_1387_),
    .A(_0026_),
    .B(_1385_),
    .C(_1386_));
 sg13g2_a21oi_1 _4317_ (.A1(_1385_),
    .A2(_1386_),
    .Y(_1388_),
    .B1(_0026_));
 sg13g2_nor3_2 _4318_ (.A(_1375_),
    .B(_1387_),
    .C(_1388_),
    .Y(_1389_));
 sg13g2_o21ai_1 _4319_ (.B1(_1375_),
    .Y(_1390_),
    .A1(_1387_),
    .A2(_1388_));
 sg13g2_nand2_1 _4320_ (.Y(_1391_),
    .A(net211),
    .B(net882));
 sg13g2_nand2_1 _4321_ (.Y(_1392_),
    .A(_0811_),
    .B(_1390_));
 sg13g2_o21ai_1 _4322_ (.B1(_1391_),
    .Y(_0163_),
    .A1(_1389_),
    .A2(_1392_));
 sg13g2_a21oi_1 _4323_ (.A1(_0026_),
    .A2(_1386_),
    .Y(_1393_),
    .B1(_1384_));
 sg13g2_a21oi_2 _4324_ (.B1(_1379_),
    .Y(_1394_),
    .A2(_1381_),
    .A1(\audio_sample_lpf[1] ));
 sg13g2_and2_1 _4325_ (.A(\bass_vol[2] ),
    .B(_1365_),
    .X(_1395_));
 sg13g2_o21ai_1 _4326_ (.B1(_1376_),
    .Y(_1396_),
    .A1(net923),
    .A2(_1395_));
 sg13g2_or3_2 _4327_ (.A(_1545_),
    .B(_1353_),
    .C(_1396_),
    .X(_1397_));
 sg13g2_o21ai_1 _4328_ (.B1(_1396_),
    .Y(_1398_),
    .A1(_1545_),
    .A2(net783));
 sg13g2_and3_1 _4329_ (.X(_1399_),
    .A(\audio_sample_lpf[2] ),
    .B(_1397_),
    .C(_1398_));
 sg13g2_nand3_1 _4330_ (.B(_1397_),
    .C(_1398_),
    .A(\audio_sample_lpf[2] ),
    .Y(_1400_));
 sg13g2_a21oi_1 _4331_ (.A1(_1397_),
    .A2(_1398_),
    .Y(_1401_),
    .B1(\audio_sample_lpf[2] ));
 sg13g2_nor3_1 _4332_ (.A(_1394_),
    .B(_1399_),
    .C(_1401_),
    .Y(_1402_));
 sg13g2_or3_1 _4333_ (.A(_1394_),
    .B(_1399_),
    .C(_1401_),
    .X(_1403_));
 sg13g2_o21ai_1 _4334_ (.B1(_1394_),
    .Y(_1404_),
    .A1(_1399_),
    .A2(_1401_));
 sg13g2_and3_1 _4335_ (.X(_1405_),
    .A(_0023_),
    .B(_1403_),
    .C(_1404_));
 sg13g2_a21oi_1 _4336_ (.A1(_1403_),
    .A2(_1404_),
    .Y(_1406_),
    .B1(_0023_));
 sg13g2_nor3_1 _4337_ (.A(_1393_),
    .B(_1405_),
    .C(_1406_),
    .Y(_1407_));
 sg13g2_o21ai_1 _4338_ (.B1(_1393_),
    .Y(_1408_),
    .A1(_1405_),
    .A2(_1406_));
 sg13g2_nor2b_1 _4339_ (.A(_1407_),
    .B_N(_1408_),
    .Y(_1409_));
 sg13g2_xnor2_1 _4340_ (.Y(_1410_),
    .A(_1389_),
    .B(_1409_));
 sg13g2_nand2_1 _4341_ (.Y(_1411_),
    .A(net200),
    .B(net882));
 sg13g2_o21ai_1 _4342_ (.B1(_1411_),
    .Y(_0164_),
    .A1(net882),
    .A2(_1410_));
 sg13g2_a21oi_1 _4343_ (.A1(_1389_),
    .A2(_1408_),
    .Y(_1412_),
    .B1(_1407_));
 sg13g2_nor2_1 _4344_ (.A(_1402_),
    .B(_1405_),
    .Y(_1413_));
 sg13g2_and2_1 _4345_ (.A(_1397_),
    .B(_1400_),
    .X(_1414_));
 sg13g2_a21oi_1 _4346_ (.A1(\bass_vol[3] ),
    .A2(_1365_),
    .Y(_1415_),
    .B1(net923));
 sg13g2_a21oi_2 _4347_ (.B1(_1415_),
    .Y(_1416_),
    .A2(net923),
    .A1(_0024_));
 sg13g2_inv_1 _4348_ (.Y(_1417_),
    .A(_1416_));
 sg13g2_nand2b_1 _4349_ (.Y(_1418_),
    .B(\sqr_vol[3] ),
    .A_N(net783));
 sg13g2_nor2_1 _4350_ (.A(_1417_),
    .B(_1418_),
    .Y(_1419_));
 sg13g2_xnor2_1 _4351_ (.Y(_1420_),
    .A(_1416_),
    .B(_1418_));
 sg13g2_xnor2_1 _4352_ (.Y(_1421_),
    .A(\audio_sample_lpf[3] ),
    .B(_1420_));
 sg13g2_nor2_1 _4353_ (.A(_1414_),
    .B(_1421_),
    .Y(_1422_));
 sg13g2_xor2_1 _4354_ (.B(_1421_),
    .A(_1414_),
    .X(_1423_));
 sg13g2_xnor2_1 _4355_ (.Y(_1424_),
    .A(_0027_),
    .B(_1423_));
 sg13g2_or2_1 _4356_ (.X(_1425_),
    .B(_1424_),
    .A(_1413_));
 sg13g2_and2_1 _4357_ (.A(_1413_),
    .B(_1424_),
    .X(_1426_));
 sg13g2_xor2_1 _4358_ (.B(_1424_),
    .A(_1413_),
    .X(_1427_));
 sg13g2_xnor2_1 _4359_ (.Y(_1428_),
    .A(_1412_),
    .B(_1427_));
 sg13g2_mux2_1 _4360_ (.A0(net269),
    .A1(_1428_),
    .S(_0811_),
    .X(_0165_));
 sg13g2_o21ai_1 _4361_ (.B1(_1425_),
    .Y(_1429_),
    .A1(_1412_),
    .A2(_1426_));
 sg13g2_a21oi_1 _4362_ (.A1(_0027_),
    .A2(_1423_),
    .Y(_1430_),
    .B1(_1422_));
 sg13g2_a21oi_2 _4363_ (.B1(_1419_),
    .Y(_1431_),
    .A2(_1420_),
    .A1(\audio_sample_lpf[3] ));
 sg13g2_a21oi_1 _4364_ (.A1(\bass_vol[4] ),
    .A2(_1365_),
    .Y(_1432_),
    .B1(net923));
 sg13g2_a21oi_2 _4365_ (.B1(_1432_),
    .Y(_1433_),
    .A2(net924),
    .A1(_0024_));
 sg13g2_inv_1 _4366_ (.Y(_1434_),
    .A(_1433_));
 sg13g2_nand2b_1 _4367_ (.Y(_1435_),
    .B(\sqr_vol[4] ),
    .A_N(net783));
 sg13g2_nor2_1 _4368_ (.A(_1434_),
    .B(_1435_),
    .Y(_1436_));
 sg13g2_xnor2_1 _4369_ (.Y(_1437_),
    .A(_1433_),
    .B(_1435_));
 sg13g2_xnor2_1 _4370_ (.Y(_1438_),
    .A(\audio_sample_lpf[4] ),
    .B(_1437_));
 sg13g2_nor2_1 _4371_ (.A(_1431_),
    .B(_1438_),
    .Y(_1439_));
 sg13g2_xor2_1 _4372_ (.B(_1438_),
    .A(_1431_),
    .X(_1440_));
 sg13g2_xnor2_1 _4373_ (.Y(_1441_),
    .A(_0028_),
    .B(_1440_));
 sg13g2_nor2_1 _4374_ (.A(_1430_),
    .B(_1441_),
    .Y(_1442_));
 sg13g2_xor2_1 _4375_ (.B(_1441_),
    .A(_1430_),
    .X(_1443_));
 sg13g2_xnor2_1 _4376_ (.Y(_1444_),
    .A(_1429_),
    .B(_1443_));
 sg13g2_nand2_1 _4377_ (.Y(_1445_),
    .A(net205),
    .B(net883));
 sg13g2_o21ai_1 _4378_ (.B1(_1445_),
    .Y(_0166_),
    .A1(net883),
    .A2(_1444_));
 sg13g2_a21oi_1 _4379_ (.A1(_1429_),
    .A2(_1443_),
    .Y(_1446_),
    .B1(_1442_));
 sg13g2_a21oi_1 _4380_ (.A1(_0028_),
    .A2(_1440_),
    .Y(_1447_),
    .B1(_1439_));
 sg13g2_a21oi_2 _4381_ (.B1(_1436_),
    .Y(_1448_),
    .A2(_1437_),
    .A1(\audio_sample_lpf[4] ));
 sg13g2_a21oi_1 _4382_ (.A1(\bass_vol[5] ),
    .A2(_1365_),
    .Y(_1449_),
    .B1(net923));
 sg13g2_a21oi_2 _4383_ (.B1(_1449_),
    .Y(_1450_),
    .A2(net923),
    .A1(_0024_));
 sg13g2_inv_1 _4384_ (.Y(_1451_),
    .A(_1450_));
 sg13g2_nand2b_1 _4385_ (.Y(_1452_),
    .B(\sqr_vol[5] ),
    .A_N(net783));
 sg13g2_nor2_1 _4386_ (.A(_1451_),
    .B(_1452_),
    .Y(_1453_));
 sg13g2_xnor2_1 _4387_ (.Y(_1454_),
    .A(_1450_),
    .B(_1452_));
 sg13g2_xnor2_1 _4388_ (.Y(_1455_),
    .A(\audio_sample_lpf[5] ),
    .B(_1454_));
 sg13g2_nor2_1 _4389_ (.A(_1448_),
    .B(_1455_),
    .Y(_1456_));
 sg13g2_xor2_1 _4390_ (.B(_1455_),
    .A(_1448_),
    .X(_1457_));
 sg13g2_xnor2_1 _4391_ (.Y(_1458_),
    .A(_0029_),
    .B(_1457_));
 sg13g2_or2_1 _4392_ (.X(_1459_),
    .B(_1458_),
    .A(_1447_));
 sg13g2_xor2_1 _4393_ (.B(_1458_),
    .A(_1447_),
    .X(_1460_));
 sg13g2_inv_1 _4394_ (.Y(_1461_),
    .A(_1460_));
 sg13g2_xnor2_1 _4395_ (.Y(_1462_),
    .A(_1446_),
    .B(_1461_));
 sg13g2_nand2_1 _4396_ (.Y(_1463_),
    .A(net228),
    .B(net882));
 sg13g2_o21ai_1 _4397_ (.B1(_1463_),
    .Y(_0167_),
    .A1(net882),
    .A2(_1462_));
 sg13g2_o21ai_1 _4398_ (.B1(_1459_),
    .Y(_1464_),
    .A1(_1446_),
    .A2(_1461_));
 sg13g2_nor2b_1 _4399_ (.A(\audio_sample_lpf[9] ),
    .B_N(\audio_sample_lpf[6] ),
    .Y(_1465_));
 sg13g2_xor2_1 _4400_ (.B(\audio_sample_lpf[9] ),
    .A(\audio_sample_lpf[6] ),
    .X(_1466_));
 sg13g2_a21oi_1 _4401_ (.A1(\audio_sample_lpf[5] ),
    .A2(_1454_),
    .Y(_1467_),
    .B1(_1453_));
 sg13g2_nor2_1 _4402_ (.A(_1466_),
    .B(_1467_),
    .Y(_1468_));
 sg13g2_xnor2_1 _4403_ (.Y(_1469_),
    .A(_1466_),
    .B(_1467_));
 sg13g2_a21oi_1 _4404_ (.A1(_0029_),
    .A2(_1457_),
    .Y(_1470_),
    .B1(_1456_));
 sg13g2_nor2_1 _4405_ (.A(_1469_),
    .B(_1470_),
    .Y(_1471_));
 sg13g2_nand2_1 _4406_ (.Y(_1472_),
    .A(_1469_),
    .B(_1470_));
 sg13g2_nand2b_1 _4407_ (.Y(_1473_),
    .B(_1472_),
    .A_N(_1471_));
 sg13g2_xnor2_1 _4408_ (.Y(_1474_),
    .A(_1464_),
    .B(_1473_));
 sg13g2_mux2_1 _4409_ (.A0(net221),
    .A1(_1474_),
    .S(_0811_),
    .X(_0168_));
 sg13g2_a21oi_1 _4410_ (.A1(_1464_),
    .A2(_1472_),
    .Y(_1475_),
    .B1(_1471_));
 sg13g2_xnor2_1 _4411_ (.Y(_1476_),
    .A(\audio_sample_lpf[7] ),
    .B(_1465_));
 sg13g2_nand2_1 _4412_ (.Y(_1477_),
    .A(_1468_),
    .B(_1476_));
 sg13g2_xnor2_1 _4413_ (.Y(_1478_),
    .A(_1468_),
    .B(_1476_));
 sg13g2_xnor2_1 _4414_ (.Y(_1479_),
    .A(_1475_),
    .B(_1478_));
 sg13g2_nand2_1 _4415_ (.Y(_1480_),
    .A(net239),
    .B(net883));
 sg13g2_o21ai_1 _4416_ (.B1(_1480_),
    .Y(_0169_),
    .A1(net883),
    .A2(_1479_));
 sg13g2_o21ai_1 _4417_ (.B1(_1477_),
    .Y(_1481_),
    .A1(_1475_),
    .A2(_1478_));
 sg13g2_nor3_1 _4418_ (.A(\audio_sample_lpf[7] ),
    .B(\audio_sample_lpf[8] ),
    .C(_1465_),
    .Y(_1482_));
 sg13g2_o21ai_1 _4419_ (.B1(net175),
    .Y(_1483_),
    .A1(\audio_sample_lpf[7] ),
    .A2(_1465_));
 sg13g2_nand2b_1 _4420_ (.Y(_1484_),
    .B(_1483_),
    .A_N(_1482_));
 sg13g2_xnor2_1 _4421_ (.Y(_1485_),
    .A(_1481_),
    .B(_1484_));
 sg13g2_nand2_1 _4422_ (.Y(_1486_),
    .A(net175),
    .B(net883));
 sg13g2_o21ai_1 _4423_ (.B1(_1486_),
    .Y(_0170_),
    .A1(net883),
    .A2(_1485_));
 sg13g2_o21ai_1 _4424_ (.B1(_0811_),
    .Y(_1487_),
    .A1(_1481_),
    .A2(_1482_));
 sg13g2_a21oi_1 _4425_ (.A1(_1481_),
    .A2(_1483_),
    .Y(_1488_),
    .B1(_1487_));
 sg13g2_xor2_1 _4426_ (.B(_1488_),
    .A(net217),
    .X(_0171_));
 sg13g2_xnor2_1 _4427_ (.Y(_0172_),
    .A(net209),
    .B(net874));
 sg13g2_a21oi_1 _4428_ (.A1(\sample_beat_ctr[0] ),
    .A2(net877),
    .Y(_1489_),
    .B1(net194));
 sg13g2_and3_1 _4429_ (.X(_1490_),
    .A(net194),
    .B(\sample_beat_ctr[0] ),
    .C(net877));
 sg13g2_nor3_1 _4430_ (.A(net864),
    .B(net195),
    .C(_1490_),
    .Y(_0173_));
 sg13g2_o21ai_1 _4431_ (.B1(_0761_),
    .Y(_1491_),
    .A1(net198),
    .A2(_1490_));
 sg13g2_inv_1 _4432_ (.Y(_0174_),
    .A(net199));
 sg13g2_nor3_1 _4433_ (.A(\sample_beat_ctr[1] ),
    .B(_0761_),
    .C(_0806_),
    .Y(_1492_));
 sg13g2_mux2_1 _4434_ (.A0(net961),
    .A1(net72),
    .S(_1492_),
    .X(_0175_));
 sg13g2_nand2_1 _4435_ (.Y(_1493_),
    .A(\hvsync_gen.vpos[0] ),
    .B(net830));
 sg13g2_nor3_1 _4436_ (.A(\hvsync_gen.vpos[8] ),
    .B(_1533_),
    .C(_0756_),
    .Y(_1494_));
 sg13g2_nand3_1 _4437_ (.B(net952),
    .C(_1494_),
    .A(\hvsync_gen.vpos[2] ),
    .Y(_1495_));
 sg13g2_nand3_1 _4438_ (.B(_0858_),
    .C(_1495_),
    .A(net1022),
    .Y(_1496_));
 sg13g2_o21ai_1 _4439_ (.B1(_1493_),
    .Y(_0176_),
    .A1(_1522_),
    .A2(_1496_));
 sg13g2_and2_1 _4440_ (.A(\hvsync_gen.vpos[0] ),
    .B(\hvsync_gen.vpos[1] ),
    .X(_1497_));
 sg13g2_nor3_1 _4441_ (.A(_0755_),
    .B(_1496_),
    .C(_1497_),
    .Y(_1498_));
 sg13g2_a21o_1 _4442_ (.A2(net830),
    .A1(net252),
    .B1(_1498_),
    .X(_0177_));
 sg13g2_nand3_1 _4443_ (.B(\hvsync_gen.vpos[1] ),
    .C(_0860_),
    .A(\hvsync_gen.vpos[0] ),
    .Y(_1499_));
 sg13g2_and2_1 _4444_ (.A(_0860_),
    .B(_1496_),
    .X(_1500_));
 sg13g2_xor2_1 _4445_ (.B(_1499_),
    .A(net960),
    .X(_1501_));
 sg13g2_nor2_1 _4446_ (.A(_1500_),
    .B(net274),
    .Y(_0178_));
 sg13g2_nand2_1 _4447_ (.Y(_1502_),
    .A(net952),
    .B(_0859_));
 sg13g2_nand3b_1 _4448_ (.B(\hvsync_gen.vpos[1] ),
    .C(\hvsync_gen.vpos[0] ),
    .Y(_1503_),
    .A_N(net276));
 sg13g2_xnor2_1 _4449_ (.Y(_1504_),
    .A(net941),
    .B(_1503_));
 sg13g2_o21ai_1 _4450_ (.B1(_1502_),
    .Y(_0179_),
    .A1(_1496_),
    .A2(_1504_));
 sg13g2_nand4_1 _4451_ (.B(\hvsync_gen.vpos[1] ),
    .C(net960),
    .A(\hvsync_gen.vpos[0] ),
    .Y(_1505_),
    .D(net952));
 sg13g2_nor2_1 _4452_ (.A(net830),
    .B(_1505_),
    .Y(_1506_));
 sg13g2_nor3_2 _4453_ (.A(_1529_),
    .B(net830),
    .C(_1505_),
    .Y(_1507_));
 sg13g2_nor2_1 _4454_ (.A(net948),
    .B(_1506_),
    .Y(_1508_));
 sg13g2_nor3_1 _4455_ (.A(_1500_),
    .B(_1507_),
    .C(_1508_),
    .Y(_0180_));
 sg13g2_nand2_1 _4456_ (.Y(_1509_),
    .A(net947),
    .B(net830));
 sg13g2_nor2_1 _4457_ (.A(net257),
    .B(_1505_),
    .Y(_1510_));
 sg13g2_xnor2_1 _4458_ (.Y(_1511_),
    .A(net947),
    .B(_1510_));
 sg13g2_o21ai_1 _4459_ (.B1(_1509_),
    .Y(_0181_),
    .A1(_1496_),
    .A2(_1511_));
 sg13g2_and2_1 _4460_ (.A(net946),
    .B(_1507_),
    .X(_1512_));
 sg13g2_nand3_1 _4461_ (.B(net950),
    .C(net944),
    .A(net946),
    .Y(_1513_));
 sg13g2_a21oi_1 _4462_ (.A1(net944),
    .A2(_1512_),
    .Y(_1514_),
    .B1(_1500_));
 sg13g2_o21ai_1 _4463_ (.B1(_1514_),
    .Y(_1515_),
    .A1(net944),
    .A2(_1512_));
 sg13g2_inv_1 _4464_ (.Y(_0182_),
    .A(_1515_));
 sg13g2_nand2_1 _4465_ (.Y(_1516_),
    .A(net943),
    .B(_1514_));
 sg13g2_or3_1 _4466_ (.A(_1496_),
    .B(_1505_),
    .C(_1513_),
    .X(_1517_));
 sg13g2_o21ai_1 _4467_ (.B1(_1516_),
    .Y(_0183_),
    .A1(net137),
    .A2(_1517_));
 sg13g2_nand3_1 _4468_ (.B(net944),
    .C(_1512_),
    .A(net943),
    .Y(_1518_));
 sg13g2_a221oi_1 _4469_ (.B2(_1532_),
    .C1(_1500_),
    .B1(_1518_),
    .A1(_0663_),
    .Y(_0184_),
    .A2(_1507_));
 sg13g2_nor2b_1 _4470_ (.A(_1500_),
    .B_N(net942),
    .Y(_1519_));
 sg13g2_o21ai_1 _4471_ (.B1(_1519_),
    .Y(_1520_),
    .A1(net189),
    .A2(_1518_));
 sg13g2_or2_1 _4472_ (.X(_1521_),
    .B(_1975_),
    .A(_1530_));
 sg13g2_o21ai_1 _4473_ (.B1(_1520_),
    .Y(_0185_),
    .A1(_1517_),
    .A2(_1521_));
 sg13g2_dfrbp_1 _4474_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net1016),
    .D(net98),
    .Q_N(\songpos[0] ),
    .Q(_0044_));
 sg13g2_dfrbp_1 _4475_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net1009),
    .D(_0060_),
    .Q_N(\songpos[1] ),
    .Q(_0045_));
 sg13g2_dfrbp_1 _4476_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net1009),
    .D(_0061_),
    .Q_N(\songpos[2] ),
    .Q(_0046_));
 sg13g2_dfrbp_1 _4477_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net1009),
    .D(_0062_),
    .Q_N(\songpos[3] ),
    .Q(_0047_));
 sg13g2_dfrbp_1 _4478_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net1009),
    .D(net89),
    .Q_N(\songpos[4] ),
    .Q(_0048_));
 sg13g2_dfrbp_1 _4479_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net1016),
    .D(_0064_),
    .Q_N(\songpos[5] ),
    .Q(_0049_));
 sg13g2_dfrbp_1 _4480_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net1016),
    .D(net110),
    .Q_N(\songpos[6] ),
    .Q(_0050_));
 sg13g2_dfrbp_1 _4481_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net1016),
    .D(_0066_),
    .Q_N(\songpos[7] ),
    .Q(_0051_));
 sg13g2_dfrbp_1 _4482_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net1009),
    .D(_0067_),
    .Q_N(\songpos[8] ),
    .Q(_0052_));
 sg13g2_dfrbp_1 _4483_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net27),
    .D(net75),
    .Q_N(_0043_),
    .Q(\kick_ctr[0] ));
 sg13g2_dfrbp_1 _4484_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net25),
    .D(_0069_),
    .Q_N(_2262_),
    .Q(\kick_ctr[1] ));
 sg13g2_dfrbp_1 _4485_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net1020),
    .D(_0000_),
    .Q_N(_2263_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _4486_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net1020),
    .D(_0001_),
    .Q_N(_2264_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _4487_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net1020),
    .D(_0002_),
    .Q_N(_2265_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _4488_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net1021),
    .D(_0003_),
    .Q_N(_2266_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _4489_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net1020),
    .D(_0004_),
    .Q_N(_2267_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _4490_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net1021),
    .D(_0005_),
    .Q_N(_2261_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _4491_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net23),
    .D(_0070_),
    .Q_N(_0042_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 _4492_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net22),
    .D(_0071_),
    .Q_N(_2260_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _4493_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net21),
    .D(_0072_),
    .Q_N(_2259_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _4494_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net20),
    .D(_0073_),
    .Q_N(_2258_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _4495_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net19),
    .D(_0074_),
    .Q_N(_2257_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _4496_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net18),
    .D(_0075_),
    .Q_N(_2256_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _4497_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net17),
    .D(_0076_),
    .Q_N(_2255_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _4498_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net16),
    .D(_0077_),
    .Q_N(_0034_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _4499_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net15),
    .D(_0078_),
    .Q_N(_0033_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _4500_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net64),
    .D(net184),
    .Q_N(_0008_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _4501_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net1016),
    .D(net71),
    .Q_N(_0041_),
    .Q(\frame_count[0] ));
 sg13g2_dfrbp_1 _4502_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net1017),
    .D(net193),
    .Q_N(_2254_),
    .Q(\frame_count[1] ));
 sg13g2_dfrbp_1 _4503_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net1017),
    .D(net180),
    .Q_N(_2253_),
    .Q(\frame_count[2] ));
 sg13g2_dfrbp_1 _4504_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net1017),
    .D(net144),
    .Q_N(_2252_),
    .Q(\frame_count[3] ));
 sg13g2_dfrbp_1 _4505_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net1020),
    .D(_0084_),
    .Q_N(_2251_),
    .Q(\frame_count[4] ));
 sg13g2_dfrbp_1 _4506_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net1020),
    .D(_0085_),
    .Q_N(_2250_),
    .Q(\frame_count[5] ));
 sg13g2_dfrbp_1 _4507_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net1020),
    .D(net178),
    .Q_N(_2249_),
    .Q(\frame_count[6] ));
 sg13g2_dfrbp_1 _4508_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net1020),
    .D(net132),
    .Q_N(_2248_),
    .Q(\frame_count[7] ));
 sg13g2_dfrbp_1 _4509_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net63),
    .D(_0088_),
    .Q_N(_2247_),
    .Q(\line_lfsr[0] ));
 sg13g2_dfrbp_1 _4510_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net61),
    .D(net155),
    .Q_N(_2246_),
    .Q(\line_lfsr[1] ));
 sg13g2_dfrbp_1 _4511_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net60),
    .D(_0090_),
    .Q_N(_2245_),
    .Q(\line_lfsr[2] ));
 sg13g2_dfrbp_1 _4512_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net58),
    .D(net163),
    .Q_N(_2244_),
    .Q(\line_lfsr[3] ));
 sg13g2_dfrbp_1 _4513_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net56),
    .D(_0092_),
    .Q_N(_2243_),
    .Q(\line_lfsr[4] ));
 sg13g2_dfrbp_1 _4514_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net54),
    .D(net169),
    .Q_N(_2242_),
    .Q(\line_lfsr[5] ));
 sg13g2_dfrbp_1 _4515_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net52),
    .D(net186),
    .Q_N(_2241_),
    .Q(\line_lfsr[6] ));
 sg13g2_dfrbp_1 _4516_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net1021),
    .D(net69),
    .Q_N(_0038_),
    .Q(\nyanframe[0] ));
 sg13g2_dfrbp_1 _4517_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net1021),
    .D(net262),
    .Q_N(_2240_),
    .Q(\nyanframe[1] ));
 sg13g2_dfrbp_1 _4518_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net1021),
    .D(net224),
    .Q_N(_0031_),
    .Q(\nyanframe[2] ));
 sg13g2_dfrbp_1 _4519_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net1012),
    .D(net102),
    .Q_N(\cos[0] ),
    .Q(_0053_));
 sg13g2_dfrbp_1 _4520_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net1012),
    .D(net128),
    .Q_N(\cos[1] ),
    .Q(_0054_));
 sg13g2_dfrbp_1 _4521_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net1012),
    .D(net117),
    .Q_N(\cos[2] ),
    .Q(_0055_));
 sg13g2_dfrbp_1 _4522_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net1012),
    .D(net107),
    .Q_N(\cos[3] ),
    .Q(_0056_));
 sg13g2_dfrbp_1 _4523_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net1011),
    .D(_0102_),
    .Q_N(\cos[4] ),
    .Q(_0057_));
 sg13g2_dfrbp_1 _4524_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net1011),
    .D(net81),
    .Q_N(\cos[5] ),
    .Q(_0058_));
 sg13g2_dfrbp_1 _4525_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net1012),
    .D(_0104_),
    .Q_N(_2239_),
    .Q(\cos[6] ));
 sg13g2_dfrbp_1 _4526_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net1011),
    .D(_0105_),
    .Q_N(_2238_),
    .Q(\sin[0] ));
 sg13g2_dfrbp_1 _4527_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net1013),
    .D(_0106_),
    .Q_N(_2237_),
    .Q(\nyan_x_offset[0] ));
 sg13g2_dfrbp_1 _4528_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net1011),
    .D(_0107_),
    .Q_N(_2236_),
    .Q(\nyan_x_offset[1] ));
 sg13g2_dfrbp_1 _4529_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net1012),
    .D(_0108_),
    .Q_N(_2235_),
    .Q(\nyan_x_offset[2] ));
 sg13g2_dfrbp_1 _4530_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net1012),
    .D(_0109_),
    .Q_N(_2234_),
    .Q(\nyan_x_offset[3] ));
 sg13g2_dfrbp_1 _4531_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net1013),
    .D(_0110_),
    .Q_N(_2233_),
    .Q(\nyan_x_offset[4] ));
 sg13g2_dfrbp_1 _4532_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net1012),
    .D(net235),
    .Q_N(_2232_),
    .Q(\sin[6] ));
 sg13g2_dfrbp_1 _4533_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net1006),
    .D(net130),
    .Q_N(_2231_),
    .Q(\bass_pha[0] ));
 sg13g2_dfrbp_1 _4534_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net1006),
    .D(_0113_),
    .Q_N(_2230_),
    .Q(\bass_pha[1] ));
 sg13g2_dfrbp_1 _4535_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net1006),
    .D(net126),
    .Q_N(_2229_),
    .Q(\bass_pha[2] ));
 sg13g2_dfrbp_1 _4536_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net1006),
    .D(_0115_),
    .Q_N(_2228_),
    .Q(\bass_pha[3] ));
 sg13g2_dfrbp_1 _4537_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net1006),
    .D(_0116_),
    .Q_N(_2227_),
    .Q(\bass_pha[4] ));
 sg13g2_dfrbp_1 _4538_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net1006),
    .D(_0117_),
    .Q_N(_2226_),
    .Q(\bass_pha[5] ));
 sg13g2_dfrbp_1 _4539_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net1006),
    .D(_0118_),
    .Q_N(_2225_),
    .Q(\bass_pha[6] ));
 sg13g2_dfrbp_1 _4540_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net1006),
    .D(_0119_),
    .Q_N(_2224_),
    .Q(\bass_pha[7] ));
 sg13g2_dfrbp_1 _4541_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net1007),
    .D(_0120_),
    .Q_N(_2223_),
    .Q(\bass_pha[8] ));
 sg13g2_dfrbp_1 _4542_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net1008),
    .D(net96),
    .Q_N(_0020_),
    .Q(\bass_pha[9] ));
 sg13g2_dfrbp_1 _4543_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net1008),
    .D(net148),
    .Q_N(_2222_),
    .Q(\bass_pha[10] ));
 sg13g2_dfrbp_1 _4544_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net1008),
    .D(net136),
    .Q_N(_2221_),
    .Q(\bass_pha[11] ));
 sg13g2_dfrbp_1 _4545_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net1008),
    .D(net100),
    .Q_N(_0021_),
    .Q(\bass_pha[12] ));
 sg13g2_dfrbp_1 _4546_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net1008),
    .D(net87),
    .Q_N(_0025_),
    .Q(\bass_pha[13] ));
 sg13g2_dfrbp_1 _4547_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net1009),
    .D(net79),
    .Q_N(_0022_),
    .Q(\bass_pha[14] ));
 sg13g2_dfrbp_1 _4548_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net1008),
    .D(net114),
    .Q_N(_0024_),
    .Q(\bass_pha[15] ));
 sg13g2_dfrbp_1 _4549_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net1008),
    .D(net158),
    .Q_N(_2220_),
    .Q(\bass_vol[0] ));
 sg13g2_dfrbp_1 _4550_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net1015),
    .D(_0129_),
    .Q_N(_2219_),
    .Q(\bass_vol[1] ));
 sg13g2_dfrbp_1 _4551_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net1008),
    .D(_0130_),
    .Q_N(_2218_),
    .Q(\bass_vol[2] ));
 sg13g2_dfrbp_1 _4552_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net1015),
    .D(net251),
    .Q_N(_2217_),
    .Q(\bass_vol[3] ));
 sg13g2_dfrbp_1 _4553_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net1015),
    .D(_0132_),
    .Q_N(_2216_),
    .Q(\bass_vol[4] ));
 sg13g2_dfrbp_1 _4554_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net1015),
    .D(net188),
    .Q_N(_2215_),
    .Q(\bass_vol[5] ));
 sg13g2_dfrbp_1 _4555_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net1013),
    .D(_0134_),
    .Q_N(_2214_),
    .Q(\sqr_pha[0] ));
 sg13g2_dfrbp_1 _4556_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net1011),
    .D(net83),
    .Q_N(_0010_),
    .Q(\sqr_pha[1] ));
 sg13g2_dfrbp_1 _4557_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net1011),
    .D(net121),
    .Q_N(_2213_),
    .Q(\sqr_pha[2] ));
 sg13g2_dfrbp_1 _4558_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net1011),
    .D(_0137_),
    .Q_N(_2212_),
    .Q(\sqr_pha[3] ));
 sg13g2_dfrbp_1 _4559_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net1011),
    .D(net150),
    .Q_N(_2211_),
    .Q(\sqr_pha[4] ));
 sg13g2_dfrbp_1 _4560_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net1007),
    .D(net123),
    .Q_N(_0011_),
    .Q(\sqr_pha[5] ));
 sg13g2_dfrbp_1 _4561_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net1007),
    .D(_0140_),
    .Q_N(_2210_),
    .Q(\sqr_pha[6] ));
 sg13g2_dfrbp_1 _4562_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net1007),
    .D(_0141_),
    .Q_N(_2209_),
    .Q(\sqr_pha[7] ));
 sg13g2_dfrbp_1 _4563_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net1010),
    .D(_0142_),
    .Q_N(_2208_),
    .Q(\sqr_pha[8] ));
 sg13g2_dfrbp_1 _4564_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net1010),
    .D(_0143_),
    .Q_N(_2207_),
    .Q(\sqr_pha[9] ));
 sg13g2_dfrbp_1 _4565_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net1007),
    .D(_0144_),
    .Q_N(_2206_),
    .Q(\sqr_pha[10] ));
 sg13g2_dfrbp_1 _4566_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net1007),
    .D(_0145_),
    .Q_N(_2205_),
    .Q(\sqr_pha[11] ));
 sg13g2_dfrbp_1 _4567_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net1007),
    .D(net105),
    .Q_N(_2204_),
    .Q(\sqr_pha[12] ));
 sg13g2_dfrbp_1 _4568_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net1015),
    .D(net152),
    .Q_N(_2203_),
    .Q(\sqr_vol[0] ));
 sg13g2_dfrbp_1 _4569_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net1015),
    .D(net256),
    .Q_N(_2202_),
    .Q(\sqr_vol[1] ));
 sg13g2_dfrbp_1 _4570_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net1018),
    .D(_0149_),
    .Q_N(_2201_),
    .Q(\sqr_vol[2] ));
 sg13g2_dfrbp_1 _4571_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net1015),
    .D(net231),
    .Q_N(_0009_),
    .Q(\sqr_vol[3] ));
 sg13g2_dfrbp_1 _4572_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net1017),
    .D(_0151_),
    .Q_N(_2200_),
    .Q(\sqr_vol[4] ));
 sg13g2_dfrbp_1 _4573_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net1017),
    .D(_0152_),
    .Q_N(_2199_),
    .Q(\sqr_vol[5] ));
 sg13g2_dfrbp_1 _4574_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net40),
    .D(_0153_),
    .Q_N(_0012_),
    .Q(\kick_osci[0] ));
 sg13g2_dfrbp_1 _4575_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net38),
    .D(net139),
    .Q_N(_0013_),
    .Q(\kick_osci[1] ));
 sg13g2_dfrbp_1 _4576_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net36),
    .D(_0155_),
    .Q_N(_0014_),
    .Q(\kick_osci[2] ));
 sg13g2_dfrbp_1 _4577_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net34),
    .D(_0156_),
    .Q_N(_0015_),
    .Q(\kick_osci[3] ));
 sg13g2_dfrbp_1 _4578_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net32),
    .D(_0157_),
    .Q_N(_0016_),
    .Q(\kick_osci[4] ));
 sg13g2_dfrbp_1 _4579_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net30),
    .D(_0158_),
    .Q_N(_0017_),
    .Q(\kick_osci[5] ));
 sg13g2_dfrbp_1 _4580_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net28),
    .D(_0159_),
    .Q_N(_0018_),
    .Q(\kick_osci[6] ));
 sg13g2_dfrbp_1 _4581_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net24),
    .D(net227),
    .Q_N(_0019_),
    .Q(\kick_osci[7] ));
 sg13g2_dfrbp_1 _4582_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net50),
    .D(net216),
    .Q_N(_2268_),
    .Q(\kick_osci[8] ));
 sg13g2_dfrbp_1 _4583_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net1018),
    .D(net85),
    .Q_N(_2269_),
    .Q(\audio_pwm_accum[0] ));
 sg13g2_dfrbp_1 _4584_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net1015),
    .D(\audio_pwm_accum_next[1] ),
    .Q_N(_2270_),
    .Q(\audio_pwm_accum[1] ));
 sg13g2_dfrbp_1 _4585_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net1019),
    .D(net243),
    .Q_N(_2271_),
    .Q(\audio_pwm_accum[2] ));
 sg13g2_dfrbp_1 _4586_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net1019),
    .D(\audio_pwm_accum_next[3] ),
    .Q_N(_2272_),
    .Q(\audio_pwm_accum[3] ));
 sg13g2_dfrbp_1 _4587_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net1022),
    .D(\audio_pwm_accum_next[4] ),
    .Q_N(_2273_),
    .Q(\audio_pwm_accum[4] ));
 sg13g2_dfrbp_1 _4588_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net1019),
    .D(net233),
    .Q_N(_2274_),
    .Q(\audio_pwm_accum[5] ));
 sg13g2_dfrbp_1 _4589_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net1019),
    .D(net268),
    .Q_N(_2275_),
    .Q(\audio_pwm_accum[6] ));
 sg13g2_dfrbp_1 _4590_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net1019),
    .D(net245),
    .Q_N(_2276_),
    .Q(\audio_pwm_accum[7] ));
 sg13g2_dfrbp_1 _4591_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net1019),
    .D(net249),
    .Q_N(_2277_),
    .Q(\audio_pwm_accum[8] ));
 sg13g2_dfrbp_1 _4592_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net1019),
    .D(\audio_pwm_accum_next[9] ),
    .Q_N(_2198_),
    .Q(\audio_pwm_accum[9] ));
 sg13g2_dfrbp_1 _4593_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net57),
    .D(net191),
    .Q_N(_2197_),
    .Q(\audio_sample_lpf[0] ));
 sg13g2_dfrbp_1 _4594_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net55),
    .D(net212),
    .Q_N(_2196_),
    .Q(\audio_sample_lpf[1] ));
 sg13g2_dfrbp_1 _4595_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net53),
    .D(net201),
    .Q_N(_2195_),
    .Q(\audio_sample_lpf[2] ));
 sg13g2_dfrbp_1 _4596_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net51),
    .D(_0165_),
    .Q_N(_2194_),
    .Q(\audio_sample_lpf[3] ));
 sg13g2_dfrbp_1 _4597_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net49),
    .D(_0166_),
    .Q_N(_0026_),
    .Q(\audio_sample_lpf[4] ));
 sg13g2_dfrbp_1 _4598_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net48),
    .D(_0167_),
    .Q_N(_0023_),
    .Q(\audio_sample_lpf[5] ));
 sg13g2_dfrbp_1 _4599_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net47),
    .D(_0168_),
    .Q_N(_0027_),
    .Q(\audio_sample_lpf[6] ));
 sg13g2_dfrbp_1 _4600_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net46),
    .D(_0169_),
    .Q_N(_0028_),
    .Q(\audio_sample_lpf[7] ));
 sg13g2_dfrbp_1 _4601_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net45),
    .D(net176),
    .Q_N(_0029_),
    .Q(\audio_sample_lpf[8] ));
 sg13g2_dfrbp_1 _4602_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net44),
    .D(net218),
    .Q_N(_2193_),
    .Q(\audio_sample_lpf[9] ));
 sg13g2_dfrbp_1 _4603_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net1017),
    .D(_0172_),
    .Q_N(_2192_),
    .Q(\sample_beat_ctr[0] ));
 sg13g2_dfrbp_1 _4604_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net1016),
    .D(net196),
    .Q_N(_2191_),
    .Q(\sample_beat_ctr[1] ));
 sg13g2_dfrbp_1 _4605_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net1016),
    .D(_0174_),
    .Q_N(_2190_),
    .Q(\sample_beat_ctr[2] ));
 sg13g2_dfrbp_1 _4606_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net1016),
    .D(net73),
    .Q_N(_2185_),
    .Q(song_loops));
 sg13g2_dfrbp_1 _4607_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net43),
    .D(_0006_),
    .Q_N(_2189_),
    .Q(hsync));
 sg13g2_dfrbp_1 _4608_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net42),
    .D(net77),
    .Q_N(_0040_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _4609_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net39),
    .D(_0177_),
    .Q_N(_0032_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _4610_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net35),
    .D(_0178_),
    .Q_N(_0030_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _4611_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net31),
    .D(_0179_),
    .Q_N(_0039_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _4612_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net26),
    .D(_0180_),
    .Q_N(_0036_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _4613_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net59),
    .D(net258),
    .Q_N(_0035_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _4614_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net37),
    .D(_0182_),
    .Q_N(_2188_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _4615_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net29),
    .D(_0183_),
    .Q_N(_2187_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _4616_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net41),
    .D(_0184_),
    .Q_N(_0037_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _4617_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net33),
    .D(_0185_),
    .Q_N(_2278_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _4618_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net62),
    .D(_0007_),
    .Q_N(_2186_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_tiehi _4498__16 (.L_HI(net16));
 sg13g2_tiehi _4497__17 (.L_HI(net17));
 sg13g2_tiehi _4496__18 (.L_HI(net18));
 sg13g2_tiehi _4495__19 (.L_HI(net19));
 sg13g2_tiehi _4494__20 (.L_HI(net20));
 sg13g2_tiehi _4493__21 (.L_HI(net21));
 sg13g2_tiehi _4492__22 (.L_HI(net22));
 sg13g2_tiehi _4491__23 (.L_HI(net23));
 sg13g2_tiehi _4581__24 (.L_HI(net24));
 sg13g2_tiehi _4484__25 (.L_HI(net25));
 sg13g2_tiehi _4612__26 (.L_HI(net26));
 sg13g2_tiehi _4483__27 (.L_HI(net27));
 sg13g2_tiehi _4580__28 (.L_HI(net28));
 sg13g2_tiehi _4615__29 (.L_HI(net29));
 sg13g2_tiehi _4579__30 (.L_HI(net30));
 sg13g2_tiehi _4611__31 (.L_HI(net31));
 sg13g2_tiehi _4578__32 (.L_HI(net32));
 sg13g2_tiehi _4617__33 (.L_HI(net33));
 sg13g2_tiehi _4577__34 (.L_HI(net34));
 sg13g2_tiehi _4610__35 (.L_HI(net35));
 sg13g2_tiehi _4576__36 (.L_HI(net36));
 sg13g2_tiehi _4614__37 (.L_HI(net37));
 sg13g2_tiehi _4575__38 (.L_HI(net38));
 sg13g2_tiehi _4609__39 (.L_HI(net39));
 sg13g2_tiehi _4574__40 (.L_HI(net40));
 sg13g2_tiehi _4616__41 (.L_HI(net41));
 sg13g2_tiehi _4608__42 (.L_HI(net42));
 sg13g2_tiehi _4607__43 (.L_HI(net43));
 sg13g2_tiehi _4602__44 (.L_HI(net44));
 sg13g2_tiehi _4601__45 (.L_HI(net45));
 sg13g2_tiehi _4600__46 (.L_HI(net46));
 sg13g2_tiehi _4599__47 (.L_HI(net47));
 sg13g2_tiehi _4598__48 (.L_HI(net48));
 sg13g2_tiehi _4597__49 (.L_HI(net49));
 sg13g2_tiehi _4582__50 (.L_HI(net50));
 sg13g2_tiehi _4596__51 (.L_HI(net51));
 sg13g2_tiehi _4515__52 (.L_HI(net52));
 sg13g2_tiehi _4595__53 (.L_HI(net53));
 sg13g2_tiehi _4514__54 (.L_HI(net54));
 sg13g2_tiehi _4594__55 (.L_HI(net55));
 sg13g2_tiehi _4513__56 (.L_HI(net56));
 sg13g2_tiehi _4593__57 (.L_HI(net57));
 sg13g2_tiehi _4512__58 (.L_HI(net58));
 sg13g2_tiehi _4613__59 (.L_HI(net59));
 sg13g2_tiehi _4511__60 (.L_HI(net60));
 sg13g2_tiehi _4510__61 (.L_HI(net61));
 sg13g2_tiehi _4618__62 (.L_HI(net62));
 sg13g2_tiehi _4509__63 (.L_HI(net63));
 sg13g2_tiehi _4500__64 (.L_HI(net64));
 sg13g2_tiehi tt_um_a1k0n_nyancat_65 (.L_HI(net65));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_a1k0n_nyancat_2 (.L_LO(net2));
 sg13g2_tielo tt_um_a1k0n_nyancat_3 (.L_LO(net3));
 sg13g2_tielo tt_um_a1k0n_nyancat_4 (.L_LO(net4));
 sg13g2_tielo tt_um_a1k0n_nyancat_5 (.L_LO(net5));
 sg13g2_tielo tt_um_a1k0n_nyancat_6 (.L_LO(net6));
 sg13g2_tielo tt_um_a1k0n_nyancat_7 (.L_LO(net7));
 sg13g2_tielo tt_um_a1k0n_nyancat_8 (.L_LO(net8));
 sg13g2_tielo tt_um_a1k0n_nyancat_9 (.L_LO(net9));
 sg13g2_tielo tt_um_a1k0n_nyancat_10 (.L_LO(net10));
 sg13g2_tielo tt_um_a1k0n_nyancat_11 (.L_LO(net11));
 sg13g2_tielo tt_um_a1k0n_nyancat_12 (.L_LO(net12));
 sg13g2_tielo tt_um_a1k0n_nyancat_13 (.L_LO(net13));
 sg13g2_tielo tt_um_a1k0n_nyancat_14 (.L_LO(net14));
 sg13g2_tiehi _4499__15 (.L_HI(net15));
 sg13g2_buf_1 _4684_ (.A(audio_pwm),
    .X(uio_out[7]));
 sg13g2_buf_1 _4685_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _4686_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout773 (.A(net774),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_0398_),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(net776),
    .X(net775));
 sg13g2_buf_1 fanout776 (.A(_2160_),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(_2058_),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(_0850_),
    .X(net778));
 sg13g2_buf_1 fanout779 (.A(_0850_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(net781),
    .X(net780));
 sg13g2_buf_1 fanout781 (.A(_0933_),
    .X(net781));
 sg13g2_buf_4 fanout782 (.X(net782),
    .A(_1658_));
 sg13g2_buf_2 fanout783 (.A(_1353_),
    .X(net783));
 sg13g2_buf_4 fanout784 (.X(net784),
    .A(_1796_));
 sg13g2_buf_2 fanout785 (.A(_1796_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(net787),
    .X(net786));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(_1721_));
 sg13g2_buf_2 fanout788 (.A(net791),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(net791),
    .X(net789));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(net791));
 sg13g2_buf_2 fanout791 (.A(_1623_),
    .X(net791));
 sg13g2_buf_4 fanout792 (.X(net792),
    .A(_1622_));
 sg13g2_buf_2 fanout793 (.A(_1622_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(net795),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_1622_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(_0487_),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_1764_));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(_1691_));
 sg13g2_buf_2 fanout799 (.A(net800),
    .X(net799));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(net804));
 sg13g2_buf_2 fanout801 (.A(net803),
    .X(net801));
 sg13g2_buf_1 fanout802 (.A(net803),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(net804),
    .X(net803));
 sg13g2_buf_1 fanout804 (.A(net808),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(net808),
    .X(net805));
 sg13g2_buf_4 fanout806 (.X(net806),
    .A(net807));
 sg13g2_buf_1 fanout807 (.A(net808),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_1647_),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(net810),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(net815),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(net815),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(net815),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(net814),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(net815),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(_1646_),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(net821),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(net820),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(net820),
    .X(net818));
 sg13g2_buf_1 fanout819 (.A(net820),
    .X(net819));
 sg13g2_buf_1 fanout820 (.A(net821),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_1646_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(net823),
    .X(net822));
 sg13g2_buf_4 fanout823 (.X(net823),
    .A(_1625_));
 sg13g2_buf_4 fanout824 (.X(net824),
    .A(net826));
 sg13g2_buf_2 fanout825 (.A(net826),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_1619_),
    .X(net826));
 sg13g2_buf_4 fanout827 (.X(net827),
    .A(net829));
 sg13g2_buf_2 fanout828 (.A(net829),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_1618_),
    .X(net829));
 sg13g2_buf_4 fanout830 (.X(net830),
    .A(_0859_));
 sg13g2_buf_4 fanout831 (.X(net831),
    .A(_1653_));
 sg13g2_buf_4 fanout832 (.X(net832),
    .A(_1651_));
 sg13g2_buf_4 fanout833 (.X(net833),
    .A(_1651_));
 sg13g2_buf_4 fanout834 (.X(net834),
    .A(net835));
 sg13g2_buf_4 fanout835 (.X(net835),
    .A(net836));
 sg13g2_buf_4 fanout836 (.X(net836),
    .A(_1635_));
 sg13g2_buf_4 fanout837 (.X(net837),
    .A(_1635_));
 sg13g2_buf_1 fanout838 (.A(_1635_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(net840),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(net842),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(net844),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(net844),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_1634_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(net853),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(net853),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(net848),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(net849),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(net853),
    .X(net849));
 sg13g2_buf_4 fanout850 (.X(net850),
    .A(net852));
 sg13g2_buf_2 fanout851 (.A(net852),
    .X(net851));
 sg13g2_buf_4 fanout852 (.X(net852),
    .A(net853));
 sg13g2_buf_1 fanout853 (.A(_1632_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(net858),
    .X(net854));
 sg13g2_buf_4 fanout855 (.X(net855),
    .A(net856));
 sg13g2_buf_4 fanout856 (.X(net856),
    .A(net857));
 sg13g2_buf_2 fanout857 (.A(net858),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_1631_),
    .X(net858));
 sg13g2_buf_4 fanout859 (.X(net859),
    .A(net861));
 sg13g2_buf_2 fanout860 (.A(net861),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_1631_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_0882_),
    .X(net862));
 sg13g2_buf_4 fanout863 (.X(net863),
    .A(_0815_));
 sg13g2_buf_2 fanout864 (.A(_0765_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_0765_),
    .X(net865));
 sg13g2_buf_4 fanout866 (.X(net866),
    .A(_1654_));
 sg13g2_buf_2 fanout867 (.A(_1654_),
    .X(net867));
 sg13g2_buf_4 fanout868 (.X(net868),
    .A(net869));
 sg13g2_buf_4 fanout869 (.X(net869),
    .A(_1641_));
 sg13g2_buf_4 fanout870 (.X(net870),
    .A(_1630_));
 sg13g2_buf_4 fanout871 (.X(net871),
    .A(net872));
 sg13g2_buf_4 fanout872 (.X(net872),
    .A(_1629_));
 sg13g2_buf_2 fanout873 (.A(net874),
    .X(net873));
 sg13g2_buf_4 fanout874 (.X(net874),
    .A(_0760_));
 sg13g2_buf_2 fanout875 (.A(net877),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(net877),
    .X(net876));
 sg13g2_buf_4 fanout877 (.X(net877),
    .A(_0759_));
 sg13g2_buf_4 fanout878 (.X(net878),
    .A(_1594_));
 sg13g2_buf_4 fanout879 (.X(net879),
    .A(net880));
 sg13g2_buf_2 fanout880 (.A(_1593_),
    .X(net880));
 sg13g2_buf_4 fanout881 (.X(net881),
    .A(_1574_));
 sg13g2_buf_4 fanout882 (.X(net882),
    .A(net883));
 sg13g2_buf_2 fanout883 (.A(_0810_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_0758_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(net886),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_0470_),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(net888),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(_1690_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(net890),
    .X(net889));
 sg13g2_buf_4 fanout890 (.X(net890),
    .A(_1689_));
 sg13g2_buf_2 fanout891 (.A(_1689_),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(net895),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(net894),
    .X(net893));
 sg13g2_buf_1 fanout894 (.A(net895),
    .X(net894));
 sg13g2_buf_1 fanout895 (.A(net896),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(_0754_),
    .X(net896));
 sg13g2_buf_4 fanout897 (.X(net897),
    .A(net898));
 sg13g2_buf_2 fanout898 (.A(net899),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(_0753_),
    .X(net899));
 sg13g2_buf_4 fanout900 (.X(net900),
    .A(_1724_));
 sg13g2_buf_2 fanout901 (.A(_1724_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(net903),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(net904),
    .X(net903));
 sg13g2_buf_4 fanout904 (.X(net904),
    .A(_1723_));
 sg13g2_buf_2 fanout905 (.A(net906),
    .X(net905));
 sg13g2_buf_4 fanout906 (.X(net906),
    .A(_1713_));
 sg13g2_buf_4 fanout907 (.X(net907),
    .A(net910));
 sg13g2_buf_4 fanout908 (.X(net908),
    .A(net909));
 sg13g2_buf_2 fanout909 (.A(net910),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(_1712_),
    .X(net910));
 sg13g2_buf_4 fanout911 (.X(net911),
    .A(_1667_));
 sg13g2_buf_2 fanout912 (.A(_1667_),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(net914),
    .X(net913));
 sg13g2_buf_4 fanout914 (.X(net914),
    .A(_1578_));
 sg13g2_buf_4 fanout915 (.X(net915),
    .A(net916));
 sg13g2_buf_4 fanout916 (.X(net916),
    .A(_1577_));
 sg13g2_buf_2 fanout917 (.A(net920),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(net920),
    .X(net918));
 sg13g2_buf_4 fanout919 (.X(net919),
    .A(net920));
 sg13g2_buf_4 fanout920 (.X(net920),
    .A(_1570_));
 sg13g2_buf_2 fanout921 (.A(net922),
    .X(net921));
 sg13g2_buf_1 fanout922 (.A(net924),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(net924),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(_0813_),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(_0787_),
    .X(net925));
 sg13g2_buf_4 fanout926 (.X(net926),
    .A(_0770_));
 sg13g2_buf_2 fanout927 (.A(_0770_),
    .X(net927));
 sg13g2_buf_4 fanout928 (.X(net928),
    .A(_0768_));
 sg13g2_buf_2 fanout929 (.A(_0768_),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(net931),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(_1666_),
    .X(net931));
 sg13g2_buf_4 fanout932 (.X(net932),
    .A(_1666_));
 sg13g2_buf_4 fanout933 (.X(net933),
    .A(net934));
 sg13g2_buf_4 fanout934 (.X(net934),
    .A(_1571_));
 sg13g2_buf_4 fanout935 (.X(net935),
    .A(net936));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(_1540_));
 sg13g2_buf_4 fanout937 (.X(net937),
    .A(_1537_));
 sg13g2_buf_4 fanout938 (.X(net938),
    .A(_1536_));
 sg13g2_buf_4 fanout939 (.X(net939),
    .A(net940));
 sg13g2_buf_4 fanout940 (.X(net940),
    .A(net941));
 sg13g2_buf_4 fanout941 (.X(net941),
    .A(_1527_));
 sg13g2_buf_2 fanout942 (.A(\hvsync_gen.vpos[9] ),
    .X(net942));
 sg13g2_buf_4 fanout943 (.X(net943),
    .A(net137));
 sg13g2_buf_2 fanout944 (.A(net945),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(\hvsync_gen.vpos[6] ),
    .X(net945));
 sg13g2_buf_4 fanout946 (.X(net946),
    .A(net947));
 sg13g2_buf_4 fanout947 (.X(net947),
    .A(\hvsync_gen.vpos[5] ));
 sg13g2_buf_4 fanout948 (.X(net948),
    .A(net950));
 sg13g2_buf_4 fanout949 (.X(net949),
    .A(net950));
 sg13g2_buf_2 fanout950 (.A(\hvsync_gen.vpos[4] ),
    .X(net950));
 sg13g2_buf_4 fanout951 (.X(net951),
    .A(net959));
 sg13g2_buf_2 fanout952 (.A(net959),
    .X(net952));
 sg13g2_buf_4 fanout953 (.X(net953),
    .A(net956));
 sg13g2_buf_2 fanout954 (.A(net956),
    .X(net954));
 sg13g2_buf_1 fanout955 (.A(net956),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(net959),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(net959),
    .X(net957));
 sg13g2_buf_1 fanout958 (.A(net959),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(\hvsync_gen.vpos[3] ),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(net273),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(song_loops),
    .X(net961));
 sg13g2_buf_4 fanout962 (.X(net962),
    .A(net963));
 sg13g2_buf_2 fanout963 (.A(net234),
    .X(net963));
 sg13g2_buf_4 fanout964 (.X(net964),
    .A(\nyanframe[0] ));
 sg13g2_buf_1 fanout965 (.A(net966),
    .X(net965));
 sg13g2_buf_4 fanout966 (.X(net966),
    .A(\nyanframe[0] ));
 sg13g2_buf_2 fanout967 (.A(net968),
    .X(net967));
 sg13g2_buf_4 fanout968 (.X(net968),
    .A(\hvsync_gen.hpos[8] ));
 sg13g2_buf_2 fanout969 (.A(\hvsync_gen.hpos[7] ),
    .X(net969));
 sg13g2_buf_4 fanout970 (.X(net970),
    .A(net275));
 sg13g2_buf_2 fanout971 (.A(\hvsync_gen.hpos[5] ),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(net973),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(\hvsync_gen.hpos[4] ),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(net976),
    .X(net974));
 sg13g2_buf_1 fanout975 (.A(net976),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(\songpos[7] ),
    .X(net976));
 sg13g2_buf_4 fanout977 (.X(net977),
    .A(\songpos[6] ));
 sg13g2_buf_4 fanout978 (.X(net978),
    .A(\songpos[5] ));
 sg13g2_buf_2 fanout979 (.A(\songpos[5] ),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(net981),
    .X(net980));
 sg13g2_buf_1 fanout981 (.A(net982),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(net984),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(net984),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(net985),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(\songpos[4] ),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(net987),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(net991),
    .X(net987));
 sg13g2_buf_4 fanout988 (.X(net988),
    .A(net991));
 sg13g2_buf_2 fanout989 (.A(net990),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(net991),
    .X(net990));
 sg13g2_buf_1 fanout991 (.A(\songpos[3] ),
    .X(net991));
 sg13g2_buf_4 fanout992 (.X(net992),
    .A(net993));
 sg13g2_buf_2 fanout993 (.A(net994),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(net996),
    .X(net994));
 sg13g2_buf_4 fanout995 (.X(net995),
    .A(net996));
 sg13g2_buf_2 fanout996 (.A(\songpos[2] ),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(net998),
    .X(net997));
 sg13g2_buf_4 fanout998 (.X(net998),
    .A(net999));
 sg13g2_buf_2 fanout999 (.A(net1000),
    .X(net999));
 sg13g2_buf_4 fanout1000 (.X(net1000),
    .A(\songpos[1] ));
 sg13g2_buf_4 fanout1001 (.X(net1001),
    .A(net1003));
 sg13g2_buf_1 fanout1002 (.A(net1003),
    .X(net1002));
 sg13g2_buf_4 fanout1003 (.X(net1003),
    .A(\songpos[0] ));
 sg13g2_buf_2 fanout1004 (.A(net1005),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(\songpos[0] ),
    .X(net1005));
 sg13g2_buf_4 fanout1006 (.X(net1006),
    .A(net1007));
 sg13g2_buf_4 fanout1007 (.X(net1007),
    .A(net1010));
 sg13g2_buf_4 fanout1008 (.X(net1008),
    .A(net1009));
 sg13g2_buf_4 fanout1009 (.X(net1009),
    .A(net1010));
 sg13g2_buf_4 fanout1010 (.X(net1010),
    .A(rst_n));
 sg13g2_buf_4 fanout1011 (.X(net1011),
    .A(net1013));
 sg13g2_buf_4 fanout1012 (.X(net1012),
    .A(net1013));
 sg13g2_buf_2 fanout1013 (.A(net1014),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(rst_n),
    .X(net1014));
 sg13g2_buf_4 fanout1015 (.X(net1015),
    .A(net1018));
 sg13g2_buf_4 fanout1016 (.X(net1016),
    .A(net1018));
 sg13g2_buf_4 fanout1017 (.X(net1017),
    .A(net1018));
 sg13g2_buf_2 fanout1018 (.A(net1019),
    .X(net1018));
 sg13g2_buf_4 fanout1019 (.X(net1019),
    .A(net1022));
 sg13g2_buf_4 fanout1020 (.X(net1020),
    .A(net1022));
 sg13g2_buf_2 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_4 fanout1022 (.X(net1022),
    .A(rst_n));
 sg13g2_tielo tt_um_a1k0n_nyancat_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0042_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0038_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0896_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0095_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0041_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0080_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold7 (.A(_2185_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0175_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0043_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0068_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0040_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0176_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold13 (.A(\bass_pha[14] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0126_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0058_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0103_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold17 (.A(\sqr_pha[1] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0135_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold19 (.A(\audio_pwm_accum[0] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold20 (.A(\audio_pwm_accum_next[0] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold21 (.A(\bass_pha[13] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0125_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0048_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0063_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0045_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0049_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0052_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0047_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold29 (.A(\sqr_pha[8] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold30 (.A(\bass_pha[9] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0121_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0044_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0059_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold34 (.A(\bass_pha[12] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0124_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0053_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0098_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0046_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold39 (.A(\sqr_pha[12] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0146_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0056_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0101_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold43 (.A(\sqr_pha[0] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0050_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0065_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold46 (.A(\sqr_pha[11] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold47 (.A(_1248_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0022_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0127_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold50 (.A(\sqr_pha[9] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0055_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0100_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold53 (.A(\sin[0] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold54 (.A(\sqr_pha[10] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold55 (.A(\sqr_pha[2] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0136_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold57 (.A(\sqr_pha[5] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0139_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0051_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold60 (.A(\bass_pha[2] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0114_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0054_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0099_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold64 (.A(\bass_pha[0] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0112_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold66 (.A(\frame_count[7] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0087_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold68 (.A(\cos[6] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold69 (.A(\bass_pha[6] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold70 (.A(\bass_pha[11] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0123_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold72 (.A(\hvsync_gen.vpos[7] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold73 (.A(\kick_osci[1] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0154_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold75 (.A(\kick_osci[2] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold76 (.A(\bass_pha[3] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold77 (.A(\frame_count[3] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0876_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0083_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold80 (.A(\bass_pha[1] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold81 (.A(\bass_pha[5] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold82 (.A(\bass_pha[10] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0122_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold84 (.A(\sqr_pha[4] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0138_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold86 (.A(\sqr_vol[0] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0147_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold88 (.A(\bass_pha[8] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold89 (.A(\line_lfsr[1] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0089_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold91 (.A(\bass_vol[0] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold92 (.A(_1076_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0128_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold94 (.A(\bass_pha[4] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold95 (.A(\bass_pha[7] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold96 (.A(\sqr_pha[6] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold97 (.A(\line_lfsr[3] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0091_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold99 (.A(\kick_osci[5] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0057_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold101 (.A(\kick_osci[0] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold102 (.A(_1299_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold103 (.A(\line_lfsr[5] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0093_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold105 (.A(\line_lfsr[2] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold106 (.A(\kick_osci[3] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold107 (.A(\sqr_pha[7] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold108 (.A(\kick_ctr[1] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0853_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold110 (.A(\audio_sample_lpf[8] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0170_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold112 (.A(\frame_count[6] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0086_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold114 (.A(\frame_count[2] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0082_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold116 (.A(\line_lfsr[4] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0890_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0033_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0079_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold120 (.A(\line_lfsr[6] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0094_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold122 (.A(\bass_vol[5] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0133_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0037_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold125 (.A(\audio_sample_lpf[0] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0162_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold127 (.A(\frame_count[1] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0081_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold129 (.A(\sample_beat_ctr[1] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold130 (.A(_1489_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0173_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold132 (.A(\bass_vol[1] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold133 (.A(\sample_beat_ctr[2] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold134 (.A(_1491_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold135 (.A(\audio_sample_lpf[2] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0164_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold137 (.A(\nyan_x_offset[1] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold138 (.A(\frame_count[5] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0878_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold140 (.A(\audio_sample_lpf[4] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold141 (.A(\audio_pwm_accum[1] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0723_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold143 (.A(\nyan_x_offset[2] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold144 (.A(\sample_beat_ctr[0] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold145 (.A(\kick_osci[4] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold146 (.A(\audio_sample_lpf[1] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0163_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold148 (.A(\bass_vol[4] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold149 (.A(\nyan_x_offset[0] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold150 (.A(\kick_osci[8] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0161_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold152 (.A(\audio_sample_lpf[9] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0171_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0009_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold155 (.A(_1296_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold156 (.A(\audio_sample_lpf[6] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold157 (.A(\nyanframe[2] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0900_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0097_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold160 (.A(\line_lfsr[0] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold161 (.A(\kick_osci[7] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0160_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold163 (.A(\audio_sample_lpf[5] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold164 (.A(\frame_count[4] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold165 (.A(\sqr_vol[3] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0150_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold167 (.A(\audio_pwm_accum[5] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold168 (.A(\audio_pwm_accum_next[5] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold169 (.A(\sin[6] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0111_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold171 (.A(\sqr_vol[2] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold172 (.A(\sqr_pha[3] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold173 (.A(\bass_vol[2] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold174 (.A(\audio_sample_lpf[7] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold175 (.A(\sqr_vol[5] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold176 (.A(_1297_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold177 (.A(\audio_pwm_accum[2] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold178 (.A(\audio_pwm_accum_next[2] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold179 (.A(\audio_pwm_accum[7] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold180 (.A(\audio_pwm_accum_next[7] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold181 (.A(\audio_pwm_accum[3] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0728_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold183 (.A(\audio_pwm_accum[8] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold184 (.A(\audio_pwm_accum_next[8] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold185 (.A(\bass_vol[3] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0131_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold187 (.A(\hvsync_gen.vpos[1] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold188 (.A(\hvsync_gen.hpos[1] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold189 (.A(\audio_pwm_accum[4] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold190 (.A(\sqr_vol[1] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0148_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0036_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0181_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold194 (.A(\audio_pwm_accum[9] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold195 (.A(\nyan_x_offset[4] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0031_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0096_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold198 (.A(\hvsync_gen.hpos[2] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0008_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold200 (.A(\audio_pwm_accum[6] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0736_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0738_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold203 (.A(\audio_pwm_accum_next[6] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold204 (.A(\audio_sample_lpf[3] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold205 (.A(\nyan_x_offset[3] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold206 (.A(\kick_osci[6] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold207 (.A(\hvsync_gen.vpos[8] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold208 (.A(\hvsync_gen.vpos[2] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold209 (.A(_1501_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold210 (.A(\hvsync_gen.hpos[6] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0030_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold212 (.A(\hvsync_gen.hpos[3] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold213 (.A(\frame_count[4] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold214 (.A(\nyan_x_offset[0] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold215 (.A(\bass_vol[2] ),
    .X(net280));
 sg13g2_antennanp ANTENNA_1 (.A(_0006_));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(_0006_));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_antennanp ANTENNA_6 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_4 FILLER_11_105 ();
 sg13g2_fill_1 FILLER_11_109 ();
 sg13g2_fill_2 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_131 ();
 sg13g2_decap_8 FILLER_11_138 ();
 sg13g2_decap_8 FILLER_11_145 ();
 sg13g2_decap_8 FILLER_11_152 ();
 sg13g2_decap_8 FILLER_11_159 ();
 sg13g2_decap_8 FILLER_11_166 ();
 sg13g2_decap_8 FILLER_11_173 ();
 sg13g2_decap_8 FILLER_11_180 ();
 sg13g2_decap_8 FILLER_11_187 ();
 sg13g2_decap_8 FILLER_11_194 ();
 sg13g2_decap_8 FILLER_11_201 ();
 sg13g2_decap_8 FILLER_11_208 ();
 sg13g2_decap_8 FILLER_11_215 ();
 sg13g2_decap_8 FILLER_11_222 ();
 sg13g2_decap_8 FILLER_11_229 ();
 sg13g2_decap_8 FILLER_11_236 ();
 sg13g2_decap_8 FILLER_11_243 ();
 sg13g2_decap_8 FILLER_11_250 ();
 sg13g2_decap_8 FILLER_11_257 ();
 sg13g2_decap_8 FILLER_11_264 ();
 sg13g2_decap_8 FILLER_11_271 ();
 sg13g2_decap_8 FILLER_11_278 ();
 sg13g2_decap_8 FILLER_11_285 ();
 sg13g2_decap_8 FILLER_11_292 ();
 sg13g2_decap_8 FILLER_11_299 ();
 sg13g2_decap_8 FILLER_11_306 ();
 sg13g2_decap_8 FILLER_11_313 ();
 sg13g2_decap_8 FILLER_11_320 ();
 sg13g2_decap_8 FILLER_11_327 ();
 sg13g2_decap_8 FILLER_11_334 ();
 sg13g2_decap_8 FILLER_11_341 ();
 sg13g2_decap_8 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_355 ();
 sg13g2_decap_8 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_369 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_4 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_43 ();
 sg13g2_decap_8 FILLER_12_50 ();
 sg13g2_decap_8 FILLER_12_57 ();
 sg13g2_decap_8 FILLER_12_64 ();
 sg13g2_decap_8 FILLER_12_71 ();
 sg13g2_decap_8 FILLER_12_78 ();
 sg13g2_decap_8 FILLER_12_85 ();
 sg13g2_decap_8 FILLER_12_92 ();
 sg13g2_fill_1 FILLER_12_99 ();
 sg13g2_fill_1 FILLER_12_110 ();
 sg13g2_decap_4 FILLER_12_123 ();
 sg13g2_decap_8 FILLER_12_144 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_8 FILLER_12_158 ();
 sg13g2_decap_8 FILLER_12_165 ();
 sg13g2_decap_8 FILLER_12_172 ();
 sg13g2_decap_8 FILLER_12_179 ();
 sg13g2_decap_8 FILLER_12_186 ();
 sg13g2_decap_8 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_214 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_4 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_32 ();
 sg13g2_fill_1 FILLER_13_38 ();
 sg13g2_decap_8 FILLER_13_52 ();
 sg13g2_decap_8 FILLER_13_59 ();
 sg13g2_decap_8 FILLER_13_66 ();
 sg13g2_decap_8 FILLER_13_73 ();
 sg13g2_decap_4 FILLER_13_80 ();
 sg13g2_fill_1 FILLER_13_84 ();
 sg13g2_fill_1 FILLER_13_125 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_fill_2 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_69 ();
 sg13g2_decap_4 FILLER_14_76 ();
 sg13g2_fill_1 FILLER_14_80 ();
 sg13g2_fill_1 FILLER_14_107 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_194 ();
 sg13g2_decap_8 FILLER_14_201 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_215 ();
 sg13g2_decap_8 FILLER_14_222 ();
 sg13g2_decap_8 FILLER_14_229 ();
 sg13g2_decap_8 FILLER_14_236 ();
 sg13g2_decap_8 FILLER_14_243 ();
 sg13g2_decap_8 FILLER_14_250 ();
 sg13g2_decap_8 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_264 ();
 sg13g2_decap_8 FILLER_14_271 ();
 sg13g2_decap_8 FILLER_14_278 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_decap_8 FILLER_14_292 ();
 sg13g2_decap_8 FILLER_14_299 ();
 sg13g2_decap_8 FILLER_14_306 ();
 sg13g2_decap_8 FILLER_14_313 ();
 sg13g2_decap_8 FILLER_14_320 ();
 sg13g2_decap_8 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_35 ();
 sg13g2_fill_2 FILLER_15_44 ();
 sg13g2_decap_8 FILLER_15_61 ();
 sg13g2_decap_8 FILLER_15_68 ();
 sg13g2_decap_4 FILLER_15_75 ();
 sg13g2_fill_1 FILLER_15_105 ();
 sg13g2_fill_2 FILLER_15_147 ();
 sg13g2_fill_1 FILLER_15_158 ();
 sg13g2_fill_2 FILLER_15_164 ();
 sg13g2_fill_1 FILLER_15_166 ();
 sg13g2_fill_1 FILLER_15_186 ();
 sg13g2_fill_2 FILLER_15_213 ();
 sg13g2_fill_1 FILLER_15_215 ();
 sg13g2_decap_8 FILLER_15_220 ();
 sg13g2_decap_8 FILLER_15_227 ();
 sg13g2_decap_8 FILLER_15_234 ();
 sg13g2_decap_8 FILLER_15_241 ();
 sg13g2_decap_8 FILLER_15_248 ();
 sg13g2_decap_8 FILLER_15_255 ();
 sg13g2_decap_8 FILLER_15_262 ();
 sg13g2_decap_8 FILLER_15_269 ();
 sg13g2_decap_8 FILLER_15_276 ();
 sg13g2_decap_8 FILLER_15_283 ();
 sg13g2_decap_8 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_297 ();
 sg13g2_decap_8 FILLER_15_304 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_23 ();
 sg13g2_fill_2 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_44 ();
 sg13g2_decap_8 FILLER_16_71 ();
 sg13g2_decap_4 FILLER_16_78 ();
 sg13g2_fill_2 FILLER_16_82 ();
 sg13g2_fill_2 FILLER_16_100 ();
 sg13g2_fill_2 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_127 ();
 sg13g2_fill_2 FILLER_16_143 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_decap_8 FILLER_16_242 ();
 sg13g2_decap_8 FILLER_16_249 ();
 sg13g2_decap_8 FILLER_16_256 ();
 sg13g2_decap_8 FILLER_16_263 ();
 sg13g2_decap_8 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_277 ();
 sg13g2_decap_8 FILLER_16_284 ();
 sg13g2_decap_8 FILLER_16_291 ();
 sg13g2_decap_8 FILLER_16_298 ();
 sg13g2_decap_8 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_312 ();
 sg13g2_decap_8 FILLER_16_319 ();
 sg13g2_decap_8 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_340 ();
 sg13g2_decap_8 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_decap_8 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_11 ();
 sg13g2_fill_1 FILLER_17_17 ();
 sg13g2_fill_1 FILLER_17_45 ();
 sg13g2_fill_1 FILLER_17_54 ();
 sg13g2_fill_2 FILLER_17_116 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_fill_2 FILLER_17_180 ();
 sg13g2_fill_2 FILLER_17_208 ();
 sg13g2_fill_1 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_236 ();
 sg13g2_decap_8 FILLER_17_243 ();
 sg13g2_decap_8 FILLER_17_250 ();
 sg13g2_decap_8 FILLER_17_257 ();
 sg13g2_decap_8 FILLER_17_264 ();
 sg13g2_decap_8 FILLER_17_271 ();
 sg13g2_decap_8 FILLER_17_278 ();
 sg13g2_decap_8 FILLER_17_285 ();
 sg13g2_decap_8 FILLER_17_292 ();
 sg13g2_decap_8 FILLER_17_299 ();
 sg13g2_decap_8 FILLER_17_306 ();
 sg13g2_decap_8 FILLER_17_313 ();
 sg13g2_decap_8 FILLER_17_320 ();
 sg13g2_decap_8 FILLER_17_327 ();
 sg13g2_decap_8 FILLER_17_334 ();
 sg13g2_decap_8 FILLER_17_341 ();
 sg13g2_decap_8 FILLER_17_348 ();
 sg13g2_decap_8 FILLER_17_355 ();
 sg13g2_decap_8 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_4 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_62 ();
 sg13g2_fill_1 FILLER_18_64 ();
 sg13g2_fill_2 FILLER_18_100 ();
 sg13g2_fill_1 FILLER_18_102 ();
 sg13g2_fill_2 FILLER_18_121 ();
 sg13g2_fill_1 FILLER_18_165 ();
 sg13g2_fill_1 FILLER_18_188 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_8 FILLER_18_232 ();
 sg13g2_decap_8 FILLER_18_239 ();
 sg13g2_decap_8 FILLER_18_246 ();
 sg13g2_decap_8 FILLER_18_253 ();
 sg13g2_decap_8 FILLER_18_260 ();
 sg13g2_decap_8 FILLER_18_267 ();
 sg13g2_decap_8 FILLER_18_274 ();
 sg13g2_decap_8 FILLER_18_281 ();
 sg13g2_decap_8 FILLER_18_288 ();
 sg13g2_decap_8 FILLER_18_295 ();
 sg13g2_decap_8 FILLER_18_302 ();
 sg13g2_decap_8 FILLER_18_309 ();
 sg13g2_decap_8 FILLER_18_316 ();
 sg13g2_decap_8 FILLER_18_323 ();
 sg13g2_decap_8 FILLER_18_330 ();
 sg13g2_decap_8 FILLER_18_337 ();
 sg13g2_decap_8 FILLER_18_344 ();
 sg13g2_decap_8 FILLER_18_351 ();
 sg13g2_decap_8 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_365 ();
 sg13g2_decap_8 FILLER_18_372 ();
 sg13g2_decap_8 FILLER_18_379 ();
 sg13g2_decap_8 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_57 ();
 sg13g2_fill_2 FILLER_19_98 ();
 sg13g2_fill_2 FILLER_19_131 ();
 sg13g2_fill_1 FILLER_19_155 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_2 FILLER_19_190 ();
 sg13g2_fill_1 FILLER_19_201 ();
 sg13g2_decap_8 FILLER_19_229 ();
 sg13g2_decap_8 FILLER_19_236 ();
 sg13g2_decap_8 FILLER_19_243 ();
 sg13g2_decap_8 FILLER_19_250 ();
 sg13g2_decap_8 FILLER_19_257 ();
 sg13g2_decap_8 FILLER_19_264 ();
 sg13g2_decap_8 FILLER_19_271 ();
 sg13g2_decap_8 FILLER_19_278 ();
 sg13g2_decap_8 FILLER_19_285 ();
 sg13g2_decap_8 FILLER_19_292 ();
 sg13g2_decap_8 FILLER_19_299 ();
 sg13g2_decap_8 FILLER_19_306 ();
 sg13g2_decap_8 FILLER_19_313 ();
 sg13g2_decap_8 FILLER_19_320 ();
 sg13g2_decap_8 FILLER_19_327 ();
 sg13g2_decap_8 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_341 ();
 sg13g2_decap_8 FILLER_19_348 ();
 sg13g2_decap_8 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_362 ();
 sg13g2_decap_8 FILLER_19_369 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_9 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_2 FILLER_20_79 ();
 sg13g2_fill_1 FILLER_20_125 ();
 sg13g2_fill_1 FILLER_20_149 ();
 sg13g2_fill_1 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_234 ();
 sg13g2_decap_8 FILLER_20_241 ();
 sg13g2_decap_8 FILLER_20_248 ();
 sg13g2_decap_8 FILLER_20_255 ();
 sg13g2_decap_8 FILLER_20_262 ();
 sg13g2_decap_8 FILLER_20_269 ();
 sg13g2_decap_8 FILLER_20_276 ();
 sg13g2_decap_8 FILLER_20_283 ();
 sg13g2_decap_8 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_297 ();
 sg13g2_decap_8 FILLER_20_304 ();
 sg13g2_decap_8 FILLER_20_311 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_8 FILLER_20_325 ();
 sg13g2_decap_8 FILLER_20_332 ();
 sg13g2_decap_8 FILLER_20_339 ();
 sg13g2_decap_8 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_353 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_11 ();
 sg13g2_fill_1 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_89 ();
 sg13g2_fill_2 FILLER_21_104 ();
 sg13g2_fill_1 FILLER_21_106 ();
 sg13g2_fill_1 FILLER_21_117 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_decap_8 FILLER_21_227 ();
 sg13g2_decap_8 FILLER_21_234 ();
 sg13g2_decap_8 FILLER_21_241 ();
 sg13g2_decap_8 FILLER_21_248 ();
 sg13g2_decap_8 FILLER_21_255 ();
 sg13g2_decap_8 FILLER_21_262 ();
 sg13g2_decap_8 FILLER_21_269 ();
 sg13g2_decap_8 FILLER_21_276 ();
 sg13g2_decap_8 FILLER_21_283 ();
 sg13g2_decap_8 FILLER_21_290 ();
 sg13g2_decap_8 FILLER_21_297 ();
 sg13g2_decap_8 FILLER_21_304 ();
 sg13g2_decap_8 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_318 ();
 sg13g2_decap_8 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_21_339 ();
 sg13g2_decap_8 FILLER_21_346 ();
 sg13g2_decap_8 FILLER_21_353 ();
 sg13g2_decap_8 FILLER_21_360 ();
 sg13g2_decap_8 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_374 ();
 sg13g2_decap_8 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_fill_1 FILLER_22_65 ();
 sg13g2_fill_2 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_107 ();
 sg13g2_fill_2 FILLER_22_116 ();
 sg13g2_fill_1 FILLER_22_118 ();
 sg13g2_fill_2 FILLER_22_128 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_fill_2 FILLER_22_204 ();
 sg13g2_decap_8 FILLER_22_214 ();
 sg13g2_decap_8 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_235 ();
 sg13g2_decap_8 FILLER_22_242 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_256 ();
 sg13g2_decap_8 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_2 FILLER_23_28 ();
 sg13g2_fill_2 FILLER_23_43 ();
 sg13g2_fill_1 FILLER_23_45 ();
 sg13g2_decap_4 FILLER_23_100 ();
 sg13g2_decap_4 FILLER_23_108 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_fill_1 FILLER_23_118 ();
 sg13g2_fill_1 FILLER_23_127 ();
 sg13g2_decap_4 FILLER_23_158 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_fill_2 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_decap_8 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_263 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_305 ();
 sg13g2_fill_1 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_23 ();
 sg13g2_decap_4 FILLER_24_30 ();
 sg13g2_fill_2 FILLER_24_34 ();
 sg13g2_fill_2 FILLER_24_64 ();
 sg13g2_fill_2 FILLER_24_88 ();
 sg13g2_decap_4 FILLER_24_95 ();
 sg13g2_fill_1 FILLER_24_104 ();
 sg13g2_fill_2 FILLER_24_115 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_1 FILLER_24_125 ();
 sg13g2_fill_2 FILLER_24_151 ();
 sg13g2_fill_1 FILLER_24_153 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_decap_8 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_256 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_284 ();
 sg13g2_decap_8 FILLER_24_291 ();
 sg13g2_decap_4 FILLER_24_298 ();
 sg13g2_decap_4 FILLER_24_307 ();
 sg13g2_fill_1 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_4 FILLER_25_26 ();
 sg13g2_fill_2 FILLER_25_83 ();
 sg13g2_fill_2 FILLER_25_90 ();
 sg13g2_fill_2 FILLER_25_97 ();
 sg13g2_fill_1 FILLER_25_109 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_fill_2 FILLER_25_177 ();
 sg13g2_fill_1 FILLER_25_188 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_4 FILLER_25_280 ();
 sg13g2_fill_2 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_327 ();
 sg13g2_decap_4 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_78 ();
 sg13g2_fill_2 FILLER_26_82 ();
 sg13g2_fill_1 FILLER_26_125 ();
 sg13g2_fill_1 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_181 ();
 sg13g2_fill_2 FILLER_26_187 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_fill_2 FILLER_26_219 ();
 sg13g2_fill_2 FILLER_26_226 ();
 sg13g2_decap_8 FILLER_26_237 ();
 sg13g2_decap_8 FILLER_26_244 ();
 sg13g2_decap_8 FILLER_26_251 ();
 sg13g2_decap_8 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_265 ();
 sg13g2_decap_8 FILLER_26_272 ();
 sg13g2_fill_2 FILLER_26_279 ();
 sg13g2_fill_2 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_299 ();
 sg13g2_fill_2 FILLER_26_315 ();
 sg13g2_fill_2 FILLER_26_325 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_36 ();
 sg13g2_fill_2 FILLER_27_68 ();
 sg13g2_fill_1 FILLER_27_70 ();
 sg13g2_fill_1 FILLER_27_76 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_95 ();
 sg13g2_fill_2 FILLER_27_117 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_fill_2 FILLER_27_148 ();
 sg13g2_fill_1 FILLER_27_150 ();
 sg13g2_fill_2 FILLER_27_185 ();
 sg13g2_fill_2 FILLER_27_216 ();
 sg13g2_decap_8 FILLER_27_223 ();
 sg13g2_decap_8 FILLER_27_230 ();
 sg13g2_decap_8 FILLER_27_237 ();
 sg13g2_decap_8 FILLER_27_244 ();
 sg13g2_decap_8 FILLER_27_251 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_260 ();
 sg13g2_fill_2 FILLER_27_314 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_fill_2 FILLER_27_323 ();
 sg13g2_fill_2 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_341 ();
 sg13g2_fill_2 FILLER_27_358 ();
 sg13g2_fill_1 FILLER_27_360 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_4 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_74 ();
 sg13g2_decap_4 FILLER_28_97 ();
 sg13g2_fill_1 FILLER_28_110 ();
 sg13g2_fill_2 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_131 ();
 sg13g2_decap_8 FILLER_28_145 ();
 sg13g2_decap_8 FILLER_28_152 ();
 sg13g2_decap_4 FILLER_28_159 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_249 ();
 sg13g2_decap_4 FILLER_28_256 ();
 sg13g2_fill_1 FILLER_28_268 ();
 sg13g2_fill_2 FILLER_28_277 ();
 sg13g2_fill_1 FILLER_28_279 ();
 sg13g2_decap_4 FILLER_28_292 ();
 sg13g2_fill_2 FILLER_28_316 ();
 sg13g2_fill_1 FILLER_28_336 ();
 sg13g2_fill_2 FILLER_28_356 ();
 sg13g2_decap_8 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_4 ();
 sg13g2_decap_4 FILLER_29_69 ();
 sg13g2_fill_2 FILLER_29_73 ();
 sg13g2_fill_1 FILLER_29_103 ();
 sg13g2_decap_8 FILLER_29_116 ();
 sg13g2_decap_4 FILLER_29_123 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_155 ();
 sg13g2_decap_4 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_166 ();
 sg13g2_decap_4 FILLER_29_172 ();
 sg13g2_fill_2 FILLER_29_176 ();
 sg13g2_fill_2 FILLER_29_187 ();
 sg13g2_fill_1 FILLER_29_189 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_fill_1 FILLER_29_208 ();
 sg13g2_decap_4 FILLER_29_226 ();
 sg13g2_decap_4 FILLER_29_243 ();
 sg13g2_decap_4 FILLER_29_251 ();
 sg13g2_fill_1 FILLER_29_255 ();
 sg13g2_decap_8 FILLER_29_276 ();
 sg13g2_fill_2 FILLER_29_283 ();
 sg13g2_decap_8 FILLER_29_298 ();
 sg13g2_decap_4 FILLER_29_318 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_fill_1 FILLER_29_343 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_2 FILLER_30_29 ();
 sg13g2_fill_2 FILLER_30_80 ();
 sg13g2_decap_8 FILLER_30_102 ();
 sg13g2_decap_4 FILLER_30_109 ();
 sg13g2_fill_1 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_170 ();
 sg13g2_decap_4 FILLER_30_177 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_fill_1 FILLER_30_246 ();
 sg13g2_fill_1 FILLER_30_289 ();
 sg13g2_fill_2 FILLER_30_304 ();
 sg13g2_fill_1 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_fill_2 FILLER_30_324 ();
 sg13g2_fill_2 FILLER_30_336 ();
 sg13g2_fill_1 FILLER_30_338 ();
 sg13g2_decap_4 FILLER_30_349 ();
 sg13g2_fill_2 FILLER_30_353 ();
 sg13g2_fill_2 FILLER_30_359 ();
 sg13g2_decap_8 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_2 ();
 sg13g2_fill_1 FILLER_31_79 ();
 sg13g2_fill_2 FILLER_31_92 ();
 sg13g2_decap_4 FILLER_31_100 ();
 sg13g2_fill_1 FILLER_31_129 ();
 sg13g2_fill_2 FILLER_31_146 ();
 sg13g2_decap_8 FILLER_31_197 ();
 sg13g2_fill_2 FILLER_31_262 ();
 sg13g2_fill_1 FILLER_31_264 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_fill_1 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_328 ();
 sg13g2_fill_1 FILLER_31_330 ();
 sg13g2_fill_2 FILLER_31_339 ();
 sg13g2_fill_2 FILLER_31_356 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_71 ();
 sg13g2_fill_1 FILLER_32_73 ();
 sg13g2_fill_2 FILLER_32_89 ();
 sg13g2_fill_1 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_167 ();
 sg13g2_fill_2 FILLER_32_178 ();
 sg13g2_fill_1 FILLER_32_180 ();
 sg13g2_decap_8 FILLER_32_201 ();
 sg13g2_decap_4 FILLER_32_208 ();
 sg13g2_fill_1 FILLER_32_212 ();
 sg13g2_decap_4 FILLER_32_217 ();
 sg13g2_fill_2 FILLER_32_261 ();
 sg13g2_fill_1 FILLER_32_279 ();
 sg13g2_fill_2 FILLER_32_353 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_32_389 ();
 sg13g2_decap_8 FILLER_32_396 ();
 sg13g2_decap_4 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_fill_2 FILLER_33_82 ();
 sg13g2_fill_2 FILLER_33_97 ();
 sg13g2_fill_1 FILLER_33_99 ();
 sg13g2_fill_2 FILLER_33_136 ();
 sg13g2_fill_1 FILLER_33_138 ();
 sg13g2_decap_8 FILLER_33_222 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_decap_4 FILLER_33_242 ();
 sg13g2_fill_2 FILLER_33_246 ();
 sg13g2_decap_4 FILLER_33_253 ();
 sg13g2_fill_2 FILLER_33_257 ();
 sg13g2_fill_2 FILLER_33_271 ();
 sg13g2_fill_1 FILLER_33_290 ();
 sg13g2_decap_4 FILLER_33_299 ();
 sg13g2_decap_8 FILLER_33_316 ();
 sg13g2_decap_4 FILLER_33_323 ();
 sg13g2_fill_1 FILLER_33_327 ();
 sg13g2_fill_1 FILLER_33_338 ();
 sg13g2_fill_2 FILLER_33_367 ();
 sg13g2_fill_1 FILLER_33_369 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_1 FILLER_34_23 ();
 sg13g2_fill_1 FILLER_34_54 ();
 sg13g2_decap_8 FILLER_34_69 ();
 sg13g2_decap_8 FILLER_34_76 ();
 sg13g2_decap_4 FILLER_34_83 ();
 sg13g2_fill_2 FILLER_34_87 ();
 sg13g2_fill_2 FILLER_34_117 ();
 sg13g2_fill_1 FILLER_34_119 ();
 sg13g2_fill_1 FILLER_34_124 ();
 sg13g2_fill_2 FILLER_34_130 ();
 sg13g2_fill_1 FILLER_34_132 ();
 sg13g2_fill_1 FILLER_34_138 ();
 sg13g2_fill_2 FILLER_34_155 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_fill_1 FILLER_34_162 ();
 sg13g2_fill_2 FILLER_34_195 ();
 sg13g2_decap_4 FILLER_34_223 ();
 sg13g2_fill_2 FILLER_34_227 ();
 sg13g2_decap_4 FILLER_34_243 ();
 sg13g2_decap_4 FILLER_34_260 ();
 sg13g2_fill_1 FILLER_34_264 ();
 sg13g2_fill_2 FILLER_34_286 ();
 sg13g2_fill_2 FILLER_34_299 ();
 sg13g2_fill_1 FILLER_34_301 ();
 sg13g2_fill_2 FILLER_34_310 ();
 sg13g2_fill_1 FILLER_34_312 ();
 sg13g2_fill_1 FILLER_34_321 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_fill_2 FILLER_35_29 ();
 sg13g2_fill_2 FILLER_35_52 ();
 sg13g2_decap_8 FILLER_35_67 ();
 sg13g2_fill_1 FILLER_35_79 ();
 sg13g2_fill_2 FILLER_35_108 ();
 sg13g2_fill_1 FILLER_35_110 ();
 sg13g2_fill_2 FILLER_35_116 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_decap_4 FILLER_35_136 ();
 sg13g2_fill_2 FILLER_35_140 ();
 sg13g2_fill_1 FILLER_35_145 ();
 sg13g2_decap_8 FILLER_35_156 ();
 sg13g2_decap_8 FILLER_35_163 ();
 sg13g2_decap_4 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_178 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_fill_2 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_decap_8 FILLER_35_264 ();
 sg13g2_fill_2 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_273 ();
 sg13g2_fill_2 FILLER_35_278 ();
 sg13g2_fill_1 FILLER_35_280 ();
 sg13g2_fill_2 FILLER_35_295 ();
 sg13g2_fill_1 FILLER_35_297 ();
 sg13g2_fill_2 FILLER_35_312 ();
 sg13g2_decap_8 FILLER_35_335 ();
 sg13g2_fill_2 FILLER_35_342 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_fill_2 FILLER_35_371 ();
 sg13g2_fill_1 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_389 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_fill_1 FILLER_36_26 ();
 sg13g2_fill_2 FILLER_36_36 ();
 sg13g2_fill_1 FILLER_36_78 ();
 sg13g2_fill_2 FILLER_36_93 ();
 sg13g2_fill_1 FILLER_36_95 ();
 sg13g2_fill_2 FILLER_36_101 ();
 sg13g2_fill_1 FILLER_36_103 ();
 sg13g2_decap_4 FILLER_36_110 ();
 sg13g2_fill_2 FILLER_36_134 ();
 sg13g2_fill_2 FILLER_36_144 ();
 sg13g2_decap_4 FILLER_36_156 ();
 sg13g2_decap_4 FILLER_36_191 ();
 sg13g2_decap_8 FILLER_36_199 ();
 sg13g2_fill_2 FILLER_36_206 ();
 sg13g2_decap_4 FILLER_36_221 ();
 sg13g2_fill_1 FILLER_36_225 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_fill_1 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_247 ();
 sg13g2_decap_4 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_258 ();
 sg13g2_decap_4 FILLER_36_274 ();
 sg13g2_fill_2 FILLER_36_310 ();
 sg13g2_fill_1 FILLER_36_312 ();
 sg13g2_decap_8 FILLER_36_326 ();
 sg13g2_decap_8 FILLER_36_333 ();
 sg13g2_decap_8 FILLER_36_346 ();
 sg13g2_fill_2 FILLER_36_353 ();
 sg13g2_fill_1 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_fill_1 FILLER_37_24 ();
 sg13g2_fill_2 FILLER_37_51 ();
 sg13g2_fill_2 FILLER_37_79 ();
 sg13g2_fill_1 FILLER_37_81 ();
 sg13g2_fill_2 FILLER_37_88 ();
 sg13g2_decap_4 FILLER_37_105 ();
 sg13g2_fill_2 FILLER_37_120 ();
 sg13g2_fill_2 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_135 ();
 sg13g2_fill_2 FILLER_37_166 ();
 sg13g2_fill_2 FILLER_37_192 ();
 sg13g2_fill_2 FILLER_37_204 ();
 sg13g2_fill_2 FILLER_37_211 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_decap_8 FILLER_37_219 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_4 FILLER_37_252 ();
 sg13g2_fill_1 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_262 ();
 sg13g2_fill_2 FILLER_37_286 ();
 sg13g2_fill_1 FILLER_37_288 ();
 sg13g2_fill_2 FILLER_37_330 ();
 sg13g2_fill_2 FILLER_37_337 ();
 sg13g2_decap_4 FILLER_37_349 ();
 sg13g2_decap_8 FILLER_37_383 ();
 sg13g2_decap_8 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_15 ();
 sg13g2_fill_1 FILLER_38_34 ();
 sg13g2_fill_2 FILLER_38_83 ();
 sg13g2_fill_1 FILLER_38_90 ();
 sg13g2_fill_2 FILLER_38_160 ();
 sg13g2_fill_2 FILLER_38_170 ();
 sg13g2_fill_2 FILLER_38_181 ();
 sg13g2_fill_2 FILLER_38_192 ();
 sg13g2_fill_1 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_211 ();
 sg13g2_fill_2 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_fill_1 FILLER_38_248 ();
 sg13g2_fill_2 FILLER_38_278 ();
 sg13g2_fill_2 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_297 ();
 sg13g2_decap_4 FILLER_38_304 ();
 sg13g2_fill_2 FILLER_38_351 ();
 sg13g2_fill_2 FILLER_38_361 ();
 sg13g2_fill_1 FILLER_38_363 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_fill_1 FILLER_39_26 ();
 sg13g2_fill_2 FILLER_39_35 ();
 sg13g2_fill_1 FILLER_39_80 ();
 sg13g2_fill_2 FILLER_39_95 ();
 sg13g2_fill_2 FILLER_39_146 ();
 sg13g2_fill_2 FILLER_39_214 ();
 sg13g2_fill_1 FILLER_39_216 ();
 sg13g2_decap_8 FILLER_39_226 ();
 sg13g2_fill_2 FILLER_39_233 ();
 sg13g2_fill_2 FILLER_39_243 ();
 sg13g2_fill_2 FILLER_39_258 ();
 sg13g2_fill_1 FILLER_39_266 ();
 sg13g2_fill_1 FILLER_39_280 ();
 sg13g2_fill_1 FILLER_39_316 ();
 sg13g2_fill_2 FILLER_39_323 ();
 sg13g2_fill_1 FILLER_39_325 ();
 sg13g2_fill_2 FILLER_39_336 ();
 sg13g2_fill_2 FILLER_39_366 ();
 sg13g2_fill_1 FILLER_39_368 ();
 sg13g2_decap_8 FILLER_39_391 ();
 sg13g2_decap_8 FILLER_39_398 ();
 sg13g2_decap_4 FILLER_39_405 ();
 sg13g2_fill_1 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_103 ();
 sg13g2_decap_4 FILLER_40_110 ();
 sg13g2_decap_4 FILLER_40_119 ();
 sg13g2_fill_2 FILLER_40_123 ();
 sg13g2_fill_2 FILLER_40_134 ();
 sg13g2_fill_2 FILLER_40_150 ();
 sg13g2_fill_1 FILLER_40_152 ();
 sg13g2_fill_2 FILLER_40_203 ();
 sg13g2_fill_1 FILLER_40_205 ();
 sg13g2_decap_4 FILLER_40_232 ();
 sg13g2_fill_2 FILLER_40_236 ();
 sg13g2_decap_8 FILLER_40_254 ();
 sg13g2_decap_4 FILLER_40_261 ();
 sg13g2_decap_4 FILLER_40_274 ();
 sg13g2_fill_1 FILLER_40_278 ();
 sg13g2_decap_4 FILLER_40_314 ();
 sg13g2_fill_2 FILLER_40_318 ();
 sg13g2_fill_2 FILLER_40_332 ();
 sg13g2_fill_1 FILLER_40_352 ();
 sg13g2_fill_2 FILLER_40_358 ();
 sg13g2_fill_2 FILLER_40_366 ();
 sg13g2_decap_8 FILLER_40_382 ();
 sg13g2_decap_8 FILLER_40_389 ();
 sg13g2_decap_8 FILLER_40_396 ();
 sg13g2_decap_4 FILLER_40_403 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_fill_2 FILLER_41_28 ();
 sg13g2_fill_1 FILLER_41_57 ();
 sg13g2_fill_2 FILLER_41_87 ();
 sg13g2_fill_2 FILLER_41_134 ();
 sg13g2_decap_8 FILLER_41_151 ();
 sg13g2_decap_8 FILLER_41_158 ();
 sg13g2_decap_4 FILLER_41_178 ();
 sg13g2_fill_2 FILLER_41_199 ();
 sg13g2_fill_2 FILLER_41_215 ();
 sg13g2_decap_8 FILLER_41_225 ();
 sg13g2_decap_8 FILLER_41_232 ();
 sg13g2_fill_2 FILLER_41_239 ();
 sg13g2_fill_1 FILLER_41_241 ();
 sg13g2_decap_8 FILLER_41_247 ();
 sg13g2_fill_2 FILLER_41_254 ();
 sg13g2_decap_4 FILLER_41_286 ();
 sg13g2_fill_1 FILLER_41_296 ();
 sg13g2_decap_4 FILLER_41_302 ();
 sg13g2_fill_1 FILLER_41_306 ();
 sg13g2_fill_1 FILLER_41_312 ();
 sg13g2_fill_2 FILLER_41_328 ();
 sg13g2_fill_1 FILLER_41_330 ();
 sg13g2_fill_2 FILLER_41_350 ();
 sg13g2_fill_1 FILLER_41_352 ();
 sg13g2_fill_2 FILLER_41_362 ();
 sg13g2_fill_1 FILLER_41_364 ();
 sg13g2_fill_1 FILLER_41_370 ();
 sg13g2_decap_8 FILLER_41_376 ();
 sg13g2_decap_8 FILLER_41_383 ();
 sg13g2_decap_8 FILLER_41_390 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_fill_1 FILLER_42_65 ();
 sg13g2_fill_2 FILLER_42_104 ();
 sg13g2_fill_2 FILLER_42_134 ();
 sg13g2_fill_1 FILLER_42_136 ();
 sg13g2_decap_4 FILLER_42_181 ();
 sg13g2_fill_1 FILLER_42_185 ();
 sg13g2_fill_2 FILLER_42_233 ();
 sg13g2_fill_1 FILLER_42_238 ();
 sg13g2_fill_2 FILLER_42_266 ();
 sg13g2_fill_1 FILLER_42_268 ();
 sg13g2_fill_1 FILLER_42_274 ();
 sg13g2_fill_1 FILLER_42_280 ();
 sg13g2_fill_2 FILLER_42_333 ();
 sg13g2_fill_2 FILLER_42_354 ();
 sg13g2_decap_8 FILLER_42_384 ();
 sg13g2_decap_8 FILLER_42_391 ();
 sg13g2_decap_8 FILLER_42_398 ();
 sg13g2_decap_4 FILLER_42_405 ();
 sg13g2_fill_2 FILLER_43_91 ();
 sg13g2_fill_1 FILLER_43_108 ();
 sg13g2_fill_1 FILLER_43_114 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_fill_2 FILLER_43_133 ();
 sg13g2_fill_1 FILLER_43_135 ();
 sg13g2_fill_1 FILLER_43_141 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_fill_2 FILLER_43_161 ();
 sg13g2_fill_1 FILLER_43_163 ();
 sg13g2_decap_4 FILLER_43_172 ();
 sg13g2_decap_4 FILLER_43_229 ();
 sg13g2_fill_2 FILLER_43_256 ();
 sg13g2_fill_2 FILLER_43_277 ();
 sg13g2_fill_1 FILLER_43_279 ();
 sg13g2_fill_2 FILLER_43_286 ();
 sg13g2_fill_1 FILLER_43_288 ();
 sg13g2_decap_8 FILLER_43_304 ();
 sg13g2_fill_2 FILLER_43_311 ();
 sg13g2_decap_8 FILLER_43_323 ();
 sg13g2_fill_2 FILLER_43_330 ();
 sg13g2_fill_1 FILLER_43_332 ();
 sg13g2_fill_2 FILLER_43_348 ();
 sg13g2_fill_1 FILLER_43_350 ();
 sg13g2_fill_2 FILLER_43_356 ();
 sg13g2_fill_1 FILLER_43_358 ();
 sg13g2_decap_8 FILLER_43_388 ();
 sg13g2_decap_8 FILLER_43_395 ();
 sg13g2_decap_8 FILLER_43_402 ();
 sg13g2_fill_2 FILLER_44_107 ();
 sg13g2_fill_1 FILLER_44_109 ();
 sg13g2_decap_8 FILLER_44_132 ();
 sg13g2_fill_1 FILLER_44_139 ();
 sg13g2_fill_2 FILLER_44_200 ();
 sg13g2_fill_1 FILLER_44_212 ();
 sg13g2_decap_8 FILLER_44_221 ();
 sg13g2_decap_8 FILLER_44_228 ();
 sg13g2_decap_8 FILLER_44_235 ();
 sg13g2_decap_8 FILLER_44_264 ();
 sg13g2_decap_4 FILLER_44_284 ();
 sg13g2_fill_2 FILLER_44_293 ();
 sg13g2_decap_8 FILLER_44_305 ();
 sg13g2_decap_8 FILLER_44_312 ();
 sg13g2_decap_8 FILLER_44_319 ();
 sg13g2_decap_4 FILLER_44_326 ();
 sg13g2_decap_8 FILLER_44_336 ();
 sg13g2_fill_2 FILLER_44_343 ();
 sg13g2_fill_2 FILLER_44_349 ();
 sg13g2_fill_1 FILLER_44_359 ();
 sg13g2_fill_2 FILLER_44_365 ();
 sg13g2_fill_1 FILLER_44_372 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_fill_2 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_fill_1 FILLER_45_4 ();
 sg13g2_fill_2 FILLER_45_9 ();
 sg13g2_fill_2 FILLER_45_41 ();
 sg13g2_fill_2 FILLER_45_75 ();
 sg13g2_fill_2 FILLER_45_99 ();
 sg13g2_fill_1 FILLER_45_101 ();
 sg13g2_fill_2 FILLER_45_133 ();
 sg13g2_fill_2 FILLER_45_158 ();
 sg13g2_fill_1 FILLER_45_160 ();
 sg13g2_decap_8 FILLER_45_179 ();
 sg13g2_fill_1 FILLER_45_186 ();
 sg13g2_decap_8 FILLER_45_192 ();
 sg13g2_decap_4 FILLER_45_199 ();
 sg13g2_decap_4 FILLER_45_215 ();
 sg13g2_fill_2 FILLER_45_219 ();
 sg13g2_decap_8 FILLER_45_232 ();
 sg13g2_decap_4 FILLER_45_239 ();
 sg13g2_decap_8 FILLER_45_251 ();
 sg13g2_fill_2 FILLER_45_258 ();
 sg13g2_fill_2 FILLER_45_282 ();
 sg13g2_fill_1 FILLER_45_284 ();
 sg13g2_fill_1 FILLER_45_293 ();
 sg13g2_fill_2 FILLER_45_302 ();
 sg13g2_fill_1 FILLER_45_304 ();
 sg13g2_fill_1 FILLER_45_316 ();
 sg13g2_decap_4 FILLER_45_331 ();
 sg13g2_fill_1 FILLER_45_335 ();
 sg13g2_decap_8 FILLER_45_356 ();
 sg13g2_decap_8 FILLER_45_363 ();
 sg13g2_fill_2 FILLER_45_370 ();
 sg13g2_fill_1 FILLER_45_372 ();
 sg13g2_decap_8 FILLER_45_387 ();
 sg13g2_decap_8 FILLER_45_394 ();
 sg13g2_decap_8 FILLER_45_401 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_16 ();
 sg13g2_fill_1 FILLER_46_22 ();
 sg13g2_fill_2 FILLER_46_96 ();
 sg13g2_fill_1 FILLER_46_98 ();
 sg13g2_fill_1 FILLER_46_143 ();
 sg13g2_fill_2 FILLER_46_157 ();
 sg13g2_fill_1 FILLER_46_159 ();
 sg13g2_decap_8 FILLER_46_164 ();
 sg13g2_decap_4 FILLER_46_171 ();
 sg13g2_fill_1 FILLER_46_189 ();
 sg13g2_decap_4 FILLER_46_194 ();
 sg13g2_fill_2 FILLER_46_198 ();
 sg13g2_fill_2 FILLER_46_243 ();
 sg13g2_fill_1 FILLER_46_245 ();
 sg13g2_fill_2 FILLER_46_251 ();
 sg13g2_fill_1 FILLER_46_253 ();
 sg13g2_fill_1 FILLER_46_292 ();
 sg13g2_fill_2 FILLER_46_326 ();
 sg13g2_fill_1 FILLER_46_328 ();
 sg13g2_fill_1 FILLER_46_335 ();
 sg13g2_decap_4 FILLER_46_342 ();
 sg13g2_fill_1 FILLER_46_346 ();
 sg13g2_decap_8 FILLER_46_352 ();
 sg13g2_fill_2 FILLER_46_359 ();
 sg13g2_fill_1 FILLER_46_370 ();
 sg13g2_decap_8 FILLER_46_389 ();
 sg13g2_decap_8 FILLER_46_396 ();
 sg13g2_decap_4 FILLER_46_403 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_36 ();
 sg13g2_fill_2 FILLER_47_103 ();
 sg13g2_fill_1 FILLER_47_105 ();
 sg13g2_fill_1 FILLER_47_111 ();
 sg13g2_fill_2 FILLER_47_142 ();
 sg13g2_decap_8 FILLER_47_149 ();
 sg13g2_fill_2 FILLER_47_156 ();
 sg13g2_decap_4 FILLER_47_162 ();
 sg13g2_fill_1 FILLER_47_166 ();
 sg13g2_fill_2 FILLER_47_191 ();
 sg13g2_decap_4 FILLER_47_204 ();
 sg13g2_decap_4 FILLER_47_214 ();
 sg13g2_fill_1 FILLER_47_222 ();
 sg13g2_fill_2 FILLER_47_231 ();
 sg13g2_fill_1 FILLER_47_233 ();
 sg13g2_fill_1 FILLER_47_239 ();
 sg13g2_decap_4 FILLER_47_255 ();
 sg13g2_fill_1 FILLER_47_264 ();
 sg13g2_fill_1 FILLER_47_272 ();
 sg13g2_fill_2 FILLER_47_358 ();
 sg13g2_decap_8 FILLER_47_391 ();
 sg13g2_decap_8 FILLER_47_398 ();
 sg13g2_decap_4 FILLER_47_405 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_46 ();
 sg13g2_fill_1 FILLER_48_70 ();
 sg13g2_fill_2 FILLER_48_98 ();
 sg13g2_fill_1 FILLER_48_100 ();
 sg13g2_fill_1 FILLER_48_111 ();
 sg13g2_decap_8 FILLER_48_145 ();
 sg13g2_fill_2 FILLER_48_152 ();
 sg13g2_fill_2 FILLER_48_159 ();
 sg13g2_decap_8 FILLER_48_211 ();
 sg13g2_fill_2 FILLER_48_218 ();
 sg13g2_fill_2 FILLER_48_226 ();
 sg13g2_fill_1 FILLER_48_266 ();
 sg13g2_fill_1 FILLER_48_285 ();
 sg13g2_decap_4 FILLER_48_305 ();
 sg13g2_fill_2 FILLER_48_324 ();
 sg13g2_fill_1 FILLER_48_326 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_fill_2 FILLER_48_406 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_32 ();
 sg13g2_fill_1 FILLER_49_40 ();
 sg13g2_fill_1 FILLER_49_71 ();
 sg13g2_fill_2 FILLER_49_113 ();
 sg13g2_fill_2 FILLER_49_124 ();
 sg13g2_fill_2 FILLER_49_197 ();
 sg13g2_fill_1 FILLER_49_232 ();
 sg13g2_decap_4 FILLER_49_261 ();
 sg13g2_fill_2 FILLER_49_265 ();
 sg13g2_fill_2 FILLER_49_272 ();
 sg13g2_decap_8 FILLER_49_279 ();
 sg13g2_decap_4 FILLER_49_286 ();
 sg13g2_fill_2 FILLER_49_290 ();
 sg13g2_fill_2 FILLER_49_300 ();
 sg13g2_decap_4 FILLER_49_307 ();
 sg13g2_fill_1 FILLER_49_316 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_fill_1 FILLER_49_336 ();
 sg13g2_fill_2 FILLER_49_361 ();
 sg13g2_decap_8 FILLER_49_376 ();
 sg13g2_decap_8 FILLER_49_383 ();
 sg13g2_decap_8 FILLER_49_390 ();
 sg13g2_decap_8 FILLER_49_397 ();
 sg13g2_decap_4 FILLER_49_404 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_fill_2 FILLER_50_66 ();
 sg13g2_fill_1 FILLER_50_103 ();
 sg13g2_fill_2 FILLER_50_130 ();
 sg13g2_fill_1 FILLER_50_132 ();
 sg13g2_fill_2 FILLER_50_188 ();
 sg13g2_decap_8 FILLER_50_223 ();
 sg13g2_fill_2 FILLER_50_230 ();
 sg13g2_fill_2 FILLER_50_244 ();
 sg13g2_decap_4 FILLER_50_251 ();
 sg13g2_fill_2 FILLER_50_255 ();
 sg13g2_decap_8 FILLER_50_262 ();
 sg13g2_decap_8 FILLER_50_278 ();
 sg13g2_decap_8 FILLER_50_285 ();
 sg13g2_fill_1 FILLER_50_305 ();
 sg13g2_fill_2 FILLER_50_317 ();
 sg13g2_decap_8 FILLER_50_323 ();
 sg13g2_decap_8 FILLER_50_330 ();
 sg13g2_decap_4 FILLER_50_337 ();
 sg13g2_decap_8 FILLER_50_349 ();
 sg13g2_fill_2 FILLER_50_356 ();
 sg13g2_fill_1 FILLER_50_358 ();
 sg13g2_decap_8 FILLER_50_388 ();
 sg13g2_decap_8 FILLER_50_395 ();
 sg13g2_decap_8 FILLER_50_402 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_69 ();
 sg13g2_fill_2 FILLER_51_82 ();
 sg13g2_fill_2 FILLER_51_122 ();
 sg13g2_fill_1 FILLER_51_130 ();
 sg13g2_fill_2 FILLER_51_147 ();
 sg13g2_fill_1 FILLER_51_149 ();
 sg13g2_fill_2 FILLER_51_163 ();
 sg13g2_decap_8 FILLER_51_177 ();
 sg13g2_decap_8 FILLER_51_184 ();
 sg13g2_fill_2 FILLER_51_191 ();
 sg13g2_fill_1 FILLER_51_193 ();
 sg13g2_decap_8 FILLER_51_215 ();
 sg13g2_decap_8 FILLER_51_222 ();
 sg13g2_decap_4 FILLER_51_229 ();
 sg13g2_fill_1 FILLER_51_233 ();
 sg13g2_fill_2 FILLER_51_238 ();
 sg13g2_fill_1 FILLER_51_240 ();
 sg13g2_decap_8 FILLER_51_249 ();
 sg13g2_fill_2 FILLER_51_256 ();
 sg13g2_fill_1 FILLER_51_258 ();
 sg13g2_fill_2 FILLER_51_265 ();
 sg13g2_fill_1 FILLER_51_267 ();
 sg13g2_fill_1 FILLER_51_277 ();
 sg13g2_fill_1 FILLER_51_283 ();
 sg13g2_decap_4 FILLER_51_289 ();
 sg13g2_decap_4 FILLER_51_308 ();
 sg13g2_fill_2 FILLER_51_338 ();
 sg13g2_fill_1 FILLER_51_340 ();
 sg13g2_fill_2 FILLER_51_364 ();
 sg13g2_fill_1 FILLER_51_366 ();
 sg13g2_fill_2 FILLER_51_371 ();
 sg13g2_decap_8 FILLER_51_390 ();
 sg13g2_decap_8 FILLER_51_397 ();
 sg13g2_decap_4 FILLER_51_404 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_fill_2 FILLER_52_49 ();
 sg13g2_fill_1 FILLER_52_72 ();
 sg13g2_decap_8 FILLER_52_104 ();
 sg13g2_fill_2 FILLER_52_111 ();
 sg13g2_decap_8 FILLER_52_144 ();
 sg13g2_fill_1 FILLER_52_151 ();
 sg13g2_decap_8 FILLER_52_161 ();
 sg13g2_fill_2 FILLER_52_168 ();
 sg13g2_fill_1 FILLER_52_170 ();
 sg13g2_fill_2 FILLER_52_180 ();
 sg13g2_decap_4 FILLER_52_187 ();
 sg13g2_fill_1 FILLER_52_191 ();
 sg13g2_fill_2 FILLER_52_196 ();
 sg13g2_fill_1 FILLER_52_198 ();
 sg13g2_decap_8 FILLER_52_207 ();
 sg13g2_decap_8 FILLER_52_214 ();
 sg13g2_fill_2 FILLER_52_221 ();
 sg13g2_fill_2 FILLER_52_241 ();
 sg13g2_fill_1 FILLER_52_243 ();
 sg13g2_decap_4 FILLER_52_259 ();
 sg13g2_fill_2 FILLER_52_288 ();
 sg13g2_fill_1 FILLER_52_320 ();
 sg13g2_fill_2 FILLER_52_358 ();
 sg13g2_fill_1 FILLER_52_360 ();
 sg13g2_fill_2 FILLER_52_376 ();
 sg13g2_decap_8 FILLER_52_386 ();
 sg13g2_decap_8 FILLER_52_393 ();
 sg13g2_decap_8 FILLER_52_400 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_fill_1 FILLER_53_58 ();
 sg13g2_fill_1 FILLER_53_78 ();
 sg13g2_fill_2 FILLER_53_84 ();
 sg13g2_fill_2 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_145 ();
 sg13g2_decap_8 FILLER_53_152 ();
 sg13g2_fill_2 FILLER_53_159 ();
 sg13g2_fill_1 FILLER_53_161 ();
 sg13g2_fill_2 FILLER_53_167 ();
 sg13g2_fill_1 FILLER_53_169 ();
 sg13g2_fill_2 FILLER_53_200 ();
 sg13g2_decap_4 FILLER_53_207 ();
 sg13g2_fill_2 FILLER_53_211 ();
 sg13g2_fill_2 FILLER_53_244 ();
 sg13g2_fill_1 FILLER_53_246 ();
 sg13g2_fill_1 FILLER_53_260 ();
 sg13g2_fill_2 FILLER_53_277 ();
 sg13g2_fill_1 FILLER_53_279 ();
 sg13g2_fill_1 FILLER_53_308 ();
 sg13g2_fill_2 FILLER_53_319 ();
 sg13g2_decap_4 FILLER_53_330 ();
 sg13g2_fill_1 FILLER_53_356 ();
 sg13g2_decap_8 FILLER_53_382 ();
 sg13g2_decap_8 FILLER_53_389 ();
 sg13g2_decap_8 FILLER_53_396 ();
 sg13g2_decap_4 FILLER_53_403 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_11 ();
 sg13g2_fill_2 FILLER_54_15 ();
 sg13g2_fill_1 FILLER_54_17 ();
 sg13g2_fill_1 FILLER_54_78 ();
 sg13g2_fill_2 FILLER_54_150 ();
 sg13g2_fill_2 FILLER_54_172 ();
 sg13g2_fill_2 FILLER_54_203 ();
 sg13g2_fill_2 FILLER_54_231 ();
 sg13g2_decap_4 FILLER_54_258 ();
 sg13g2_fill_1 FILLER_54_262 ();
 sg13g2_decap_4 FILLER_54_273 ();
 sg13g2_fill_2 FILLER_54_277 ();
 sg13g2_fill_2 FILLER_54_291 ();
 sg13g2_fill_2 FILLER_54_301 ();
 sg13g2_fill_2 FILLER_54_309 ();
 sg13g2_fill_1 FILLER_54_311 ();
 sg13g2_fill_1 FILLER_54_335 ();
 sg13g2_fill_1 FILLER_54_342 ();
 sg13g2_fill_1 FILLER_54_353 ();
 sg13g2_fill_2 FILLER_54_358 ();
 sg13g2_fill_1 FILLER_54_360 ();
 sg13g2_decap_8 FILLER_54_374 ();
 sg13g2_decap_8 FILLER_54_381 ();
 sg13g2_decap_8 FILLER_54_388 ();
 sg13g2_decap_8 FILLER_54_395 ();
 sg13g2_decap_8 FILLER_54_402 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_4 FILLER_55_14 ();
 sg13g2_fill_1 FILLER_55_18 ();
 sg13g2_decap_8 FILLER_55_23 ();
 sg13g2_decap_4 FILLER_55_45 ();
 sg13g2_fill_1 FILLER_55_56 ();
 sg13g2_fill_1 FILLER_55_79 ();
 sg13g2_fill_1 FILLER_55_108 ();
 sg13g2_fill_2 FILLER_55_173 ();
 sg13g2_fill_1 FILLER_55_175 ();
 sg13g2_fill_2 FILLER_55_184 ();
 sg13g2_fill_1 FILLER_55_186 ();
 sg13g2_decap_8 FILLER_55_207 ();
 sg13g2_fill_2 FILLER_55_214 ();
 sg13g2_fill_1 FILLER_55_221 ();
 sg13g2_decap_8 FILLER_55_248 ();
 sg13g2_fill_2 FILLER_55_263 ();
 sg13g2_fill_1 FILLER_55_279 ();
 sg13g2_fill_1 FILLER_55_297 ();
 sg13g2_fill_2 FILLER_55_322 ();
 sg13g2_fill_2 FILLER_55_341 ();
 sg13g2_decap_4 FILLER_55_351 ();
 sg13g2_fill_2 FILLER_55_355 ();
 sg13g2_decap_4 FILLER_55_365 ();
 sg13g2_decap_8 FILLER_55_383 ();
 sg13g2_decap_8 FILLER_55_390 ();
 sg13g2_decap_8 FILLER_55_397 ();
 sg13g2_decap_4 FILLER_55_404 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_2 ();
 sg13g2_fill_1 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_21 ();
 sg13g2_fill_1 FILLER_56_43 ();
 sg13g2_fill_1 FILLER_56_87 ();
 sg13g2_fill_2 FILLER_56_117 ();
 sg13g2_fill_1 FILLER_56_119 ();
 sg13g2_fill_2 FILLER_56_130 ();
 sg13g2_fill_2 FILLER_56_178 ();
 sg13g2_fill_2 FILLER_56_188 ();
 sg13g2_fill_1 FILLER_56_196 ();
 sg13g2_decap_8 FILLER_56_203 ();
 sg13g2_fill_2 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_253 ();
 sg13g2_fill_1 FILLER_56_260 ();
 sg13g2_fill_1 FILLER_56_265 ();
 sg13g2_fill_1 FILLER_56_276 ();
 sg13g2_fill_1 FILLER_56_326 ();
 sg13g2_fill_1 FILLER_56_341 ();
 sg13g2_fill_2 FILLER_56_352 ();
 sg13g2_fill_1 FILLER_56_354 ();
 sg13g2_decap_8 FILLER_56_373 ();
 sg13g2_decap_8 FILLER_56_380 ();
 sg13g2_decap_8 FILLER_56_387 ();
 sg13g2_decap_8 FILLER_56_394 ();
 sg13g2_decap_8 FILLER_56_401 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_fill_2 FILLER_57_31 ();
 sg13g2_fill_1 FILLER_57_68 ();
 sg13g2_fill_2 FILLER_57_84 ();
 sg13g2_decap_4 FILLER_57_167 ();
 sg13g2_fill_2 FILLER_57_171 ();
 sg13g2_decap_8 FILLER_57_178 ();
 sg13g2_decap_4 FILLER_57_185 ();
 sg13g2_fill_1 FILLER_57_189 ();
 sg13g2_decap_4 FILLER_57_211 ();
 sg13g2_fill_2 FILLER_57_235 ();
 sg13g2_fill_1 FILLER_57_237 ();
 sg13g2_decap_4 FILLER_57_266 ();
 sg13g2_fill_2 FILLER_57_276 ();
 sg13g2_fill_1 FILLER_57_278 ();
 sg13g2_fill_1 FILLER_57_283 ();
 sg13g2_decap_8 FILLER_57_306 ();
 sg13g2_fill_1 FILLER_57_313 ();
 sg13g2_decap_8 FILLER_57_319 ();
 sg13g2_fill_2 FILLER_57_326 ();
 sg13g2_fill_1 FILLER_57_328 ();
 sg13g2_fill_2 FILLER_57_344 ();
 sg13g2_decap_4 FILLER_57_357 ();
 sg13g2_decap_8 FILLER_57_390 ();
 sg13g2_decap_8 FILLER_57_397 ();
 sg13g2_decap_4 FILLER_57_404 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_fill_2 FILLER_58_26 ();
 sg13g2_fill_1 FILLER_58_40 ();
 sg13g2_fill_2 FILLER_58_65 ();
 sg13g2_fill_1 FILLER_58_93 ();
 sg13g2_decap_8 FILLER_58_176 ();
 sg13g2_decap_8 FILLER_58_183 ();
 sg13g2_fill_2 FILLER_58_208 ();
 sg13g2_fill_2 FILLER_58_221 ();
 sg13g2_fill_1 FILLER_58_233 ();
 sg13g2_fill_2 FILLER_58_254 ();
 sg13g2_fill_2 FILLER_58_261 ();
 sg13g2_fill_1 FILLER_58_263 ();
 sg13g2_decap_8 FILLER_58_273 ();
 sg13g2_decap_4 FILLER_58_280 ();
 sg13g2_decap_4 FILLER_58_301 ();
 sg13g2_fill_1 FILLER_58_305 ();
 sg13g2_fill_1 FILLER_58_332 ();
 sg13g2_fill_1 FILLER_58_344 ();
 sg13g2_decap_8 FILLER_58_393 ();
 sg13g2_decap_8 FILLER_58_400 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_19 ();
 sg13g2_fill_1 FILLER_59_46 ();
 sg13g2_fill_2 FILLER_59_117 ();
 sg13g2_fill_2 FILLER_59_164 ();
 sg13g2_fill_1 FILLER_59_166 ();
 sg13g2_fill_2 FILLER_59_187 ();
 sg13g2_decap_4 FILLER_59_205 ();
 sg13g2_fill_2 FILLER_59_209 ();
 sg13g2_decap_8 FILLER_59_223 ();
 sg13g2_decap_4 FILLER_59_230 ();
 sg13g2_decap_8 FILLER_59_246 ();
 sg13g2_decap_8 FILLER_59_253 ();
 sg13g2_decap_8 FILLER_59_260 ();
 sg13g2_decap_4 FILLER_59_267 ();
 sg13g2_fill_1 FILLER_59_271 ();
 sg13g2_decap_8 FILLER_59_280 ();
 sg13g2_fill_2 FILLER_59_287 ();
 sg13g2_fill_1 FILLER_59_289 ();
 sg13g2_fill_1 FILLER_59_294 ();
 sg13g2_decap_8 FILLER_59_303 ();
 sg13g2_fill_1 FILLER_59_310 ();
 sg13g2_fill_2 FILLER_59_315 ();
 sg13g2_fill_1 FILLER_59_317 ();
 sg13g2_fill_1 FILLER_59_323 ();
 sg13g2_decap_8 FILLER_59_328 ();
 sg13g2_fill_2 FILLER_59_359 ();
 sg13g2_fill_1 FILLER_59_361 ();
 sg13g2_decap_8 FILLER_59_384 ();
 sg13g2_decap_8 FILLER_59_391 ();
 sg13g2_decap_8 FILLER_59_398 ();
 sg13g2_decap_4 FILLER_59_405 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_36 ();
 sg13g2_fill_1 FILLER_60_76 ();
 sg13g2_fill_2 FILLER_60_86 ();
 sg13g2_fill_2 FILLER_60_101 ();
 sg13g2_fill_1 FILLER_60_108 ();
 sg13g2_fill_2 FILLER_60_161 ();
 sg13g2_fill_2 FILLER_60_177 ();
 sg13g2_fill_1 FILLER_60_179 ();
 sg13g2_fill_2 FILLER_60_195 ();
 sg13g2_decap_4 FILLER_60_219 ();
 sg13g2_fill_1 FILLER_60_223 ();
 sg13g2_fill_1 FILLER_60_233 ();
 sg13g2_decap_8 FILLER_60_242 ();
 sg13g2_fill_2 FILLER_60_249 ();
 sg13g2_fill_1 FILLER_60_251 ();
 sg13g2_fill_1 FILLER_60_269 ();
 sg13g2_fill_2 FILLER_60_289 ();
 sg13g2_fill_2 FILLER_60_296 ();
 sg13g2_fill_1 FILLER_60_298 ();
 sg13g2_fill_2 FILLER_60_335 ();
 sg13g2_fill_1 FILLER_60_337 ();
 sg13g2_fill_1 FILLER_60_368 ();
 sg13g2_decap_8 FILLER_60_374 ();
 sg13g2_decap_8 FILLER_60_381 ();
 sg13g2_decap_8 FILLER_60_388 ();
 sg13g2_decap_8 FILLER_60_395 ();
 sg13g2_decap_8 FILLER_60_402 ();
 sg13g2_fill_2 FILLER_61_92 ();
 sg13g2_fill_2 FILLER_61_139 ();
 sg13g2_fill_1 FILLER_61_156 ();
 sg13g2_fill_2 FILLER_61_183 ();
 sg13g2_fill_1 FILLER_61_185 ();
 sg13g2_fill_2 FILLER_61_197 ();
 sg13g2_fill_1 FILLER_61_199 ();
 sg13g2_fill_2 FILLER_61_209 ();
 sg13g2_fill_2 FILLER_61_279 ();
 sg13g2_fill_1 FILLER_61_281 ();
 sg13g2_fill_1 FILLER_61_363 ();
 sg13g2_decap_8 FILLER_61_378 ();
 sg13g2_decap_8 FILLER_61_385 ();
 sg13g2_decap_8 FILLER_61_392 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_2 FILLER_62_15 ();
 sg13g2_fill_2 FILLER_62_46 ();
 sg13g2_fill_2 FILLER_62_56 ();
 sg13g2_fill_2 FILLER_62_116 ();
 sg13g2_fill_1 FILLER_62_143 ();
 sg13g2_fill_2 FILLER_62_164 ();
 sg13g2_fill_1 FILLER_62_166 ();
 sg13g2_fill_2 FILLER_62_203 ();
 sg13g2_fill_2 FILLER_62_210 ();
 sg13g2_fill_1 FILLER_62_212 ();
 sg13g2_fill_1 FILLER_62_221 ();
 sg13g2_fill_2 FILLER_62_240 ();
 sg13g2_fill_1 FILLER_62_242 ();
 sg13g2_fill_1 FILLER_62_251 ();
 sg13g2_fill_2 FILLER_62_335 ();
 sg13g2_fill_1 FILLER_62_337 ();
 sg13g2_decap_8 FILLER_62_386 ();
 sg13g2_decap_8 FILLER_62_393 ();
 sg13g2_decap_8 FILLER_62_400 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_fill_1 FILLER_63_37 ();
 sg13g2_fill_2 FILLER_63_43 ();
 sg13g2_fill_2 FILLER_63_107 ();
 sg13g2_fill_1 FILLER_63_173 ();
 sg13g2_fill_1 FILLER_63_186 ();
 sg13g2_fill_2 FILLER_63_197 ();
 sg13g2_decap_4 FILLER_63_230 ();
 sg13g2_fill_1 FILLER_63_234 ();
 sg13g2_decap_4 FILLER_63_251 ();
 sg13g2_fill_2 FILLER_63_255 ();
 sg13g2_decap_8 FILLER_63_264 ();
 sg13g2_fill_2 FILLER_63_271 ();
 sg13g2_fill_1 FILLER_63_278 ();
 sg13g2_decap_4 FILLER_63_288 ();
 sg13g2_fill_2 FILLER_63_296 ();
 sg13g2_decap_8 FILLER_63_307 ();
 sg13g2_decap_8 FILLER_63_314 ();
 sg13g2_decap_8 FILLER_63_321 ();
 sg13g2_fill_2 FILLER_63_328 ();
 sg13g2_fill_2 FILLER_63_338 ();
 sg13g2_fill_1 FILLER_63_340 ();
 sg13g2_fill_2 FILLER_63_354 ();
 sg13g2_fill_2 FILLER_63_361 ();
 sg13g2_fill_1 FILLER_63_368 ();
 sg13g2_decap_8 FILLER_63_382 ();
 sg13g2_decap_8 FILLER_63_389 ();
 sg13g2_decap_8 FILLER_63_396 ();
 sg13g2_decap_4 FILLER_63_403 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_60 ();
 sg13g2_fill_2 FILLER_64_89 ();
 sg13g2_fill_1 FILLER_64_117 ();
 sg13g2_fill_2 FILLER_64_132 ();
 sg13g2_fill_1 FILLER_64_142 ();
 sg13g2_fill_1 FILLER_64_163 ();
 sg13g2_decap_4 FILLER_64_175 ();
 sg13g2_fill_2 FILLER_64_191 ();
 sg13g2_fill_2 FILLER_64_197 ();
 sg13g2_fill_1 FILLER_64_203 ();
 sg13g2_fill_2 FILLER_64_213 ();
 sg13g2_decap_8 FILLER_64_224 ();
 sg13g2_fill_2 FILLER_64_231 ();
 sg13g2_decap_8 FILLER_64_247 ();
 sg13g2_decap_8 FILLER_64_254 ();
 sg13g2_decap_4 FILLER_64_270 ();
 sg13g2_fill_2 FILLER_64_274 ();
 sg13g2_fill_2 FILLER_64_281 ();
 sg13g2_fill_1 FILLER_64_283 ();
 sg13g2_decap_8 FILLER_64_288 ();
 sg13g2_decap_8 FILLER_64_295 ();
 sg13g2_decap_8 FILLER_64_302 ();
 sg13g2_fill_1 FILLER_64_314 ();
 sg13g2_fill_2 FILLER_64_324 ();
 sg13g2_decap_8 FILLER_64_331 ();
 sg13g2_fill_1 FILLER_64_338 ();
 sg13g2_decap_8 FILLER_64_362 ();
 sg13g2_decap_8 FILLER_64_369 ();
 sg13g2_decap_8 FILLER_64_376 ();
 sg13g2_decap_8 FILLER_64_383 ();
 sg13g2_decap_8 FILLER_64_390 ();
 sg13g2_decap_8 FILLER_64_397 ();
 sg13g2_decap_4 FILLER_64_404 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_22 ();
 sg13g2_fill_1 FILLER_65_40 ();
 sg13g2_fill_1 FILLER_65_76 ();
 sg13g2_fill_2 FILLER_65_81 ();
 sg13g2_fill_2 FILLER_65_136 ();
 sg13g2_decap_4 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_168 ();
 sg13g2_fill_2 FILLER_65_175 ();
 sg13g2_fill_2 FILLER_65_195 ();
 sg13g2_fill_1 FILLER_65_197 ();
 sg13g2_fill_2 FILLER_65_208 ();
 sg13g2_fill_1 FILLER_65_210 ();
 sg13g2_fill_2 FILLER_65_248 ();
 sg13g2_fill_2 FILLER_65_273 ();
 sg13g2_fill_2 FILLER_65_291 ();
 sg13g2_fill_1 FILLER_65_293 ();
 sg13g2_fill_2 FILLER_65_310 ();
 sg13g2_decap_8 FILLER_65_377 ();
 sg13g2_decap_8 FILLER_65_384 ();
 sg13g2_decap_8 FILLER_65_391 ();
 sg13g2_decap_8 FILLER_65_398 ();
 sg13g2_decap_4 FILLER_65_405 ();
 sg13g2_fill_1 FILLER_66_26 ();
 sg13g2_fill_2 FILLER_66_96 ();
 sg13g2_fill_1 FILLER_66_98 ();
 sg13g2_fill_1 FILLER_66_104 ();
 sg13g2_fill_1 FILLER_66_173 ();
 sg13g2_fill_1 FILLER_66_201 ();
 sg13g2_fill_2 FILLER_66_207 ();
 sg13g2_fill_1 FILLER_66_209 ();
 sg13g2_fill_2 FILLER_66_227 ();
 sg13g2_decap_8 FILLER_66_237 ();
 sg13g2_decap_8 FILLER_66_244 ();
 sg13g2_decap_8 FILLER_66_251 ();
 sg13g2_decap_8 FILLER_66_258 ();
 sg13g2_fill_1 FILLER_66_265 ();
 sg13g2_fill_2 FILLER_66_278 ();
 sg13g2_fill_1 FILLER_66_280 ();
 sg13g2_fill_1 FILLER_66_310 ();
 sg13g2_fill_1 FILLER_66_321 ();
 sg13g2_fill_2 FILLER_66_352 ();
 sg13g2_decap_8 FILLER_66_366 ();
 sg13g2_decap_8 FILLER_66_373 ();
 sg13g2_decap_8 FILLER_66_380 ();
 sg13g2_decap_8 FILLER_66_387 ();
 sg13g2_decap_8 FILLER_66_394 ();
 sg13g2_decap_8 FILLER_66_401 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_2 ();
 sg13g2_fill_1 FILLER_67_12 ();
 sg13g2_fill_2 FILLER_67_47 ();
 sg13g2_fill_1 FILLER_67_100 ();
 sg13g2_fill_2 FILLER_67_152 ();
 sg13g2_fill_1 FILLER_67_162 ();
 sg13g2_fill_1 FILLER_67_207 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_8 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_238 ();
 sg13g2_decap_4 FILLER_67_245 ();
 sg13g2_fill_1 FILLER_67_249 ();
 sg13g2_fill_2 FILLER_67_269 ();
 sg13g2_fill_2 FILLER_67_317 ();
 sg13g2_fill_1 FILLER_67_319 ();
 sg13g2_decap_8 FILLER_67_366 ();
 sg13g2_decap_8 FILLER_67_373 ();
 sg13g2_decap_8 FILLER_67_380 ();
 sg13g2_decap_8 FILLER_67_387 ();
 sg13g2_decap_8 FILLER_67_394 ();
 sg13g2_decap_8 FILLER_67_401 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_4 ();
 sg13g2_fill_2 FILLER_68_19 ();
 sg13g2_fill_2 FILLER_68_52 ();
 sg13g2_fill_2 FILLER_68_79 ();
 sg13g2_fill_1 FILLER_68_81 ();
 sg13g2_fill_2 FILLER_68_108 ();
 sg13g2_fill_1 FILLER_68_202 ();
 sg13g2_fill_2 FILLER_68_211 ();
 sg13g2_fill_1 FILLER_68_213 ();
 sg13g2_fill_1 FILLER_68_221 ();
 sg13g2_fill_2 FILLER_68_261 ();
 sg13g2_fill_2 FILLER_68_274 ();
 sg13g2_decap_8 FILLER_68_324 ();
 sg13g2_decap_4 FILLER_68_341 ();
 sg13g2_decap_4 FILLER_68_351 ();
 sg13g2_decap_8 FILLER_68_373 ();
 sg13g2_decap_8 FILLER_68_380 ();
 sg13g2_decap_8 FILLER_68_387 ();
 sg13g2_decap_8 FILLER_68_394 ();
 sg13g2_decap_8 FILLER_68_401 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_fill_2 FILLER_69_26 ();
 sg13g2_fill_1 FILLER_69_28 ();
 sg13g2_fill_2 FILLER_69_44 ();
 sg13g2_fill_1 FILLER_69_61 ();
 sg13g2_fill_1 FILLER_69_84 ();
 sg13g2_fill_2 FILLER_69_152 ();
 sg13g2_fill_2 FILLER_69_196 ();
 sg13g2_fill_1 FILLER_69_198 ();
 sg13g2_fill_1 FILLER_69_234 ();
 sg13g2_fill_1 FILLER_69_258 ();
 sg13g2_fill_2 FILLER_69_263 ();
 sg13g2_fill_1 FILLER_69_265 ();
 sg13g2_decap_4 FILLER_69_283 ();
 sg13g2_fill_1 FILLER_69_287 ();
 sg13g2_fill_2 FILLER_69_292 ();
 sg13g2_fill_1 FILLER_69_294 ();
 sg13g2_fill_2 FILLER_69_300 ();
 sg13g2_fill_1 FILLER_69_302 ();
 sg13g2_decap_4 FILLER_69_311 ();
 sg13g2_decap_8 FILLER_69_319 ();
 sg13g2_decap_4 FILLER_69_326 ();
 sg13g2_fill_2 FILLER_69_330 ();
 sg13g2_fill_1 FILLER_69_342 ();
 sg13g2_fill_2 FILLER_69_348 ();
 sg13g2_decap_8 FILLER_69_365 ();
 sg13g2_decap_8 FILLER_69_372 ();
 sg13g2_decap_8 FILLER_69_379 ();
 sg13g2_decap_8 FILLER_69_386 ();
 sg13g2_decap_8 FILLER_69_393 ();
 sg13g2_decap_8 FILLER_69_400 ();
 sg13g2_fill_2 FILLER_69_407 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_7 ();
 sg13g2_fill_1 FILLER_70_9 ();
 sg13g2_fill_2 FILLER_70_22 ();
 sg13g2_fill_1 FILLER_70_24 ();
 sg13g2_fill_1 FILLER_70_83 ();
 sg13g2_fill_2 FILLER_70_92 ();
 sg13g2_fill_1 FILLER_70_94 ();
 sg13g2_fill_2 FILLER_70_143 ();
 sg13g2_fill_1 FILLER_70_145 ();
 sg13g2_fill_2 FILLER_70_154 ();
 sg13g2_fill_1 FILLER_70_174 ();
 sg13g2_fill_1 FILLER_70_180 ();
 sg13g2_fill_1 FILLER_70_207 ();
 sg13g2_fill_2 FILLER_70_217 ();
 sg13g2_fill_1 FILLER_70_238 ();
 sg13g2_fill_1 FILLER_70_244 ();
 sg13g2_decap_4 FILLER_70_249 ();
 sg13g2_decap_4 FILLER_70_262 ();
 sg13g2_fill_1 FILLER_70_266 ();
 sg13g2_decap_4 FILLER_70_284 ();
 sg13g2_fill_1 FILLER_70_288 ();
 sg13g2_fill_1 FILLER_70_294 ();
 sg13g2_fill_2 FILLER_70_300 ();
 sg13g2_fill_1 FILLER_70_302 ();
 sg13g2_fill_2 FILLER_70_309 ();
 sg13g2_fill_2 FILLER_70_331 ();
 sg13g2_fill_1 FILLER_70_343 ();
 sg13g2_decap_8 FILLER_70_362 ();
 sg13g2_decap_8 FILLER_70_369 ();
 sg13g2_decap_8 FILLER_70_376 ();
 sg13g2_decap_8 FILLER_70_383 ();
 sg13g2_decap_8 FILLER_70_390 ();
 sg13g2_decap_8 FILLER_70_397 ();
 sg13g2_decap_4 FILLER_70_404 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_27 ();
 sg13g2_fill_1 FILLER_71_36 ();
 sg13g2_fill_2 FILLER_71_70 ();
 sg13g2_fill_1 FILLER_71_80 ();
 sg13g2_fill_1 FILLER_71_120 ();
 sg13g2_fill_1 FILLER_71_130 ();
 sg13g2_fill_1 FILLER_71_188 ();
 sg13g2_fill_1 FILLER_71_228 ();
 sg13g2_decap_8 FILLER_71_260 ();
 sg13g2_fill_2 FILLER_71_267 ();
 sg13g2_decap_4 FILLER_71_274 ();
 sg13g2_fill_2 FILLER_71_344 ();
 sg13g2_fill_1 FILLER_71_346 ();
 sg13g2_decap_8 FILLER_71_359 ();
 sg13g2_decap_8 FILLER_71_366 ();
 sg13g2_decap_8 FILLER_71_373 ();
 sg13g2_decap_8 FILLER_71_380 ();
 sg13g2_decap_8 FILLER_71_387 ();
 sg13g2_decap_8 FILLER_71_394 ();
 sg13g2_decap_8 FILLER_71_401 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_14 ();
 sg13g2_fill_1 FILLER_72_16 ();
 sg13g2_fill_1 FILLER_72_66 ();
 sg13g2_fill_2 FILLER_72_109 ();
 sg13g2_fill_2 FILLER_72_189 ();
 sg13g2_fill_1 FILLER_72_191 ();
 sg13g2_fill_2 FILLER_72_196 ();
 sg13g2_fill_1 FILLER_72_198 ();
 sg13g2_fill_2 FILLER_72_243 ();
 sg13g2_fill_1 FILLER_72_245 ();
 sg13g2_fill_1 FILLER_72_280 ();
 sg13g2_fill_1 FILLER_72_293 ();
 sg13g2_fill_1 FILLER_72_336 ();
 sg13g2_decap_8 FILLER_72_353 ();
 sg13g2_decap_8 FILLER_72_360 ();
 sg13g2_decap_8 FILLER_72_367 ();
 sg13g2_decap_8 FILLER_72_374 ();
 sg13g2_decap_8 FILLER_72_381 ();
 sg13g2_decap_8 FILLER_72_388 ();
 sg13g2_decap_8 FILLER_72_395 ();
 sg13g2_decap_8 FILLER_72_402 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_fill_2 FILLER_73_21 ();
 sg13g2_fill_2 FILLER_73_134 ();
 sg13g2_fill_2 FILLER_73_158 ();
 sg13g2_fill_1 FILLER_73_160 ();
 sg13g2_fill_2 FILLER_73_166 ();
 sg13g2_fill_2 FILLER_73_176 ();
 sg13g2_decap_8 FILLER_73_194 ();
 sg13g2_decap_8 FILLER_73_201 ();
 sg13g2_fill_2 FILLER_73_208 ();
 sg13g2_decap_8 FILLER_73_213 ();
 sg13g2_fill_2 FILLER_73_220 ();
 sg13g2_fill_1 FILLER_73_222 ();
 sg13g2_fill_1 FILLER_73_238 ();
 sg13g2_decap_8 FILLER_73_294 ();
 sg13g2_fill_2 FILLER_73_301 ();
 sg13g2_fill_2 FILLER_73_310 ();
 sg13g2_fill_1 FILLER_73_312 ();
 sg13g2_fill_1 FILLER_73_327 ();
 sg13g2_decap_8 FILLER_73_341 ();
 sg13g2_decap_8 FILLER_73_348 ();
 sg13g2_decap_8 FILLER_73_355 ();
 sg13g2_decap_8 FILLER_73_362 ();
 sg13g2_decap_8 FILLER_73_369 ();
 sg13g2_decap_8 FILLER_73_376 ();
 sg13g2_decap_8 FILLER_73_383 ();
 sg13g2_decap_8 FILLER_73_390 ();
 sg13g2_decap_8 FILLER_73_397 ();
 sg13g2_decap_4 FILLER_73_404 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_4 FILLER_74_14 ();
 sg13g2_fill_1 FILLER_74_18 ();
 sg13g2_fill_2 FILLER_74_38 ();
 sg13g2_fill_2 FILLER_74_45 ();
 sg13g2_fill_1 FILLER_74_56 ();
 sg13g2_fill_1 FILLER_74_77 ();
 sg13g2_fill_2 FILLER_74_88 ();
 sg13g2_fill_1 FILLER_74_142 ();
 sg13g2_fill_1 FILLER_74_209 ();
 sg13g2_fill_1 FILLER_74_225 ();
 sg13g2_fill_2 FILLER_74_266 ();
 sg13g2_decap_8 FILLER_74_300 ();
 sg13g2_decap_8 FILLER_74_307 ();
 sg13g2_decap_8 FILLER_74_314 ();
 sg13g2_decap_8 FILLER_74_321 ();
 sg13g2_fill_1 FILLER_74_328 ();
 sg13g2_decap_8 FILLER_74_333 ();
 sg13g2_decap_8 FILLER_74_340 ();
 sg13g2_decap_8 FILLER_74_347 ();
 sg13g2_decap_8 FILLER_74_354 ();
 sg13g2_decap_8 FILLER_74_361 ();
 sg13g2_decap_8 FILLER_74_368 ();
 sg13g2_decap_8 FILLER_74_375 ();
 sg13g2_decap_8 FILLER_74_382 ();
 sg13g2_decap_8 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_74_396 ();
 sg13g2_decap_4 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_fill_1 FILLER_75_28 ();
 sg13g2_fill_1 FILLER_75_39 ();
 sg13g2_fill_1 FILLER_75_53 ();
 sg13g2_fill_2 FILLER_75_98 ();
 sg13g2_fill_1 FILLER_75_173 ();
 sg13g2_decap_8 FILLER_75_221 ();
 sg13g2_fill_2 FILLER_75_228 ();
 sg13g2_fill_2 FILLER_75_240 ();
 sg13g2_fill_2 FILLER_75_247 ();
 sg13g2_fill_2 FILLER_75_254 ();
 sg13g2_fill_1 FILLER_75_256 ();
 sg13g2_decap_8 FILLER_75_317 ();
 sg13g2_decap_8 FILLER_75_324 ();
 sg13g2_decap_8 FILLER_75_331 ();
 sg13g2_decap_8 FILLER_75_338 ();
 sg13g2_decap_8 FILLER_75_345 ();
 sg13g2_decap_8 FILLER_75_352 ();
 sg13g2_decap_8 FILLER_75_359 ();
 sg13g2_decap_8 FILLER_75_366 ();
 sg13g2_decap_8 FILLER_75_373 ();
 sg13g2_decap_8 FILLER_75_380 ();
 sg13g2_decap_8 FILLER_75_387 ();
 sg13g2_decap_8 FILLER_75_394 ();
 sg13g2_decap_8 FILLER_75_401 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_fill_2 FILLER_76_21 ();
 sg13g2_fill_1 FILLER_76_23 ();
 sg13g2_fill_2 FILLER_76_63 ();
 sg13g2_fill_1 FILLER_76_92 ();
 sg13g2_fill_1 FILLER_76_171 ();
 sg13g2_fill_1 FILLER_76_209 ();
 sg13g2_fill_2 FILLER_76_220 ();
 sg13g2_fill_2 FILLER_76_250 ();
 sg13g2_fill_1 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_392 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_fill_2 FILLER_76_406 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_fill_2 FILLER_77_128 ();
 sg13g2_fill_1 FILLER_77_130 ();
 sg13g2_fill_2 FILLER_77_140 ();
 sg13g2_fill_2 FILLER_77_151 ();
 sg13g2_fill_2 FILLER_77_231 ();
 sg13g2_fill_2 FILLER_77_245 ();
 sg13g2_decap_8 FILLER_77_287 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_decap_8 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_364 ();
 sg13g2_decap_8 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_fill_2 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_fill_2 FILLER_78_35 ();
 sg13g2_fill_1 FILLER_78_72 ();
 sg13g2_fill_2 FILLER_78_125 ();
 sg13g2_fill_2 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_279 ();
 sg13g2_decap_8 FILLER_78_286 ();
 sg13g2_decap_8 FILLER_78_293 ();
 sg13g2_decap_8 FILLER_78_300 ();
 sg13g2_decap_8 FILLER_78_307 ();
 sg13g2_decap_8 FILLER_78_314 ();
 sg13g2_decap_8 FILLER_78_321 ();
 sg13g2_decap_8 FILLER_78_328 ();
 sg13g2_decap_8 FILLER_78_335 ();
 sg13g2_decap_8 FILLER_78_342 ();
 sg13g2_decap_8 FILLER_78_349 ();
 sg13g2_decap_8 FILLER_78_356 ();
 sg13g2_decap_8 FILLER_78_363 ();
 sg13g2_decap_8 FILLER_78_370 ();
 sg13g2_decap_8 FILLER_78_377 ();
 sg13g2_decap_8 FILLER_78_384 ();
 sg13g2_decap_8 FILLER_78_391 ();
 sg13g2_decap_8 FILLER_78_398 ();
 sg13g2_decap_4 FILLER_78_405 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_fill_2 FILLER_79_28 ();
 sg13g2_fill_1 FILLER_79_30 ();
 sg13g2_fill_1 FILLER_79_105 ();
 sg13g2_fill_2 FILLER_79_111 ();
 sg13g2_fill_2 FILLER_79_122 ();
 sg13g2_fill_1 FILLER_79_124 ();
 sg13g2_fill_1 FILLER_79_156 ();
 sg13g2_fill_1 FILLER_79_183 ();
 sg13g2_fill_1 FILLER_79_241 ();
 sg13g2_decap_8 FILLER_79_268 ();
 sg13g2_decap_8 FILLER_79_275 ();
 sg13g2_decap_8 FILLER_79_282 ();
 sg13g2_decap_8 FILLER_79_289 ();
 sg13g2_decap_8 FILLER_79_296 ();
 sg13g2_decap_8 FILLER_79_303 ();
 sg13g2_decap_8 FILLER_79_310 ();
 sg13g2_decap_8 FILLER_79_317 ();
 sg13g2_decap_8 FILLER_79_324 ();
 sg13g2_decap_8 FILLER_79_331 ();
 sg13g2_decap_8 FILLER_79_338 ();
 sg13g2_decap_8 FILLER_79_345 ();
 sg13g2_decap_8 FILLER_79_352 ();
 sg13g2_decap_8 FILLER_79_359 ();
 sg13g2_decap_8 FILLER_79_366 ();
 sg13g2_decap_8 FILLER_79_373 ();
 sg13g2_decap_8 FILLER_79_380 ();
 sg13g2_decap_8 FILLER_79_387 ();
 sg13g2_decap_8 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_401 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_fill_2 FILLER_80_21 ();
 sg13g2_fill_1 FILLER_80_23 ();
 sg13g2_fill_2 FILLER_80_85 ();
 sg13g2_fill_1 FILLER_80_87 ();
 sg13g2_fill_2 FILLER_80_96 ();
 sg13g2_fill_1 FILLER_80_126 ();
 sg13g2_fill_1 FILLER_80_175 ();
 sg13g2_fill_1 FILLER_80_189 ();
 sg13g2_fill_2 FILLER_80_202 ();
 sg13g2_fill_1 FILLER_80_204 ();
 sg13g2_fill_1 FILLER_80_209 ();
 sg13g2_decap_8 FILLER_80_218 ();
 sg13g2_decap_8 FILLER_80_225 ();
 sg13g2_decap_8 FILLER_80_232 ();
 sg13g2_fill_1 FILLER_80_239 ();
 sg13g2_decap_4 FILLER_80_245 ();
 sg13g2_fill_1 FILLER_80_249 ();
 sg13g2_fill_2 FILLER_80_255 ();
 sg13g2_decap_8 FILLER_80_261 ();
 sg13g2_decap_8 FILLER_80_268 ();
 sg13g2_decap_8 FILLER_80_275 ();
 sg13g2_decap_8 FILLER_80_282 ();
 sg13g2_decap_8 FILLER_80_289 ();
 sg13g2_decap_8 FILLER_80_296 ();
 sg13g2_decap_8 FILLER_80_303 ();
 sg13g2_decap_8 FILLER_80_310 ();
 sg13g2_decap_8 FILLER_80_317 ();
 sg13g2_decap_8 FILLER_80_324 ();
 sg13g2_decap_8 FILLER_80_331 ();
 sg13g2_decap_8 FILLER_80_338 ();
 sg13g2_decap_8 FILLER_80_345 ();
 sg13g2_decap_8 FILLER_80_352 ();
 sg13g2_decap_8 FILLER_80_359 ();
 sg13g2_decap_8 FILLER_80_366 ();
 sg13g2_decap_8 FILLER_80_373 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net65;
 assign uio_out[0] = net8;
 assign uio_out[1] = net9;
 assign uio_out[2] = net10;
 assign uio_out[3] = net11;
 assign uio_out[4] = net12;
 assign uio_out[5] = net13;
 assign uio_out[6] = net14;
endmodule

module tt_um_systolicLif (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire net26;
 wire net27;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire \first.enable_Reg ;
 wire \first.out_data[3] ;
 wire \first.out_data[4] ;
 wire \first.out_data[5] ;
 wire \first.out_data[6] ;
 wire \four.spike ;
 wire \four.state[2] ;
 wire \four.state[3] ;
 wire \four.state[4] ;
 wire \four.state[5] ;
 wire \four.state[6] ;
 wire \four.state[7] ;
 wire \fourth.accumulate[1] ;
 wire \fourth.accumulate[2] ;
 wire \fourth.accumulate[3] ;
 wire \fourth.accumulate[4] ;
 wire \fourth.accumulate[5] ;
 wire \fourth.accumulate[6] ;
 wire \fourth.enable_Reg ;
 wire \fourth.out_data[0] ;
 wire \fourth.out_data[1] ;
 wire \fourth.out_data[2] ;
 wire \fourth.out_data[3] ;
 wire \fourth.out_data[4] ;
 wire \fourth.out_data[5] ;
 wire \fourth.out_data[6] ;
 wire \mac_Out_two[2] ;
 wire \mac_Out_two[3] ;
 wire \mac_Out_two[4] ;
 wire \mac_Out_two[5] ;
 wire \mac_Out_two[6] ;
 wire \one.spike ;
 wire \one.state[3] ;
 wire \one.state[4] ;
 wire \one.state[5] ;
 wire \one.state[6] ;
 wire \one.state[7] ;
 wire \second.enable_Reg ;
 wire \third.enable_Reg ;
 wire \three.spike ;
 wire \three.state[3] ;
 wire \three.state[4] ;
 wire \three.state[5] ;
 wire \three.state[6] ;
 wire \three.state[7] ;
 wire \two.spike ;
 wire \two.state[3] ;
 wire \two.state[4] ;
 wire \two.state[5] ;
 wire \two.state[6] ;
 wire \two.state[7] ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_0_clk;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;

 sg13g2_inv_2 _336_ (.Y(_047_),
    .A(net33));
 sg13g2_inv_2 _337_ (.Y(_048_),
    .A(net4));
 sg13g2_inv_2 _338_ (.Y(_049_),
    .A(net5));
 sg13g2_inv_1 _339_ (.Y(_050_),
    .A(\mac_Out_two[3] ));
 sg13g2_inv_1 _340_ (.Y(_051_),
    .A(net85));
 sg13g2_inv_1 _341_ (.Y(_052_),
    .A(\fourth.out_data[1] ));
 sg13g2_inv_1 _342_ (.Y(_053_),
    .A(\fourth.out_data[0] ));
 sg13g2_inv_1 _343_ (.Y(_054_),
    .A(\fourth.out_data[2] ));
 sg13g2_nand2_2 _344_ (.Y(_055_),
    .A(\three.state[7] ),
    .B(\three.state[6] ));
 sg13g2_nor3_1 _345_ (.A(\three.state[3] ),
    .B(\three.state[4] ),
    .C(\three.state[5] ),
    .Y(_056_));
 sg13g2_or2_1 _346_ (.X(_057_),
    .B(_056_),
    .A(_055_));
 sg13g2_inv_1 _347_ (.Y(\three.spike ),
    .A(_057_));
 sg13g2_nand2_1 _348_ (.Y(_058_),
    .A(\four.state[7] ),
    .B(\four.state[6] ));
 sg13g2_nor3_1 _349_ (.A(\four.state[3] ),
    .B(\four.state[4] ),
    .C(\four.state[5] ),
    .Y(_059_));
 sg13g2_or2_1 _350_ (.X(_060_),
    .B(_059_),
    .A(_058_));
 sg13g2_inv_1 _351_ (.Y(\four.spike ),
    .A(net30));
 sg13g2_or3_1 _352_ (.A(\one.state[3] ),
    .B(\one.state[4] ),
    .C(\one.state[5] ),
    .X(_061_));
 sg13g2_nand3_1 _353_ (.B(\one.state[6] ),
    .C(_061_),
    .A(net134),
    .Y(_062_));
 sg13g2_inv_1 _354_ (.Y(\one.spike ),
    .A(_062_));
 sg13g2_or3_1 _355_ (.A(\two.state[3] ),
    .B(\two.state[4] ),
    .C(\two.state[5] ),
    .X(_063_));
 sg13g2_nand3_1 _356_ (.B(\two.state[6] ),
    .C(_063_),
    .A(\two.state[7] ),
    .Y(_064_));
 sg13g2_inv_1 _357_ (.Y(\two.spike ),
    .A(_064_));
 sg13g2_nor2_1 _358_ (.A(net32),
    .B(\one.spike ),
    .Y(_065_));
 sg13g2_and2_1 _359_ (.A(net82),
    .B(_065_),
    .X(_000_));
 sg13g2_nand2_1 _360_ (.Y(_066_),
    .A(net3),
    .B(\mac_Out_two[6] ));
 sg13g2_and2_1 _361_ (.A(net2),
    .B(\mac_Out_two[5] ),
    .X(_067_));
 sg13g2_and2_1 _362_ (.A(net1),
    .B(net86),
    .X(_068_));
 sg13g2_xor2_1 _363_ (.B(net114),
    .A(net2),
    .X(_069_));
 sg13g2_a21oi_1 _364_ (.A1(_068_),
    .A2(_069_),
    .Y(_070_),
    .B1(_067_));
 sg13g2_xnor2_1 _365_ (.Y(_071_),
    .A(net3),
    .B(net116));
 sg13g2_o21ai_1 _366_ (.B1(_066_),
    .Y(_072_),
    .A1(_070_),
    .A2(_071_));
 sg13g2_nand2_1 _367_ (.Y(_073_),
    .A(net4),
    .B(_072_));
 sg13g2_xnor2_1 _368_ (.Y(_074_),
    .A(_048_),
    .B(_072_));
 sg13g2_xor2_1 _369_ (.B(_071_),
    .A(_070_),
    .X(_075_));
 sg13g2_xnor2_1 _370_ (.Y(_076_),
    .A(_068_),
    .B(_069_));
 sg13g2_xnor2_1 _371_ (.Y(_077_),
    .A(net1),
    .B(net86));
 sg13g2_nand2_1 _372_ (.Y(_078_),
    .A(net129),
    .B(net85));
 sg13g2_nand3_1 _373_ (.B(_077_),
    .C(_078_),
    .A(_076_),
    .Y(_079_));
 sg13g2_nand3_1 _374_ (.B(_075_),
    .C(_079_),
    .A(_074_),
    .Y(_080_));
 sg13g2_xnor2_1 _375_ (.Y(_081_),
    .A(_049_),
    .B(_073_));
 sg13g2_nand2_1 _376_ (.Y(_082_),
    .A(_080_),
    .B(_081_));
 sg13g2_and4_1 _377_ (.A(net128),
    .B(\fourth.accumulate[1] ),
    .C(_055_),
    .D(net29),
    .X(_083_));
 sg13g2_nand4_1 _378_ (.B(net91),
    .C(_055_),
    .A(net103),
    .Y(_084_),
    .D(net29));
 sg13g2_nand2_1 _379_ (.Y(_085_),
    .A(\three.state[4] ),
    .B(_055_));
 sg13g2_inv_1 _380_ (.Y(_086_),
    .A(_085_));
 sg13g2_and3_1 _381_ (.X(_087_),
    .A(net87),
    .B(net29),
    .C(_086_));
 sg13g2_a21o_1 _382_ (.A2(net29),
    .A1(net87),
    .B1(_086_),
    .X(_088_));
 sg13g2_nand2b_1 _383_ (.Y(_089_),
    .B(_088_),
    .A_N(_087_));
 sg13g2_o21ai_1 _384_ (.B1(net33),
    .Y(_090_),
    .A1(_084_),
    .A2(_089_));
 sg13g2_a21oi_1 _385_ (.A1(net104),
    .A2(_089_),
    .Y(_001_),
    .B1(_090_));
 sg13g2_and2_1 _386_ (.A(\three.state[5] ),
    .B(_055_),
    .X(_091_));
 sg13g2_nand3_1 _387_ (.B(net29),
    .C(_091_),
    .A(net89),
    .Y(_092_));
 sg13g2_a21o_1 _388_ (.A2(net29),
    .A1(net89),
    .B1(_091_),
    .X(_093_));
 sg13g2_nand2_1 _389_ (.Y(_094_),
    .A(_092_),
    .B(_093_));
 sg13g2_a21oi_1 _390_ (.A1(_083_),
    .A2(_088_),
    .Y(_095_),
    .B1(_087_));
 sg13g2_o21ai_1 _391_ (.B1(net33),
    .Y(_096_),
    .A1(_094_),
    .A2(_095_));
 sg13g2_a21oi_1 _392_ (.A1(_094_),
    .A2(_095_),
    .Y(_002_),
    .B1(_096_));
 sg13g2_o21ai_1 _393_ (.B1(_092_),
    .Y(_097_),
    .A1(_094_),
    .A2(_095_));
 sg13g2_nand2_1 _394_ (.Y(_098_),
    .A(\fourth.accumulate[4] ),
    .B(_082_));
 sg13g2_nand2_1 _395_ (.Y(_099_),
    .A(net132),
    .B(_057_));
 sg13g2_nor2_1 _396_ (.A(_098_),
    .B(_099_),
    .Y(_100_));
 sg13g2_xor2_1 _397_ (.B(_099_),
    .A(_098_),
    .X(_101_));
 sg13g2_o21ai_1 _398_ (.B1(net33),
    .Y(_102_),
    .A1(_097_),
    .A2(_101_));
 sg13g2_a21oi_1 _399_ (.A1(_097_),
    .A2(_101_),
    .Y(_003_),
    .B1(_102_));
 sg13g2_a21oi_1 _400_ (.A1(_097_),
    .A2(_101_),
    .Y(_103_),
    .B1(net133));
 sg13g2_and2_1 _401_ (.A(\fourth.accumulate[5] ),
    .B(net29),
    .X(_104_));
 sg13g2_nand3_1 _402_ (.B(_057_),
    .C(_104_),
    .A(net123),
    .Y(_105_));
 sg13g2_a21o_1 _403_ (.A2(_057_),
    .A1(net123),
    .B1(_104_),
    .X(_106_));
 sg13g2_nand2_1 _404_ (.Y(_107_),
    .A(_105_),
    .B(_106_));
 sg13g2_o21ai_1 _405_ (.B1(net33),
    .Y(_108_),
    .A1(_103_),
    .A2(_107_));
 sg13g2_a21oi_1 _406_ (.A1(_103_),
    .A2(_107_),
    .Y(_004_),
    .B1(_108_));
 sg13g2_and2_1 _407_ (.A(net112),
    .B(net29),
    .X(_109_));
 sg13g2_o21ai_1 _408_ (.B1(_105_),
    .Y(_110_),
    .A1(_103_),
    .A2(_107_));
 sg13g2_o21ai_1 _409_ (.B1(net33),
    .Y(_111_),
    .A1(_109_),
    .A2(_110_));
 sg13g2_a21oi_1 _410_ (.A1(_109_),
    .A2(_110_),
    .Y(_005_),
    .B1(_111_));
 sg13g2_and2_1 _411_ (.A(net3),
    .B(\fourth.accumulate[6] ),
    .X(_112_));
 sg13g2_nand2_1 _412_ (.Y(_113_),
    .A(net2),
    .B(\fourth.accumulate[5] ));
 sg13g2_nand2_1 _413_ (.Y(_114_),
    .A(net1),
    .B(net110));
 sg13g2_xnor2_1 _414_ (.Y(_115_),
    .A(net2),
    .B(\fourth.accumulate[5] ));
 sg13g2_o21ai_1 _415_ (.B1(_113_),
    .Y(_116_),
    .A1(_114_),
    .A2(_115_));
 sg13g2_xor2_1 _416_ (.B(\fourth.accumulate[6] ),
    .A(net3),
    .X(_117_));
 sg13g2_a21oi_2 _417_ (.B1(net113),
    .Y(_118_),
    .A2(_117_),
    .A1(_116_));
 sg13g2_nor3_1 _418_ (.A(_048_),
    .B(_049_),
    .C(_118_),
    .Y(_119_));
 sg13g2_nand3b_1 _419_ (.B(net5),
    .C(net4),
    .Y(_120_),
    .A_N(_118_));
 sg13g2_xnor2_1 _420_ (.Y(_121_),
    .A(_116_),
    .B(_117_));
 sg13g2_xnor2_1 _421_ (.Y(_122_),
    .A(_114_),
    .B(_115_));
 sg13g2_o21ai_1 _422_ (.B1(\fourth.accumulate[3] ),
    .Y(_123_),
    .A1(\fourth.accumulate[2] ),
    .A2(\fourth.accumulate[1] ));
 sg13g2_xnor2_1 _423_ (.Y(_124_),
    .A(net1),
    .B(net110));
 sg13g2_and2_1 _424_ (.A(_123_),
    .B(_124_),
    .X(_125_));
 sg13g2_a221oi_1 _425_ (.B2(_125_),
    .C1(_121_),
    .B1(_122_),
    .A1(_048_),
    .Y(_126_),
    .A2(_118_));
 sg13g2_o21ai_1 _426_ (.B1(_049_),
    .Y(_127_),
    .A1(_048_),
    .A2(_118_));
 sg13g2_nor2_1 _427_ (.A(_126_),
    .B(_127_),
    .Y(_128_));
 sg13g2_xnor2_1 _428_ (.Y(_129_),
    .A(_048_),
    .B(_118_));
 sg13g2_nor2_1 _429_ (.A(_119_),
    .B(_128_),
    .Y(_130_));
 sg13g2_o21ai_1 _430_ (.B1(_120_),
    .Y(_131_),
    .A1(_126_),
    .A2(_127_));
 sg13g2_nand2_1 _431_ (.Y(_132_),
    .A(\four.state[2] ),
    .B(net30));
 sg13g2_nor3_1 _432_ (.A(_053_),
    .B(_131_),
    .C(_132_),
    .Y(_133_));
 sg13g2_nand4_1 _433_ (.B(\fourth.out_data[0] ),
    .C(net30),
    .A(net97),
    .Y(_134_),
    .D(net28));
 sg13g2_nand2_1 _434_ (.Y(_135_),
    .A(\four.state[3] ),
    .B(_058_));
 sg13g2_nor3_1 _435_ (.A(_052_),
    .B(_131_),
    .C(_135_),
    .Y(_136_));
 sg13g2_o21ai_1 _436_ (.B1(_135_),
    .Y(_137_),
    .A1(_052_),
    .A2(_131_));
 sg13g2_nand2b_1 _437_ (.Y(_138_),
    .B(_137_),
    .A_N(_136_));
 sg13g2_o21ai_1 _438_ (.B1(net35),
    .Y(_139_),
    .A1(net98),
    .A2(_138_));
 sg13g2_a21oi_1 _439_ (.A1(net98),
    .A2(_138_),
    .Y(_006_),
    .B1(_139_));
 sg13g2_nor2_1 _440_ (.A(_054_),
    .B(_131_),
    .Y(_140_));
 sg13g2_nand2_1 _441_ (.Y(_141_),
    .A(net136),
    .B(_058_));
 sg13g2_nand3_1 _442_ (.B(net30),
    .C(_140_),
    .A(net126),
    .Y(_142_));
 sg13g2_xor2_1 _443_ (.B(_141_),
    .A(_140_),
    .X(_143_));
 sg13g2_a21oi_1 _444_ (.A1(_133_),
    .A2(_137_),
    .Y(_144_),
    .B1(_136_));
 sg13g2_and2_1 _445_ (.A(_143_),
    .B(_144_),
    .X(_145_));
 sg13g2_nor2_1 _446_ (.A(_143_),
    .B(_144_),
    .Y(_146_));
 sg13g2_nor3_1 _447_ (.A(_047_),
    .B(_145_),
    .C(_146_),
    .Y(_007_));
 sg13g2_o21ai_1 _448_ (.B1(_142_),
    .Y(_147_),
    .A1(_143_),
    .A2(_144_));
 sg13g2_and4_1 _449_ (.A(\four.state[5] ),
    .B(\fourth.out_data[3] ),
    .C(net30),
    .D(net28),
    .X(_148_));
 sg13g2_nand4_1 _450_ (.B(\fourth.out_data[3] ),
    .C(net30),
    .A(\four.state[5] ),
    .Y(_149_),
    .D(net28));
 sg13g2_a22oi_1 _451_ (.Y(_150_),
    .B1(net28),
    .B2(\fourth.out_data[3] ),
    .A2(net30),
    .A1(\four.state[5] ));
 sg13g2_nor2_1 _452_ (.A(_148_),
    .B(_150_),
    .Y(_151_));
 sg13g2_o21ai_1 _453_ (.B1(net35),
    .Y(_152_),
    .A1(_147_),
    .A2(_151_));
 sg13g2_a21oi_1 _454_ (.A1(_147_),
    .A2(_151_),
    .Y(_008_),
    .B1(_152_));
 sg13g2_a21oi_1 _455_ (.A1(_142_),
    .A2(_149_),
    .Y(_153_),
    .B1(_150_));
 sg13g2_a21oi_1 _456_ (.A1(_146_),
    .A2(_151_),
    .Y(_154_),
    .B1(_153_));
 sg13g2_and4_1 _457_ (.A(\four.state[6] ),
    .B(\fourth.out_data[4] ),
    .C(_060_),
    .D(_130_),
    .X(_155_));
 sg13g2_a22oi_1 _458_ (.Y(_156_),
    .B1(net28),
    .B2(net119),
    .A2(_060_),
    .A1(\four.state[6] ));
 sg13g2_or2_1 _459_ (.X(_157_),
    .B(net120),
    .A(_155_));
 sg13g2_or2_1 _460_ (.X(_158_),
    .B(_157_),
    .A(_154_));
 sg13g2_nand2_1 _461_ (.Y(_159_),
    .A(net34),
    .B(_158_));
 sg13g2_a21oi_1 _462_ (.A1(_154_),
    .A2(_157_),
    .Y(_009_),
    .B1(_159_));
 sg13g2_nand2b_1 _463_ (.Y(_160_),
    .B(_158_),
    .A_N(_155_));
 sg13g2_a22oi_1 _464_ (.Y(_161_),
    .B1(net28),
    .B2(net130),
    .A2(_060_),
    .A1(\four.state[7] ));
 sg13g2_and4_1 _465_ (.A(\four.state[7] ),
    .B(\fourth.out_data[5] ),
    .C(net30),
    .D(net28),
    .X(_162_));
 sg13g2_nor2_1 _466_ (.A(net131),
    .B(_162_),
    .Y(_163_));
 sg13g2_inv_1 _467_ (.Y(_164_),
    .A(_163_));
 sg13g2_o21ai_1 _468_ (.B1(net34),
    .Y(_165_),
    .A1(_160_),
    .A2(_163_));
 sg13g2_a21oi_1 _469_ (.A1(_160_),
    .A2(_163_),
    .Y(_010_),
    .B1(_165_));
 sg13g2_and2_1 _470_ (.A(net107),
    .B(net28),
    .X(_166_));
 sg13g2_nor2_1 _471_ (.A(_155_),
    .B(_162_),
    .Y(_167_));
 sg13g2_or2_1 _472_ (.X(_168_),
    .B(_167_),
    .A(_161_));
 sg13g2_o21ai_1 _473_ (.B1(_168_),
    .Y(_169_),
    .A1(_158_),
    .A2(_164_));
 sg13g2_o21ai_1 _474_ (.B1(net34),
    .Y(_170_),
    .A1(_166_),
    .A2(_169_));
 sg13g2_a21oi_1 _475_ (.A1(_166_),
    .A2(_169_),
    .Y(_011_),
    .B1(_170_));
 sg13g2_nor2_1 _476_ (.A(_047_),
    .B(net81),
    .Y(_171_));
 sg13g2_and2_1 _477_ (.A(net1),
    .B(_171_),
    .X(_012_));
 sg13g2_and2_1 _478_ (.A(net2),
    .B(_171_),
    .X(_013_));
 sg13g2_and2_1 _479_ (.A(net3),
    .B(_171_),
    .X(_014_));
 sg13g2_nor3_1 _480_ (.A(net32),
    .B(_048_),
    .C(net81),
    .Y(_015_));
 sg13g2_or2_1 _481_ (.X(_172_),
    .B(net2),
    .A(net1));
 sg13g2_nand3_1 _482_ (.B(net4),
    .C(_172_),
    .A(net3),
    .Y(_173_));
 sg13g2_nand2_2 _483_ (.Y(_174_),
    .A(_049_),
    .B(_173_));
 sg13g2_a22oi_1 _484_ (.Y(_175_),
    .B1(_174_),
    .B2(net93),
    .A2(net135),
    .A1(net95));
 sg13g2_nand4_1 _485_ (.B(net93),
    .C(_062_),
    .A(net95),
    .Y(_176_),
    .D(_174_));
 sg13g2_nand2_1 _486_ (.Y(_177_),
    .A(net34),
    .B(_176_));
 sg13g2_nor2_1 _487_ (.A(_175_),
    .B(_177_),
    .Y(_016_));
 sg13g2_nand2_1 _488_ (.Y(_178_),
    .A(net101),
    .B(_174_));
 sg13g2_nand2_1 _489_ (.Y(_179_),
    .A(net105),
    .B(_062_));
 sg13g2_xnor2_1 _490_ (.Y(_180_),
    .A(_178_),
    .B(_179_));
 sg13g2_or2_1 _491_ (.X(_181_),
    .B(_180_),
    .A(_176_));
 sg13g2_nand2_1 _492_ (.Y(_182_),
    .A(net34),
    .B(_181_));
 sg13g2_a21oi_1 _493_ (.A1(_176_),
    .A2(_180_),
    .Y(_017_),
    .B1(_182_));
 sg13g2_nand2_1 _494_ (.Y(_183_),
    .A(\first.out_data[5] ),
    .B(_174_));
 sg13g2_nand2_1 _495_ (.Y(_184_),
    .A(net125),
    .B(_062_));
 sg13g2_or2_1 _496_ (.X(_185_),
    .B(_184_),
    .A(_183_));
 sg13g2_xor2_1 _497_ (.B(_184_),
    .A(_183_),
    .X(_186_));
 sg13g2_o21ai_1 _498_ (.B1(_181_),
    .Y(_187_),
    .A1(_178_),
    .A2(_179_));
 sg13g2_nand2_1 _499_ (.Y(_188_),
    .A(_186_),
    .B(_187_));
 sg13g2_o21ai_1 _500_ (.B1(net35),
    .Y(_189_),
    .A1(_186_),
    .A2(_187_));
 sg13g2_nor2b_1 _501_ (.A(_189_),
    .B_N(_188_),
    .Y(_018_));
 sg13g2_nand2_1 _502_ (.Y(_190_),
    .A(net106),
    .B(_174_));
 sg13g2_a21oi_1 _503_ (.A1(_185_),
    .A2(_188_),
    .Y(_191_),
    .B1(_190_));
 sg13g2_nand3_1 _504_ (.B(_188_),
    .C(_190_),
    .A(_185_),
    .Y(_192_));
 sg13g2_nand2_1 _505_ (.Y(_193_),
    .A(net35),
    .B(_192_));
 sg13g2_nor2_1 _506_ (.A(_191_),
    .B(_193_),
    .Y(_019_));
 sg13g2_a21oi_1 _507_ (.A1(_049_),
    .A2(_173_),
    .Y(_020_),
    .B1(net32));
 sg13g2_and2_1 _508_ (.A(net3),
    .B(\first.out_data[6] ),
    .X(_194_));
 sg13g2_nand2_1 _509_ (.Y(_195_),
    .A(net2),
    .B(\first.out_data[5] ));
 sg13g2_nand2_1 _510_ (.Y(_196_),
    .A(net1),
    .B(net101));
 sg13g2_xnor2_1 _511_ (.Y(_197_),
    .A(net2),
    .B(\first.out_data[5] ));
 sg13g2_o21ai_1 _512_ (.B1(_195_),
    .Y(_198_),
    .A1(_196_),
    .A2(_197_));
 sg13g2_xor2_1 _513_ (.B(net106),
    .A(net3),
    .X(_199_));
 sg13g2_a21o_1 _514_ (.A2(_199_),
    .A1(_198_),
    .B1(_194_),
    .X(_200_));
 sg13g2_xnor2_1 _515_ (.Y(_201_),
    .A(_048_),
    .B(_200_));
 sg13g2_xnor2_1 _516_ (.Y(_202_),
    .A(net1),
    .B(net101));
 sg13g2_xnor2_1 _517_ (.Y(_203_),
    .A(_196_),
    .B(_197_));
 sg13g2_xnor2_1 _518_ (.Y(_204_),
    .A(_198_),
    .B(_199_));
 sg13g2_a21oi_1 _519_ (.A1(_202_),
    .A2(_203_),
    .Y(_205_),
    .B1(_204_));
 sg13g2_and2_1 _520_ (.A(_201_),
    .B(_205_),
    .X(_206_));
 sg13g2_nand3_1 _521_ (.B(net5),
    .C(_200_),
    .A(net4),
    .Y(_207_));
 sg13g2_a21o_1 _522_ (.A2(_200_),
    .A1(net4),
    .B1(net5),
    .X(_208_));
 sg13g2_a22oi_1 _523_ (.Y(_209_),
    .B1(_207_),
    .B2(_208_),
    .A2(_205_),
    .A1(_201_));
 sg13g2_a21o_1 _524_ (.A2(_208_),
    .A1(_207_),
    .B1(_206_),
    .X(_210_));
 sg13g2_nor2_1 _525_ (.A(net32),
    .B(_209_),
    .Y(_021_));
 sg13g2_a21oi_1 _526_ (.A1(_080_),
    .A2(_081_),
    .Y(_022_),
    .B1(net31));
 sg13g2_nand2_1 _527_ (.Y(_211_),
    .A(net100),
    .B(_064_));
 sg13g2_a22oi_1 _528_ (.Y(_212_),
    .B1(_210_),
    .B2(net85),
    .A2(_064_),
    .A1(net100));
 sg13g2_nor3_1 _529_ (.A(_051_),
    .B(_209_),
    .C(_211_),
    .Y(_213_));
 sg13g2_nor3_1 _530_ (.A(net31),
    .B(_212_),
    .C(_213_),
    .Y(_023_));
 sg13g2_nand2_1 _531_ (.Y(_214_),
    .A(net117),
    .B(_064_));
 sg13g2_or3_1 _532_ (.A(_050_),
    .B(_209_),
    .C(_214_),
    .X(_215_));
 sg13g2_o21ai_1 _533_ (.B1(_214_),
    .Y(_216_),
    .A1(_050_),
    .A2(_209_));
 sg13g2_a21oi_1 _534_ (.A1(_215_),
    .A2(net118),
    .Y(_217_),
    .B1(_213_));
 sg13g2_nand3_1 _535_ (.B(_215_),
    .C(_216_),
    .A(_213_),
    .Y(_218_));
 sg13g2_nand2_1 _536_ (.Y(_219_),
    .A(net33),
    .B(_218_));
 sg13g2_nor2_1 _537_ (.A(_217_),
    .B(_219_),
    .Y(_024_));
 sg13g2_nand2_1 _538_ (.Y(_220_),
    .A(net86),
    .B(_210_));
 sg13g2_nand2_1 _539_ (.Y(_221_),
    .A(net124),
    .B(_064_));
 sg13g2_nor2_1 _540_ (.A(_220_),
    .B(_221_),
    .Y(_222_));
 sg13g2_xor2_1 _541_ (.B(_221_),
    .A(_220_),
    .X(_223_));
 sg13g2_and2_1 _542_ (.A(_215_),
    .B(_218_),
    .X(_224_));
 sg13g2_nor2b_1 _543_ (.A(_223_),
    .B_N(_224_),
    .Y(_225_));
 sg13g2_nor2b_1 _544_ (.A(_224_),
    .B_N(_223_),
    .Y(_226_));
 sg13g2_nor3_1 _545_ (.A(net31),
    .B(_225_),
    .C(_226_),
    .Y(_025_));
 sg13g2_nor2_1 _546_ (.A(_222_),
    .B(_226_),
    .Y(_227_));
 sg13g2_nand2_1 _547_ (.Y(_228_),
    .A(net114),
    .B(_210_));
 sg13g2_nand2_1 _548_ (.Y(_229_),
    .A(net122),
    .B(_064_));
 sg13g2_or2_1 _549_ (.X(_230_),
    .B(_229_),
    .A(_228_));
 sg13g2_xnor2_1 _550_ (.Y(_231_),
    .A(_228_),
    .B(_229_));
 sg13g2_or2_1 _551_ (.X(_232_),
    .B(_231_),
    .A(_227_));
 sg13g2_nand2_1 _552_ (.Y(_233_),
    .A(net34),
    .B(_232_));
 sg13g2_a21oi_1 _553_ (.A1(_227_),
    .A2(_231_),
    .Y(_026_),
    .B1(_233_));
 sg13g2_nand2_1 _554_ (.Y(_234_),
    .A(net115),
    .B(_210_));
 sg13g2_a21oi_1 _555_ (.A1(_230_),
    .A2(_232_),
    .Y(_235_),
    .B1(_234_));
 sg13g2_and3_1 _556_ (.X(_236_),
    .A(_230_),
    .B(_232_),
    .C(_234_));
 sg13g2_nor3_1 _557_ (.A(net31),
    .B(_235_),
    .C(_236_),
    .Y(_027_));
 sg13g2_nor2_1 _558_ (.A(net32),
    .B(_131_),
    .Y(_028_));
 sg13g2_nor2_1 _559_ (.A(net32),
    .B(\fourth.enable_Reg ),
    .Y(_237_));
 sg13g2_nand2b_1 _560_ (.Y(_238_),
    .B(net34),
    .A_N(net108));
 sg13g2_and2_1 _561_ (.A(net91),
    .B(_237_),
    .X(_029_));
 sg13g2_and2_1 _562_ (.A(net87),
    .B(_237_),
    .X(_030_));
 sg13g2_and2_1 _563_ (.A(net89),
    .B(_237_),
    .X(_031_));
 sg13g2_nor2_1 _564_ (.A(_124_),
    .B(_238_),
    .Y(_032_));
 sg13g2_nor2_1 _565_ (.A(net111),
    .B(_238_),
    .Y(_033_));
 sg13g2_nor2_1 _566_ (.A(_121_),
    .B(_238_),
    .Y(_034_));
 sg13g2_nor2_1 _567_ (.A(_129_),
    .B(_238_),
    .Y(_035_));
 sg13g2_nor2_1 _568_ (.A(net31),
    .B(net83),
    .Y(_239_));
 sg13g2_nor3_1 _569_ (.A(net31),
    .B(_051_),
    .C(net83),
    .Y(_036_));
 sg13g2_nor3_1 _570_ (.A(net31),
    .B(_050_),
    .C(net83),
    .Y(_037_));
 sg13g2_nor3_1 _571_ (.A(net31),
    .B(net83),
    .C(_077_),
    .Y(_038_));
 sg13g2_nor2b_1 _572_ (.A(_076_),
    .B_N(_239_),
    .Y(_039_));
 sg13g2_and2_1 _573_ (.A(_075_),
    .B(_239_),
    .X(_040_));
 sg13g2_and2_1 _574_ (.A(_074_),
    .B(_239_),
    .X(_041_));
 sg13g2_nor2_1 _575_ (.A(net32),
    .B(net96),
    .Y(_240_));
 sg13g2_nand2b_1 _576_ (.Y(_241_),
    .B(net33),
    .A_N(net96));
 sg13g2_and2_1 _577_ (.A(net93),
    .B(_240_),
    .X(_042_));
 sg13g2_nor2_1 _578_ (.A(_202_),
    .B(_241_),
    .Y(_043_));
 sg13g2_nor2_1 _579_ (.A(net102),
    .B(_241_),
    .Y(_044_));
 sg13g2_nor2_1 _580_ (.A(_204_),
    .B(_241_),
    .Y(_045_));
 sg13g2_and2_1 _581_ (.A(_201_),
    .B(_240_),
    .X(_046_));
 sg13g2_dfrbp_1 _582_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net73),
    .D(_000_),
    .Q_N(_288_),
    .Q(\one.state[3] ));
 sg13g2_dfrbp_1 _583_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net72),
    .D(_001_),
    .Q_N(_287_),
    .Q(\three.state[3] ));
 sg13g2_dfrbp_1 _584_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net71),
    .D(_002_),
    .Q_N(_286_),
    .Q(\three.state[4] ));
 sg13g2_dfrbp_1 _585_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net70),
    .D(_003_),
    .Q_N(_285_),
    .Q(\three.state[5] ));
 sg13g2_dfrbp_1 _586_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net69),
    .D(_004_),
    .Q_N(_284_),
    .Q(\three.state[6] ));
 sg13g2_dfrbp_1 _587_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net68),
    .D(_005_),
    .Q_N(_283_),
    .Q(\three.state[7] ));
 sg13g2_dfrbp_1 _588_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net67),
    .D(net99),
    .Q_N(_282_),
    .Q(\four.state[2] ));
 sg13g2_dfrbp_1 _589_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net66),
    .D(_007_),
    .Q_N(_281_),
    .Q(\four.state[3] ));
 sg13g2_dfrbp_1 _590_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net65),
    .D(net127),
    .Q_N(_280_),
    .Q(\four.state[4] ));
 sg13g2_dfrbp_1 _591_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net64),
    .D(net121),
    .Q_N(_279_),
    .Q(\four.state[5] ));
 sg13g2_dfrbp_1 _592_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net63),
    .D(_010_),
    .Q_N(_278_),
    .Q(\four.state[6] ));
 sg13g2_dfrbp_1 _593_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net62),
    .D(_011_),
    .Q_N(_277_),
    .Q(\four.state[7] ));
 sg13g2_dfrbp_1 _594_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net61),
    .D(_012_),
    .Q_N(_276_),
    .Q(\first.out_data[3] ));
 sg13g2_dfrbp_1 _595_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net60),
    .D(_013_),
    .Q_N(_275_),
    .Q(\first.out_data[4] ));
 sg13g2_dfrbp_1 _596_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net59),
    .D(_014_),
    .Q_N(_274_),
    .Q(\first.out_data[5] ));
 sg13g2_dfrbp_1 _597_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net58),
    .D(_015_),
    .Q_N(_273_),
    .Q(\first.out_data[6] ));
 sg13g2_dfrbp_1 _598_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net57),
    .D(_016_),
    .Q_N(_272_),
    .Q(\one.state[4] ));
 sg13g2_dfrbp_1 _599_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net56),
    .D(_017_),
    .Q_N(_271_),
    .Q(\one.state[5] ));
 sg13g2_dfrbp_1 _600_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net55),
    .D(_018_),
    .Q_N(_270_),
    .Q(\one.state[6] ));
 sg13g2_dfrbp_1 _601_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net54),
    .D(_019_),
    .Q_N(_269_),
    .Q(\one.state[7] ));
 sg13g2_dfrbp_1 _602_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net53),
    .D(_020_),
    .Q_N(_268_),
    .Q(\first.enable_Reg ));
 sg13g2_dfrbp_1 _603_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net52),
    .D(_021_),
    .Q_N(_267_),
    .Q(\second.enable_Reg ));
 sg13g2_dfrbp_1 _604_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net51),
    .D(_022_),
    .Q_N(_266_),
    .Q(\third.enable_Reg ));
 sg13g2_dfrbp_1 _605_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net50),
    .D(_023_),
    .Q_N(_265_),
    .Q(\two.state[3] ));
 sg13g2_dfrbp_1 _606_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net49),
    .D(_024_),
    .Q_N(_264_),
    .Q(\two.state[4] ));
 sg13g2_dfrbp_1 _607_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net48),
    .D(_025_),
    .Q_N(_263_),
    .Q(\two.state[5] ));
 sg13g2_dfrbp_1 _608_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net47),
    .D(_026_),
    .Q_N(_262_),
    .Q(\two.state[6] ));
 sg13g2_dfrbp_1 _609_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net46),
    .D(_027_),
    .Q_N(_261_),
    .Q(\two.state[7] ));
 sg13g2_dfrbp_1 _610_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net45),
    .D(_028_),
    .Q_N(_260_),
    .Q(\fourth.enable_Reg ));
 sg13g2_dfrbp_1 _611_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net44),
    .D(net92),
    .Q_N(_259_),
    .Q(\fourth.out_data[0] ));
 sg13g2_dfrbp_1 _612_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net43),
    .D(net88),
    .Q_N(_258_),
    .Q(\fourth.out_data[1] ));
 sg13g2_dfrbp_1 _613_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net42),
    .D(net90),
    .Q_N(_257_),
    .Q(\fourth.out_data[2] ));
 sg13g2_dfrbp_1 _614_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net41),
    .D(_032_),
    .Q_N(_256_),
    .Q(\fourth.out_data[3] ));
 sg13g2_dfrbp_1 _615_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net40),
    .D(_033_),
    .Q_N(_255_),
    .Q(\fourth.out_data[4] ));
 sg13g2_dfrbp_1 _616_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net39),
    .D(net109),
    .Q_N(_254_),
    .Q(\fourth.out_data[5] ));
 sg13g2_dfrbp_1 _617_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net38),
    .D(_035_),
    .Q_N(_253_),
    .Q(\fourth.out_data[6] ));
 sg13g2_dfrbp_1 _618_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net37),
    .D(_036_),
    .Q_N(_252_),
    .Q(\fourth.accumulate[1] ));
 sg13g2_dfrbp_1 _619_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net36),
    .D(net84),
    .Q_N(_251_),
    .Q(\fourth.accumulate[2] ));
 sg13g2_dfrbp_1 _620_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net27),
    .D(_038_),
    .Q_N(_250_),
    .Q(\fourth.accumulate[3] ));
 sg13g2_dfrbp_1 _621_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net26),
    .D(_039_),
    .Q_N(_249_),
    .Q(\fourth.accumulate[4] ));
 sg13g2_dfrbp_1 _622_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net25),
    .D(_040_),
    .Q_N(_248_),
    .Q(\fourth.accumulate[5] ));
 sg13g2_dfrbp_1 _623_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net79),
    .D(_041_),
    .Q_N(_247_),
    .Q(\fourth.accumulate[6] ));
 sg13g2_dfrbp_1 _624_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net78),
    .D(net94),
    .Q_N(_246_),
    .Q(\mac_Out_two[2] ));
 sg13g2_dfrbp_1 _625_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net77),
    .D(_043_),
    .Q_N(_245_),
    .Q(\mac_Out_two[3] ));
 sg13g2_dfrbp_1 _626_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net76),
    .D(_044_),
    .Q_N(_244_),
    .Q(\mac_Out_two[4] ));
 sg13g2_dfrbp_1 _627_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net75),
    .D(_045_),
    .Q_N(_243_),
    .Q(\mac_Out_two[5] ));
 sg13g2_dfrbp_1 _628_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net74),
    .D(_046_),
    .Q_N(_242_),
    .Q(\mac_Out_two[6] ));
 sg13g2_tiehi _621__26 (.L_HI(net26));
 sg13g2_tiehi _620__27 (.L_HI(net27));
 sg13g2_tiehi _619__28 (.L_HI(net36));
 sg13g2_tiehi _618__29 (.L_HI(net37));
 sg13g2_tiehi _617__30 (.L_HI(net38));
 sg13g2_tiehi _616__31 (.L_HI(net39));
 sg13g2_tiehi _615__32 (.L_HI(net40));
 sg13g2_tiehi _614__33 (.L_HI(net41));
 sg13g2_tiehi _613__34 (.L_HI(net42));
 sg13g2_tiehi _612__35 (.L_HI(net43));
 sg13g2_tiehi _611__36 (.L_HI(net44));
 sg13g2_tiehi _610__37 (.L_HI(net45));
 sg13g2_tiehi _609__38 (.L_HI(net46));
 sg13g2_tiehi _608__39 (.L_HI(net47));
 sg13g2_tiehi _607__40 (.L_HI(net48));
 sg13g2_tiehi _606__41 (.L_HI(net49));
 sg13g2_tiehi _605__42 (.L_HI(net50));
 sg13g2_tiehi _604__43 (.L_HI(net51));
 sg13g2_tiehi _603__44 (.L_HI(net52));
 sg13g2_tiehi _602__45 (.L_HI(net53));
 sg13g2_tiehi _601__46 (.L_HI(net54));
 sg13g2_tiehi _600__47 (.L_HI(net55));
 sg13g2_tiehi _599__48 (.L_HI(net56));
 sg13g2_tiehi _598__49 (.L_HI(net57));
 sg13g2_tiehi _597__50 (.L_HI(net58));
 sg13g2_tiehi _596__51 (.L_HI(net59));
 sg13g2_tiehi _595__52 (.L_HI(net60));
 sg13g2_tiehi _594__53 (.L_HI(net61));
 sg13g2_tiehi _593__54 (.L_HI(net62));
 sg13g2_tiehi _592__55 (.L_HI(net63));
 sg13g2_tiehi _591__56 (.L_HI(net64));
 sg13g2_tiehi _590__57 (.L_HI(net65));
 sg13g2_tiehi _589__58 (.L_HI(net66));
 sg13g2_tiehi _588__59 (.L_HI(net67));
 sg13g2_tiehi _587__60 (.L_HI(net68));
 sg13g2_tiehi _586__61 (.L_HI(net69));
 sg13g2_tiehi _585__62 (.L_HI(net70));
 sg13g2_tiehi _584__63 (.L_HI(net71));
 sg13g2_tiehi _583__64 (.L_HI(net72));
 sg13g2_tiehi _582__65 (.L_HI(net73));
 sg13g2_tiehi _628__66 (.L_HI(net74));
 sg13g2_tiehi _627__67 (.L_HI(net75));
 sg13g2_tiehi _626__68 (.L_HI(net76));
 sg13g2_tiehi _625__69 (.L_HI(net77));
 sg13g2_tiehi _624__70 (.L_HI(net78));
 sg13g2_tiehi _623__71 (.L_HI(net79));
 sg13g2_tiehi tt_um_systolicLif_72 (.L_HI(net80));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_systolicLif_7 (.L_LO(net7));
 sg13g2_tielo tt_um_systolicLif_8 (.L_LO(net8));
 sg13g2_tielo tt_um_systolicLif_9 (.L_LO(net9));
 sg13g2_tielo tt_um_systolicLif_10 (.L_LO(net10));
 sg13g2_tielo tt_um_systolicLif_11 (.L_LO(net11));
 sg13g2_tielo tt_um_systolicLif_12 (.L_LO(net12));
 sg13g2_tielo tt_um_systolicLif_13 (.L_LO(net13));
 sg13g2_tielo tt_um_systolicLif_14 (.L_LO(net14));
 sg13g2_tielo tt_um_systolicLif_15 (.L_LO(net15));
 sg13g2_tielo tt_um_systolicLif_16 (.L_LO(net16));
 sg13g2_tielo tt_um_systolicLif_17 (.L_LO(net17));
 sg13g2_tielo tt_um_systolicLif_18 (.L_LO(net18));
 sg13g2_tielo tt_um_systolicLif_19 (.L_LO(net19));
 sg13g2_tielo tt_um_systolicLif_20 (.L_LO(net20));
 sg13g2_tielo tt_um_systolicLif_21 (.L_LO(net21));
 sg13g2_tielo tt_um_systolicLif_22 (.L_LO(net22));
 sg13g2_tielo tt_um_systolicLif_23 (.L_LO(net23));
 sg13g2_tielo tt_um_systolicLif_24 (.L_LO(net24));
 sg13g2_tiehi _622__25 (.L_HI(net25));
 sg13g2_buf_2 _696_ (.A(\four.spike ),
    .X(uo_out[4]));
 sg13g2_buf_2 _697_ (.A(\three.spike ),
    .X(uo_out[5]));
 sg13g2_buf_1 _698_ (.A(\two.spike ),
    .X(uo_out[6]));
 sg13g2_buf_1 _699_ (.A(\one.spike ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout28 (.A(_130_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_082_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_060_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(net32),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_047_),
    .X(net32));
 sg13g2_buf_4 fanout33 (.X(net33),
    .A(net34));
 sg13g2_buf_4 fanout34 (.X(net34),
    .A(rst_n));
 sg13g2_buf_2 fanout35 (.A(rst_n),
    .X(net35));
 sg13g2_buf_4 input1 (.X(net1),
    .A(ui_in[0]));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[1]));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[2]));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_tielo tt_um_systolicLif_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\first.enable_Reg ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold2 (.A(\one.state[4] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold3 (.A(\third.enable_Reg ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold4 (.A(_037_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mac_Out_two[2] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mac_Out_two[4] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold7 (.A(\fourth.accumulate[2] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold8 (.A(_030_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold9 (.A(\fourth.accumulate[3] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold10 (.A(_031_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold11 (.A(\fourth.accumulate[1] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold12 (.A(_029_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold13 (.A(\first.out_data[3] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold14 (.A(_042_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold15 (.A(\one.state[5] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold16 (.A(\second.enable_Reg ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold17 (.A(\four.state[2] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold18 (.A(_134_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold19 (.A(_006_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold20 (.A(\two.state[4] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold21 (.A(\first.out_data[4] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold22 (.A(_203_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold23 (.A(\three.state[3] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold24 (.A(_084_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold25 (.A(\one.state[6] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold26 (.A(\first.out_data[6] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold27 (.A(\fourth.out_data[6] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold28 (.A(\fourth.enable_Reg ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold29 (.A(_034_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold30 (.A(\fourth.accumulate[4] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold31 (.A(_122_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold32 (.A(\fourth.accumulate[6] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold33 (.A(_112_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold34 (.A(\mac_Out_two[5] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold35 (.A(\mac_Out_two[6] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mac_Out_two[6] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold37 (.A(\two.state[5] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold38 (.A(_216_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold39 (.A(\fourth.out_data[4] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold40 (.A(_156_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold41 (.A(_009_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold42 (.A(\two.state[7] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold43 (.A(\three.state[7] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold44 (.A(\two.state[6] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold45 (.A(\one.state[7] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold46 (.A(\four.state[4] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold47 (.A(_008_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold48 (.A(\three.state[3] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold49 (.A(\mac_Out_two[3] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold50 (.A(\fourth.out_data[5] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold51 (.A(_161_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold52 (.A(\three.state[6] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold53 (.A(_100_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold54 (.A(\one.state[7] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold55 (.A(_062_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold56 (.A(\four.state[4] ),
    .X(net136));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_4 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_254 ();
 sg13g2_fill_2 FILLER_21_261 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_fill_2 FILLER_21_268 ();
 sg13g2_fill_1 FILLER_21_270 ();
 sg13g2_decap_8 FILLER_21_297 ();
 sg13g2_decap_8 FILLER_21_304 ();
 sg13g2_decap_8 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_318 ();
 sg13g2_decap_8 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_21_339 ();
 sg13g2_decap_8 FILLER_21_346 ();
 sg13g2_decap_8 FILLER_21_353 ();
 sg13g2_decap_8 FILLER_21_360 ();
 sg13g2_decap_8 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_374 ();
 sg13g2_decap_8 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_fill_2 FILLER_22_236 ();
 sg13g2_fill_1 FILLER_22_238 ();
 sg13g2_decap_4 FILLER_22_243 ();
 sg13g2_fill_2 FILLER_22_252 ();
 sg13g2_fill_2 FILLER_22_280 ();
 sg13g2_fill_2 FILLER_22_286 ();
 sg13g2_fill_1 FILLER_22_288 ();
 sg13g2_fill_1 FILLER_22_293 ();
 sg13g2_decap_8 FILLER_22_302 ();
 sg13g2_decap_8 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_decap_8 FILLER_22_323 ();
 sg13g2_decap_8 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_fill_1 FILLER_23_210 ();
 sg13g2_fill_2 FILLER_23_237 ();
 sg13g2_fill_1 FILLER_23_239 ();
 sg13g2_decap_4 FILLER_23_280 ();
 sg13g2_fill_1 FILLER_23_284 ();
 sg13g2_fill_1 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_decap_8 FILLER_23_335 ();
 sg13g2_decap_8 FILLER_23_342 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_23_363 ();
 sg13g2_decap_4 FILLER_23_370 ();
 sg13g2_fill_1 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_fill_2 FILLER_24_168 ();
 sg13g2_fill_1 FILLER_24_170 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_fill_2 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_217 ();
 sg13g2_fill_2 FILLER_24_279 ();
 sg13g2_fill_1 FILLER_24_281 ();
 sg13g2_decap_4 FILLER_24_323 ();
 sg13g2_fill_2 FILLER_24_327 ();
 sg13g2_decap_8 FILLER_24_333 ();
 sg13g2_decap_8 FILLER_24_340 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_fill_2 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_4 FILLER_25_154 ();
 sg13g2_fill_2 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_193 ();
 sg13g2_fill_2 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_4 FILLER_25_231 ();
 sg13g2_fill_2 FILLER_25_235 ();
 sg13g2_fill_2 FILLER_25_284 ();
 sg13g2_fill_1 FILLER_25_286 ();
 sg13g2_fill_1 FILLER_25_318 ();
 sg13g2_decap_4 FILLER_25_345 ();
 sg13g2_fill_1 FILLER_25_352 ();
 sg13g2_fill_1 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_4 FILLER_26_119 ();
 sg13g2_fill_2 FILLER_26_123 ();
 sg13g2_decap_4 FILLER_26_159 ();
 sg13g2_fill_1 FILLER_26_163 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_194 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_fill_1 FILLER_26_255 ();
 sg13g2_decap_8 FILLER_26_275 ();
 sg13g2_fill_2 FILLER_26_282 ();
 sg13g2_fill_2 FILLER_26_289 ();
 sg13g2_fill_2 FILLER_26_296 ();
 sg13g2_fill_2 FILLER_26_342 ();
 sg13g2_decap_4 FILLER_26_359 ();
 sg13g2_fill_2 FILLER_26_377 ();
 sg13g2_fill_2 FILLER_26_388 ();
 sg13g2_fill_1 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_fill_2 FILLER_27_126 ();
 sg13g2_fill_1 FILLER_27_128 ();
 sg13g2_fill_1 FILLER_27_146 ();
 sg13g2_fill_1 FILLER_27_154 ();
 sg13g2_fill_1 FILLER_27_176 ();
 sg13g2_fill_1 FILLER_27_192 ();
 sg13g2_decap_8 FILLER_27_233 ();
 sg13g2_fill_2 FILLER_27_240 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_262 ();
 sg13g2_decap_8 FILLER_27_267 ();
 sg13g2_fill_1 FILLER_27_309 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_decap_4 FILLER_27_348 ();
 sg13g2_fill_1 FILLER_27_352 ();
 sg13g2_fill_1 FILLER_27_358 ();
 sg13g2_fill_2 FILLER_27_364 ();
 sg13g2_fill_2 FILLER_27_371 ();
 sg13g2_fill_1 FILLER_27_373 ();
 sg13g2_fill_1 FILLER_27_379 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_172 ();
 sg13g2_fill_2 FILLER_28_198 ();
 sg13g2_fill_1 FILLER_28_220 ();
 sg13g2_fill_1 FILLER_28_230 ();
 sg13g2_fill_1 FILLER_28_251 ();
 sg13g2_decap_4 FILLER_28_278 ();
 sg13g2_fill_2 FILLER_28_282 ();
 sg13g2_fill_2 FILLER_28_288 ();
 sg13g2_decap_4 FILLER_28_331 ();
 sg13g2_fill_2 FILLER_28_335 ();
 sg13g2_decap_4 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_fill_2 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_4 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_130 ();
 sg13g2_decap_8 FILLER_29_135 ();
 sg13g2_fill_2 FILLER_29_142 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_170 ();
 sg13g2_decap_4 FILLER_29_177 ();
 sg13g2_decap_4 FILLER_29_211 ();
 sg13g2_fill_1 FILLER_29_215 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_fill_2 FILLER_29_231 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_decap_8 FILLER_29_239 ();
 sg13g2_fill_2 FILLER_29_246 ();
 sg13g2_fill_1 FILLER_29_248 ();
 sg13g2_decap_4 FILLER_29_345 ();
 sg13g2_fill_2 FILLER_29_349 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_119 ();
 sg13g2_fill_2 FILLER_30_159 ();
 sg13g2_fill_1 FILLER_30_161 ();
 sg13g2_fill_1 FILLER_30_167 ();
 sg13g2_decap_8 FILLER_30_178 ();
 sg13g2_decap_8 FILLER_30_185 ();
 sg13g2_fill_2 FILLER_30_209 ();
 sg13g2_fill_1 FILLER_30_234 ();
 sg13g2_fill_1 FILLER_30_251 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_327 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_338 ();
 sg13g2_decap_8 FILLER_30_345 ();
 sg13g2_fill_1 FILLER_30_352 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_fill_2 FILLER_31_119 ();
 sg13g2_fill_1 FILLER_31_121 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_fill_1 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_214 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_fill_1 FILLER_31_251 ();
 sg13g2_fill_1 FILLER_31_268 ();
 sg13g2_fill_2 FILLER_31_315 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_166 ();
 sg13g2_fill_1 FILLER_32_179 ();
 sg13g2_decap_4 FILLER_32_224 ();
 sg13g2_fill_2 FILLER_32_241 ();
 sg13g2_decap_4 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_268 ();
 sg13g2_fill_2 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_309 ();
 sg13g2_fill_2 FILLER_32_345 ();
 sg13g2_fill_1 FILLER_32_347 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_fill_1 FILLER_33_174 ();
 sg13g2_fill_2 FILLER_33_216 ();
 sg13g2_fill_1 FILLER_33_218 ();
 sg13g2_fill_2 FILLER_33_255 ();
 sg13g2_fill_2 FILLER_33_262 ();
 sg13g2_fill_1 FILLER_33_264 ();
 sg13g2_fill_2 FILLER_33_270 ();
 sg13g2_fill_1 FILLER_33_272 ();
 sg13g2_fill_2 FILLER_33_278 ();
 sg13g2_decap_4 FILLER_33_326 ();
 sg13g2_decap_4 FILLER_33_334 ();
 sg13g2_fill_2 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_369 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_4 FILLER_34_154 ();
 sg13g2_fill_2 FILLER_34_330 ();
 sg13g2_fill_1 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_4 FILLER_35_168 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_fill_1 FILLER_35_187 ();
 sg13g2_decap_8 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_decap_4 FILLER_35_214 ();
 sg13g2_fill_2 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_233 ();
 sg13g2_fill_1 FILLER_35_235 ();
 sg13g2_fill_2 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_278 ();
 sg13g2_decap_8 FILLER_35_293 ();
 sg13g2_decap_8 FILLER_35_300 ();
 sg13g2_decap_4 FILLER_35_307 ();
 sg13g2_fill_1 FILLER_35_336 ();
 sg13g2_fill_2 FILLER_35_360 ();
 sg13g2_fill_1 FILLER_35_383 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_4 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_198 ();
 sg13g2_decap_8 FILLER_36_205 ();
 sg13g2_decap_8 FILLER_36_212 ();
 sg13g2_decap_8 FILLER_36_219 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_decap_4 FILLER_36_242 ();
 sg13g2_decap_4 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_289 ();
 sg13g2_decap_8 FILLER_36_296 ();
 sg13g2_decap_4 FILLER_36_303 ();
 sg13g2_fill_1 FILLER_36_307 ();
 sg13g2_fill_2 FILLER_36_323 ();
 sg13g2_fill_1 FILLER_36_330 ();
 sg13g2_fill_2 FILLER_36_380 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_fill_2 FILLER_37_301 ();
 sg13g2_fill_1 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_decap_4 FILLER_38_220 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_decap_4 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_244 ();
 sg13g2_decap_8 FILLER_38_251 ();
 sg13g2_decap_8 FILLER_38_258 ();
 sg13g2_decap_8 FILLER_38_265 ();
 sg13g2_decap_8 FILLER_38_272 ();
 sg13g2_decap_8 FILLER_38_279 ();
 sg13g2_decap_8 FILLER_38_286 ();
 sg13g2_decap_8 FILLER_38_293 ();
 sg13g2_decap_8 FILLER_38_300 ();
 sg13g2_decap_8 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_314 ();
 sg13g2_fill_1 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_351 ();
 sg13g2_fill_2 FILLER_38_368 ();
 sg13g2_fill_1 FILLER_38_370 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net8;
 assign uio_oe[3] = net9;
 assign uio_oe[4] = net10;
 assign uio_oe[5] = net11;
 assign uio_oe[6] = net12;
 assign uio_oe[7] = net80;
 assign uio_out[0] = net13;
 assign uio_out[1] = net14;
 assign uio_out[2] = net15;
 assign uio_out[3] = net16;
 assign uio_out[4] = net17;
 assign uio_out[5] = net18;
 assign uio_out[6] = net19;
 assign uio_out[7] = net20;
 assign uo_out[0] = net21;
 assign uo_out[1] = net22;
 assign uo_out[2] = net23;
 assign uo_out[3] = net24;
endmodule

module tt_um_algofoogle_vga (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire \clock_color_offset[0] ;
 wire \clock_color_offset[1] ;
 wire \clock_color_offset[2] ;
 wire \clock_hrs_d[0] ;
 wire \clock_hrs_d[1] ;
 wire \clock_hrs_u[0] ;
 wire \clock_hrs_u[1] ;
 wire \clock_hrs_u[2] ;
 wire \clock_hrs_u[3] ;
 wire \clock_min_d[0] ;
 wire \clock_min_d[1] ;
 wire \clock_min_d[2] ;
 wire \clock_min_u[0] ;
 wire \clock_min_u[1] ;
 wire \clock_min_u[2] ;
 wire \clock_min_u[3] ;
 wire \clock_sec_d[0] ;
 wire \clock_sec_d[1] ;
 wire \clock_sec_d[2] ;
 wire \clock_sec_u[0] ;
 wire \clock_sec_u[1] ;
 wire \clock_sec_u[2] ;
 wire \clock_sec_u[3] ;
 wire dx;
 wire \h[0] ;
 wire \h[1] ;
 wire \h[2] ;
 wire \h[3] ;
 wire \h[4] ;
 wire \h[5] ;
 wire \h[6] ;
 wire \h[7] ;
 wire \h[8] ;
 wire \h[9] ;
 wire hblank;
 wire hmax;
 wire \matt_venn_clock.pulse_hrs.comp[0] ;
 wire \matt_venn_clock.pulse_hrs.comp[1] ;
 wire \matt_venn_clock.pulse_hrs.comp[2] ;
 wire \matt_venn_clock.pulse_hrs.comp[3] ;
 wire \matt_venn_clock.pulse_hrs.comp[4] ;
 wire \matt_venn_clock.pulse_hrs.count[0] ;
 wire \matt_venn_clock.pulse_hrs.count[1] ;
 wire \matt_venn_clock.pulse_hrs.count[2] ;
 wire \matt_venn_clock.pulse_hrs.count[3] ;
 wire \matt_venn_clock.pulse_hrs.count[4] ;
 wire \matt_venn_clock.pulse_min.comp[0] ;
 wire \matt_venn_clock.pulse_min.comp[1] ;
 wire \matt_venn_clock.pulse_min.comp[2] ;
 wire \matt_venn_clock.pulse_min.comp[3] ;
 wire \matt_venn_clock.pulse_min.comp[4] ;
 wire \matt_venn_clock.pulse_min.count[0] ;
 wire \matt_venn_clock.pulse_min.count[1] ;
 wire \matt_venn_clock.pulse_min.count[2] ;
 wire \matt_venn_clock.pulse_min.count[3] ;
 wire \matt_venn_clock.pulse_min.count[4] ;
 wire \matt_venn_clock.pulse_sec.comp[0] ;
 wire \matt_venn_clock.pulse_sec.comp[1] ;
 wire \matt_venn_clock.pulse_sec.comp[2] ;
 wire \matt_venn_clock.pulse_sec.comp[3] ;
 wire \matt_venn_clock.pulse_sec.comp[4] ;
 wire \matt_venn_clock.pulse_sec.count[0] ;
 wire \matt_venn_clock.pulse_sec.count[1] ;
 wire \matt_venn_clock.pulse_sec.count[2] ;
 wire \matt_venn_clock.pulse_sec.count[3] ;
 wire \matt_venn_clock.pulse_sec.count[4] ;
 wire \matt_venn_clock.sec_counter[0] ;
 wire \matt_venn_clock.sec_counter[10] ;
 wire \matt_venn_clock.sec_counter[11] ;
 wire \matt_venn_clock.sec_counter[12] ;
 wire \matt_venn_clock.sec_counter[13] ;
 wire \matt_venn_clock.sec_counter[14] ;
 wire \matt_venn_clock.sec_counter[15] ;
 wire \matt_venn_clock.sec_counter[16] ;
 wire \matt_venn_clock.sec_counter[17] ;
 wire \matt_venn_clock.sec_counter[18] ;
 wire \matt_venn_clock.sec_counter[19] ;
 wire \matt_venn_clock.sec_counter[1] ;
 wire \matt_venn_clock.sec_counter[20] ;
 wire \matt_venn_clock.sec_counter[21] ;
 wire \matt_venn_clock.sec_counter[22] ;
 wire \matt_venn_clock.sec_counter[23] ;
 wire \matt_venn_clock.sec_counter[24] ;
 wire \matt_venn_clock.sec_counter[2] ;
 wire \matt_venn_clock.sec_counter[3] ;
 wire \matt_venn_clock.sec_counter[4] ;
 wire \matt_venn_clock.sec_counter[5] ;
 wire \matt_venn_clock.sec_counter[6] ;
 wire \matt_venn_clock.sec_counter[7] ;
 wire \matt_venn_clock.sec_counter[8] ;
 wire \matt_venn_clock.sec_counter[9] ;
 wire \matt_venn_vga.activevideo ;
 wire \matt_venn_vga.col_index[0] ;
 wire \matt_venn_vga.col_index[1] ;
 wire \matt_venn_vga.col_index_q[0] ;
 wire \matt_venn_vga.col_index_q[1] ;
 wire \matt_venn_vga.color[0] ;
 wire \matt_venn_vga.color[1] ;
 wire \matt_venn_vga.color[2] ;
 wire \matt_venn_vga.color[3] ;
 wire \matt_venn_vga.color[4] ;
 wire \matt_venn_vga.color[5] ;
 wire \matt_venn_vga.digit_0.char[0] ;
 wire \matt_venn_vga.digit_0.digit_index[0] ;
 wire \matt_venn_vga.digit_0.digit_index[1] ;
 wire \matt_venn_vga.digit_0.digit_index[2] ;
 wire \matt_venn_vga.digit_0.digit_index[3] ;
 wire \matt_venn_vga.digit_0.digit_index[4] ;
 wire \matt_venn_vga.digit_0.digit_index[5] ;
 wire \matt_venn_vga.draw ;
 wire \matt_venn_vga.font_0.dout[1] ;
 wire \matt_venn_vga.font_0.dout[2] ;
 wire \matt_venn_vga.font_0.dout[3] ;
 wire \matt_venn_vga.x_block_q[5] ;
 wire \matt_venn_vga.y_block_q[0] ;
 wire \matt_venn_vga.y_block_q[1] ;
 wire \matt_venn_vga.y_block_q[2] ;
 wire \matt_venn_vga.y_block_q[3] ;
 wire \matt_venn_vga.y_block_q[4] ;
 wire \matt_venn_vga.y_block_q[5] ;
 wire \matt_venn_vga.y_px[0] ;
 wire \matt_venn_vga.y_px[1] ;
 wire \matt_venn_vga.y_px[2] ;
 wire \matt_venn_vga.y_px[3] ;
 wire \matt_venn_vga.y_px[4] ;
 wire \matt_venn_vga.y_px[5] ;
 wire \matt_venn_vga.y_px[6] ;
 wire \matt_venn_vga.y_px[7] ;
 wire \matt_venn_vga.y_px[8] ;
 wire \matt_venn_vga.y_px[9] ;
 wire \matt_venn_vga_shadow.col_index[0] ;
 wire \matt_venn_vga_shadow.col_index[1] ;
 wire \matt_venn_vga_shadow.col_index_q[0] ;
 wire \matt_venn_vga_shadow.col_index_q[1] ;
 wire \matt_venn_vga_shadow.color[0] ;
 wire \matt_venn_vga_shadow.color[1] ;
 wire \matt_venn_vga_shadow.color[2] ;
 wire \matt_venn_vga_shadow.color[3] ;
 wire \matt_venn_vga_shadow.color[4] ;
 wire \matt_venn_vga_shadow.color[5] ;
 wire \matt_venn_vga_shadow.digit_0.digit_index[0] ;
 wire \matt_venn_vga_shadow.digit_0.digit_index[1] ;
 wire \matt_venn_vga_shadow.digit_0.digit_index[2] ;
 wire \matt_venn_vga_shadow.digit_0.digit_index[3] ;
 wire \matt_venn_vga_shadow.digit_0.digit_index[4] ;
 wire \matt_venn_vga_shadow.digit_0.digit_index[5] ;
 wire \matt_venn_vga_shadow.draw ;
 wire \matt_venn_vga_shadow.font_0.dout[1] ;
 wire \matt_venn_vga_shadow.font_0.dout[2] ;
 wire \matt_venn_vga_shadow.font_0.dout[3] ;
 wire \matt_venn_vga_shadow.x_block_q[5] ;
 wire \matt_venn_vga_shadow.y_block_q[0] ;
 wire \matt_venn_vga_shadow.y_block_q[1] ;
 wire \matt_venn_vga_shadow.y_block_q[2] ;
 wire \matt_venn_vga_shadow.y_block_q[3] ;
 wire \matt_venn_vga_shadow.y_block_q[4] ;
 wire \matt_venn_vga_shadow.y_block_q[5] ;
 wire \product_comp[10] ;
 wire \product_comp[1] ;
 wire \product_comp[2] ;
 wire \product_comp[3] ;
 wire \product_comp[4] ;
 wire \product_comp[5] ;
 wire \product_comp[6] ;
 wire \product_comp[7] ;
 wire \product_comp[8] ;
 wire \product_comp[9] ;
 wire product_comp_dir;
 wire \px[0] ;
 wire \px[1] ;
 wire \px[2] ;
 wire \px[3] ;
 wire \px[4] ;
 wire \px[5] ;
 wire \px[6] ;
 wire \px[7] ;
 wire \px[8] ;
 wire \px[9] ;
 wire \pxm[0] ;
 wire \pxm[1] ;
 wire \py[0] ;
 wire \py[1] ;
 wire \py[2] ;
 wire \py[3] ;
 wire \py[4] ;
 wire \py[5] ;
 wire \py[6] ;
 wire \py[7] ;
 wire \py[8] ;
 wire \py[9] ;
 wire \pym[10] ;
 wire \pym[11] ;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire clknet_0_clk;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire vblank;
 wire \vga_sync.hsync ;
 wire \vga_sync.o_vmax ;
 wire \vga_sync.vsync ;
 wire \ydelta[0] ;
 wire \ydelta[1] ;
 wire \ydelta[2] ;
 wire \ydelta[3] ;
 wire \ydelta[4] ;
 wire \ydelta[5] ;
 wire \ydelta[6] ;
 wire \ydelta[7] ;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;

 sg13g2_inv_1 _2044_ (.Y(_1176_),
    .A(\product_comp[10] ));
 sg13g2_inv_1 _2045_ (.Y(_1177_),
    .A(\product_comp[9] ));
 sg13g2_inv_1 _2046_ (.Y(_1178_),
    .A(\product_comp[8] ));
 sg13g2_inv_1 _2047_ (.Y(_1179_),
    .A(net230));
 sg13g2_inv_1 _2048_ (.Y(_1180_),
    .A(net375));
 sg13g2_inv_2 _2049_ (.Y(_1181_),
    .A(net497));
 sg13g2_inv_1 _2050_ (.Y(_1182_),
    .A(\clock_min_d[0] ));
 sg13g2_inv_1 _2051_ (.Y(_1183_),
    .A(\clock_hrs_d[0] ));
 sg13g2_inv_1 _2052_ (.Y(_1184_),
    .A(net221));
 sg13g2_inv_1 _2053_ (.Y(_1185_),
    .A(net268));
 sg13g2_inv_1 _2054_ (.Y(_1186_),
    .A(net487));
 sg13g2_inv_1 _2055_ (.Y(_1187_),
    .A(net451));
 sg13g2_inv_1 _2056_ (.Y(_1188_),
    .A(net530));
 sg13g2_inv_1 _2057_ (.Y(_1189_),
    .A(net493));
 sg13g2_inv_1 _2058_ (.Y(_1190_),
    .A(\matt_venn_clock.pulse_min.comp[4] ));
 sg13g2_inv_1 _2059_ (.Y(_1191_),
    .A(net397));
 sg13g2_inv_1 _2060_ (.Y(_1192_),
    .A(net440));
 sg13g2_inv_1 _2061_ (.Y(_1193_),
    .A(net269));
 sg13g2_inv_1 _2062_ (.Y(_1194_),
    .A(net443));
 sg13g2_inv_1 _2063_ (.Y(_1195_),
    .A(net524));
 sg13g2_inv_1 _2064_ (.Y(_1196_),
    .A(net475));
 sg13g2_inv_1 _2065_ (.Y(_1197_),
    .A(net319));
 sg13g2_inv_2 _2066_ (.Y(_1198_),
    .A(net321));
 sg13g2_inv_1 _2067_ (.Y(_1199_),
    .A(net327));
 sg13g2_inv_1 _2068_ (.Y(_1200_),
    .A(\matt_venn_vga.y_px[1] ));
 sg13g2_inv_2 _2069_ (.Y(_1201_),
    .A(net335));
 sg13g2_inv_2 _2070_ (.Y(_1202_),
    .A(net337));
 sg13g2_inv_2 _2071_ (.Y(_1203_),
    .A(\py[6] ));
 sg13g2_inv_2 _2072_ (.Y(_1204_),
    .A(net507));
 sg13g2_inv_1 _2073_ (.Y(_1205_),
    .A(net343));
 sg13g2_inv_1 _2074_ (.Y(_1206_),
    .A(net344));
 sg13g2_inv_1 _2075_ (.Y(_1207_),
    .A(net503));
 sg13g2_inv_1 _2076_ (.Y(_1208_),
    .A(net417));
 sg13g2_inv_1 _2077_ (.Y(_1209_),
    .A(net349));
 sg13g2_inv_1 _2078_ (.Y(_1210_),
    .A(net468));
 sg13g2_inv_1 _2079_ (.Y(_1211_),
    .A(net472));
 sg13g2_inv_1 _2080_ (.Y(_1212_),
    .A(net476));
 sg13g2_inv_1 _2081_ (.Y(_1213_),
    .A(net309));
 sg13g2_inv_1 _2082_ (.Y(_1214_),
    .A(_0051_));
 sg13g2_inv_2 _2083_ (.Y(_1215_),
    .A(net313));
 sg13g2_inv_2 _2084_ (.Y(_1216_),
    .A(\h[3] ));
 sg13g2_inv_2 _2085_ (.Y(_1217_),
    .A(\h[9] ));
 sg13g2_inv_1 _2086_ (.Y(_1218_),
    .A(net316));
 sg13g2_inv_1 _2087_ (.Y(_1219_),
    .A(net364));
 sg13g2_inv_1 _2088_ (.Y(_1220_),
    .A(net1));
 sg13g2_inv_2 _2089_ (.Y(_1221_),
    .A(_0057_));
 sg13g2_inv_2 _2090_ (.Y(_1222_),
    .A(_0023_));
 sg13g2_inv_1 _2091_ (.Y(_1223_),
    .A(_0024_));
 sg13g2_inv_1 _2092_ (.Y(_1224_),
    .A(_0028_));
 sg13g2_inv_1 _2093_ (.Y(_1225_),
    .A(_0029_));
 sg13g2_inv_1 _2094_ (.Y(_1226_),
    .A(\matt_venn_vga.color[3] ));
 sg13g2_inv_1 _2095_ (.Y(_1227_),
    .A(\matt_venn_vga.color[4] ));
 sg13g2_inv_1 _2096_ (.Y(_1228_),
    .A(net356));
 sg13g2_inv_1 _2097_ (.Y(_1229_),
    .A(_0035_));
 sg13g2_inv_1 _2098_ (.Y(_1230_),
    .A(_0038_));
 sg13g2_inv_1 _2099_ (.Y(_1231_),
    .A(_0036_));
 sg13g2_inv_1 _2100_ (.Y(_1232_),
    .A(\matt_venn_vga.font_0.dout[2] ));
 sg13g2_inv_1 _2101_ (.Y(_1233_),
    .A(\matt_venn_vga.col_index_q[1] ));
 sg13g2_inv_1 _2102_ (.Y(_1234_),
    .A(\matt_venn_vga_shadow.font_0.dout[2] ));
 sg13g2_inv_1 _2103_ (.Y(_1235_),
    .A(\matt_venn_vga_shadow.col_index_q[1] ));
 sg13g2_and2_2 _2104_ (.A(\h[0] ),
    .B(net505),
    .X(_1236_));
 sg13g2_nor2_1 _2105_ (.A(_0050_),
    .B(net311),
    .Y(_1237_));
 sg13g2_nand4_1 _2106_ (.B(\h[3] ),
    .C(_1236_),
    .A(net314),
    .Y(_1238_),
    .D(_1237_));
 sg13g2_or2_1 _2107_ (.X(_1239_),
    .B(net354),
    .A(net307));
 sg13g2_o21ai_1 _2108_ (.B1(_1239_),
    .Y(_1240_),
    .A1(net315),
    .A2(net305));
 sg13g2_a22oi_1 _2109_ (.Y(_1241_),
    .B1(net354),
    .B2(net307),
    .A2(\h[9] ),
    .A1(\h[2] ));
 sg13g2_inv_1 _2110_ (.Y(_1242_),
    .A(_1241_));
 sg13g2_nor2_2 _2111_ (.A(net307),
    .B(net310),
    .Y(_1243_));
 sg13g2_nand2_2 _2112_ (.Y(_1244_),
    .A(net307),
    .B(net309));
 sg13g2_inv_1 _2113_ (.Y(_1245_),
    .A(_1244_));
 sg13g2_nand2b_2 _2114_ (.Y(_1246_),
    .B(_1244_),
    .A_N(_1243_));
 sg13g2_nand3_1 _2115_ (.B(_1242_),
    .C(_1246_),
    .A(_1240_),
    .Y(_1247_));
 sg13g2_nor2_2 _2116_ (.A(_1238_),
    .B(_1247_),
    .Y(hmax));
 sg13g2_nand2_2 _2117_ (.Y(_1248_),
    .A(net319),
    .B(net320));
 sg13g2_nor3_1 _2118_ (.A(net328),
    .B(net330),
    .C(_1248_),
    .Y(_1249_));
 sg13g2_nand4_1 _2119_ (.B(net333),
    .C(net354),
    .A(\matt_venn_vga.y_px[1] ),
    .Y(_1250_),
    .D(_1249_));
 sg13g2_nand2_1 _2120_ (.Y(_1251_),
    .A(net325),
    .B(_1250_));
 sg13g2_nand2_2 _2121_ (.Y(_1252_),
    .A(net328),
    .B(net329));
 sg13g2_inv_1 _2122_ (.Y(_1253_),
    .A(_1252_));
 sg13g2_or2_1 _2123_ (.X(_1254_),
    .B(net333),
    .A(\matt_venn_vga.y_px[1] ));
 sg13g2_or2_1 _2124_ (.X(_1255_),
    .B(_1254_),
    .A(_1252_));
 sg13g2_nor4_1 _2125_ (.A(net319),
    .B(net320),
    .C(net355),
    .D(_1255_),
    .Y(_1256_));
 sg13g2_or2_1 _2126_ (.X(_1257_),
    .B(_1256_),
    .A(net325));
 sg13g2_nor3_1 _2127_ (.A(net322),
    .B(net326),
    .C(_0052_),
    .Y(_1258_));
 sg13g2_and3_2 _2128_ (.X(\vga_sync.o_vmax ),
    .A(_1251_),
    .B(_1257_),
    .C(_1258_));
 sg13g2_a21oi_1 _2129_ (.A1(net305),
    .A2(_1239_),
    .Y(_1259_),
    .B1(\h[8] ));
 sg13g2_nand2_1 _2130_ (.Y(_1260_),
    .A(_1215_),
    .B(_1216_));
 sg13g2_nand4_1 _2131_ (.B(\h[5] ),
    .C(net354),
    .A(net309),
    .Y(_1261_),
    .D(_1260_));
 sg13g2_a21oi_1 _2132_ (.A1(net307),
    .A2(net354),
    .Y(_1262_),
    .B1(\h[9] ));
 sg13g2_a21o_1 _2133_ (.A2(_1262_),
    .A1(_1261_),
    .B1(_1259_),
    .X(_1263_));
 sg13g2_inv_1 _2134_ (.Y(hblank),
    .A(_1263_));
 sg13g2_nand2_1 _2135_ (.Y(_1264_),
    .A(net321),
    .B(net323));
 sg13g2_nor2_2 _2136_ (.A(_1197_),
    .B(net326),
    .Y(_1265_));
 sg13g2_nor2b_1 _2137_ (.A(net317),
    .B_N(net325),
    .Y(_1266_));
 sg13g2_nand4_1 _2138_ (.B(net322),
    .C(_1265_),
    .A(net320),
    .Y(_1267_),
    .D(_1266_));
 sg13g2_or4_1 _2139_ (.A(net328),
    .B(net329),
    .C(_1254_),
    .D(_1267_),
    .X(_1268_));
 sg13g2_nand4_1 _2140_ (.B(net320),
    .C(net322),
    .A(net319),
    .Y(_1269_),
    .D(_1221_));
 sg13g2_a21oi_1 _2141_ (.A1(_1268_),
    .A2(_1269_),
    .Y(_1270_),
    .B1(net355));
 sg13g2_or2_2 _2142_ (.X(_1271_),
    .B(net328),
    .A(net326));
 sg13g2_nor3_2 _2143_ (.A(net322),
    .B(net325),
    .C(_1271_),
    .Y(_1272_));
 sg13g2_nor2b_1 _2144_ (.A(net329),
    .B_N(_1272_),
    .Y(_1273_));
 sg13g2_o21ai_1 _2145_ (.B1(net355),
    .Y(_1274_),
    .A1(_1248_),
    .A2(_1273_));
 sg13g2_o21ai_1 _2146_ (.B1(_1274_),
    .Y(_1275_),
    .A1(net318),
    .A2(_1270_));
 sg13g2_inv_1 _2147_ (.Y(vblank),
    .A(_1275_));
 sg13g2_nor2_2 _2148_ (.A(hblank),
    .B(vblank),
    .Y(\matt_venn_vga.activevideo ));
 sg13g2_nand2_2 _2149_ (.Y(_1276_),
    .A(_1228_),
    .B(\matt_venn_vga.activevideo ));
 sg13g2_nor3_2 _2150_ (.A(_1198_),
    .B(net322),
    .C(net325),
    .Y(_1277_));
 sg13g2_nor2b_1 _2151_ (.A(net317),
    .B_N(_1277_),
    .Y(_1278_));
 sg13g2_nor2_1 _2152_ (.A(_1200_),
    .B(net333),
    .Y(_1279_));
 sg13g2_nand4_1 _2153_ (.B(net329),
    .C(_1278_),
    .A(net319),
    .Y(_1280_),
    .D(_1279_));
 sg13g2_nand2_2 _2154_ (.Y(_1281_),
    .A(net326),
    .B(net327));
 sg13g2_nor2_1 _2155_ (.A(_1280_),
    .B(_1281_),
    .Y(_1282_));
 sg13g2_a21oi_1 _2156_ (.A1(_1277_),
    .A2(_1281_),
    .Y(_1283_),
    .B1(_1248_));
 sg13g2_nor2_1 _2157_ (.A(net317),
    .B(_1283_),
    .Y(_1284_));
 sg13g2_or2_1 _2158_ (.X(_1285_),
    .B(_1283_),
    .A(net317));
 sg13g2_nand3_1 _2159_ (.B(net331),
    .C(net333),
    .A(net329),
    .Y(_1286_));
 sg13g2_nand3_1 _2160_ (.B(_1278_),
    .C(_1286_),
    .A(net326),
    .Y(_1287_));
 sg13g2_a21oi_1 _2161_ (.A1(_1285_),
    .A2(_1287_),
    .Y(_1288_),
    .B1(_1282_));
 sg13g2_inv_1 _2162_ (.Y(_1289_),
    .A(_1288_));
 sg13g2_a21oi_1 _2163_ (.A1(_1272_),
    .A2(_1286_),
    .Y(_1290_),
    .B1(_1248_));
 sg13g2_nor2_1 _2164_ (.A(net317),
    .B(_1290_),
    .Y(_1291_));
 sg13g2_o21ai_1 _2165_ (.B1(_1291_),
    .Y(_1292_),
    .A1(_1271_),
    .A2(_1280_));
 sg13g2_nand2_1 _2166_ (.Y(_1293_),
    .A(_1265_),
    .B(_1277_));
 sg13g2_nor4_1 _2167_ (.A(net327),
    .B(net329),
    .C(_1254_),
    .D(_1293_),
    .Y(_1294_));
 sg13g2_nor2_1 _2168_ (.A(net317),
    .B(_1294_),
    .Y(_1295_));
 sg13g2_o21ai_1 _2169_ (.B1(_1295_),
    .Y(_1296_),
    .A1(_1197_),
    .A2(_0031_));
 sg13g2_or2_1 _2170_ (.X(_1297_),
    .B(_1296_),
    .A(_1292_));
 sg13g2_nand3_1 _2171_ (.B(net5),
    .C(\matt_venn_vga.activevideo ),
    .A(\matt_venn_vga.draw ),
    .Y(_1298_));
 sg13g2_nand4_1 _2172_ (.B(\matt_venn_vga.color[5] ),
    .C(net5),
    .A(\matt_venn_vga.draw ),
    .Y(_1299_),
    .D(\matt_venn_vga.activevideo ));
 sg13g2_nor2_1 _2173_ (.A(net340),
    .B(\py[0] ),
    .Y(_1300_));
 sg13g2_nor3_1 _2174_ (.A(\py[2] ),
    .B(net340),
    .C(net341),
    .Y(_1301_));
 sg13g2_nor2b_1 _2175_ (.A(\py[3] ),
    .B_N(_1301_),
    .Y(_1302_));
 sg13g2_nor2b_1 _2176_ (.A(\py[4] ),
    .B_N(_1302_),
    .Y(_1303_));
 sg13g2_nor2b_1 _2177_ (.A(\py[5] ),
    .B_N(_1303_),
    .Y(_1304_));
 sg13g2_nand2_1 _2178_ (.Y(_1305_),
    .A(_1203_),
    .B(_1304_));
 sg13g2_nand3_1 _2179_ (.B(\py[7] ),
    .C(_1305_),
    .A(\py[8] ),
    .Y(_1306_));
 sg13g2_a21o_1 _2180_ (.A2(_1305_),
    .A1(\py[7] ),
    .B1(\py[8] ),
    .X(_1307_));
 sg13g2_and2_1 _2181_ (.A(_1306_),
    .B(_1307_),
    .X(_1308_));
 sg13g2_inv_1 _2182_ (.Y(_1309_),
    .A(_1308_));
 sg13g2_xnor2_1 _2183_ (.Y(_1310_),
    .A(\py[6] ),
    .B(_1304_));
 sg13g2_inv_1 _2184_ (.Y(_1311_),
    .A(_1310_));
 sg13g2_xnor2_1 _2185_ (.Y(_1312_),
    .A(\py[5] ),
    .B(_1303_));
 sg13g2_nand2b_1 _2186_ (.Y(_1313_),
    .B(net324),
    .A_N(_1312_));
 sg13g2_xnor2_1 _2187_ (.Y(_1314_),
    .A(net339),
    .B(_1302_));
 sg13g2_nand2_1 _2188_ (.Y(_1315_),
    .A(_0025_),
    .B(_1314_));
 sg13g2_nor2_1 _2189_ (.A(net331),
    .B(net340),
    .Y(_1316_));
 sg13g2_nand2_1 _2190_ (.Y(_1317_),
    .A(net332),
    .B(net341));
 sg13g2_a22oi_1 _2191_ (.Y(_1318_),
    .B1(net341),
    .B2(net332),
    .A2(net340),
    .A1(net331));
 sg13g2_nor2_1 _2192_ (.A(_1316_),
    .B(_1318_),
    .Y(_1319_));
 sg13g2_or2_1 _2193_ (.X(_1320_),
    .B(_1319_),
    .A(_1300_));
 sg13g2_xor2_1 _2194_ (.B(_1300_),
    .A(\py[2] ),
    .X(_1321_));
 sg13g2_xnor2_1 _2195_ (.Y(_1322_),
    .A(_0026_),
    .B(_1321_));
 sg13g2_a22oi_1 _2196_ (.Y(_1323_),
    .B1(_1322_),
    .B2(_1320_),
    .A2(_1321_),
    .A1(net330));
 sg13g2_xnor2_1 _2197_ (.Y(_1324_),
    .A(\py[3] ),
    .B(_1301_));
 sg13g2_xnor2_1 _2198_ (.Y(_1325_),
    .A(_1199_),
    .B(_1324_));
 sg13g2_nor2_1 _2199_ (.A(_0025_),
    .B(_1314_),
    .Y(_1326_));
 sg13g2_or2_1 _2200_ (.X(_1327_),
    .B(_1324_),
    .A(_0027_));
 sg13g2_o21ai_1 _2201_ (.B1(_1327_),
    .Y(_1328_),
    .A1(_1323_),
    .A2(_1325_));
 sg13g2_a21oi_1 _2202_ (.A1(_1315_),
    .A2(_1328_),
    .Y(_1329_),
    .B1(_1326_));
 sg13g2_nand2_1 _2203_ (.Y(_1330_),
    .A(_1221_),
    .B(_1312_));
 sg13g2_xnor2_1 _2204_ (.Y(_1331_),
    .A(_0057_),
    .B(_1312_));
 sg13g2_o21ai_1 _2205_ (.B1(_1313_),
    .Y(_1332_),
    .A1(_1329_),
    .A2(_1331_));
 sg13g2_xnor2_1 _2206_ (.Y(_1333_),
    .A(_1223_),
    .B(_1310_));
 sg13g2_a22oi_1 _2207_ (.Y(_1334_),
    .B1(_1332_),
    .B2(_1333_),
    .A2(_1311_),
    .A1(net323));
 sg13g2_xor2_1 _2208_ (.B(_1305_),
    .A(_0022_),
    .X(_1335_));
 sg13g2_inv_1 _2209_ (.Y(_1336_),
    .A(_1335_));
 sg13g2_a21oi_1 _2210_ (.A1(_1198_),
    .A2(_1335_),
    .Y(_1337_),
    .B1(_1334_));
 sg13g2_a221oi_1 _2211_ (.B2(net321),
    .C1(_1337_),
    .B1(_1336_),
    .A1(_1222_),
    .Y(_1338_),
    .A2(_1308_));
 sg13g2_a21oi_1 _2212_ (.A1(_0023_),
    .A2(_1309_),
    .Y(_1339_),
    .B1(_1338_));
 sg13g2_nand2_1 _2213_ (.Y(_1340_),
    .A(\px[6] ),
    .B(net517));
 sg13g2_nor2_1 _2214_ (.A(_0059_),
    .B(_1340_),
    .Y(_1341_));
 sg13g2_xnor2_1 _2215_ (.Y(_1342_),
    .A(_1204_),
    .B(_1341_));
 sg13g2_nor2b_1 _2216_ (.A(_1342_),
    .B_N(\h[8] ),
    .Y(_1343_));
 sg13g2_xnor2_1 _2217_ (.Y(_1344_),
    .A(\px[6] ),
    .B(net344));
 sg13g2_xnor2_1 _2218_ (.Y(_1345_),
    .A(\matt_venn_vga.digit_0.char[0] ),
    .B(_1344_));
 sg13g2_nor2b_2 _2219_ (.A(\h[0] ),
    .B_N(\px[0] ),
    .Y(_1346_));
 sg13g2_nor2b_1 _2220_ (.A(net346),
    .B_N(net316),
    .Y(_1347_));
 sg13g2_nor2b_1 _2221_ (.A(net316),
    .B_N(net346),
    .Y(_1348_));
 sg13g2_xnor2_1 _2222_ (.Y(_1349_),
    .A(net346),
    .B(net316));
 sg13g2_inv_1 _2223_ (.Y(_1350_),
    .A(_1349_));
 sg13g2_nand2b_1 _2224_ (.Y(_1351_),
    .B(_1349_),
    .A_N(_1346_));
 sg13g2_nand2b_1 _2225_ (.Y(_1352_),
    .B(net315),
    .A_N(\px[2] ));
 sg13g2_xor2_1 _2226_ (.B(net315),
    .A(\px[2] ),
    .X(_1353_));
 sg13g2_nor3_1 _2227_ (.A(net346),
    .B(_1218_),
    .C(_1353_),
    .Y(_1354_));
 sg13g2_xnor2_1 _2228_ (.Y(_1355_),
    .A(_1347_),
    .B(_1353_));
 sg13g2_nor4_1 _2229_ (.A(_1346_),
    .B(_1347_),
    .C(_1348_),
    .D(_1353_),
    .Y(_1356_));
 sg13g2_nor2_1 _2230_ (.A(\px[3] ),
    .B(_1216_),
    .Y(_1357_));
 sg13g2_xnor2_1 _2231_ (.Y(_1358_),
    .A(\px[3] ),
    .B(\h[3] ));
 sg13g2_nor2b_1 _2232_ (.A(_1352_),
    .B_N(_1358_),
    .Y(_1359_));
 sg13g2_xnor2_1 _2233_ (.Y(_1360_),
    .A(_1352_),
    .B(_1358_));
 sg13g2_a221oi_1 _2234_ (.B2(_1356_),
    .C1(_1359_),
    .B1(_1360_),
    .A1(_1354_),
    .Y(_1361_),
    .A2(_1358_));
 sg13g2_a21oi_1 _2235_ (.A1(_1207_),
    .A2(net313),
    .Y(_1362_),
    .B1(_1357_));
 sg13g2_a22oi_1 _2236_ (.Y(_1363_),
    .B1(_1361_),
    .B2(_1362_),
    .A2(_1215_),
    .A1(\px[4] ));
 sg13g2_a21oi_1 _2237_ (.A1(net344),
    .A2(net312),
    .Y(_1364_),
    .B1(_1363_));
 sg13g2_o21ai_1 _2238_ (.B1(_1345_),
    .Y(_1365_),
    .A1(net344),
    .A2(net312));
 sg13g2_xnor2_1 _2239_ (.Y(_1366_),
    .A(_0059_),
    .B(_1340_));
 sg13g2_a22oi_1 _2240_ (.Y(_1367_),
    .B1(_1366_),
    .B2(net308),
    .A2(_1344_),
    .A1(net309));
 sg13g2_o21ai_1 _2241_ (.B1(_1367_),
    .Y(_1368_),
    .A1(_1364_),
    .A2(_1365_));
 sg13g2_xor2_1 _2242_ (.B(_1342_),
    .A(_0050_),
    .X(_1369_));
 sg13g2_o21ai_1 _2243_ (.B1(_1368_),
    .Y(_1370_),
    .A1(net308),
    .A2(_1366_));
 sg13g2_inv_1 _2244_ (.Y(_1371_),
    .A(_1370_));
 sg13g2_a21oi_1 _2245_ (.A1(_1369_),
    .A2(_1371_),
    .Y(_1372_),
    .B1(_1343_));
 sg13g2_nor2_1 _2246_ (.A(\px[9] ),
    .B(_1217_),
    .Y(_1373_));
 sg13g2_nand2_1 _2247_ (.Y(_1374_),
    .A(\px[9] ),
    .B(_1217_));
 sg13g2_nand4_1 _2248_ (.B(\px[7] ),
    .C(net343),
    .A(\px[8] ),
    .Y(_1375_),
    .D(net344));
 sg13g2_a21oi_1 _2249_ (.A1(_1374_),
    .A2(_1375_),
    .Y(_1376_),
    .B1(_1373_));
 sg13g2_nor2_1 _2250_ (.A(_1372_),
    .B(_1376_),
    .Y(_1377_));
 sg13g2_nor2_1 _2251_ (.A(_1310_),
    .B(_1312_),
    .Y(_1378_));
 sg13g2_nor2b_1 _2252_ (.A(_1335_),
    .B_N(_1378_),
    .Y(_1379_));
 sg13g2_xnor2_1 _2253_ (.Y(_1380_),
    .A(_1335_),
    .B(_1378_));
 sg13g2_nor2_1 _2254_ (.A(net321),
    .B(_1380_),
    .Y(_1381_));
 sg13g2_a21oi_1 _2255_ (.A1(_1203_),
    .A2(_1312_),
    .Y(_1382_),
    .B1(_1378_));
 sg13g2_xnor2_1 _2256_ (.Y(_1383_),
    .A(net324),
    .B(_1312_));
 sg13g2_o21ai_1 _2257_ (.B1(_1330_),
    .Y(_1384_),
    .A1(_1329_),
    .A2(_1383_));
 sg13g2_xnor2_1 _2258_ (.Y(_1385_),
    .A(_0024_),
    .B(_1382_));
 sg13g2_a22oi_1 _2259_ (.Y(_1386_),
    .B1(_1384_),
    .B2(_1385_),
    .A2(_1382_),
    .A1(net323));
 sg13g2_nor2_1 _2260_ (.A(_1381_),
    .B(_1386_),
    .Y(_1387_));
 sg13g2_nor2_1 _2261_ (.A(_1308_),
    .B(_1379_),
    .Y(_1388_));
 sg13g2_nand2_1 _2262_ (.Y(_1389_),
    .A(_1308_),
    .B(_1379_));
 sg13g2_nor2_1 _2263_ (.A(_0023_),
    .B(_1388_),
    .Y(_1390_));
 sg13g2_a221oi_1 _2264_ (.B2(_1390_),
    .C1(_1387_),
    .B1(_1389_),
    .A1(net321),
    .Y(_1391_),
    .A2(_1380_));
 sg13g2_a21oi_1 _2265_ (.A1(_1204_),
    .A2(\h[8] ),
    .Y(_1392_),
    .B1(_1373_));
 sg13g2_inv_1 _2266_ (.Y(_1393_),
    .A(_1392_));
 sg13g2_nor2b_1 _2267_ (.A(net342),
    .B_N(net308),
    .Y(_1394_));
 sg13g2_nor2_1 _2268_ (.A(net309),
    .B(_1394_),
    .Y(_1395_));
 sg13g2_o21ai_1 _2269_ (.B1(_1363_),
    .Y(_1396_),
    .A1(_1206_),
    .A2(net312));
 sg13g2_a221oi_1 _2270_ (.B2(_1206_),
    .C1(_1394_),
    .B1(net312),
    .A1(_1205_),
    .Y(_1397_),
    .A2(net309));
 sg13g2_nand2b_1 _2271_ (.Y(_1398_),
    .B(\px[8] ),
    .A_N(\h[8] ));
 sg13g2_nand2b_1 _2272_ (.Y(_1399_),
    .B(net342),
    .A_N(net308));
 sg13g2_nand3_1 _2273_ (.B(_1398_),
    .C(_1399_),
    .A(_1392_),
    .Y(_1400_));
 sg13g2_a221oi_1 _2274_ (.B2(_1397_),
    .C1(_1400_),
    .B1(_1396_),
    .A1(net343),
    .Y(_1401_),
    .A2(_1395_));
 sg13g2_nor2_1 _2275_ (.A(net318),
    .B(\py[9] ),
    .Y(_1402_));
 sg13g2_nand3_1 _2276_ (.B(_1374_),
    .C(_1402_),
    .A(_0052_),
    .Y(_1403_));
 sg13g2_a21oi_1 _2277_ (.A1(_1373_),
    .A2(_1375_),
    .Y(_1404_),
    .B1(_1403_));
 sg13g2_nand3_1 _2278_ (.B(_1389_),
    .C(_1404_),
    .A(_1306_),
    .Y(_1405_));
 sg13g2_a21oi_1 _2279_ (.A1(_0023_),
    .A2(_1388_),
    .Y(_1406_),
    .B1(_1405_));
 sg13g2_o21ai_1 _2280_ (.B1(_1406_),
    .Y(_1407_),
    .A1(_1393_),
    .A2(_1401_));
 sg13g2_nor4_2 _2281_ (.A(_1339_),
    .B(_1377_),
    .C(_1391_),
    .Y(_1408_),
    .D(_1407_));
 sg13g2_xnor2_1 _2282_ (.Y(_1409_),
    .A(\px[0] ),
    .B(\h[0] ));
 sg13g2_xor2_1 _2283_ (.B(\h[0] ),
    .A(\px[0] ),
    .X(_1410_));
 sg13g2_xnor2_1 _2284_ (.Y(_1411_),
    .A(_1351_),
    .B(_1355_));
 sg13g2_inv_2 _2285_ (.Y(_1412_),
    .A(_1411_));
 sg13g2_nor2_1 _2286_ (.A(_1354_),
    .B(_1356_),
    .Y(_1413_));
 sg13g2_xnor2_1 _2287_ (.Y(_1414_),
    .A(_1360_),
    .B(_1413_));
 sg13g2_inv_1 _2288_ (.Y(_1415_),
    .A(_1414_));
 sg13g2_and2_1 _2289_ (.A(_1411_),
    .B(_1414_),
    .X(_1416_));
 sg13g2_nand2_1 _2290_ (.Y(_1417_),
    .A(_1411_),
    .B(_1414_));
 sg13g2_xnor2_1 _2291_ (.Y(_1418_),
    .A(_1412_),
    .B(_1414_));
 sg13g2_nand2_1 _2292_ (.Y(_1419_),
    .A(net304),
    .B(_1418_));
 sg13g2_xor2_1 _2293_ (.B(net341),
    .A(net332),
    .X(_1420_));
 sg13g2_xnor2_1 _2294_ (.Y(_1421_),
    .A(net332),
    .B(net341));
 sg13g2_nand2_1 _2295_ (.Y(_1422_),
    .A(net330),
    .B(\py[2] ));
 sg13g2_xnor2_1 _2296_ (.Y(_1423_),
    .A(net330),
    .B(\py[2] ));
 sg13g2_nor3_1 _2297_ (.A(_1316_),
    .B(_1318_),
    .C(_1423_),
    .Y(_1424_));
 sg13g2_nand2_1 _2298_ (.Y(_1425_),
    .A(net327),
    .B(\py[3] ));
 sg13g2_xnor2_1 _2299_ (.Y(_1426_),
    .A(net327),
    .B(\py[3] ));
 sg13g2_nor2_1 _2300_ (.A(_1422_),
    .B(_1426_),
    .Y(_1427_));
 sg13g2_xor2_1 _2301_ (.B(_1426_),
    .A(_1422_),
    .X(_1428_));
 sg13g2_xnor2_1 _2302_ (.Y(_1429_),
    .A(_1424_),
    .B(_1428_));
 sg13g2_nor2_1 _2303_ (.A(_1421_),
    .B(_1429_),
    .Y(_1430_));
 sg13g2_nand3_1 _2304_ (.B(_1414_),
    .C(_1430_),
    .A(net304),
    .Y(_1431_));
 sg13g2_a21o_1 _2305_ (.A2(_1414_),
    .A1(net304),
    .B1(_1430_),
    .X(_1432_));
 sg13g2_and2_1 _2306_ (.A(_1431_),
    .B(_1432_),
    .X(_1433_));
 sg13g2_nand2b_1 _2307_ (.Y(_1434_),
    .B(_1433_),
    .A_N(_1419_));
 sg13g2_o21ai_1 _2308_ (.B1(_1434_),
    .Y(_1435_),
    .A1(_1409_),
    .A2(_1417_));
 sg13g2_xor2_1 _2309_ (.B(net313),
    .A(\px[4] ),
    .X(_1436_));
 sg13g2_xnor2_1 _2310_ (.Y(_1437_),
    .A(_1357_),
    .B(_1436_));
 sg13g2_xnor2_1 _2311_ (.Y(_1438_),
    .A(_1361_),
    .B(_1437_));
 sg13g2_nor2_1 _2312_ (.A(net304),
    .B(net300),
    .Y(_1439_));
 sg13g2_xnor2_1 _2313_ (.Y(_1440_),
    .A(_1346_),
    .B(_1349_));
 sg13g2_nand2_1 _2314_ (.Y(_1441_),
    .A(_1355_),
    .B(_1440_));
 sg13g2_a21oi_1 _2315_ (.A1(_1424_),
    .A2(_1428_),
    .Y(_1442_),
    .B1(_1427_));
 sg13g2_xor2_1 _2316_ (.B(net339),
    .A(net326),
    .X(_1443_));
 sg13g2_xnor2_1 _2317_ (.Y(_1444_),
    .A(_1425_),
    .B(_1443_));
 sg13g2_xor2_1 _2318_ (.B(_1444_),
    .A(_1442_),
    .X(_1445_));
 sg13g2_inv_1 _2319_ (.Y(_1446_),
    .A(net298));
 sg13g2_xor2_1 _2320_ (.B(net298),
    .A(_1441_),
    .X(_1447_));
 sg13g2_xnor2_1 _2321_ (.Y(_1448_),
    .A(_1439_),
    .B(_1447_));
 sg13g2_xnor2_1 _2322_ (.Y(_1449_),
    .A(_1412_),
    .B(_1448_));
 sg13g2_nand2_1 _2323_ (.Y(_1450_),
    .A(_1435_),
    .B(_1449_));
 sg13g2_xnor2_1 _2324_ (.Y(_1451_),
    .A(_1435_),
    .B(_1449_));
 sg13g2_xor2_1 _2325_ (.B(net340),
    .A(net331),
    .X(_1452_));
 sg13g2_xor2_1 _2326_ (.B(_1452_),
    .A(_1317_),
    .X(_1453_));
 sg13g2_xnor2_1 _2327_ (.Y(_1454_),
    .A(_1317_),
    .B(_1452_));
 sg13g2_xnor2_1 _2328_ (.Y(_1455_),
    .A(_1319_),
    .B(_1423_));
 sg13g2_nand2_1 _2329_ (.Y(_1456_),
    .A(_1454_),
    .B(net302));
 sg13g2_nor2_2 _2330_ (.A(_1429_),
    .B(_1453_),
    .Y(_1457_));
 sg13g2_nor2_2 _2331_ (.A(_1421_),
    .B(_1446_),
    .Y(_1458_));
 sg13g2_nand2_2 _2332_ (.Y(_1459_),
    .A(_1420_),
    .B(_1445_));
 sg13g2_nor2_2 _2333_ (.A(net299),
    .B(_1459_),
    .Y(_1460_));
 sg13g2_xnor2_1 _2334_ (.Y(_1461_),
    .A(_1439_),
    .B(_1459_));
 sg13g2_xnor2_1 _2335_ (.Y(_1462_),
    .A(_1457_),
    .B(_1461_));
 sg13g2_or2_1 _2336_ (.X(_1463_),
    .B(_1462_),
    .A(_1431_));
 sg13g2_xnor2_1 _2337_ (.Y(_1464_),
    .A(_1431_),
    .B(_1462_));
 sg13g2_xnor2_1 _2338_ (.Y(_1465_),
    .A(_1456_),
    .B(_1464_));
 sg13g2_o21ai_1 _2339_ (.B1(_1450_),
    .Y(_1466_),
    .A1(_1451_),
    .A2(_1465_));
 sg13g2_a22oi_1 _2340_ (.Y(_1467_),
    .B1(_1448_),
    .B2(_1411_),
    .A2(_1440_),
    .A1(_1355_));
 sg13g2_nand2_2 _2341_ (.Y(_1468_),
    .A(net304),
    .B(_1440_));
 sg13g2_o21ai_1 _2342_ (.B1(_1468_),
    .Y(_1469_),
    .A1(_1350_),
    .A2(net304));
 sg13g2_nor2_2 _2343_ (.A(_1415_),
    .B(net299),
    .Y(_1470_));
 sg13g2_nor2_1 _2344_ (.A(net299),
    .B(_1469_),
    .Y(_1471_));
 sg13g2_xnor2_1 _2345_ (.Y(_1472_),
    .A(_1416_),
    .B(_1471_));
 sg13g2_a21o_1 _2346_ (.A2(_1446_),
    .A1(_1409_),
    .B1(net300),
    .X(_1473_));
 sg13g2_nor2_1 _2347_ (.A(_1472_),
    .B(_1473_),
    .Y(_1474_));
 sg13g2_nand2_1 _2348_ (.Y(_1475_),
    .A(_1472_),
    .B(_1473_));
 sg13g2_xnor2_1 _2349_ (.Y(_1476_),
    .A(_1472_),
    .B(_1473_));
 sg13g2_nor2_1 _2350_ (.A(net300),
    .B(_1440_),
    .Y(_1477_));
 sg13g2_and2_1 _2351_ (.A(_1416_),
    .B(_1477_),
    .X(_1478_));
 sg13g2_xnor2_1 _2352_ (.Y(_1479_),
    .A(_1417_),
    .B(_1477_));
 sg13g2_xnor2_1 _2353_ (.Y(_1480_),
    .A(_1459_),
    .B(_1479_));
 sg13g2_xnor2_1 _2354_ (.Y(_1481_),
    .A(_1476_),
    .B(_1480_));
 sg13g2_nor2b_1 _2355_ (.A(_1467_),
    .B_N(_1481_),
    .Y(_1482_));
 sg13g2_xnor2_1 _2356_ (.Y(_1483_),
    .A(_1467_),
    .B(_1481_));
 sg13g2_a22oi_1 _2357_ (.Y(_1484_),
    .B1(_1461_),
    .B2(_1457_),
    .A2(_1460_),
    .A1(_1409_));
 sg13g2_nand2_1 _2358_ (.Y(_1485_),
    .A(net298),
    .B(_1454_));
 sg13g2_inv_1 _2359_ (.Y(_1486_),
    .A(_1485_));
 sg13g2_nand2_1 _2360_ (.Y(_1487_),
    .A(_1414_),
    .B(_1440_));
 sg13g2_or2_1 _2361_ (.X(_1488_),
    .B(_1487_),
    .A(_1485_));
 sg13g2_xor2_1 _2362_ (.B(_1487_),
    .A(_1485_),
    .X(_1489_));
 sg13g2_nand2b_1 _2363_ (.Y(_1490_),
    .B(_1489_),
    .A_N(_1484_));
 sg13g2_xnor2_1 _2364_ (.Y(_1491_),
    .A(_1484_),
    .B(_1489_));
 sg13g2_xor2_1 _2365_ (.B(_1491_),
    .A(_1483_),
    .X(_1492_));
 sg13g2_and2_1 _2366_ (.A(_1466_),
    .B(_1492_),
    .X(_1493_));
 sg13g2_or2_1 _2367_ (.X(_1494_),
    .B(_1492_),
    .A(_1466_));
 sg13g2_xnor2_1 _2368_ (.Y(_1495_),
    .A(_1466_),
    .B(_1492_));
 sg13g2_xor2_1 _2369_ (.B(_1457_),
    .A(net302),
    .X(_1496_));
 sg13g2_nand3_1 _2370_ (.B(_1445_),
    .C(_1496_),
    .A(_1421_),
    .Y(_1497_));
 sg13g2_o21ai_1 _2371_ (.B1(_1497_),
    .Y(_1498_),
    .A1(_1429_),
    .A2(_1456_));
 sg13g2_o21ai_1 _2372_ (.B1(_1463_),
    .Y(_1499_),
    .A1(_1456_),
    .A2(_1464_));
 sg13g2_nand2_1 _2373_ (.Y(_1500_),
    .A(net298),
    .B(_1453_));
 sg13g2_nor3_1 _2374_ (.A(_1446_),
    .B(_1454_),
    .C(_1463_),
    .Y(_1501_));
 sg13g2_xor2_1 _2375_ (.B(_1500_),
    .A(_1499_),
    .X(_1502_));
 sg13g2_inv_1 _2376_ (.Y(_1503_),
    .A(_1502_));
 sg13g2_xnor2_1 _2377_ (.Y(_1504_),
    .A(_1498_),
    .B(_1502_));
 sg13g2_a21oi_1 _2378_ (.A1(_1494_),
    .A2(_1504_),
    .Y(_1505_),
    .B1(_1493_));
 sg13g2_or2_1 _2379_ (.X(_1506_),
    .B(net302),
    .A(_1446_));
 sg13g2_a21oi_2 _2380_ (.B1(_1506_),
    .Y(_1507_),
    .A2(_1490_),
    .A1(_1488_));
 sg13g2_nand3_1 _2381_ (.B(_1490_),
    .C(_1506_),
    .A(_1488_),
    .Y(_1508_));
 sg13g2_nor2b_1 _2382_ (.A(_1507_),
    .B_N(_1508_),
    .Y(_1509_));
 sg13g2_a21oi_1 _2383_ (.A1(_1483_),
    .A2(_1491_),
    .Y(_1510_),
    .B1(_1482_));
 sg13g2_a21oi_1 _2384_ (.A1(_1475_),
    .A2(_1480_),
    .Y(_1511_),
    .B1(_1474_));
 sg13g2_nor2_1 _2385_ (.A(net299),
    .B(_1468_),
    .Y(_1512_));
 sg13g2_nor3_2 _2386_ (.A(_1412_),
    .B(net299),
    .C(_1468_),
    .Y(_1513_));
 sg13g2_a21oi_1 _2387_ (.A1(_1412_),
    .A2(_1469_),
    .Y(_1514_),
    .B1(net299));
 sg13g2_o21ai_1 _2388_ (.B1(_1514_),
    .Y(_1515_),
    .A1(_1412_),
    .A2(_1469_));
 sg13g2_a21oi_1 _2389_ (.A1(_1416_),
    .A2(_1471_),
    .Y(_1516_),
    .B1(_1512_));
 sg13g2_a21oi_1 _2390_ (.A1(_1515_),
    .A2(_1516_),
    .Y(_1517_),
    .B1(_1513_));
 sg13g2_nand2_1 _2391_ (.Y(_1518_),
    .A(_1414_),
    .B(net300));
 sg13g2_o21ai_1 _2392_ (.B1(_1518_),
    .Y(_1519_),
    .A1(_1418_),
    .A2(net299));
 sg13g2_xnor2_1 _2393_ (.Y(_1520_),
    .A(_1459_),
    .B(_1519_));
 sg13g2_xor2_1 _2394_ (.B(_1520_),
    .A(_1517_),
    .X(_1521_));
 sg13g2_nor2b_1 _2395_ (.A(_1511_),
    .B_N(_1521_),
    .Y(_1522_));
 sg13g2_xnor2_1 _2396_ (.Y(_1523_),
    .A(_1511_),
    .B(_1521_));
 sg13g2_nand2_2 _2397_ (.Y(_1524_),
    .A(_1428_),
    .B(_1455_));
 sg13g2_a21o_1 _2398_ (.A2(_1479_),
    .A1(_1458_),
    .B1(_1478_),
    .X(_1525_));
 sg13g2_xnor2_1 _2399_ (.Y(_1526_),
    .A(_1454_),
    .B(net302));
 sg13g2_nand2b_1 _2400_ (.Y(_1527_),
    .B(net298),
    .A_N(_1526_));
 sg13g2_nor2_1 _2401_ (.A(_1429_),
    .B(_1527_),
    .Y(_1528_));
 sg13g2_and2_1 _2402_ (.A(_1429_),
    .B(_1527_),
    .X(_1529_));
 sg13g2_nor2_1 _2403_ (.A(_1528_),
    .B(_1529_),
    .Y(_1530_));
 sg13g2_nand2_1 _2404_ (.Y(_1531_),
    .A(_1525_),
    .B(_1530_));
 sg13g2_xnor2_1 _2405_ (.Y(_1532_),
    .A(_1525_),
    .B(_1530_));
 sg13g2_xor2_1 _2406_ (.B(_1532_),
    .A(_1524_),
    .X(_1533_));
 sg13g2_xnor2_1 _2407_ (.Y(_1534_),
    .A(_1523_),
    .B(_1533_));
 sg13g2_nor2_1 _2408_ (.A(_1510_),
    .B(_1534_),
    .Y(_1535_));
 sg13g2_xor2_1 _2409_ (.B(_1534_),
    .A(_1510_),
    .X(_1536_));
 sg13g2_xnor2_1 _2410_ (.Y(_1537_),
    .A(_1509_),
    .B(_1536_));
 sg13g2_or2_1 _2411_ (.X(_1538_),
    .B(_1537_),
    .A(_1505_));
 sg13g2_a21oi_1 _2412_ (.A1(_1498_),
    .A2(_1503_),
    .Y(_1539_),
    .B1(_1501_));
 sg13g2_and2_1 _2413_ (.A(_1505_),
    .B(_1537_),
    .X(_1540_));
 sg13g2_xor2_1 _2414_ (.B(_1537_),
    .A(_1505_),
    .X(_1541_));
 sg13g2_o21ai_1 _2415_ (.B1(_1538_),
    .Y(_1542_),
    .A1(_1539_),
    .A2(_1540_));
 sg13g2_a21oi_1 _2416_ (.A1(_1509_),
    .A2(_1536_),
    .Y(_1543_),
    .B1(_1535_));
 sg13g2_o21ai_1 _2417_ (.B1(_1531_),
    .Y(_1544_),
    .A1(_1524_),
    .A2(_1532_));
 sg13g2_nand2_1 _2418_ (.Y(_1545_),
    .A(_1429_),
    .B(net298));
 sg13g2_nand2b_1 _2419_ (.Y(_1546_),
    .B(_1544_),
    .A_N(_1545_));
 sg13g2_xor2_1 _2420_ (.B(_1545_),
    .A(_1544_),
    .X(_1547_));
 sg13g2_a21oi_1 _2421_ (.A1(_1523_),
    .A2(_1533_),
    .Y(_1548_),
    .B1(_1522_));
 sg13g2_a21oi_1 _2422_ (.A1(_1517_),
    .A2(_1520_),
    .Y(_1549_),
    .B1(_1513_));
 sg13g2_xor2_1 _2423_ (.B(_1459_),
    .A(net299),
    .X(_1550_));
 sg13g2_mux2_2 _2424_ (.A0(_1514_),
    .A1(_1412_),
    .S(_1512_),
    .X(_1551_));
 sg13g2_xor2_1 _2425_ (.B(_1551_),
    .A(_1550_),
    .X(_1552_));
 sg13g2_nand2b_1 _2426_ (.Y(_1553_),
    .B(_1552_),
    .A_N(_1549_));
 sg13g2_xor2_1 _2427_ (.B(_1552_),
    .A(_1549_),
    .X(_1554_));
 sg13g2_a21oi_2 _2428_ (.B1(_1528_),
    .Y(_1555_),
    .A2(_1486_),
    .A1(net302));
 sg13g2_a21oi_1 _2429_ (.A1(net298),
    .A2(_1526_),
    .Y(_1556_),
    .B1(_1429_));
 sg13g2_nor2_2 _2430_ (.A(_1529_),
    .B(_1556_),
    .Y(_1557_));
 sg13g2_a22oi_1 _2431_ (.Y(_1558_),
    .B1(_1519_),
    .B2(_1458_),
    .A2(_1470_),
    .A1(_1412_));
 sg13g2_nand2b_1 _2432_ (.Y(_1559_),
    .B(_1557_),
    .A_N(_1558_));
 sg13g2_xnor2_1 _2433_ (.Y(_1560_),
    .A(_1557_),
    .B(_1558_));
 sg13g2_nand2b_1 _2434_ (.Y(_1561_),
    .B(_1560_),
    .A_N(_1555_));
 sg13g2_xnor2_1 _2435_ (.Y(_1562_),
    .A(_1555_),
    .B(_1560_));
 sg13g2_nand2b_1 _2436_ (.Y(_1563_),
    .B(_1562_),
    .A_N(_1554_));
 sg13g2_xnor2_1 _2437_ (.Y(_1564_),
    .A(_1554_),
    .B(_1562_));
 sg13g2_nand2b_1 _2438_ (.Y(_1565_),
    .B(_1564_),
    .A_N(_1548_));
 sg13g2_xnor2_1 _2439_ (.Y(_1566_),
    .A(_1548_),
    .B(_1564_));
 sg13g2_nand2b_1 _2440_ (.Y(_1567_),
    .B(_1566_),
    .A_N(_1547_));
 sg13g2_xnor2_1 _2441_ (.Y(_1568_),
    .A(_1547_),
    .B(_1566_));
 sg13g2_nor2b_1 _2442_ (.A(_1543_),
    .B_N(_1568_),
    .Y(_1569_));
 sg13g2_xnor2_1 _2443_ (.Y(_1570_),
    .A(_1543_),
    .B(_1568_));
 sg13g2_xor2_1 _2444_ (.B(_1570_),
    .A(_1507_),
    .X(_1571_));
 sg13g2_nor2_1 _2445_ (.A(_1542_),
    .B(_1571_),
    .Y(_1572_));
 sg13g2_nand2_1 _2446_ (.Y(_1573_),
    .A(_1542_),
    .B(_1571_));
 sg13g2_xor2_1 _2447_ (.B(_1571_),
    .A(_1542_),
    .X(_1574_));
 sg13g2_nand2_1 _2448_ (.Y(_1575_),
    .A(_1420_),
    .B(_1455_));
 sg13g2_nor2_2 _2449_ (.A(_1349_),
    .B(net304),
    .Y(_1576_));
 sg13g2_nand3_1 _2450_ (.B(net302),
    .C(_1576_),
    .A(_1420_),
    .Y(_1577_));
 sg13g2_nand2_1 _2451_ (.Y(_1578_),
    .A(_1468_),
    .B(_1577_));
 sg13g2_xnor2_1 _2452_ (.Y(_1579_),
    .A(_1419_),
    .B(_1433_));
 sg13g2_and2_1 _2453_ (.A(_1420_),
    .B(_1452_),
    .X(_1580_));
 sg13g2_nand2_1 _2454_ (.Y(_1581_),
    .A(net302),
    .B(_1580_));
 sg13g2_nor2_1 _2455_ (.A(_1429_),
    .B(_1581_),
    .Y(_1582_));
 sg13g2_nor2b_1 _2456_ (.A(_1430_),
    .B_N(_1581_),
    .Y(_1583_));
 sg13g2_nor2_1 _2457_ (.A(_1582_),
    .B(_1583_),
    .Y(_1584_));
 sg13g2_xnor2_1 _2458_ (.Y(_1585_),
    .A(_1578_),
    .B(_1579_));
 sg13g2_nor3_1 _2459_ (.A(_1582_),
    .B(_1583_),
    .C(_1585_),
    .Y(_1586_));
 sg13g2_a21o_1 _2460_ (.A2(_1579_),
    .A1(_1578_),
    .B1(_1586_),
    .X(_1587_));
 sg13g2_xor2_1 _2461_ (.B(_1465_),
    .A(_1451_),
    .X(_1588_));
 sg13g2_nand2_1 _2462_ (.Y(_1589_),
    .A(_1587_),
    .B(_1588_));
 sg13g2_a21o_1 _2463_ (.A2(net298),
    .A1(_1421_),
    .B1(_1496_),
    .X(_1590_));
 sg13g2_a21oi_1 _2464_ (.A1(_1497_),
    .A2(_1590_),
    .Y(_1591_),
    .B1(_1582_));
 sg13g2_xnor2_1 _2465_ (.Y(_1592_),
    .A(_1587_),
    .B(_1588_));
 sg13g2_o21ai_1 _2466_ (.B1(_1589_),
    .Y(_1593_),
    .A1(_1591_),
    .A2(_1592_));
 sg13g2_xnor2_1 _2467_ (.Y(_1594_),
    .A(_1495_),
    .B(_1504_));
 sg13g2_nand2_1 _2468_ (.Y(_1595_),
    .A(_1593_),
    .B(_1594_));
 sg13g2_xnor2_1 _2469_ (.Y(_1596_),
    .A(_1539_),
    .B(_1541_));
 sg13g2_nand2b_1 _2470_ (.Y(_1597_),
    .B(_1596_),
    .A_N(_1595_));
 sg13g2_xnor2_1 _2471_ (.Y(_1598_),
    .A(_1595_),
    .B(_1596_));
 sg13g2_xor2_1 _2472_ (.B(_1596_),
    .A(_1595_),
    .X(_1599_));
 sg13g2_xor2_1 _2473_ (.B(_1592_),
    .A(_1591_),
    .X(_1600_));
 sg13g2_xnor2_1 _2474_ (.Y(_1601_),
    .A(_1584_),
    .B(_1585_));
 sg13g2_a22oi_1 _2475_ (.Y(_1602_),
    .B1(_1580_),
    .B2(net302),
    .A2(_1575_),
    .A1(_1453_));
 sg13g2_xnor2_1 _2476_ (.Y(_1603_),
    .A(_1575_),
    .B(_1576_));
 sg13g2_nand2_1 _2477_ (.Y(_1604_),
    .A(_1602_),
    .B(_1603_));
 sg13g2_and3_1 _2478_ (.X(_1605_),
    .A(_1601_),
    .B(_1602_),
    .C(_1603_));
 sg13g2_nand2_1 _2479_ (.Y(_1606_),
    .A(_1600_),
    .B(_1605_));
 sg13g2_xor2_1 _2480_ (.B(_1594_),
    .A(_1593_),
    .X(_1607_));
 sg13g2_nor2b_1 _2481_ (.A(_1606_),
    .B_N(_1607_),
    .Y(_1608_));
 sg13g2_xnor2_1 _2482_ (.Y(_1609_),
    .A(_1601_),
    .B(_1604_));
 sg13g2_xor2_1 _2483_ (.B(_1603_),
    .A(_1602_),
    .X(_1610_));
 sg13g2_and2_1 _2484_ (.A(_1580_),
    .B(_1610_),
    .X(_1611_));
 sg13g2_and2_1 _2485_ (.A(_1609_),
    .B(_1611_),
    .X(_1612_));
 sg13g2_and2_1 _2486_ (.A(_1600_),
    .B(_1612_),
    .X(_1613_));
 sg13g2_xnor2_1 _2487_ (.Y(_1614_),
    .A(_1606_),
    .B(_1607_));
 sg13g2_a21oi_2 _2488_ (.B1(_1608_),
    .Y(_1615_),
    .A2(_1614_),
    .A1(_1613_));
 sg13g2_o21ai_1 _2489_ (.B1(_1597_),
    .Y(_1616_),
    .A1(_1599_),
    .A2(_1615_));
 sg13g2_xnor2_1 _2490_ (.Y(_1617_),
    .A(_1574_),
    .B(_1616_));
 sg13g2_xor2_1 _2491_ (.B(_1616_),
    .A(_1574_),
    .X(_1618_));
 sg13g2_xnor2_1 _2492_ (.Y(_1619_),
    .A(_1598_),
    .B(_1615_));
 sg13g2_nor2b_1 _2493_ (.A(_1619_),
    .B_N(\product_comp[6] ),
    .Y(_1620_));
 sg13g2_nand2b_1 _2494_ (.Y(_1621_),
    .B(_1619_),
    .A_N(\product_comp[6] ));
 sg13g2_xor2_1 _2495_ (.B(_1614_),
    .A(_1613_),
    .X(_1622_));
 sg13g2_nand2b_1 _2496_ (.Y(_1623_),
    .B(\product_comp[5] ),
    .A_N(_1622_));
 sg13g2_nor2b_1 _2497_ (.A(\product_comp[5] ),
    .B_N(_1622_),
    .Y(_1624_));
 sg13g2_nor2_1 _2498_ (.A(_1605_),
    .B(_1612_),
    .Y(_1625_));
 sg13g2_xor2_1 _2499_ (.B(_1625_),
    .A(_1600_),
    .X(_1626_));
 sg13g2_nor2_1 _2500_ (.A(_1410_),
    .B(_1420_),
    .Y(_1627_));
 sg13g2_inv_1 _2501_ (.Y(_1628_),
    .A(_1627_));
 sg13g2_xnor2_1 _2502_ (.Y(_1629_),
    .A(net304),
    .B(_1420_));
 sg13g2_o21ai_1 _2503_ (.B1(\product_comp[2] ),
    .Y(_1630_),
    .A1(\product_comp[1] ),
    .A2(_1629_));
 sg13g2_nor2b_1 _2504_ (.A(_1611_),
    .B_N(_1630_),
    .Y(_1631_));
 sg13g2_o21ai_1 _2505_ (.B1(_1631_),
    .Y(_1632_),
    .A1(_1580_),
    .A2(_1610_));
 sg13g2_or3_1 _2506_ (.A(\product_comp[2] ),
    .B(\product_comp[1] ),
    .C(_1627_),
    .X(_1633_));
 sg13g2_xor2_1 _2507_ (.B(_1611_),
    .A(_1609_),
    .X(_1634_));
 sg13g2_nor2_1 _2508_ (.A(_0030_),
    .B(_1634_),
    .Y(_1635_));
 sg13g2_a21oi_1 _2509_ (.A1(_1632_),
    .A2(_1633_),
    .Y(_1636_),
    .B1(_1635_));
 sg13g2_a21oi_1 _2510_ (.A1(_0030_),
    .A2(_1634_),
    .Y(_1637_),
    .B1(_1636_));
 sg13g2_a21o_1 _2511_ (.A2(_1637_),
    .A1(_1626_),
    .B1(\product_comp[4] ),
    .X(_1638_));
 sg13g2_o21ai_1 _2512_ (.B1(_1638_),
    .Y(_1639_),
    .A1(_1626_),
    .A2(_1637_));
 sg13g2_a21oi_1 _2513_ (.A1(_1623_),
    .A2(_1639_),
    .Y(_1640_),
    .B1(_1624_));
 sg13g2_a221oi_1 _2514_ (.B2(_1640_),
    .C1(_1620_),
    .B1(_1621_),
    .A1(_1225_),
    .Y(_1641_),
    .A2(_1617_));
 sg13g2_a21oi_1 _2515_ (.A1(_1507_),
    .A2(_1570_),
    .Y(_1642_),
    .B1(_1569_));
 sg13g2_nand2_1 _2516_ (.Y(_1643_),
    .A(_1565_),
    .B(_1567_));
 sg13g2_nand2_1 _2517_ (.Y(_1644_),
    .A(_1559_),
    .B(_1561_));
 sg13g2_nand2_1 _2518_ (.Y(_1645_),
    .A(_1553_),
    .B(_1563_));
 sg13g2_xor2_1 _2519_ (.B(_1557_),
    .A(_1460_),
    .X(_1646_));
 sg13g2_nor2b_1 _2520_ (.A(_1555_),
    .B_N(_1646_),
    .Y(_1647_));
 sg13g2_xnor2_1 _2521_ (.Y(_1648_),
    .A(_1555_),
    .B(_1646_));
 sg13g2_a21oi_1 _2522_ (.A1(_1550_),
    .A2(_1551_),
    .Y(_1649_),
    .B1(_1513_));
 sg13g2_nand2_1 _2523_ (.Y(_1650_),
    .A(_1458_),
    .B(_1470_));
 sg13g2_xnor2_1 _2524_ (.Y(_1651_),
    .A(_1459_),
    .B(_1470_));
 sg13g2_xnor2_1 _2525_ (.Y(_1652_),
    .A(_1551_),
    .B(_1651_));
 sg13g2_nor2_1 _2526_ (.A(_1649_),
    .B(_1652_),
    .Y(_1653_));
 sg13g2_xor2_1 _2527_ (.B(_1652_),
    .A(_1649_),
    .X(_1654_));
 sg13g2_xnor2_1 _2528_ (.Y(_1655_),
    .A(_1648_),
    .B(_1654_));
 sg13g2_inv_1 _2529_ (.Y(_1656_),
    .A(_1655_));
 sg13g2_xnor2_1 _2530_ (.Y(_1657_),
    .A(_1645_),
    .B(_1656_));
 sg13g2_nor2b_1 _2531_ (.A(_1657_),
    .B_N(_1644_),
    .Y(_1658_));
 sg13g2_xor2_1 _2532_ (.B(_1657_),
    .A(_1644_),
    .X(_1659_));
 sg13g2_nand2b_1 _2533_ (.Y(_1660_),
    .B(_1643_),
    .A_N(_1659_));
 sg13g2_xor2_1 _2534_ (.B(_1659_),
    .A(_1643_),
    .X(_1661_));
 sg13g2_xor2_1 _2535_ (.B(_1661_),
    .A(_1546_),
    .X(_1662_));
 sg13g2_nor2b_1 _2536_ (.A(_1642_),
    .B_N(_1662_),
    .Y(_1663_));
 sg13g2_xor2_1 _2537_ (.B(_1662_),
    .A(_1642_),
    .X(_1664_));
 sg13g2_nand3b_1 _2538_ (.B(_1598_),
    .C(_1574_),
    .Y(_1665_),
    .A_N(_1615_));
 sg13g2_a21o_1 _2539_ (.A2(_1597_),
    .A1(_1573_),
    .B1(_1572_),
    .X(_1666_));
 sg13g2_nand2_1 _2540_ (.Y(_1667_),
    .A(_1665_),
    .B(_1666_));
 sg13g2_a21oi_1 _2541_ (.A1(_1665_),
    .A2(_1666_),
    .Y(_1668_),
    .B1(_1664_));
 sg13g2_xnor2_1 _2542_ (.Y(_1669_),
    .A(_1664_),
    .B(_1667_));
 sg13g2_xor2_1 _2543_ (.B(_1667_),
    .A(_1664_),
    .X(_1670_));
 sg13g2_a221oi_1 _2544_ (.B2(_1178_),
    .C1(_1641_),
    .B1(_1669_),
    .A1(_0029_),
    .Y(_1671_),
    .A2(_1618_));
 sg13g2_a21oi_1 _2545_ (.A1(_1645_),
    .A2(_1656_),
    .Y(_1672_),
    .B1(_1658_));
 sg13g2_a21oi_1 _2546_ (.A1(_1648_),
    .A2(_1654_),
    .Y(_1673_),
    .B1(_1653_));
 sg13g2_a21oi_1 _2547_ (.A1(_1460_),
    .A2(_1557_),
    .Y(_1674_),
    .B1(_1647_));
 sg13g2_xnor2_1 _2548_ (.Y(_1675_),
    .A(_1557_),
    .B(_1650_));
 sg13g2_xnor2_1 _2549_ (.Y(_1676_),
    .A(_1555_),
    .B(_1675_));
 sg13g2_nor3_1 _2550_ (.A(_1513_),
    .B(_1551_),
    .C(_1651_),
    .Y(_1677_));
 sg13g2_a21oi_1 _2551_ (.A1(_1513_),
    .A2(_1651_),
    .Y(_1678_),
    .B1(_1677_));
 sg13g2_xnor2_1 _2552_ (.Y(_1679_),
    .A(_1676_),
    .B(_1678_));
 sg13g2_xnor2_1 _2553_ (.Y(_1680_),
    .A(_1673_),
    .B(_1679_));
 sg13g2_xnor2_1 _2554_ (.Y(_1681_),
    .A(_1674_),
    .B(_1680_));
 sg13g2_xnor2_1 _2555_ (.Y(_1682_),
    .A(_1672_),
    .B(_1681_));
 sg13g2_o21ai_1 _2556_ (.B1(_1660_),
    .Y(_1683_),
    .A1(_1546_),
    .A2(_1661_));
 sg13g2_or2_1 _2557_ (.X(_1684_),
    .B(_1683_),
    .A(_1682_));
 sg13g2_o21ai_1 _2558_ (.B1(_1684_),
    .Y(_1685_),
    .A1(_1663_),
    .A2(_1668_));
 sg13g2_and2_1 _2559_ (.A(_1224_),
    .B(_1685_),
    .X(_1686_));
 sg13g2_nor2_1 _2560_ (.A(_1178_),
    .B(_1669_),
    .Y(_1687_));
 sg13g2_nor3_1 _2561_ (.A(_1671_),
    .B(_1686_),
    .C(_1687_),
    .Y(_1688_));
 sg13g2_nor2_1 _2562_ (.A(_1224_),
    .B(_1685_),
    .Y(_1689_));
 sg13g2_o21ai_1 _2563_ (.B1(_1176_),
    .Y(_1690_),
    .A1(_1688_),
    .A2(_1689_));
 sg13g2_nor3_1 _2564_ (.A(_1609_),
    .B(_1610_),
    .C(_1628_),
    .Y(_1691_));
 sg13g2_nor2_1 _2565_ (.A(_1626_),
    .B(_1691_),
    .Y(_1692_));
 sg13g2_nand4_1 _2566_ (.B(_1619_),
    .C(_1622_),
    .A(_1618_),
    .Y(_1693_),
    .D(_1692_));
 sg13g2_nor4_2 _2567_ (.A(_1339_),
    .B(_1377_),
    .C(_1391_),
    .Y(_1694_),
    .D(_1407_));
 sg13g2_nand4_1 _2568_ (.B(_1685_),
    .C(_1693_),
    .A(_1670_),
    .Y(_0240_),
    .D(_1694_));
 sg13g2_inv_1 _2569_ (.Y(_0241_),
    .A(_0240_));
 sg13g2_a21oi_2 _2570_ (.B1(_0241_),
    .Y(_0242_),
    .A2(_1694_),
    .A1(_1690_));
 sg13g2_or4_1 _2571_ (.A(\product_comp[10] ),
    .B(_1671_),
    .C(_1686_),
    .D(_1687_),
    .X(_0243_));
 sg13g2_nand2_1 _2572_ (.Y(_0244_),
    .A(_1176_),
    .B(_1689_));
 sg13g2_nand3_1 _2573_ (.B(_0243_),
    .C(_0244_),
    .A(_1408_),
    .Y(_0245_));
 sg13g2_a21oi_1 _2574_ (.A1(_1299_),
    .A2(_0242_),
    .Y(_0246_),
    .B1(_1297_));
 sg13g2_nor2_1 _2575_ (.A(_1289_),
    .B(_0246_),
    .Y(_0247_));
 sg13g2_nand2_1 _2576_ (.Y(_0248_),
    .A(_0058_),
    .B(net356));
 sg13g2_o21ai_1 _2577_ (.B1(_0248_),
    .Y(uo_out[0]),
    .A1(_1276_),
    .A2(_0247_));
 sg13g2_nor2_1 _2578_ (.A(\matt_venn_vga.color[5] ),
    .B(\matt_venn_vga.color[0] ),
    .Y(_0249_));
 sg13g2_nor4_1 _2579_ (.A(\matt_venn_vga.color[1] ),
    .B(\matt_venn_vga.color[2] ),
    .C(\matt_venn_vga.color[3] ),
    .D(\matt_venn_vga.color[4] ),
    .Y(_0250_));
 sg13g2_a21oi_2 _2580_ (.B1(_1298_),
    .Y(_0251_),
    .A2(_0250_),
    .A1(_0249_));
 sg13g2_inv_1 _2581_ (.Y(_0252_),
    .A(_0251_));
 sg13g2_nor2_1 _2582_ (.A(\matt_venn_vga_shadow.color[0] ),
    .B(\matt_venn_vga_shadow.color[1] ),
    .Y(_0253_));
 sg13g2_nor4_1 _2583_ (.A(\matt_venn_vga_shadow.color[2] ),
    .B(\matt_venn_vga_shadow.color[3] ),
    .C(\matt_venn_vga_shadow.color[4] ),
    .D(\matt_venn_vga_shadow.color[5] ),
    .Y(_0254_));
 sg13g2_nand2_1 _2584_ (.Y(_0255_),
    .A(_0253_),
    .B(_0254_));
 sg13g2_nand4_1 _2585_ (.B(\matt_venn_vga_shadow.draw ),
    .C(\matt_venn_vga.activevideo ),
    .A(net5),
    .Y(_0256_),
    .D(_0255_));
 sg13g2_nor2_1 _2586_ (.A(_0251_),
    .B(_0256_),
    .Y(_0257_));
 sg13g2_xor2_1 _2587_ (.B(net316),
    .A(net331),
    .X(_0258_));
 sg13g2_xnor2_1 _2588_ (.Y(_0259_),
    .A(_0027_),
    .B(_0258_));
 sg13g2_xor2_1 _2589_ (.B(\h[0] ),
    .A(net332),
    .X(_0260_));
 sg13g2_xor2_1 _2590_ (.B(_0260_),
    .A(net330),
    .X(_0261_));
 sg13g2_nor2_2 _2591_ (.A(_0259_),
    .B(_0261_),
    .Y(_0262_));
 sg13g2_nor3_1 _2592_ (.A(net324),
    .B(_1223_),
    .C(_1271_),
    .Y(_0263_));
 sg13g2_a22oi_1 _2593_ (.Y(_0264_),
    .B1(_0263_),
    .B2(_0260_),
    .A2(_0262_),
    .A1(net315));
 sg13g2_nor2b_1 _2594_ (.A(net315),
    .B_N(net330),
    .Y(_0265_));
 sg13g2_o21ai_1 _2595_ (.B1(_0262_),
    .Y(_0266_),
    .A1(_0057_),
    .A2(_0265_));
 sg13g2_o21ai_1 _2596_ (.B1(_0266_),
    .Y(_0267_),
    .A1(net330),
    .A2(_0264_));
 sg13g2_nor4_2 _2597_ (.A(net318),
    .B(net319),
    .C(net320),
    .Y(_0268_),
    .D(net322));
 sg13g2_nand3_1 _2598_ (.B(_0267_),
    .C(_0268_),
    .A(_0252_),
    .Y(_0269_));
 sg13g2_nand2b_1 _2599_ (.Y(_0270_),
    .B(_0269_),
    .A_N(_0257_));
 sg13g2_a21oi_1 _2600_ (.A1(_1226_),
    .A2(_0251_),
    .Y(_0271_),
    .B1(_0270_));
 sg13g2_a21o_1 _2601_ (.A2(_0271_),
    .A1(_0242_),
    .B1(_1297_),
    .X(_0272_));
 sg13g2_nand2_1 _2602_ (.Y(_0273_),
    .A(_1292_),
    .B(_0262_));
 sg13g2_nand3_1 _2603_ (.B(_0272_),
    .C(_0273_),
    .A(_1284_),
    .Y(_0274_));
 sg13g2_xnor2_1 _2604_ (.Y(_0275_),
    .A(net355),
    .B(\vga_sync.vsync ));
 sg13g2_nand2_1 _2605_ (.Y(_0276_),
    .A(net356),
    .B(_0275_));
 sg13g2_o21ai_1 _2606_ (.B1(_0276_),
    .Y(uo_out[1]),
    .A1(_1276_),
    .A2(_0274_));
 sg13g2_nor2_1 _2607_ (.A(_1297_),
    .B(_0257_),
    .Y(_0277_));
 sg13g2_inv_1 _2608_ (.Y(_0278_),
    .A(_0277_));
 sg13g2_and2_1 _2609_ (.A(_0242_),
    .B(_0277_),
    .X(_0279_));
 sg13g2_o21ai_1 _2610_ (.B1(_0279_),
    .Y(_0280_),
    .A1(\matt_venn_vga.color[1] ),
    .A2(_0252_));
 sg13g2_nand2b_1 _2611_ (.Y(_0281_),
    .B(_0251_),
    .A_N(\matt_venn_vga.color[0] ));
 sg13g2_nand2_1 _2612_ (.Y(_0282_),
    .A(_0279_),
    .B(_0281_));
 sg13g2_nand3_1 _2613_ (.B(_0279_),
    .C(_0281_),
    .A(net4),
    .Y(_0283_));
 sg13g2_o21ai_1 _2614_ (.B1(_0283_),
    .Y(uo_out[2]),
    .A1(_1276_),
    .A2(_0280_));
 sg13g2_nor2_1 _2615_ (.A(net356),
    .B(_0275_),
    .Y(_0284_));
 sg13g2_a21oi_2 _2616_ (.B1(_0284_),
    .Y(uo_out[3]),
    .A2(_0280_),
    .A1(net356));
 sg13g2_a21oi_1 _2617_ (.A1(_1227_),
    .A2(_0251_),
    .Y(_0285_),
    .B1(_0270_));
 sg13g2_a21oi_1 _2618_ (.A1(_0240_),
    .A2(_0285_),
    .Y(_0286_),
    .B1(_1296_));
 sg13g2_a21oi_1 _2619_ (.A1(_0245_),
    .A2(_0286_),
    .Y(_0287_),
    .B1(_1292_));
 sg13g2_o21ai_1 _2620_ (.B1(_1288_),
    .Y(_0288_),
    .A1(_1285_),
    .A2(_0287_));
 sg13g2_or2_1 _2621_ (.X(_0289_),
    .B(_0288_),
    .A(_1276_));
 sg13g2_and2_1 _2622_ (.A(_1297_),
    .B(_0262_),
    .X(_0290_));
 sg13g2_nand2_1 _2623_ (.Y(_0291_),
    .A(\matt_venn_vga.color[2] ),
    .B(_0251_));
 sg13g2_a21oi_1 _2624_ (.A1(_0269_),
    .A2(_0291_),
    .Y(_0292_),
    .B1(_0278_));
 sg13g2_a21o_1 _2625_ (.A2(_0292_),
    .A1(_0242_),
    .B1(_0290_),
    .X(_0293_));
 sg13g2_a21oi_1 _2626_ (.A1(_1284_),
    .A2(_0293_),
    .Y(_0294_),
    .B1(_1289_));
 sg13g2_o21ai_1 _2627_ (.B1(_0289_),
    .Y(uo_out[4]),
    .A1(_1228_),
    .A2(_0294_));
 sg13g2_nand4_1 _2628_ (.B(_1284_),
    .C(_0272_),
    .A(net356),
    .Y(_0295_),
    .D(_0273_));
 sg13g2_o21ai_1 _2629_ (.B1(_0295_),
    .Y(uo_out[5]),
    .A1(_1276_),
    .A2(_0294_));
 sg13g2_or2_1 _2630_ (.X(_0296_),
    .B(_0288_),
    .A(_1228_));
 sg13g2_o21ai_1 _2631_ (.B1(_0296_),
    .Y(uo_out[6]),
    .A1(_1276_),
    .A2(_0282_));
 sg13g2_nor2_1 _2632_ (.A(_0058_),
    .B(net356),
    .Y(_0297_));
 sg13g2_a21oi_2 _2633_ (.B1(_0297_),
    .Y(uo_out[7]),
    .A2(_0247_),
    .A1(net356));
 sg13g2_nor3_1 _2634_ (.A(net306),
    .B(_1213_),
    .C(net305),
    .Y(_0298_));
 sg13g2_nor2_2 _2635_ (.A(net305),
    .B(_1243_),
    .Y(_0299_));
 sg13g2_and2_1 _2636_ (.A(_0050_),
    .B(_0299_),
    .X(_0300_));
 sg13g2_nand2_2 _2637_ (.Y(_0301_),
    .A(_0050_),
    .B(_0299_));
 sg13g2_nor2_2 _2638_ (.A(net306),
    .B(_0301_),
    .Y(_0302_));
 sg13g2_inv_1 _2639_ (.Y(_0303_),
    .A(_0302_));
 sg13g2_nand2_1 _2640_ (.Y(_0304_),
    .A(\h[8] ),
    .B(_1217_));
 sg13g2_xor2_1 _2641_ (.B(net305),
    .A(\h[8] ),
    .X(_0305_));
 sg13g2_a21oi_2 _2642_ (.B1(_0299_),
    .Y(_0306_),
    .A2(_0305_),
    .A1(_1243_));
 sg13g2_xnor2_1 _2643_ (.Y(_0307_),
    .A(_0050_),
    .B(_1243_));
 sg13g2_nor2b_1 _2644_ (.A(net301),
    .B_N(_0307_),
    .Y(_0308_));
 sg13g2_and2_1 _2645_ (.A(net306),
    .B(_0308_),
    .X(_0309_));
 sg13g2_nand2_1 _2646_ (.Y(_0310_),
    .A(_1245_),
    .B(_0308_));
 sg13g2_nor2_1 _2647_ (.A(_0062_),
    .B(_0310_),
    .Y(_0311_));
 sg13g2_nor2_2 _2648_ (.A(net301),
    .B(_0307_),
    .Y(_0312_));
 sg13g2_inv_1 _2649_ (.Y(_0313_),
    .A(_0312_));
 sg13g2_nor2_2 _2650_ (.A(_0298_),
    .B(_0312_),
    .Y(_0314_));
 sg13g2_nor2b_1 _2651_ (.A(net301),
    .B_N(_0032_),
    .Y(_0315_));
 sg13g2_o21ai_1 _2652_ (.B1(_0314_),
    .Y(_0316_),
    .A1(_0309_),
    .A2(_0315_));
 sg13g2_nand2_1 _2653_ (.Y(_0317_),
    .A(_0298_),
    .B(_0313_));
 sg13g2_inv_1 _2654_ (.Y(_0318_),
    .A(_0317_));
 sg13g2_o21ai_1 _2655_ (.B1(_0301_),
    .Y(_0319_),
    .A1(\clock_min_u[0] ),
    .A2(_0317_));
 sg13g2_a21oi_1 _2656_ (.A1(_1182_),
    .A2(_0312_),
    .Y(_0320_),
    .B1(_0319_));
 sg13g2_o21ai_1 _2657_ (.B1(_0320_),
    .Y(_0321_),
    .A1(_0311_),
    .A2(_0316_));
 sg13g2_nor2_2 _2658_ (.A(_1245_),
    .B(_0301_),
    .Y(_0322_));
 sg13g2_a21oi_1 _2659_ (.A1(\clock_hrs_u[0] ),
    .A2(_0322_),
    .Y(_0323_),
    .B1(_0302_));
 sg13g2_a22oi_1 _2660_ (.Y(_0324_),
    .B1(_0321_),
    .B2(_0323_),
    .A2(_0302_),
    .A1(_1183_));
 sg13g2_nand2_1 _2661_ (.Y(_0325_),
    .A(net537),
    .B(_0322_));
 sg13g2_nor3_1 _2662_ (.A(_1229_),
    .B(net301),
    .C(_0309_),
    .Y(_0326_));
 sg13g2_nand2_1 _2663_ (.Y(_0327_),
    .A(_0310_),
    .B(_0314_));
 sg13g2_nor2_1 _2664_ (.A(_0326_),
    .B(_0327_),
    .Y(_0328_));
 sg13g2_o21ai_1 _2665_ (.B1(_0301_),
    .Y(_0329_),
    .A1(_0034_),
    .A2(_0317_));
 sg13g2_o21ai_1 _2666_ (.B1(_0325_),
    .Y(_0330_),
    .A1(_0328_),
    .A2(_0329_));
 sg13g2_nor3_1 _2667_ (.A(_0040_),
    .B(net301),
    .C(_0309_),
    .Y(_0331_));
 sg13g2_o21ai_1 _2668_ (.B1(_0314_),
    .Y(_0332_),
    .A1(_0039_),
    .A2(_0310_));
 sg13g2_or2_1 _2669_ (.X(_0333_),
    .B(_0332_),
    .A(_0331_));
 sg13g2_a221oi_1 _2670_ (.B2(_0038_),
    .C1(_0300_),
    .B1(_0318_),
    .A1(_0037_),
    .Y(_0334_),
    .A2(_0312_));
 sg13g2_a22oi_1 _2671_ (.Y(_0335_),
    .B1(_0333_),
    .B2(_0334_),
    .A2(_0322_),
    .A1(_1231_));
 sg13g2_nor2_1 _2672_ (.A(_0302_),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_nand2b_1 _2673_ (.Y(_0337_),
    .B(_0303_),
    .A_N(_0330_));
 sg13g2_inv_1 _2674_ (.Y(_0338_),
    .A(_0337_));
 sg13g2_or2_1 _2675_ (.X(_0339_),
    .B(_0337_),
    .A(_0335_));
 sg13g2_and2_1 _2676_ (.A(_0324_),
    .B(_0339_),
    .X(_0000_));
 sg13g2_or3_1 _2677_ (.A(\clock_sec_u[1] ),
    .B(net301),
    .C(_0309_),
    .X(_0340_));
 sg13g2_o21ai_1 _2678_ (.B1(_0340_),
    .Y(_0341_),
    .A1(\clock_sec_d[1] ),
    .A2(_0310_));
 sg13g2_nor2_1 _2679_ (.A(\clock_min_d[1] ),
    .B(_0313_),
    .Y(_0342_));
 sg13g2_a221oi_1 _2680_ (.B2(_0314_),
    .C1(_0342_),
    .B1(_0341_),
    .A1(_1181_),
    .Y(_0343_),
    .A2(_0318_));
 sg13g2_a21oi_1 _2681_ (.A1(_0042_),
    .A2(_0322_),
    .Y(_0344_),
    .B1(_0302_));
 sg13g2_o21ai_1 _2682_ (.B1(_0344_),
    .Y(_0345_),
    .A1(_0300_),
    .A2(_0343_));
 sg13g2_o21ai_1 _2683_ (.B1(_0345_),
    .Y(_0346_),
    .A1(net527),
    .A2(_0303_));
 sg13g2_and2_1 _2684_ (.A(_0339_),
    .B(_0346_),
    .X(_0001_));
 sg13g2_nand2_1 _2685_ (.Y(_0347_),
    .A(_0330_),
    .B(_0336_));
 sg13g2_mux2_1 _2686_ (.A0(_0347_),
    .A1(_0336_),
    .S(_0324_),
    .X(_0348_));
 sg13g2_inv_1 _2687_ (.Y(_0002_),
    .A(_0348_));
 sg13g2_a21oi_1 _2688_ (.A1(_0324_),
    .A2(_0336_),
    .Y(_0349_),
    .B1(_0338_));
 sg13g2_nor2b_1 _2689_ (.A(_0346_),
    .B_N(_0339_),
    .Y(_0350_));
 sg13g2_mux2_1 _2690_ (.A0(_0350_),
    .A1(_0346_),
    .S(_0349_),
    .X(_0003_));
 sg13g2_nand2_1 _2691_ (.Y(_0351_),
    .A(_0324_),
    .B(_0346_));
 sg13g2_nand2b_1 _2692_ (.Y(_0352_),
    .B(_0351_),
    .A_N(_0347_));
 sg13g2_nand2_1 _2693_ (.Y(_0353_),
    .A(_0335_),
    .B(_0338_));
 sg13g2_nand3_1 _2694_ (.B(_0338_),
    .C(_0346_),
    .A(_0335_),
    .Y(_0354_));
 sg13g2_nand2_1 _2695_ (.Y(_0004_),
    .A(_0352_),
    .B(_0354_));
 sg13g2_o21ai_1 _2696_ (.B1(_0353_),
    .Y(_0005_),
    .A1(_0347_),
    .A2(_0351_));
 sg13g2_nor2_2 _2697_ (.A(\h[3] ),
    .B(\h[2] ),
    .Y(_0355_));
 sg13g2_nand2_2 _2698_ (.Y(_0356_),
    .A(_1215_),
    .B(_0355_));
 sg13g2_nor2_1 _2699_ (.A(net311),
    .B(_0356_),
    .Y(_0357_));
 sg13g2_o21ai_1 _2700_ (.B1(net310),
    .Y(_0358_),
    .A1(net311),
    .A2(_0356_));
 sg13g2_nor2b_2 _2701_ (.A(net306),
    .B_N(_0358_),
    .Y(_0359_));
 sg13g2_xnor2_1 _2702_ (.Y(_0360_),
    .A(net306),
    .B(_0358_));
 sg13g2_inv_1 _2703_ (.Y(_0361_),
    .A(_0360_));
 sg13g2_nor2_2 _2704_ (.A(_0313_),
    .B(_0361_),
    .Y(_0362_));
 sg13g2_nor2_1 _2705_ (.A(net305),
    .B(_0359_),
    .Y(_0363_));
 sg13g2_a21o_2 _2706_ (.A2(_0359_),
    .A1(_0305_),
    .B1(_0363_),
    .X(_0364_));
 sg13g2_a21oi_2 _2707_ (.B1(_0363_),
    .Y(_0365_),
    .A2(_0359_),
    .A1(_0305_));
 sg13g2_xnor2_1 _2708_ (.Y(_0366_),
    .A(_0050_),
    .B(_0359_));
 sg13g2_nor2_2 _2709_ (.A(_0365_),
    .B(_0366_),
    .Y(_0367_));
 sg13g2_nand2_1 _2710_ (.Y(_0368_),
    .A(_1213_),
    .B(_0357_));
 sg13g2_and2_2 _2711_ (.A(_0358_),
    .B(_0368_),
    .X(_0369_));
 sg13g2_nor3_2 _2712_ (.A(_0361_),
    .B(_0365_),
    .C(_0369_),
    .Y(_0370_));
 sg13g2_nor2_1 _2713_ (.A(net305),
    .B(_0361_),
    .Y(_0371_));
 sg13g2_nor3_2 _2714_ (.A(_0367_),
    .B(_0370_),
    .C(_0371_),
    .Y(_0372_));
 sg13g2_nor2b_1 _2715_ (.A(_0369_),
    .B_N(_0308_),
    .Y(_0373_));
 sg13g2_nand2b_1 _2716_ (.Y(_0374_),
    .B(_0308_),
    .A_N(_0369_));
 sg13g2_nor2_1 _2717_ (.A(_0039_),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_nor3_1 _2718_ (.A(_0040_),
    .B(_0365_),
    .C(_0373_),
    .Y(_0376_));
 sg13g2_o21ai_1 _2719_ (.B1(_0372_),
    .Y(_0377_),
    .A1(_0375_),
    .A2(_0376_));
 sg13g2_a21oi_1 _2720_ (.A1(_1230_),
    .A2(_0370_),
    .Y(_0378_),
    .B1(_0367_));
 sg13g2_a21oi_2 _2721_ (.B1(_0313_),
    .Y(_0379_),
    .A2(_0368_),
    .A1(_0359_));
 sg13g2_a221oi_1 _2722_ (.B2(_0378_),
    .C1(_0379_),
    .B1(_0377_),
    .A1(_0037_),
    .Y(_0380_),
    .A2(_0367_));
 sg13g2_a21oi_2 _2723_ (.B1(_0380_),
    .Y(_0381_),
    .A2(_0362_),
    .A1(_1231_));
 sg13g2_o21ai_1 _2724_ (.B1(_0374_),
    .Y(_0382_),
    .A1(_1229_),
    .A2(_0365_));
 sg13g2_a221oi_1 _2725_ (.B2(_0382_),
    .C1(_0367_),
    .B1(_0372_),
    .A1(_0034_),
    .Y(_0383_),
    .A2(_0370_));
 sg13g2_nand2b_2 _2726_ (.Y(_0384_),
    .B(_0322_),
    .A_N(_0369_));
 sg13g2_o21ai_1 _2727_ (.B1(_0384_),
    .Y(_0385_),
    .A1(_0379_),
    .A2(_0383_));
 sg13g2_a21oi_2 _2728_ (.B1(_0385_),
    .Y(_0386_),
    .A2(_0362_),
    .A1(net535));
 sg13g2_nor2b_1 _2729_ (.A(_0381_),
    .B_N(_0386_),
    .Y(_0387_));
 sg13g2_and2_1 _2730_ (.A(_0032_),
    .B(_0374_),
    .X(_0388_));
 sg13g2_a22oi_1 _2731_ (.Y(_0389_),
    .B1(_0388_),
    .B2(_0364_),
    .A2(_0373_),
    .A1(_0062_));
 sg13g2_a221oi_1 _2732_ (.B2(_0389_),
    .C1(_0367_),
    .B1(_0372_),
    .A1(\clock_min_u[0] ),
    .Y(_0390_),
    .A2(_0370_));
 sg13g2_a21oi_1 _2733_ (.A1(_1182_),
    .A2(_0367_),
    .Y(_0391_),
    .B1(_0379_));
 sg13g2_nand2b_1 _2734_ (.Y(_0392_),
    .B(_0391_),
    .A_N(_0390_));
 sg13g2_nand2_1 _2735_ (.Y(_0393_),
    .A(\clock_hrs_u[0] ),
    .B(_0362_));
 sg13g2_nand3_1 _2736_ (.B(_0392_),
    .C(_0393_),
    .A(_0384_),
    .Y(_0394_));
 sg13g2_o21ai_1 _2737_ (.B1(_0394_),
    .Y(_0395_),
    .A1(\clock_hrs_d[0] ),
    .A2(_0384_));
 sg13g2_nor2_1 _2738_ (.A(_0387_),
    .B(_0395_),
    .Y(_0011_));
 sg13g2_nor2_1 _2739_ (.A(\clock_sec_d[1] ),
    .B(_0374_),
    .Y(_0396_));
 sg13g2_nor3_1 _2740_ (.A(\clock_sec_u[1] ),
    .B(_0365_),
    .C(_0373_),
    .Y(_0397_));
 sg13g2_o21ai_1 _2741_ (.B1(_0372_),
    .Y(_0398_),
    .A1(_0396_),
    .A2(_0397_));
 sg13g2_a21oi_1 _2742_ (.A1(_1181_),
    .A2(_0370_),
    .Y(_0399_),
    .B1(_0367_));
 sg13g2_a221oi_1 _2743_ (.B2(_0399_),
    .C1(_0379_),
    .B1(_0398_),
    .A1(\clock_min_d[1] ),
    .Y(_0400_),
    .A2(_0367_));
 sg13g2_a21oi_1 _2744_ (.A1(_0042_),
    .A2(_0362_),
    .Y(_0401_),
    .B1(_0400_));
 sg13g2_nand2_1 _2745_ (.Y(_0402_),
    .A(_0384_),
    .B(_0401_));
 sg13g2_o21ai_1 _2746_ (.B1(_0402_),
    .Y(_0403_),
    .A1(net547),
    .A2(_0384_));
 sg13g2_nor2b_1 _2747_ (.A(_0387_),
    .B_N(_0403_),
    .Y(_0012_));
 sg13g2_nand2b_2 _2748_ (.Y(_0404_),
    .B(_0384_),
    .A_N(_0381_));
 sg13g2_nor2_1 _2749_ (.A(_0395_),
    .B(_0404_),
    .Y(_0405_));
 sg13g2_or2_1 _2750_ (.X(_0406_),
    .B(_0404_),
    .A(_0386_));
 sg13g2_a21oi_1 _2751_ (.A1(_0395_),
    .A2(_0406_),
    .Y(_0013_),
    .B1(_0405_));
 sg13g2_nor2_1 _2752_ (.A(_0386_),
    .B(_0405_),
    .Y(_0407_));
 sg13g2_nor3_1 _2753_ (.A(_0387_),
    .B(_0403_),
    .C(_0407_),
    .Y(_0408_));
 sg13g2_a21o_1 _2754_ (.A2(_0407_),
    .A1(_0403_),
    .B1(_0408_),
    .X(_0014_));
 sg13g2_nand2_1 _2755_ (.Y(_0409_),
    .A(_0381_),
    .B(_0386_));
 sg13g2_nand2b_1 _2756_ (.Y(_0410_),
    .B(_0403_),
    .A_N(_0409_));
 sg13g2_nor2b_1 _2757_ (.A(_0395_),
    .B_N(_0403_),
    .Y(_0411_));
 sg13g2_o21ai_1 _2758_ (.B1(_0410_),
    .Y(_0015_),
    .A1(_0406_),
    .A2(_0411_));
 sg13g2_nand2b_1 _2759_ (.Y(_0412_),
    .B(_0411_),
    .A_N(_0406_));
 sg13g2_nand2_1 _2760_ (.Y(_0016_),
    .A(_0409_),
    .B(_0412_));
 sg13g2_o21ai_1 _2761_ (.B1(net322),
    .Y(_0413_),
    .A1(net324),
    .A2(_1271_));
 sg13g2_nor2_1 _2762_ (.A(_1198_),
    .B(_0413_),
    .Y(_0414_));
 sg13g2_xnor2_1 _2763_ (.Y(_0415_),
    .A(net320),
    .B(_0413_));
 sg13g2_nor2b_2 _2764_ (.A(_1272_),
    .B_N(_0413_),
    .Y(_0416_));
 sg13g2_xnor2_1 _2765_ (.Y(_0417_),
    .A(_1221_),
    .B(_1271_));
 sg13g2_nand2_1 _2766_ (.Y(_0418_),
    .A(\matt_venn_vga.digit_0.digit_index[1] ),
    .B(_0417_));
 sg13g2_nand2_2 _2767_ (.Y(_0419_),
    .A(_1271_),
    .B(_1281_));
 sg13g2_nand2_1 _2768_ (.Y(_0420_),
    .A(\matt_venn_vga.digit_0.digit_index[0] ),
    .B(_0419_));
 sg13g2_xnor2_1 _2769_ (.Y(_0421_),
    .A(\matt_venn_vga.digit_0.digit_index[1] ),
    .B(_0417_));
 sg13g2_o21ai_1 _2770_ (.B1(_0418_),
    .Y(_0422_),
    .A1(_0420_),
    .A2(_0421_));
 sg13g2_xnor2_1 _2771_ (.Y(_0423_),
    .A(\matt_venn_vga.digit_0.digit_index[2] ),
    .B(_0416_));
 sg13g2_nor2b_1 _2772_ (.A(_0423_),
    .B_N(_0422_),
    .Y(_0424_));
 sg13g2_a21o_1 _2773_ (.A2(_0416_),
    .A1(\matt_venn_vga.digit_0.digit_index[2] ),
    .B1(_0424_),
    .X(_0425_));
 sg13g2_xnor2_1 _2774_ (.Y(_0426_),
    .A(\matt_venn_vga.digit_0.digit_index[3] ),
    .B(_0415_));
 sg13g2_nor2b_1 _2775_ (.A(_0426_),
    .B_N(_0425_),
    .Y(_0427_));
 sg13g2_a21oi_1 _2776_ (.A1(\matt_venn_vga.digit_0.digit_index[3] ),
    .A2(_0415_),
    .Y(_0428_),
    .B1(_0427_));
 sg13g2_xnor2_1 _2777_ (.Y(_0429_),
    .A(\matt_venn_vga.y_px[8] ),
    .B(_0414_));
 sg13g2_nand2_1 _2778_ (.Y(_0430_),
    .A(\matt_venn_vga.digit_0.digit_index[4] ),
    .B(_0429_));
 sg13g2_xnor2_1 _2779_ (.Y(_0431_),
    .A(\matt_venn_vga.digit_0.digit_index[4] ),
    .B(_0429_));
 sg13g2_xor2_1 _2780_ (.B(_0431_),
    .A(_0428_),
    .X(_0432_));
 sg13g2_xor2_1 _2781_ (.B(_0423_),
    .A(_0422_),
    .X(_0433_));
 sg13g2_inv_1 _2782_ (.Y(_0434_),
    .A(net297));
 sg13g2_xnor2_1 _2783_ (.Y(_0435_),
    .A(_0425_),
    .B(_0426_));
 sg13g2_nand2_1 _2784_ (.Y(_0436_),
    .A(_0434_),
    .B(net285));
 sg13g2_xor2_1 _2785_ (.B(_0419_),
    .A(\matt_venn_vga.digit_0.digit_index[0] ),
    .X(_0437_));
 sg13g2_nand2_1 _2786_ (.Y(_0438_),
    .A(_0421_),
    .B(_0437_));
 sg13g2_nand3_1 _2787_ (.B(net286),
    .C(_0438_),
    .A(_0434_),
    .Y(_0439_));
 sg13g2_xor2_1 _2788_ (.B(_0421_),
    .A(_0420_),
    .X(_0440_));
 sg13g2_nor2_2 _2789_ (.A(_0437_),
    .B(_0440_),
    .Y(_0441_));
 sg13g2_inv_1 _2790_ (.Y(_0442_),
    .A(_0441_));
 sg13g2_o21ai_1 _2791_ (.B1(_0430_),
    .Y(_0443_),
    .A1(_0428_),
    .A2(_0431_));
 sg13g2_a21oi_1 _2792_ (.A1(_1197_),
    .A2(_0414_),
    .Y(_0444_),
    .B1(_1222_));
 sg13g2_xnor2_1 _2793_ (.Y(_0445_),
    .A(_0052_),
    .B(_0444_));
 sg13g2_xor2_1 _2794_ (.B(_0445_),
    .A(\matt_venn_vga.digit_0.digit_index[5] ),
    .X(_0446_));
 sg13g2_xnor2_1 _2795_ (.Y(_0447_),
    .A(_0443_),
    .B(_0446_));
 sg13g2_xor2_1 _2796_ (.B(_0446_),
    .A(_0443_),
    .X(_0448_));
 sg13g2_nand3_1 _2797_ (.B(_0441_),
    .C(_0447_),
    .A(net286),
    .Y(_0449_));
 sg13g2_o21ai_1 _2798_ (.B1(_0449_),
    .Y(_0450_),
    .A1(_0433_),
    .A2(_0441_));
 sg13g2_a21oi_1 _2799_ (.A1(_0439_),
    .A2(_0450_),
    .Y(_0451_),
    .B1(net282));
 sg13g2_nor2_1 _2800_ (.A(_0434_),
    .B(net286),
    .Y(_0452_));
 sg13g2_nand2b_1 _2801_ (.Y(_0453_),
    .B(_0452_),
    .A_N(_0440_));
 sg13g2_nand3_1 _2802_ (.B(_0448_),
    .C(_0453_),
    .A(_0436_),
    .Y(_0454_));
 sg13g2_nand2_1 _2803_ (.Y(_0455_),
    .A(net297),
    .B(_0437_));
 sg13g2_nand3_1 _2804_ (.B(_0440_),
    .C(_0455_),
    .A(net286),
    .Y(_0456_));
 sg13g2_a21o_1 _2805_ (.A2(_0456_),
    .A1(net282),
    .B1(_0448_),
    .X(_0457_));
 sg13g2_a21o_1 _2806_ (.A2(_0457_),
    .A1(_0454_),
    .B1(_0451_),
    .X(_0008_));
 sg13g2_o21ai_1 _2807_ (.B1(_0437_),
    .Y(_0458_),
    .A1(_0421_),
    .A2(net297));
 sg13g2_a21oi_1 _2808_ (.A1(_0421_),
    .A2(net297),
    .Y(_0459_),
    .B1(_0458_));
 sg13g2_nand2b_1 _2809_ (.Y(_0460_),
    .B(_0459_),
    .A_N(net285));
 sg13g2_nand3_1 _2810_ (.B(_0436_),
    .C(_0460_),
    .A(net282),
    .Y(_0461_));
 sg13g2_xnor2_1 _2811_ (.Y(_0462_),
    .A(net297),
    .B(_0438_));
 sg13g2_nand2b_1 _2812_ (.Y(_0463_),
    .B(_0440_),
    .A_N(_0437_));
 sg13g2_o21ai_1 _2813_ (.B1(_0455_),
    .Y(_0464_),
    .A1(net297),
    .A2(_0463_));
 sg13g2_nor2_1 _2814_ (.A(net285),
    .B(_0462_),
    .Y(_0465_));
 sg13g2_a21oi_1 _2815_ (.A1(net286),
    .A2(_0464_),
    .Y(_0466_),
    .B1(_0465_));
 sg13g2_o21ai_1 _2816_ (.B1(_0461_),
    .Y(_0467_),
    .A1(net282),
    .A2(_0466_));
 sg13g2_a221oi_1 _2817_ (.B2(net285),
    .C1(net282),
    .B1(_0459_),
    .A1(_0442_),
    .Y(_0468_),
    .A2(_0452_));
 sg13g2_o21ai_1 _2818_ (.B1(net282),
    .Y(_0469_),
    .A1(net285),
    .A2(_0464_));
 sg13g2_a21oi_1 _2819_ (.A1(net286),
    .A2(_0458_),
    .Y(_0470_),
    .B1(_0469_));
 sg13g2_nor3_1 _2820_ (.A(_0448_),
    .B(_0468_),
    .C(_0470_),
    .Y(_0471_));
 sg13g2_a21oi_1 _2821_ (.A1(_0448_),
    .A2(_0467_),
    .Y(_0009_),
    .B1(_0471_));
 sg13g2_nor2_1 _2822_ (.A(net297),
    .B(_0437_),
    .Y(_0472_));
 sg13g2_nor2_1 _2823_ (.A(net285),
    .B(_0472_),
    .Y(_0473_));
 sg13g2_a22oi_1 _2824_ (.Y(_0474_),
    .B1(_0458_),
    .B2(_0473_),
    .A2(_0441_),
    .A1(net286));
 sg13g2_nand3_1 _2825_ (.B(_0438_),
    .C(_0463_),
    .A(net297),
    .Y(_0475_));
 sg13g2_a21oi_1 _2826_ (.A1(_0434_),
    .A2(_0440_),
    .Y(_0476_),
    .B1(net285));
 sg13g2_a21oi_1 _2827_ (.A1(net285),
    .A2(_0475_),
    .Y(_0477_),
    .B1(_0476_));
 sg13g2_o21ai_1 _2828_ (.B1(_0447_),
    .Y(_0478_),
    .A1(net282),
    .A2(_0477_));
 sg13g2_a21oi_1 _2829_ (.A1(net282),
    .A2(_0474_),
    .Y(_0479_),
    .B1(_0478_));
 sg13g2_nor2_1 _2830_ (.A(_0433_),
    .B(_0440_),
    .Y(_0480_));
 sg13g2_o21ai_1 _2831_ (.B1(_0436_),
    .Y(_0481_),
    .A1(_0432_),
    .A2(_0480_));
 sg13g2_nor2_1 _2832_ (.A(_0447_),
    .B(_0481_),
    .Y(_0482_));
 sg13g2_nor2_1 _2833_ (.A(_0479_),
    .B(_0482_),
    .Y(_0010_));
 sg13g2_nand2_1 _2834_ (.Y(_0483_),
    .A(_0025_),
    .B(_1252_));
 sg13g2_xnor2_1 _2835_ (.Y(_0484_),
    .A(_1221_),
    .B(_0483_));
 sg13g2_nand2_1 _2836_ (.Y(_0485_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[1] ),
    .B(_0484_));
 sg13g2_xor2_1 _2837_ (.B(_1252_),
    .A(\matt_venn_vga.y_px[4] ),
    .X(_0486_));
 sg13g2_nand2_1 _2838_ (.Y(_0487_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[0] ),
    .B(_0486_));
 sg13g2_xnor2_1 _2839_ (.Y(_0488_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[1] ),
    .B(_0484_));
 sg13g2_o21ai_1 _2840_ (.B1(_0485_),
    .Y(_0489_),
    .A1(_0487_),
    .A2(_0488_));
 sg13g2_nor3_2 _2841_ (.A(net324),
    .B(\matt_venn_vga.y_px[4] ),
    .C(_1253_),
    .Y(_0490_));
 sg13g2_nor2b_2 _2842_ (.A(_0490_),
    .B_N(net323),
    .Y(_0491_));
 sg13g2_xnor2_1 _2843_ (.Y(_0492_),
    .A(net322),
    .B(_0490_));
 sg13g2_xnor2_1 _2844_ (.Y(_0493_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[2] ),
    .B(_0492_));
 sg13g2_nor2b_1 _2845_ (.A(_0493_),
    .B_N(_0489_),
    .Y(_0494_));
 sg13g2_xnor2_1 _2846_ (.Y(_0495_),
    .A(_0489_),
    .B(_0493_));
 sg13g2_xor2_1 _2847_ (.B(_0493_),
    .A(_0489_),
    .X(_0496_));
 sg13g2_a21oi_1 _2848_ (.A1(\matt_venn_vga_shadow.digit_0.digit_index[2] ),
    .A2(_0492_),
    .Y(_0497_),
    .B1(_0494_));
 sg13g2_xnor2_1 _2849_ (.Y(_0498_),
    .A(net533),
    .B(_0491_));
 sg13g2_nand2_1 _2850_ (.Y(_0499_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[3] ),
    .B(_0498_));
 sg13g2_xnor2_1 _2851_ (.Y(_0500_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[3] ),
    .B(_0498_));
 sg13g2_xnor2_1 _2852_ (.Y(_0501_),
    .A(_0497_),
    .B(_0500_));
 sg13g2_or2_1 _2853_ (.X(_0502_),
    .B(net283),
    .A(net295));
 sg13g2_nand2_1 _2854_ (.Y(_0503_),
    .A(net321),
    .B(_0491_));
 sg13g2_xnor2_1 _2855_ (.Y(_0504_),
    .A(_1222_),
    .B(_0503_));
 sg13g2_nor2b_1 _2856_ (.A(_0504_),
    .B_N(\matt_venn_vga_shadow.digit_0.digit_index[4] ),
    .Y(_0505_));
 sg13g2_xnor2_1 _2857_ (.Y(_0506_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[4] ),
    .B(_0504_));
 sg13g2_o21ai_1 _2858_ (.B1(_0499_),
    .Y(_0507_),
    .A1(_0497_),
    .A2(_0500_));
 sg13g2_a21o_1 _2859_ (.A2(_0507_),
    .A1(_0506_),
    .B1(_0505_),
    .X(_0508_));
 sg13g2_a21oi_1 _2860_ (.A1(net321),
    .A2(_0491_),
    .Y(_0509_),
    .B1(net319));
 sg13g2_xnor2_1 _2861_ (.Y(_0510_),
    .A(_0052_),
    .B(_0509_));
 sg13g2_xnor2_1 _2862_ (.Y(_0511_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[5] ),
    .B(_0510_));
 sg13g2_xnor2_1 _2863_ (.Y(_0512_),
    .A(_0508_),
    .B(_0511_));
 sg13g2_xor2_1 _2864_ (.B(_0507_),
    .A(_0506_),
    .X(_0513_));
 sg13g2_inv_1 _2865_ (.Y(_0514_),
    .A(net281));
 sg13g2_xor2_1 _2866_ (.B(_0486_),
    .A(\matt_venn_vga_shadow.digit_0.digit_index[0] ),
    .X(_0515_));
 sg13g2_and2_1 _2867_ (.A(_0488_),
    .B(_0515_),
    .X(_0516_));
 sg13g2_xnor2_1 _2868_ (.Y(_0517_),
    .A(_0487_),
    .B(_0488_));
 sg13g2_nand2_1 _2869_ (.Y(_0518_),
    .A(_0501_),
    .B(_0517_));
 sg13g2_nor2b_1 _2870_ (.A(_0515_),
    .B_N(_0517_),
    .Y(_0519_));
 sg13g2_o21ai_1 _2871_ (.B1(_0514_),
    .Y(_0520_),
    .A1(net295),
    .A2(_0519_));
 sg13g2_o21ai_1 _2872_ (.B1(_0520_),
    .Y(_0521_),
    .A1(_0495_),
    .A2(_0518_));
 sg13g2_nand2_1 _2873_ (.Y(_0522_),
    .A(net295),
    .B(_0515_));
 sg13g2_a21oi_1 _2874_ (.A1(net295),
    .A2(_0515_),
    .Y(_0523_),
    .B1(_0517_));
 sg13g2_nor2_1 _2875_ (.A(_0514_),
    .B(_0523_),
    .Y(_0524_));
 sg13g2_o21ai_1 _2876_ (.B1(_0501_),
    .Y(_0525_),
    .A1(net281),
    .A2(_0519_));
 sg13g2_nor3_1 _2877_ (.A(_0495_),
    .B(net281),
    .C(_0519_),
    .Y(_0526_));
 sg13g2_nor2b_1 _2878_ (.A(_0521_),
    .B_N(_0502_),
    .Y(_0527_));
 sg13g2_nor2b_1 _2879_ (.A(_0512_),
    .B_N(_0525_),
    .Y(_0528_));
 sg13g2_nor3_1 _2880_ (.A(_0502_),
    .B(net281),
    .C(_0516_),
    .Y(_0529_));
 sg13g2_nor3_1 _2881_ (.A(_0524_),
    .B(_0526_),
    .C(_0529_),
    .Y(_0530_));
 sg13g2_a22oi_1 _2882_ (.Y(_0019_),
    .B1(_0528_),
    .B2(_0530_),
    .A2(_0527_),
    .A1(_0512_));
 sg13g2_nand2_1 _2883_ (.Y(_0531_),
    .A(_0495_),
    .B(_0516_));
 sg13g2_o21ai_1 _2884_ (.B1(_0531_),
    .Y(_0532_),
    .A1(_0488_),
    .A2(_0522_));
 sg13g2_inv_1 _2885_ (.Y(_0533_),
    .A(_0532_));
 sg13g2_nand2_1 _2886_ (.Y(_0534_),
    .A(_0502_),
    .B(net281));
 sg13g2_xnor2_1 _2887_ (.Y(_0535_),
    .A(_0496_),
    .B(_0516_));
 sg13g2_or2_1 _2888_ (.X(_0536_),
    .B(_0517_),
    .A(_0515_));
 sg13g2_o21ai_1 _2889_ (.B1(_0522_),
    .Y(_0537_),
    .A1(_0496_),
    .A2(_0536_));
 sg13g2_inv_1 _2890_ (.Y(_0538_),
    .A(_0537_));
 sg13g2_mux4_1 _2891_ (.S0(net283),
    .A0(_0537_),
    .A1(_0535_),
    .A2(net295),
    .A3(_0533_),
    .S1(net281),
    .X(_0539_));
 sg13g2_o21ai_1 _2892_ (.B1(_0515_),
    .Y(_0540_),
    .A1(_0488_),
    .A2(net295));
 sg13g2_a21oi_1 _2893_ (.A1(net281),
    .A2(_0540_),
    .Y(_0541_),
    .B1(net283));
 sg13g2_o21ai_1 _2894_ (.B1(_0541_),
    .Y(_0542_),
    .A1(net281),
    .A2(_0533_));
 sg13g2_a21oi_1 _2895_ (.A1(_0513_),
    .A2(_0538_),
    .Y(_0543_),
    .B1(_0526_));
 sg13g2_a21oi_1 _2896_ (.A1(net283),
    .A2(_0543_),
    .Y(_0544_),
    .B1(_0512_));
 sg13g2_a22oi_1 _2897_ (.Y(_0020_),
    .B1(_0542_),
    .B2(_0544_),
    .A2(_0539_),
    .A1(_0512_));
 sg13g2_o21ai_1 _2898_ (.B1(_0540_),
    .Y(_0545_),
    .A1(net295),
    .A2(_0515_));
 sg13g2_nand2b_1 _2899_ (.Y(_0546_),
    .B(net283),
    .A_N(_0545_));
 sg13g2_nand2b_1 _2900_ (.Y(_0547_),
    .B(_0519_),
    .A_N(net283));
 sg13g2_nand3_1 _2901_ (.B(_0546_),
    .C(_0547_),
    .A(_0513_),
    .Y(_0548_));
 sg13g2_nor2_1 _2902_ (.A(net295),
    .B(_0517_),
    .Y(_0549_));
 sg13g2_nor3_1 _2903_ (.A(_0495_),
    .B(net283),
    .C(_0516_),
    .Y(_0550_));
 sg13g2_a22oi_1 _2904_ (.Y(_0551_),
    .B1(_0550_),
    .B2(_0536_),
    .A2(_0549_),
    .A1(net283));
 sg13g2_a21oi_1 _2905_ (.A1(_0514_),
    .A2(_0551_),
    .Y(_0552_),
    .B1(_0512_));
 sg13g2_o21ai_1 _2906_ (.B1(_0534_),
    .Y(_0553_),
    .A1(_0496_),
    .A2(_0518_));
 sg13g2_a22oi_1 _2907_ (.Y(_0021_),
    .B1(_0553_),
    .B2(_0512_),
    .A2(_0552_),
    .A1(_0548_));
 sg13g2_nand2_1 _2908_ (.Y(_0554_),
    .A(\clock_color_offset[0] ),
    .B(_0369_));
 sg13g2_xor2_1 _2909_ (.B(_0369_),
    .A(\clock_color_offset[0] ),
    .X(_0555_));
 sg13g2_xnor2_1 _2910_ (.Y(_0556_),
    .A(net544),
    .B(_0360_));
 sg13g2_nand2_1 _2911_ (.Y(_0557_),
    .A(_0555_),
    .B(_0556_));
 sg13g2_nand2b_1 _2912_ (.Y(_0558_),
    .B(_0556_),
    .A_N(_0554_));
 sg13g2_o21ai_1 _2913_ (.B1(_0558_),
    .Y(_0559_),
    .A1(_0051_),
    .A2(_0360_));
 sg13g2_xnor2_1 _2914_ (.Y(_0560_),
    .A(\clock_color_offset[2] ),
    .B(_0366_));
 sg13g2_xnor2_1 _2915_ (.Y(_0561_),
    .A(_0559_),
    .B(_0560_));
 sg13g2_inv_1 _2916_ (.Y(_0562_),
    .A(_0561_));
 sg13g2_xor2_1 _2917_ (.B(_0556_),
    .A(_0554_),
    .X(_0563_));
 sg13g2_a22oi_1 _2918_ (.Y(_0017_),
    .B1(_0561_),
    .B2(_0563_),
    .A2(_0556_),
    .A1(_0555_));
 sg13g2_mux2_1 _2919_ (.A0(_0557_),
    .A1(_0555_),
    .S(_0561_),
    .X(_0018_));
 sg13g2_nor2b_1 _2920_ (.A(net310),
    .B_N(\clock_color_offset[0] ),
    .Y(_0564_));
 sg13g2_xnor2_1 _2921_ (.Y(_0565_),
    .A(\clock_color_offset[0] ),
    .B(net310));
 sg13g2_xor2_1 _2922_ (.B(_1246_),
    .A(net549),
    .X(_0566_));
 sg13g2_nand2_1 _2923_ (.Y(_0567_),
    .A(_0565_),
    .B(_0566_));
 sg13g2_xnor2_1 _2924_ (.Y(_0568_),
    .A(_0564_),
    .B(_0566_));
 sg13g2_a22oi_1 _2925_ (.Y(_0569_),
    .B1(_0564_),
    .B2(_0566_),
    .A2(_1246_),
    .A1(_1214_));
 sg13g2_xor2_1 _2926_ (.B(_0307_),
    .A(\clock_color_offset[2] ),
    .X(_0570_));
 sg13g2_xnor2_1 _2927_ (.Y(_0571_),
    .A(_0569_),
    .B(_0570_));
 sg13g2_inv_1 _2928_ (.Y(_0572_),
    .A(_0571_));
 sg13g2_a22oi_1 _2929_ (.Y(_0006_),
    .B1(_0568_),
    .B2(_0571_),
    .A2(_0566_),
    .A1(_0565_));
 sg13g2_mux2_1 _2930_ (.A0(_0567_),
    .A1(_0565_),
    .S(_0571_),
    .X(_0007_));
 sg13g2_nand2b_1 _2931_ (.Y(_0573_),
    .B(_0563_),
    .A_N(_0555_));
 sg13g2_nor2b_1 _2932_ (.A(_0561_),
    .B_N(_0573_),
    .Y(_0068_));
 sg13g2_a21oi_1 _2933_ (.A1(_0557_),
    .A2(_0573_),
    .Y(_0069_),
    .B1(_0562_));
 sg13g2_and2_1 _2934_ (.A(_0557_),
    .B(_0561_),
    .X(_0070_));
 sg13g2_and2_2 _2935_ (.A(hmax),
    .B(\vga_sync.o_vmax ),
    .X(_0574_));
 sg13g2_nand2_2 _2936_ (.Y(_0575_),
    .A(hmax),
    .B(\vga_sync.o_vmax ));
 sg13g2_nand3b_1 _2937_ (.B(net313),
    .C(_1236_),
    .Y(_0576_),
    .A_N(net311));
 sg13g2_nor4_1 _2938_ (.A(_0050_),
    .B(_1216_),
    .C(_1241_),
    .D(_0576_),
    .Y(_0577_));
 sg13g2_nand3_1 _2939_ (.B(_1246_),
    .C(_0577_),
    .A(_1240_),
    .Y(_0578_));
 sg13g2_nand4_1 _2940_ (.B(_1246_),
    .C(\vga_sync.o_vmax ),
    .A(_1240_),
    .Y(_0579_),
    .D(_0577_));
 sg13g2_inv_2 _2941_ (.Y(_0580_),
    .A(_0579_));
 sg13g2_and4_2 _2942_ (.A(hmax),
    .B(_1251_),
    .C(_1257_),
    .D(_1258_),
    .X(_0581_));
 sg13g2_a21oi_1 _2943_ (.A1(\ydelta[0] ),
    .A2(_0579_),
    .Y(_0582_),
    .B1(net351));
 sg13g2_nor2_1 _2944_ (.A(\ydelta[1] ),
    .B(\ydelta[0] ),
    .Y(_0583_));
 sg13g2_nor3_2 _2945_ (.A(\ydelta[2] ),
    .B(\ydelta[1] ),
    .C(\ydelta[0] ),
    .Y(_0584_));
 sg13g2_nand2b_2 _2946_ (.Y(_0585_),
    .B(_0584_),
    .A_N(\ydelta[3] ));
 sg13g2_nor3_2 _2947_ (.A(\ydelta[5] ),
    .B(\ydelta[4] ),
    .C(_0585_),
    .Y(_0586_));
 sg13g2_nor2b_2 _2948_ (.A(\ydelta[6] ),
    .B_N(_0586_),
    .Y(_0587_));
 sg13g2_o21ai_1 _2949_ (.B1(_0022_),
    .Y(_0588_),
    .A1(_1209_),
    .A2(_0587_));
 sg13g2_xor2_1 _2950_ (.B(_0586_),
    .A(\ydelta[6] ),
    .X(_0589_));
 sg13g2_inv_1 _2951_ (.Y(_0590_),
    .A(_0589_));
 sg13g2_xor2_1 _2952_ (.B(net349),
    .A(\py[7] ),
    .X(_0591_));
 sg13g2_xor2_1 _2953_ (.B(_0591_),
    .A(_0587_),
    .X(_0592_));
 sg13g2_o21ai_1 _2954_ (.B1(_0592_),
    .Y(_0593_),
    .A1(_1203_),
    .A2(_0590_));
 sg13g2_xnor2_1 _2955_ (.Y(_0594_),
    .A(net339),
    .B(\ydelta[4] ));
 sg13g2_nand2_1 _2956_ (.Y(_0595_),
    .A(\py[2] ),
    .B(\ydelta[2] ));
 sg13g2_xor2_1 _2957_ (.B(\ydelta[2] ),
    .A(\py[2] ),
    .X(_0596_));
 sg13g2_xnor2_1 _2958_ (.Y(_0597_),
    .A(_0583_),
    .B(_0596_));
 sg13g2_nor2_1 _2959_ (.A(\py[3] ),
    .B(\ydelta[3] ),
    .Y(_0598_));
 sg13g2_xor2_1 _2960_ (.B(\ydelta[3] ),
    .A(\py[3] ),
    .X(_0599_));
 sg13g2_xnor2_1 _2961_ (.Y(_0600_),
    .A(_0584_),
    .B(_0599_));
 sg13g2_nor2_1 _2962_ (.A(_0597_),
    .B(_0600_),
    .Y(_0601_));
 sg13g2_nand2_1 _2963_ (.Y(_0602_),
    .A(net340),
    .B(\ydelta[1] ));
 sg13g2_nand2_1 _2964_ (.Y(_0603_),
    .A(net341),
    .B(\ydelta[0] ));
 sg13g2_xnor2_1 _2965_ (.Y(_0604_),
    .A(net340),
    .B(\ydelta[1] ));
 sg13g2_o21ai_1 _2966_ (.B1(_0602_),
    .Y(_0605_),
    .A1(_0603_),
    .A2(_0604_));
 sg13g2_nor2_1 _2967_ (.A(_0595_),
    .B(_0598_),
    .Y(_0606_));
 sg13g2_a221oi_1 _2968_ (.B2(_0605_),
    .C1(_0606_),
    .B1(_0601_),
    .A1(\py[3] ),
    .Y(_0607_),
    .A2(\ydelta[3] ));
 sg13g2_nor2_1 _2969_ (.A(_0594_),
    .B(_0607_),
    .Y(_0608_));
 sg13g2_xnor2_1 _2970_ (.Y(_0609_),
    .A(_0594_),
    .B(_0607_));
 sg13g2_xor2_1 _2971_ (.B(\ydelta[0] ),
    .A(\ydelta[1] ),
    .X(_0610_));
 sg13g2_xnor2_1 _2972_ (.Y(_0611_),
    .A(net341),
    .B(\ydelta[0] ));
 sg13g2_xnor2_1 _2973_ (.Y(_0612_),
    .A(net340),
    .B(_0610_));
 sg13g2_nand3_1 _2974_ (.B(_0611_),
    .C(_0612_),
    .A(_0601_),
    .Y(_0613_));
 sg13g2_xnor2_1 _2975_ (.Y(_0614_),
    .A(\ydelta[4] ),
    .B(_0585_));
 sg13g2_o21ai_1 _2976_ (.B1(\ydelta[5] ),
    .Y(_0615_),
    .A1(\ydelta[4] ),
    .A2(_0585_));
 sg13g2_nor2b_1 _2977_ (.A(_0586_),
    .B_N(_0615_),
    .Y(_0616_));
 sg13g2_nand2b_1 _2978_ (.Y(_0617_),
    .B(\py[5] ),
    .A_N(_0616_));
 sg13g2_nor2_1 _2979_ (.A(\py[6] ),
    .B(_0589_),
    .Y(_0618_));
 sg13g2_nand2b_1 _2980_ (.Y(_0619_),
    .B(_0616_),
    .A_N(\py[5] ));
 sg13g2_a22oi_1 _2981_ (.Y(_0620_),
    .B1(_0614_),
    .B2(net339),
    .A2(_0613_),
    .A1(_0609_));
 sg13g2_o21ai_1 _2982_ (.B1(_0619_),
    .Y(_0621_),
    .A1(net339),
    .A2(_0614_));
 sg13g2_o21ai_1 _2983_ (.B1(_0617_),
    .Y(_0622_),
    .A1(_0620_),
    .A2(_0621_));
 sg13g2_nor2b_1 _2984_ (.A(_0618_),
    .B_N(_0622_),
    .Y(_0623_));
 sg13g2_o21ai_1 _2985_ (.B1(_0588_),
    .Y(_0624_),
    .A1(_0593_),
    .A2(_0623_));
 sg13g2_nor2_1 _2986_ (.A(\pym[11] ),
    .B(\pym[10] ),
    .Y(_0625_));
 sg13g2_nor3_1 _2987_ (.A(\py[9] ),
    .B(\py[8] ),
    .C(net393),
    .Y(_0626_));
 sg13g2_nand3_1 _2988_ (.B(_0625_),
    .C(_0626_),
    .A(_0624_),
    .Y(_0627_));
 sg13g2_a21oi_2 _2989_ (.B1(_0627_),
    .Y(_0628_),
    .A2(_0587_),
    .A1(_1209_));
 sg13g2_nor2b_1 _2990_ (.A(net235),
    .B_N(_0628_),
    .Y(_0629_));
 sg13g2_o21ai_1 _2991_ (.B1(_0574_),
    .Y(_0630_),
    .A1(_0044_),
    .A2(_0628_));
 sg13g2_o21ai_1 _2992_ (.B1(_0582_),
    .Y(_0071_),
    .A1(_0629_),
    .A2(_0630_));
 sg13g2_nor2_1 _2993_ (.A(net473),
    .B(net296),
    .Y(_0631_));
 sg13g2_xor2_1 _2994_ (.B(net347),
    .A(net345),
    .X(_0632_));
 sg13g2_o21ai_1 _2995_ (.B1(net296),
    .Y(_0633_),
    .A1(_0610_),
    .A2(_0628_));
 sg13g2_a21oi_1 _2996_ (.A1(_0628_),
    .A2(_0632_),
    .Y(_0634_),
    .B1(_0633_));
 sg13g2_nor3_1 _2997_ (.A(net351),
    .B(_0631_),
    .C(_0634_),
    .Y(_0072_));
 sg13g2_nor2_1 _2998_ (.A(net353),
    .B(net296),
    .Y(_0635_));
 sg13g2_nand2_2 _2999_ (.Y(_0636_),
    .A(net360),
    .B(net294));
 sg13g2_xnor2_1 _3000_ (.Y(_0637_),
    .A(_1211_),
    .B(_0583_));
 sg13g2_nand2b_1 _3001_ (.Y(_0638_),
    .B(_0637_),
    .A_N(_0628_));
 sg13g2_nor2_2 _3002_ (.A(net351),
    .B(net294),
    .Y(_0639_));
 sg13g2_nand2_2 _3003_ (.Y(_0640_),
    .A(net361),
    .B(_0574_));
 sg13g2_nand2b_1 _3004_ (.Y(_0641_),
    .B(_0639_),
    .A_N(_0628_));
 sg13g2_nand4_1 _3005_ (.B(net345),
    .C(net347),
    .A(\px[2] ),
    .Y(_0642_),
    .D(_0639_));
 sg13g2_and2_1 _3006_ (.A(net279),
    .B(_0642_),
    .X(_0643_));
 sg13g2_a21o_1 _3007_ (.A2(net347),
    .A1(net345),
    .B1(\px[2] ),
    .X(_0644_));
 sg13g2_o21ai_1 _3008_ (.B1(_0643_),
    .Y(_0645_),
    .A1(_0640_),
    .A2(_0644_));
 sg13g2_nand3b_1 _3009_ (.B(_0580_),
    .C(net361),
    .Y(_0646_),
    .A_N(_0628_));
 sg13g2_nand2_2 _3010_ (.Y(_0647_),
    .A(net357),
    .B(net296));
 sg13g2_a22oi_1 _3011_ (.Y(_0073_),
    .B1(_0638_),
    .B2(_0645_),
    .A2(net290),
    .A1(_1211_));
 sg13g2_nand2_1 _3012_ (.Y(_0648_),
    .A(net433),
    .B(net290));
 sg13g2_xor2_1 _3013_ (.B(_0584_),
    .A(net433),
    .X(_0649_));
 sg13g2_nor2_1 _3014_ (.A(_0628_),
    .B(_0649_),
    .Y(_0650_));
 sg13g2_o21ai_1 _3015_ (.B1(_0648_),
    .Y(_0074_),
    .A1(_0643_),
    .A2(_0650_));
 sg13g2_nor2_1 _3016_ (.A(_0614_),
    .B(net279),
    .Y(_0651_));
 sg13g2_a21oi_1 _3017_ (.A1(_1210_),
    .A2(net290),
    .Y(_0075_),
    .B1(_0651_));
 sg13g2_nand2_1 _3018_ (.Y(_0652_),
    .A(net399),
    .B(net289));
 sg13g2_o21ai_1 _3019_ (.B1(_0652_),
    .Y(_0076_),
    .A1(_0616_),
    .A2(net279));
 sg13g2_nand2_1 _3020_ (.Y(_0653_),
    .A(net424),
    .B(net289));
 sg13g2_o21ai_1 _3021_ (.B1(_0653_),
    .Y(_0077_),
    .A1(_0590_),
    .A2(net280));
 sg13g2_nand2_1 _3022_ (.Y(_0654_),
    .A(net349),
    .B(net288));
 sg13g2_xor2_1 _3023_ (.B(_0587_),
    .A(net393),
    .X(_0655_));
 sg13g2_o21ai_1 _3024_ (.B1(_0654_),
    .Y(_0078_),
    .A1(net280),
    .A2(_0655_));
 sg13g2_a22oi_1 _3025_ (.Y(_0656_),
    .B1(_0639_),
    .B2(net228),
    .A2(net287),
    .A1(\pxm[0] ));
 sg13g2_inv_1 _3026_ (.Y(_0079_),
    .A(net229));
 sg13g2_nand2_1 _3027_ (.Y(_0657_),
    .A(net250),
    .B(net287));
 sg13g2_nor2b_1 _3028_ (.A(net334),
    .B_N(\pxm[1] ),
    .Y(_0658_));
 sg13g2_nand2b_1 _3029_ (.Y(_0659_),
    .B(net334),
    .A_N(\pxm[1] ));
 sg13g2_nand2b_1 _3030_ (.Y(_0660_),
    .B(_0659_),
    .A_N(_0658_));
 sg13g2_xnor2_1 _3031_ (.Y(_0661_),
    .A(net228),
    .B(_0660_));
 sg13g2_o21ai_1 _3032_ (.B1(_0657_),
    .Y(_0080_),
    .A1(_0640_),
    .A2(_0661_));
 sg13g2_nand2_1 _3033_ (.Y(_0662_),
    .A(net347),
    .B(net287));
 sg13g2_nand2_1 _3034_ (.Y(_0663_),
    .A(_1201_),
    .B(net347));
 sg13g2_xor2_1 _3035_ (.B(net347),
    .A(net334),
    .X(_0664_));
 sg13g2_o21ai_1 _3036_ (.B1(_0659_),
    .Y(_0665_),
    .A1(\pxm[0] ),
    .A2(_0658_));
 sg13g2_xnor2_1 _3037_ (.Y(_0666_),
    .A(_0664_),
    .B(_0665_));
 sg13g2_o21ai_1 _3038_ (.B1(_0662_),
    .Y(_0081_),
    .A1(_0640_),
    .A2(_0666_));
 sg13g2_nand2_1 _3039_ (.Y(_0667_),
    .A(net345),
    .B(net287));
 sg13g2_xor2_1 _3040_ (.B(net345),
    .A(net334),
    .X(_0668_));
 sg13g2_o21ai_1 _3041_ (.B1(_0663_),
    .Y(_0669_),
    .A1(_0664_),
    .A2(_0665_));
 sg13g2_xnor2_1 _3042_ (.Y(_0670_),
    .A(_0668_),
    .B(_0669_));
 sg13g2_o21ai_1 _3043_ (.B1(_0667_),
    .Y(_0082_),
    .A1(_0640_),
    .A2(_0670_));
 sg13g2_nand2_1 _3044_ (.Y(_0671_),
    .A(net474),
    .B(net287));
 sg13g2_xor2_1 _3045_ (.B(\px[2] ),
    .A(net334),
    .X(_0672_));
 sg13g2_o21ai_1 _3046_ (.B1(net345),
    .Y(_0673_),
    .A1(net334),
    .A2(net347));
 sg13g2_o21ai_1 _3047_ (.B1(_0673_),
    .Y(_0674_),
    .A1(_0664_),
    .A2(_0665_));
 sg13g2_o21ai_1 _3048_ (.B1(_0674_),
    .Y(_0675_),
    .A1(net334),
    .A2(net345));
 sg13g2_nor2_1 _3049_ (.A(_0672_),
    .B(_0675_),
    .Y(_0676_));
 sg13g2_xnor2_1 _3050_ (.Y(_0677_),
    .A(_0672_),
    .B(_0675_));
 sg13g2_o21ai_1 _3051_ (.B1(_0671_),
    .Y(_0083_),
    .A1(_0640_),
    .A2(_0677_));
 sg13g2_xor2_1 _3052_ (.B(\px[3] ),
    .A(net335),
    .X(_0678_));
 sg13g2_a21oi_1 _3053_ (.A1(_1201_),
    .A2(\px[2] ),
    .Y(_0679_),
    .B1(_0676_));
 sg13g2_a21oi_1 _3054_ (.A1(_0678_),
    .A2(_0679_),
    .Y(_0680_),
    .B1(_0640_));
 sg13g2_o21ai_1 _3055_ (.B1(_0680_),
    .Y(_0681_),
    .A1(_0678_),
    .A2(_0679_));
 sg13g2_o21ai_1 _3056_ (.B1(_0681_),
    .Y(_0084_),
    .A1(_1208_),
    .A2(_0636_));
 sg13g2_xor2_1 _3057_ (.B(\px[4] ),
    .A(net336),
    .X(_0682_));
 sg13g2_or3_1 _3058_ (.A(_0672_),
    .B(_0675_),
    .C(_0678_),
    .X(_0683_));
 sg13g2_nor2_1 _3059_ (.A(\px[3] ),
    .B(\px[2] ),
    .Y(_0684_));
 sg13g2_or2_1 _3060_ (.X(_0685_),
    .B(_0684_),
    .A(net335));
 sg13g2_and3_1 _3061_ (.X(_0686_),
    .A(_0682_),
    .B(_0683_),
    .C(_0685_));
 sg13g2_a21oi_1 _3062_ (.A1(_0683_),
    .A2(_0685_),
    .Y(_0687_),
    .B1(_0682_));
 sg13g2_or3_1 _3063_ (.A(_0647_),
    .B(_0686_),
    .C(_0687_),
    .X(_0688_));
 sg13g2_o21ai_1 _3064_ (.B1(_0688_),
    .Y(_0085_),
    .A1(_1207_),
    .A2(_0636_));
 sg13g2_xor2_1 _3065_ (.B(net344),
    .A(net335),
    .X(_0689_));
 sg13g2_a21oi_1 _3066_ (.A1(_1201_),
    .A2(\px[4] ),
    .Y(_0690_),
    .B1(_0687_));
 sg13g2_a21oi_1 _3067_ (.A1(_0689_),
    .A2(_0690_),
    .Y(_0691_),
    .B1(_0640_));
 sg13g2_o21ai_1 _3068_ (.B1(_0691_),
    .Y(_0692_),
    .A1(_0689_),
    .A2(_0690_));
 sg13g2_o21ai_1 _3069_ (.B1(_0692_),
    .Y(_0086_),
    .A1(_1206_),
    .A2(_0636_));
 sg13g2_xnor2_1 _3070_ (.Y(_0693_),
    .A(net334),
    .B(net343));
 sg13g2_nor3_1 _3071_ (.A(_0682_),
    .B(_0683_),
    .C(_0689_),
    .Y(_0694_));
 sg13g2_o21ai_1 _3072_ (.B1(_1201_),
    .Y(_0695_),
    .A1(net344),
    .A2(\px[4] ));
 sg13g2_nand2_1 _3073_ (.Y(_0696_),
    .A(_0685_),
    .B(_0695_));
 sg13g2_nor2_1 _3074_ (.A(_0694_),
    .B(_0696_),
    .Y(_0697_));
 sg13g2_nor3_1 _3075_ (.A(_0693_),
    .B(_0694_),
    .C(_0696_),
    .Y(_0698_));
 sg13g2_nor2b_2 _3076_ (.A(_0697_),
    .B_N(_0693_),
    .Y(_0699_));
 sg13g2_nor3_1 _3077_ (.A(_0647_),
    .B(_0698_),
    .C(_0699_),
    .Y(_0700_));
 sg13g2_a21o_1 _3078_ (.A2(net287),
    .A1(net343),
    .B1(_0700_),
    .X(_0087_));
 sg13g2_nand2_1 _3079_ (.Y(_0701_),
    .A(net342),
    .B(net288));
 sg13g2_nand2b_1 _3080_ (.Y(_0702_),
    .B(net335),
    .A_N(net342));
 sg13g2_nor2b_1 _3081_ (.A(net335),
    .B_N(net342),
    .Y(_0703_));
 sg13g2_xor2_1 _3082_ (.B(net342),
    .A(net336),
    .X(_0704_));
 sg13g2_a21oi_1 _3083_ (.A1(_1201_),
    .A2(net343),
    .Y(_0705_),
    .B1(_0699_));
 sg13g2_xnor2_1 _3084_ (.Y(_0706_),
    .A(_0704_),
    .B(_0705_));
 sg13g2_o21ai_1 _3085_ (.B1(_0701_),
    .Y(_0088_),
    .A1(_0647_),
    .A2(_0706_));
 sg13g2_a221oi_1 _3086_ (.B2(_0702_),
    .C1(_0703_),
    .B1(_0699_),
    .A1(_1201_),
    .Y(_0707_),
    .A2(net343));
 sg13g2_nor2_1 _3087_ (.A(net335),
    .B(_1204_),
    .Y(_0708_));
 sg13g2_xor2_1 _3088_ (.B(\px[8] ),
    .A(net335),
    .X(_0709_));
 sg13g2_a21oi_1 _3089_ (.A1(_0707_),
    .A2(_0709_),
    .Y(_0710_),
    .B1(_0640_));
 sg13g2_o21ai_1 _3090_ (.B1(_0710_),
    .Y(_0711_),
    .A1(_0707_),
    .A2(_0709_));
 sg13g2_o21ai_1 _3091_ (.B1(_0711_),
    .Y(_0089_),
    .A1(_1204_),
    .A2(_0636_));
 sg13g2_a21oi_1 _3092_ (.A1(net342),
    .A2(_0699_),
    .Y(_0712_),
    .B1(_1201_));
 sg13g2_o21ai_1 _3093_ (.B1(_0580_),
    .Y(_0713_),
    .A1(\px[8] ),
    .A2(_0707_));
 sg13g2_nor3_1 _3094_ (.A(_0708_),
    .B(_0712_),
    .C(_0713_),
    .Y(_0714_));
 sg13g2_o21ai_1 _3095_ (.B1(net357),
    .Y(_0715_),
    .A1(net377),
    .A2(_0714_));
 sg13g2_a21oi_1 _3096_ (.A1(net377),
    .A2(_0714_),
    .Y(_0090_),
    .B1(_0715_));
 sg13g2_nand2_1 _3097_ (.Y(_0716_),
    .A(net341),
    .B(net290));
 sg13g2_o21ai_1 _3098_ (.B1(_0716_),
    .Y(_0091_),
    .A1(_0611_),
    .A2(net280));
 sg13g2_nand2_1 _3099_ (.Y(_0717_),
    .A(net237),
    .B(net290));
 sg13g2_xnor2_1 _3100_ (.Y(_0718_),
    .A(_0603_),
    .B(_0604_));
 sg13g2_o21ai_1 _3101_ (.B1(_0717_),
    .Y(_0092_),
    .A1(net279),
    .A2(_0718_));
 sg13g2_nand2_1 _3102_ (.Y(_0719_),
    .A(net492),
    .B(net290));
 sg13g2_nand2_1 _3103_ (.Y(_0720_),
    .A(_0596_),
    .B(_0605_));
 sg13g2_xnor2_1 _3104_ (.Y(_0721_),
    .A(_0596_),
    .B(_0605_));
 sg13g2_o21ai_1 _3105_ (.B1(_0719_),
    .Y(_0093_),
    .A1(net279),
    .A2(_0721_));
 sg13g2_nand2_1 _3106_ (.Y(_0722_),
    .A(net514),
    .B(net290));
 sg13g2_nand2_1 _3107_ (.Y(_0723_),
    .A(_0595_),
    .B(_0720_));
 sg13g2_xnor2_1 _3108_ (.Y(_0724_),
    .A(_0599_),
    .B(_0723_));
 sg13g2_o21ai_1 _3109_ (.B1(_0722_),
    .Y(_0094_),
    .A1(net279),
    .A2(_0724_));
 sg13g2_nand2_1 _3110_ (.Y(_0725_),
    .A(net339),
    .B(net290));
 sg13g2_o21ai_1 _3111_ (.B1(_0725_),
    .Y(_0095_),
    .A1(_0609_),
    .A2(net279));
 sg13g2_nand2_1 _3112_ (.Y(_0726_),
    .A(net500),
    .B(net293));
 sg13g2_a21oi_1 _3113_ (.A1(net339),
    .A2(\ydelta[4] ),
    .Y(_0727_),
    .B1(_0608_));
 sg13g2_xor2_1 _3114_ (.B(\ydelta[5] ),
    .A(\py[5] ),
    .X(_0728_));
 sg13g2_xor2_1 _3115_ (.B(_0728_),
    .A(_0727_),
    .X(_0729_));
 sg13g2_o21ai_1 _3116_ (.B1(_0726_),
    .Y(_0096_),
    .A1(net279),
    .A2(_0729_));
 sg13g2_nand2_1 _3117_ (.Y(_0730_),
    .A(net504),
    .B(net289));
 sg13g2_nor2_1 _3118_ (.A(\py[6] ),
    .B(\ydelta[6] ),
    .Y(_0731_));
 sg13g2_nand2_1 _3119_ (.Y(_0732_),
    .A(\py[6] ),
    .B(\ydelta[6] ));
 sg13g2_nand2b_1 _3120_ (.Y(_0733_),
    .B(_0732_),
    .A_N(_0731_));
 sg13g2_nand2_1 _3121_ (.Y(_0734_),
    .A(_0608_),
    .B(_0728_));
 sg13g2_and3_1 _3122_ (.X(_0735_),
    .A(net339),
    .B(\ydelta[4] ),
    .C(_0728_));
 sg13g2_a21oi_1 _3123_ (.A1(\py[5] ),
    .A2(\ydelta[5] ),
    .Y(_0736_),
    .B1(_0735_));
 sg13g2_and2_1 _3124_ (.A(_0734_),
    .B(_0736_),
    .X(_0737_));
 sg13g2_xnor2_1 _3125_ (.Y(_0738_),
    .A(_0733_),
    .B(_0737_));
 sg13g2_o21ai_1 _3126_ (.B1(_0730_),
    .Y(_0097_),
    .A1(net280),
    .A2(_0738_));
 sg13g2_nand2_1 _3127_ (.Y(_0739_),
    .A(net463),
    .B(net288));
 sg13g2_o21ai_1 _3128_ (.B1(_0732_),
    .Y(_0740_),
    .A1(_0731_),
    .A2(_0737_));
 sg13g2_xnor2_1 _3129_ (.Y(_0741_),
    .A(_0591_),
    .B(_0740_));
 sg13g2_o21ai_1 _3130_ (.B1(_0739_),
    .Y(_0098_),
    .A1(net280),
    .A2(_0741_));
 sg13g2_nand2_1 _3131_ (.Y(_0742_),
    .A(net469),
    .B(net287));
 sg13g2_and2_1 _3132_ (.A(\py[8] ),
    .B(net348),
    .X(_0743_));
 sg13g2_xor2_1 _3133_ (.B(net348),
    .A(\py[8] ),
    .X(_0744_));
 sg13g2_nor3_1 _3134_ (.A(_0593_),
    .B(_0618_),
    .C(_0734_),
    .Y(_0745_));
 sg13g2_a22oi_1 _3135_ (.Y(_0746_),
    .B1(\ydelta[6] ),
    .B2(\py[6] ),
    .A2(net349),
    .A1(\py[7] ));
 sg13g2_o21ai_1 _3136_ (.B1(_0746_),
    .Y(_0747_),
    .A1(_0731_),
    .A2(_0736_));
 sg13g2_o21ai_1 _3137_ (.B1(_0747_),
    .Y(_0748_),
    .A1(\py[7] ),
    .A2(net349));
 sg13g2_nand2b_1 _3138_ (.Y(_0749_),
    .B(_0748_),
    .A_N(_0745_));
 sg13g2_xnor2_1 _3139_ (.Y(_0750_),
    .A(_0744_),
    .B(_0749_));
 sg13g2_o21ai_1 _3140_ (.B1(_0742_),
    .Y(_0099_),
    .A1(net280),
    .A2(_0750_));
 sg13g2_nand2_1 _3141_ (.Y(_0751_),
    .A(net483),
    .B(net287));
 sg13g2_xor2_1 _3142_ (.B(net348),
    .A(\py[9] ),
    .X(_0752_));
 sg13g2_a21o_1 _3143_ (.A2(_0749_),
    .A1(_0744_),
    .B1(_0743_),
    .X(_0753_));
 sg13g2_xnor2_1 _3144_ (.Y(_0754_),
    .A(_0752_),
    .B(_0753_));
 sg13g2_o21ai_1 _3145_ (.B1(_0751_),
    .Y(_0100_),
    .A1(net280),
    .A2(_0754_));
 sg13g2_nand2_1 _3146_ (.Y(_0755_),
    .A(net382),
    .B(net289));
 sg13g2_xnor2_1 _3147_ (.Y(_0756_),
    .A(\pym[10] ),
    .B(net348));
 sg13g2_a21o_1 _3148_ (.A2(net348),
    .A1(\py[9] ),
    .B1(_0753_),
    .X(_0757_));
 sg13g2_o21ai_1 _3149_ (.B1(_0757_),
    .Y(_0758_),
    .A1(\py[9] ),
    .A2(net348));
 sg13g2_xnor2_1 _3150_ (.Y(_0759_),
    .A(_0756_),
    .B(_0758_));
 sg13g2_o21ai_1 _3151_ (.B1(_0755_),
    .Y(_0101_),
    .A1(_0646_),
    .A2(_0759_));
 sg13g2_nand2_1 _3152_ (.Y(_0760_),
    .A(net369),
    .B(net289));
 sg13g2_nand2_1 _3153_ (.Y(_0761_),
    .A(net546),
    .B(net348));
 sg13g2_o21ai_1 _3154_ (.B1(_0761_),
    .Y(_0762_),
    .A1(_0756_),
    .A2(_0758_));
 sg13g2_xor2_1 _3155_ (.B(net348),
    .A(net369),
    .X(_0763_));
 sg13g2_xnor2_1 _3156_ (.Y(_0764_),
    .A(_0762_),
    .B(_0763_));
 sg13g2_o21ai_1 _3157_ (.B1(_0760_),
    .Y(_0102_),
    .A1(_0646_),
    .A2(_0764_));
 sg13g2_nor3_1 _3158_ (.A(\product_comp[5] ),
    .B(\product_comp[4] ),
    .C(\product_comp[3] ),
    .Y(_0765_));
 sg13g2_nand2_1 _3159_ (.Y(_0766_),
    .A(\product_comp[7] ),
    .B(\product_comp[6] ));
 sg13g2_nor2_1 _3160_ (.A(_0765_),
    .B(_0766_),
    .Y(_0767_));
 sg13g2_nor4_2 _3161_ (.A(net387),
    .B(net411),
    .C(\product_comp[8] ),
    .Y(_0768_),
    .D(_0767_));
 sg13g2_o21ai_1 _3162_ (.B1(net337),
    .Y(_0769_),
    .A1(net294),
    .A2(_0768_));
 sg13g2_o21ai_1 _3163_ (.B1(\product_comp[4] ),
    .Y(_0770_),
    .A1(\product_comp[3] ),
    .A2(\product_comp[2] ));
 sg13g2_nor4_1 _3164_ (.A(\product_comp[9] ),
    .B(\product_comp[8] ),
    .C(\product_comp[7] ),
    .D(\product_comp[6] ),
    .Y(_0771_));
 sg13g2_nor2_1 _3165_ (.A(\product_comp[5] ),
    .B(net337),
    .Y(_0772_));
 sg13g2_nand4_1 _3166_ (.B(_0770_),
    .C(_0771_),
    .A(net453),
    .Y(_0773_),
    .D(_0772_));
 sg13g2_o21ai_1 _3167_ (.B1(net360),
    .Y(_0774_),
    .A1(net294),
    .A2(_0773_));
 sg13g2_nand2b_1 _3168_ (.Y(_0103_),
    .B(_0769_),
    .A_N(_0774_));
 sg13g2_nor4_1 _3169_ (.A(net343),
    .B(net344),
    .C(net345),
    .D(net347),
    .Y(_0775_));
 sg13g2_nor3_1 _3170_ (.A(\px[8] ),
    .B(net342),
    .C(\px[4] ),
    .Y(_0776_));
 sg13g2_nand3_1 _3171_ (.B(_0775_),
    .C(_0776_),
    .A(_0684_),
    .Y(_0777_));
 sg13g2_a21o_1 _3172_ (.A2(_0777_),
    .A1(_1201_),
    .B1(net377),
    .X(_0778_));
 sg13g2_nand3b_1 _3173_ (.B(_1340_),
    .C(_1204_),
    .Y(_0779_),
    .A_N(_0702_));
 sg13g2_nand3_1 _3174_ (.B(_0778_),
    .C(_0779_),
    .A(net357),
    .Y(_0104_));
 sg13g2_nor3_1 _3175_ (.A(_0565_),
    .B(_0568_),
    .C(_0571_),
    .Y(_0105_));
 sg13g2_nor2_1 _3176_ (.A(\h[0] ),
    .B(net316),
    .Y(_0780_));
 sg13g2_or2_1 _3177_ (.X(_0781_),
    .B(net316),
    .A(\h[0] ));
 sg13g2_nand2b_1 _3178_ (.Y(_0782_),
    .B(_0355_),
    .A_N(net354));
 sg13g2_nor4_1 _3179_ (.A(\h[8] ),
    .B(_1217_),
    .C(_0781_),
    .D(_0782_),
    .Y(_0783_));
 sg13g2_xnor2_1 _3180_ (.Y(_0784_),
    .A(net314),
    .B(_0355_));
 sg13g2_nand3b_1 _3181_ (.B(\h[3] ),
    .C(net315),
    .Y(_0785_),
    .A_N(net306));
 sg13g2_nand4_1 _3182_ (.B(net311),
    .C(net314),
    .A(net309),
    .Y(_0786_),
    .D(net354));
 sg13g2_nor4_1 _3183_ (.A(_0304_),
    .B(_0781_),
    .C(_0785_),
    .D(_0786_),
    .Y(_0787_));
 sg13g2_nor2_1 _3184_ (.A(net309),
    .B(\h[5] ),
    .Y(_0788_));
 sg13g2_and4_1 _3185_ (.A(net306),
    .B(_0783_),
    .C(_0784_),
    .D(_0788_),
    .X(_0789_));
 sg13g2_nor3_1 _3186_ (.A(net420),
    .B(_0787_),
    .C(_0789_),
    .Y(_0790_));
 sg13g2_nand4_1 _3187_ (.B(net313),
    .C(_1245_),
    .A(net311),
    .Y(_0791_),
    .D(_0783_));
 sg13g2_nand4_1 _3188_ (.B(net311),
    .C(net316),
    .A(net306),
    .Y(_0792_),
    .D(net354));
 sg13g2_or4_1 _3189_ (.A(net310),
    .B(\h[0] ),
    .C(_0304_),
    .D(_0356_),
    .X(_0793_));
 sg13g2_o21ai_1 _3190_ (.B1(_0791_),
    .Y(_0794_),
    .A1(_0792_),
    .A2(_0793_));
 sg13g2_nor3_1 _3191_ (.A(net350),
    .B(net421),
    .C(_0794_),
    .Y(_0106_));
 sg13g2_nor2_1 _3192_ (.A(net332),
    .B(hmax),
    .Y(_0795_));
 sg13g2_and2_1 _3193_ (.A(net332),
    .B(hmax),
    .X(_0796_));
 sg13g2_nor3_1 _3194_ (.A(_0636_),
    .B(_0795_),
    .C(_0796_),
    .Y(_0107_));
 sg13g2_o21ai_1 _3195_ (.B1(net364),
    .Y(_0797_),
    .A1(net331),
    .A2(_0796_));
 sg13g2_nand2_2 _3196_ (.Y(_0798_),
    .A(net331),
    .B(_0796_));
 sg13g2_nor2b_1 _3197_ (.A(_0797_),
    .B_N(_0798_),
    .Y(_0108_));
 sg13g2_a21oi_1 _3198_ (.A1(net331),
    .A2(_0796_),
    .Y(_0799_),
    .B1(net329));
 sg13g2_nor2_1 _3199_ (.A(_1286_),
    .B(_0578_),
    .Y(_0800_));
 sg13g2_nor3_1 _3200_ (.A(_0636_),
    .B(net510),
    .C(_0800_),
    .Y(_0109_));
 sg13g2_nor2_1 _3201_ (.A(net405),
    .B(_0798_),
    .Y(_0801_));
 sg13g2_o21ai_1 _3202_ (.B1(net291),
    .Y(_0802_),
    .A1(net327),
    .A2(_0801_));
 sg13g2_a21oi_1 _3203_ (.A1(net327),
    .A2(_0801_),
    .Y(_0110_),
    .B1(_0802_));
 sg13g2_nor2_1 _3204_ (.A(_1252_),
    .B(_0798_),
    .Y(_0803_));
 sg13g2_xnor2_1 _3205_ (.Y(_0804_),
    .A(net326),
    .B(_0803_));
 sg13g2_nor2_1 _3206_ (.A(net353),
    .B(_0804_),
    .Y(_0111_));
 sg13g2_nor3_1 _3207_ (.A(_0025_),
    .B(_1252_),
    .C(_0798_),
    .Y(_0805_));
 sg13g2_o21ai_1 _3208_ (.B1(net291),
    .Y(_0806_),
    .A1(net324),
    .A2(_0805_));
 sg13g2_a21oi_1 _3209_ (.A1(net324),
    .A2(_0805_),
    .Y(_0112_),
    .B1(_0806_));
 sg13g2_nand3_1 _3210_ (.B(net326),
    .C(_0803_),
    .A(net324),
    .Y(_0807_));
 sg13g2_xor2_1 _3211_ (.B(_0807_),
    .A(net323),
    .X(_0808_));
 sg13g2_nor2_1 _3212_ (.A(net351),
    .B(_0808_),
    .Y(_0113_));
 sg13g2_nor2_2 _3213_ (.A(net480),
    .B(_0807_),
    .Y(_0809_));
 sg13g2_o21ai_1 _3214_ (.B1(net291),
    .Y(_0810_),
    .A1(net320),
    .A2(_0809_));
 sg13g2_a21oi_1 _3215_ (.A1(net320),
    .A2(_0809_),
    .Y(_0114_),
    .B1(_0810_));
 sg13g2_nor2_1 _3216_ (.A(_1264_),
    .B(_0807_),
    .Y(_0811_));
 sg13g2_xnor2_1 _3217_ (.Y(_0812_),
    .A(net319),
    .B(_0811_));
 sg13g2_nor2_1 _3218_ (.A(_0636_),
    .B(_0812_),
    .Y(_0115_));
 sg13g2_nor3_1 _3219_ (.A(_0023_),
    .B(_1264_),
    .C(_0807_),
    .Y(_0813_));
 sg13g2_o21ai_1 _3220_ (.B1(net291),
    .Y(_0814_),
    .A1(net318),
    .A2(_0813_));
 sg13g2_a21oi_1 _3221_ (.A1(net318),
    .A2(_0813_),
    .Y(_0116_),
    .B1(_0814_));
 sg13g2_o21ai_1 _3222_ (.B1(net364),
    .Y(_0815_),
    .A1(_1255_),
    .A2(_1267_));
 sg13g2_nand2b_1 _3223_ (.Y(_0816_),
    .B(net327),
    .A_N(net329));
 sg13g2_nor4_1 _3224_ (.A(_1200_),
    .B(net332),
    .C(_1267_),
    .D(_0816_),
    .Y(_0817_));
 sg13g2_nor3_1 _3225_ (.A(net355),
    .B(_0815_),
    .C(_0817_),
    .Y(_0818_));
 sg13g2_nand4_1 _3226_ (.B(net330),
    .C(_1200_),
    .A(_1199_),
    .Y(_0819_),
    .D(net333));
 sg13g2_nor2_1 _3227_ (.A(_1254_),
    .B(_0816_),
    .Y(_0820_));
 sg13g2_o21ai_1 _3228_ (.B1(_0819_),
    .Y(_0821_),
    .A1(_1254_),
    .A2(_0816_));
 sg13g2_nand4_1 _3229_ (.B(_1265_),
    .C(_1277_),
    .A(net317),
    .Y(_0822_),
    .D(_0821_));
 sg13g2_nand3_1 _3230_ (.B(net364),
    .C(_0822_),
    .A(net355),
    .Y(_0823_));
 sg13g2_nor2b_1 _3231_ (.A(_0818_),
    .B_N(_0823_),
    .Y(_0824_));
 sg13g2_nand4_1 _3232_ (.B(_1265_),
    .C(_1277_),
    .A(net317),
    .Y(_0825_),
    .D(_0820_));
 sg13g2_nand2b_1 _3233_ (.Y(_0826_),
    .B(_0825_),
    .A_N(_0815_));
 sg13g2_nor2_1 _3234_ (.A(net253),
    .B(_0824_),
    .Y(_0827_));
 sg13g2_a21oi_1 _3235_ (.A1(_0824_),
    .A2(_0826_),
    .Y(_0117_),
    .B1(_0827_));
 sg13g2_nand2_2 _3236_ (.Y(_0118_),
    .A(_0364_),
    .B(_0784_));
 sg13g2_xor2_1 _3237_ (.B(_0356_),
    .A(net312),
    .X(_0828_));
 sg13g2_nand2_2 _3238_ (.Y(_0119_),
    .A(_0364_),
    .B(_0828_));
 sg13g2_nor3_1 _3239_ (.A(_0555_),
    .B(_0561_),
    .C(_0563_),
    .Y(_0120_));
 sg13g2_nand2_2 _3240_ (.Y(_0829_),
    .A(net357),
    .B(_0578_));
 sg13g2_and3_1 _3241_ (.X(_0121_),
    .A(net357),
    .B(net220),
    .C(_0578_));
 sg13g2_nor3_1 _3242_ (.A(net351),
    .B(_1236_),
    .C(_0780_),
    .Y(_0122_));
 sg13g2_and2_1 _3243_ (.A(net315),
    .B(_1236_),
    .X(_0830_));
 sg13g2_nor2_1 _3244_ (.A(net315),
    .B(_1236_),
    .Y(_0831_));
 sg13g2_nor3_1 _3245_ (.A(_0829_),
    .B(_0830_),
    .C(_0831_),
    .Y(_0123_));
 sg13g2_and2_1 _3246_ (.A(\h[3] ),
    .B(_0830_),
    .X(_0832_));
 sg13g2_nor2_1 _3247_ (.A(net508),
    .B(_0830_),
    .Y(_0833_));
 sg13g2_nor3_1 _3248_ (.A(_0829_),
    .B(_0832_),
    .C(_0833_),
    .Y(_0124_));
 sg13g2_xnor2_1 _3249_ (.Y(_0834_),
    .A(net313),
    .B(_0832_));
 sg13g2_nor2_1 _3250_ (.A(_0829_),
    .B(_0834_),
    .Y(_0125_));
 sg13g2_nand3_1 _3251_ (.B(net313),
    .C(_0832_),
    .A(net312),
    .Y(_0835_));
 sg13g2_inv_1 _3252_ (.Y(_0836_),
    .A(_0835_));
 sg13g2_a21oi_1 _3253_ (.A1(net313),
    .A2(_0832_),
    .Y(_0837_),
    .B1(net312));
 sg13g2_nor3_1 _3254_ (.A(_0829_),
    .B(_0836_),
    .C(_0837_),
    .Y(_0126_));
 sg13g2_xnor2_1 _3255_ (.Y(_0838_),
    .A(_1213_),
    .B(_0835_));
 sg13g2_nor2_1 _3256_ (.A(_0829_),
    .B(_0838_),
    .Y(_0127_));
 sg13g2_nor2_1 _3257_ (.A(net481),
    .B(_0835_),
    .Y(_0839_));
 sg13g2_xnor2_1 _3258_ (.Y(_0840_),
    .A(net308),
    .B(_0839_));
 sg13g2_nor2_1 _3259_ (.A(_0829_),
    .B(net482),
    .Y(_0128_));
 sg13g2_nor2_1 _3260_ (.A(_1244_),
    .B(_0835_),
    .Y(_0841_));
 sg13g2_xnor2_1 _3261_ (.Y(_0842_),
    .A(net521),
    .B(_0841_));
 sg13g2_nor2_1 _3262_ (.A(_0829_),
    .B(_0842_),
    .Y(_0129_));
 sg13g2_nor3_1 _3263_ (.A(net536),
    .B(_1244_),
    .C(_0835_),
    .Y(_0843_));
 sg13g2_xnor2_1 _3264_ (.Y(_0844_),
    .A(net305),
    .B(_0843_));
 sg13g2_nor2_1 _3265_ (.A(_0829_),
    .B(_0844_),
    .Y(_0130_));
 sg13g2_nor3_1 _3266_ (.A(\matt_venn_clock.pulse_hrs.count[3] ),
    .B(\matt_venn_clock.pulse_hrs.count[1] ),
    .C(\matt_venn_clock.pulse_hrs.count[0] ),
    .Y(_0845_));
 sg13g2_nand3b_1 _3267_ (.B(_0056_),
    .C(_0845_),
    .Y(_0846_),
    .A_N(\matt_venn_clock.pulse_hrs.count[2] ));
 sg13g2_nor3_1 _3268_ (.A(\matt_venn_clock.pulse_hrs.comp[4] ),
    .B(\matt_venn_clock.pulse_hrs.comp[3] ),
    .C(\matt_venn_clock.pulse_hrs.comp[2] ),
    .Y(_0847_));
 sg13g2_or2_1 _3269_ (.X(_0848_),
    .B(_0847_),
    .A(_0846_));
 sg13g2_nand2_2 _3270_ (.Y(_0849_),
    .A(net1),
    .B(_0574_));
 sg13g2_inv_1 _3271_ (.Y(_0850_),
    .A(_0849_));
 sg13g2_nor2_1 _3272_ (.A(_0579_),
    .B(_0848_),
    .Y(_0851_));
 sg13g2_nand2_1 _3273_ (.Y(_0852_),
    .A(net1),
    .B(_0848_));
 sg13g2_o21ai_1 _3274_ (.B1(net475),
    .Y(_0853_),
    .A1(_0848_),
    .A2(_0849_));
 sg13g2_nand3_1 _3275_ (.B(_0581_),
    .C(_0852_),
    .A(_1196_),
    .Y(_0854_));
 sg13g2_nand3_1 _3276_ (.B(_0853_),
    .C(_0854_),
    .A(net366),
    .Y(_0131_));
 sg13g2_nand2_1 _3277_ (.Y(_0855_),
    .A(net456),
    .B(_0854_));
 sg13g2_o21ai_1 _3278_ (.B1(net366),
    .Y(_0856_),
    .A1(net1),
    .A2(net294));
 sg13g2_or2_1 _3279_ (.X(_0857_),
    .B(_0854_),
    .A(net456));
 sg13g2_nand3b_1 _3280_ (.B(_0857_),
    .C(_0855_),
    .Y(_0132_),
    .A_N(_0856_));
 sg13g2_nand2_1 _3281_ (.Y(_0858_),
    .A(net464),
    .B(_0857_));
 sg13g2_nor3_1 _3282_ (.A(\matt_venn_clock.pulse_hrs.comp[2] ),
    .B(net456),
    .C(net475),
    .Y(_0859_));
 sg13g2_a22oi_1 _3283_ (.Y(_0860_),
    .B1(_0851_),
    .B2(_0859_),
    .A2(_0580_),
    .A1(_1220_));
 sg13g2_nand3_1 _3284_ (.B(_0858_),
    .C(_0860_),
    .A(net364),
    .Y(_0133_));
 sg13g2_nor2_2 _3285_ (.A(_0846_),
    .B(_0849_),
    .Y(_0861_));
 sg13g2_or2_2 _3286_ (.X(_0862_),
    .B(_0849_),
    .A(_0846_));
 sg13g2_a21o_1 _3287_ (.A2(_0861_),
    .A1(_0859_),
    .B1(_1195_),
    .X(_0863_));
 sg13g2_or2_1 _3288_ (.X(_0864_),
    .B(_0860_),
    .A(net524));
 sg13g2_nand3_1 _3289_ (.B(_0863_),
    .C(_0864_),
    .A(net364),
    .Y(_0134_));
 sg13g2_nor4_1 _3290_ (.A(net418),
    .B(\matt_venn_clock.pulse_hrs.comp[3] ),
    .C(\matt_venn_clock.pulse_hrs.comp[2] ),
    .D(_0857_),
    .Y(_0865_));
 sg13g2_a21oi_1 _3291_ (.A1(net418),
    .A2(_0864_),
    .Y(_0866_),
    .B1(_0865_));
 sg13g2_nor2_1 _3292_ (.A(_0856_),
    .B(net419),
    .Y(_0135_));
 sg13g2_xor2_1 _3293_ (.B(\matt_venn_clock.pulse_hrs.comp[2] ),
    .A(\matt_venn_clock.pulse_hrs.count[2] ),
    .X(_0867_));
 sg13g2_a22oi_1 _3294_ (.Y(_0868_),
    .B1(_1196_),
    .B2(\matt_venn_clock.pulse_hrs.count[0] ),
    .A2(\matt_venn_clock.pulse_hrs.comp[3] ),
    .A1(_1193_));
 sg13g2_xnor2_1 _3295_ (.Y(_0869_),
    .A(\matt_venn_clock.pulse_hrs.count[4] ),
    .B(\matt_venn_clock.pulse_hrs.comp[4] ));
 sg13g2_xnor2_1 _3296_ (.Y(_0870_),
    .A(\matt_venn_clock.pulse_hrs.count[1] ),
    .B(\matt_venn_clock.pulse_hrs.comp[1] ));
 sg13g2_a221oi_1 _3297_ (.B2(_1194_),
    .C1(_0867_),
    .B1(\matt_venn_clock.pulse_hrs.comp[0] ),
    .A1(\matt_venn_clock.pulse_hrs.count[3] ),
    .Y(_0871_),
    .A2(_1195_));
 sg13g2_nand4_1 _3298_ (.B(_0869_),
    .C(_0870_),
    .A(_0868_),
    .Y(_0872_),
    .D(_0871_));
 sg13g2_a21oi_1 _3299_ (.A1(_0850_),
    .A2(_0872_),
    .Y(_0873_),
    .B1(net443));
 sg13g2_o21ai_1 _3300_ (.B1(net364),
    .Y(_0874_),
    .A1(_1194_),
    .A2(net294));
 sg13g2_nor2_1 _3301_ (.A(_0873_),
    .B(_0874_),
    .Y(_0136_));
 sg13g2_nand2_1 _3302_ (.Y(_0875_),
    .A(net436),
    .B(net291));
 sg13g2_xnor2_1 _3303_ (.Y(_0876_),
    .A(net436),
    .B(\matt_venn_clock.pulse_hrs.count[0] ));
 sg13g2_nand3_1 _3304_ (.B(_0850_),
    .C(_0872_),
    .A(net364),
    .Y(_0877_));
 sg13g2_o21ai_1 _3305_ (.B1(_0875_),
    .Y(_0137_),
    .A1(_0876_),
    .A2(_0877_));
 sg13g2_nand2_1 _3306_ (.Y(_0878_),
    .A(net395),
    .B(net291));
 sg13g2_nand3_1 _3307_ (.B(\matt_venn_clock.pulse_hrs.count[1] ),
    .C(\matt_venn_clock.pulse_hrs.count[0] ),
    .A(\matt_venn_clock.pulse_hrs.count[2] ),
    .Y(_0879_));
 sg13g2_a21o_1 _3308_ (.A2(\matt_venn_clock.pulse_hrs.count[0] ),
    .A1(\matt_venn_clock.pulse_hrs.count[1] ),
    .B1(net395),
    .X(_0880_));
 sg13g2_nand2_1 _3309_ (.Y(_0881_),
    .A(_0879_),
    .B(_0880_));
 sg13g2_o21ai_1 _3310_ (.B1(_0878_),
    .Y(_0138_),
    .A1(_0877_),
    .A2(_0881_));
 sg13g2_nand2_1 _3311_ (.Y(_0882_),
    .A(net269),
    .B(net291));
 sg13g2_or2_1 _3312_ (.X(_0883_),
    .B(_0879_),
    .A(_1193_));
 sg13g2_xnor2_1 _3313_ (.Y(_0884_),
    .A(_1193_),
    .B(_0879_));
 sg13g2_o21ai_1 _3314_ (.B1(_0882_),
    .Y(_0139_),
    .A1(_0877_),
    .A2(_0884_));
 sg13g2_nand2_1 _3315_ (.Y(_0885_),
    .A(net254),
    .B(net291));
 sg13g2_xnor2_1 _3316_ (.Y(_0886_),
    .A(_0056_),
    .B(_0883_));
 sg13g2_o21ai_1 _3317_ (.B1(_0885_),
    .Y(_0140_),
    .A1(_0877_),
    .A2(_0886_));
 sg13g2_nor3_2 _3318_ (.A(net414),
    .B(net545),
    .C(\matt_venn_clock.pulse_min.comp[2] ),
    .Y(_0887_));
 sg13g2_nor3_1 _3319_ (.A(\matt_venn_clock.pulse_min.count[3] ),
    .B(\matt_venn_clock.pulse_min.count[1] ),
    .C(\matt_venn_clock.pulse_min.count[0] ),
    .Y(_0888_));
 sg13g2_nand3b_1 _3320_ (.B(_0055_),
    .C(_0888_),
    .Y(_0889_),
    .A_N(\matt_venn_clock.pulse_min.count[2] ));
 sg13g2_inv_1 _3321_ (.Y(_0890_),
    .A(_0889_));
 sg13g2_nand3_1 _3322_ (.B(_0574_),
    .C(_0890_),
    .A(net2),
    .Y(_0891_));
 sg13g2_nor3_1 _3323_ (.A(_0579_),
    .B(_0887_),
    .C(_0889_),
    .Y(_0892_));
 sg13g2_o21ai_1 _3324_ (.B1(net2),
    .Y(_0893_),
    .A1(_0887_),
    .A2(_0889_));
 sg13g2_o21ai_1 _3325_ (.B1(net440),
    .Y(_0894_),
    .A1(_0887_),
    .A2(_0891_));
 sg13g2_nand3_1 _3326_ (.B(_0581_),
    .C(_0893_),
    .A(_1192_),
    .Y(_0895_));
 sg13g2_nor2_1 _3327_ (.A(net2),
    .B(_0579_),
    .Y(_0896_));
 sg13g2_nand3_1 _3328_ (.B(_0894_),
    .C(_0895_),
    .A(net365),
    .Y(_0141_));
 sg13g2_nand2_1 _3329_ (.Y(_0897_),
    .A(net397),
    .B(_0895_));
 sg13g2_o21ai_1 _3330_ (.B1(net365),
    .Y(_0898_),
    .A1(net2),
    .A2(_0575_));
 sg13g2_nand2b_1 _3331_ (.Y(_0899_),
    .B(_1191_),
    .A_N(_0895_));
 sg13g2_nand3b_1 _3332_ (.B(_0899_),
    .C(_0897_),
    .Y(_0142_),
    .A_N(_0898_));
 sg13g2_nand2_1 _3333_ (.Y(_0900_),
    .A(net462),
    .B(_0899_));
 sg13g2_nor3_1 _3334_ (.A(\matt_venn_clock.pulse_min.comp[2] ),
    .B(net397),
    .C(net440),
    .Y(_0901_));
 sg13g2_a21oi_1 _3335_ (.A1(_0892_),
    .A2(_0901_),
    .Y(_0902_),
    .B1(_0896_));
 sg13g2_nand3_1 _3336_ (.B(_0900_),
    .C(_0902_),
    .A(net365),
    .Y(_0143_));
 sg13g2_nand4_1 _3337_ (.B(net296),
    .C(_0890_),
    .A(net2),
    .Y(_0903_),
    .D(_0901_));
 sg13g2_or2_1 _3338_ (.X(_0904_),
    .B(_0902_),
    .A(net452));
 sg13g2_a21oi_1 _3339_ (.A1(net452),
    .A2(_0903_),
    .Y(_0905_),
    .B1(net352));
 sg13g2_nand2_1 _3340_ (.Y(_0144_),
    .A(_0904_),
    .B(_0905_));
 sg13g2_nand2_1 _3341_ (.Y(_0906_),
    .A(net414),
    .B(_0904_));
 sg13g2_nand4_1 _3342_ (.B(_1192_),
    .C(_0887_),
    .A(_1191_),
    .Y(_0907_),
    .D(_0896_));
 sg13g2_a21oi_1 _3343_ (.A1(_0906_),
    .A2(_0907_),
    .Y(_0145_),
    .B1(_0898_));
 sg13g2_nand2b_1 _3344_ (.Y(_0908_),
    .B(\matt_venn_clock.pulse_min.comp[2] ),
    .A_N(\matt_venn_clock.pulse_min.count[2] ));
 sg13g2_nor2_1 _3345_ (.A(\matt_venn_clock.pulse_min.count[4] ),
    .B(_1190_),
    .Y(_0909_));
 sg13g2_nor2b_1 _3346_ (.A(\matt_venn_clock.pulse_min.comp[2] ),
    .B_N(\matt_venn_clock.pulse_min.count[2] ),
    .Y(_0910_));
 sg13g2_o21ai_1 _3347_ (.B1(_0908_),
    .Y(_0911_),
    .A1(\matt_venn_clock.pulse_min.count[1] ),
    .A2(_1191_));
 sg13g2_xor2_1 _3348_ (.B(\matt_venn_clock.pulse_min.comp[3] ),
    .A(\matt_venn_clock.pulse_min.count[3] ),
    .X(_0912_));
 sg13g2_a221oi_1 _3349_ (.B2(_1189_),
    .C1(_0912_),
    .B1(\matt_venn_clock.pulse_min.comp[0] ),
    .A1(\matt_venn_clock.pulse_min.count[4] ),
    .Y(_0913_),
    .A2(_1190_));
 sg13g2_nor3_1 _3350_ (.A(_0909_),
    .B(_0910_),
    .C(_0911_),
    .Y(_0914_));
 sg13g2_a22oi_1 _3351_ (.Y(_0915_),
    .B1(_1192_),
    .B2(\matt_venn_clock.pulse_min.count[0] ),
    .A2(_1191_),
    .A1(\matt_venn_clock.pulse_min.count[1] ));
 sg13g2_nand3_1 _3352_ (.B(_0914_),
    .C(_0915_),
    .A(_0913_),
    .Y(_0916_));
 sg13g2_nand3_1 _3353_ (.B(_0574_),
    .C(_0916_),
    .A(net2),
    .Y(_0917_));
 sg13g2_o21ai_1 _3354_ (.B1(net365),
    .Y(_0918_),
    .A1(_1189_),
    .A2(_0575_));
 sg13g2_a21oi_1 _3355_ (.A1(_1189_),
    .A2(_0917_),
    .Y(_0146_),
    .B1(_0918_));
 sg13g2_nand2_1 _3356_ (.Y(_0919_),
    .A(net447),
    .B(net292));
 sg13g2_xnor2_1 _3357_ (.Y(_0920_),
    .A(net447),
    .B(\matt_venn_clock.pulse_min.count[0] ));
 sg13g2_or2_1 _3358_ (.X(_0921_),
    .B(_0917_),
    .A(net352));
 sg13g2_o21ai_1 _3359_ (.B1(_0919_),
    .Y(_0147_),
    .A1(_0920_),
    .A2(_0921_));
 sg13g2_nand2_1 _3360_ (.Y(_0922_),
    .A(net422),
    .B(net292));
 sg13g2_a21oi_1 _3361_ (.A1(\matt_venn_clock.pulse_min.count[1] ),
    .A2(\matt_venn_clock.pulse_min.count[0] ),
    .Y(_0923_),
    .B1(net422));
 sg13g2_nand3_1 _3362_ (.B(\matt_venn_clock.pulse_min.count[1] ),
    .C(\matt_venn_clock.pulse_min.count[0] ),
    .A(\matt_venn_clock.pulse_min.count[2] ),
    .Y(_0924_));
 sg13g2_nand2b_1 _3363_ (.Y(_0925_),
    .B(_0924_),
    .A_N(_0923_));
 sg13g2_o21ai_1 _3364_ (.B1(_0922_),
    .Y(_0148_),
    .A1(_0921_),
    .A2(_0925_));
 sg13g2_nand2_1 _3365_ (.Y(_0926_),
    .A(net425),
    .B(net292));
 sg13g2_nand4_1 _3366_ (.B(\matt_venn_clock.pulse_min.count[2] ),
    .C(\matt_venn_clock.pulse_min.count[1] ),
    .A(\matt_venn_clock.pulse_min.count[3] ),
    .Y(_0927_),
    .D(\matt_venn_clock.pulse_min.count[0] ));
 sg13g2_xor2_1 _3367_ (.B(_0924_),
    .A(net425),
    .X(_0928_));
 sg13g2_o21ai_1 _3368_ (.B1(_0926_),
    .Y(_0149_),
    .A1(_0921_),
    .A2(_0928_));
 sg13g2_nand2_1 _3369_ (.Y(_0929_),
    .A(net251),
    .B(net292));
 sg13g2_xnor2_1 _3370_ (.Y(_0930_),
    .A(_0055_),
    .B(_0927_));
 sg13g2_o21ai_1 _3371_ (.B1(_0929_),
    .Y(_0150_),
    .A1(_0921_),
    .A2(_0930_));
 sg13g2_nor3_1 _3372_ (.A(net383),
    .B(\matt_venn_clock.pulse_sec.comp[3] ),
    .C(\matt_venn_clock.pulse_sec.comp[2] ),
    .Y(_0931_));
 sg13g2_nor3_1 _3373_ (.A(\matt_venn_clock.pulse_sec.count[3] ),
    .B(\matt_venn_clock.pulse_sec.count[1] ),
    .C(\matt_venn_clock.pulse_sec.count[0] ),
    .Y(_0932_));
 sg13g2_nand3b_1 _3374_ (.B(_0054_),
    .C(_0932_),
    .Y(_0933_),
    .A_N(\matt_venn_clock.pulse_sec.count[2] ));
 sg13g2_nor3_1 _3375_ (.A(_0579_),
    .B(_0931_),
    .C(_0933_),
    .Y(_0934_));
 sg13g2_o21ai_1 _3376_ (.B1(net3),
    .Y(_0935_),
    .A1(_0931_),
    .A2(_0933_));
 sg13g2_a21o_1 _3377_ (.A2(_0934_),
    .A1(net3),
    .B1(_1188_),
    .X(_0936_));
 sg13g2_nand3_1 _3378_ (.B(net296),
    .C(_0935_),
    .A(_1188_),
    .Y(_0937_));
 sg13g2_nor2_1 _3379_ (.A(net3),
    .B(_0579_),
    .Y(_0938_));
 sg13g2_nand3_1 _3380_ (.B(_0936_),
    .C(_0937_),
    .A(net366),
    .Y(_0151_));
 sg13g2_nand2_1 _3381_ (.Y(_0939_),
    .A(net451),
    .B(_0937_));
 sg13g2_o21ai_1 _3382_ (.B1(net366),
    .Y(_0940_),
    .A1(net3),
    .A2(net294));
 sg13g2_nand2b_1 _3383_ (.Y(_0941_),
    .B(_1187_),
    .A_N(_0937_));
 sg13g2_nand3b_1 _3384_ (.B(_0941_),
    .C(_0939_),
    .Y(_0152_),
    .A_N(_0940_));
 sg13g2_nand2_1 _3385_ (.Y(_0942_),
    .A(net441),
    .B(_0941_));
 sg13g2_nor3_1 _3386_ (.A(\matt_venn_clock.pulse_sec.comp[2] ),
    .B(net451),
    .C(\matt_venn_clock.pulse_sec.comp[0] ),
    .Y(_0943_));
 sg13g2_a21oi_1 _3387_ (.A1(_0934_),
    .A2(_0943_),
    .Y(_0944_),
    .B1(_0938_));
 sg13g2_nand3_1 _3388_ (.B(_0942_),
    .C(_0944_),
    .A(net365),
    .Y(_0153_));
 sg13g2_nand2_1 _3389_ (.Y(_0945_),
    .A(net3),
    .B(net296));
 sg13g2_nor2_2 _3390_ (.A(_0933_),
    .B(_0945_),
    .Y(_0946_));
 sg13g2_nand2_1 _3391_ (.Y(_0947_),
    .A(_0943_),
    .B(_0946_));
 sg13g2_or2_1 _3392_ (.X(_0948_),
    .B(_0944_),
    .A(net470));
 sg13g2_a21oi_1 _3393_ (.A1(net470),
    .A2(_0947_),
    .Y(_0949_),
    .B1(net352));
 sg13g2_nand2_1 _3394_ (.Y(_0154_),
    .A(_0948_),
    .B(net471));
 sg13g2_nand2_1 _3395_ (.Y(_0950_),
    .A(net383),
    .B(_0948_));
 sg13g2_nand4_1 _3396_ (.B(_1188_),
    .C(_0931_),
    .A(_1187_),
    .Y(_0951_),
    .D(_0938_));
 sg13g2_a21oi_1 _3397_ (.A1(net384),
    .A2(_0951_),
    .Y(_0155_),
    .B1(_0940_));
 sg13g2_xnor2_1 _3398_ (.Y(_0952_),
    .A(net246),
    .B(\matt_venn_clock.pulse_sec.comp[4] ));
 sg13g2_xnor2_1 _3399_ (.Y(_0953_),
    .A(\matt_venn_clock.pulse_sec.count[2] ),
    .B(\matt_venn_clock.pulse_sec.comp[2] ));
 sg13g2_a22oi_1 _3400_ (.Y(_0954_),
    .B1(_1188_),
    .B2(\matt_venn_clock.pulse_sec.count[0] ),
    .A2(\matt_venn_clock.pulse_sec.comp[3] ),
    .A1(_1185_));
 sg13g2_a22oi_1 _3401_ (.Y(_0955_),
    .B1(\matt_venn_clock.pulse_sec.comp[0] ),
    .B2(_1186_),
    .A2(_1187_),
    .A1(\matt_venn_clock.pulse_sec.count[1] ));
 sg13g2_nand2b_1 _3402_ (.Y(_0956_),
    .B(\matt_venn_clock.pulse_sec.comp[1] ),
    .A_N(\matt_venn_clock.pulse_sec.count[1] ));
 sg13g2_nand2b_1 _3403_ (.Y(_0957_),
    .B(\matt_venn_clock.pulse_sec.count[3] ),
    .A_N(\matt_venn_clock.pulse_sec.comp[3] ));
 sg13g2_and4_1 _3404_ (.A(_0954_),
    .B(_0955_),
    .C(_0956_),
    .D(_0957_),
    .X(_0958_));
 sg13g2_nand3_1 _3405_ (.B(_0953_),
    .C(_0958_),
    .A(_0952_),
    .Y(_0959_));
 sg13g2_nand3_1 _3406_ (.B(_0574_),
    .C(_0959_),
    .A(net3),
    .Y(_0960_));
 sg13g2_o21ai_1 _3407_ (.B1(net365),
    .Y(_0961_),
    .A1(_1186_),
    .A2(net294));
 sg13g2_a21oi_1 _3408_ (.A1(_1186_),
    .A2(_0960_),
    .Y(_0156_),
    .B1(_0961_));
 sg13g2_nand2_1 _3409_ (.Y(_0962_),
    .A(net445),
    .B(net292));
 sg13g2_xnor2_1 _3410_ (.Y(_0963_),
    .A(net445),
    .B(\matt_venn_clock.pulse_sec.count[0] ));
 sg13g2_or2_1 _3411_ (.X(_0964_),
    .B(_0960_),
    .A(net352));
 sg13g2_o21ai_1 _3412_ (.B1(_0962_),
    .Y(_0157_),
    .A1(_0963_),
    .A2(_0964_));
 sg13g2_nand2_1 _3413_ (.Y(_0965_),
    .A(net429),
    .B(net292));
 sg13g2_a21oi_1 _3414_ (.A1(\matt_venn_clock.pulse_sec.count[1] ),
    .A2(\matt_venn_clock.pulse_sec.count[0] ),
    .Y(_0966_),
    .B1(net429));
 sg13g2_nand3_1 _3415_ (.B(\matt_venn_clock.pulse_sec.count[1] ),
    .C(\matt_venn_clock.pulse_sec.count[0] ),
    .A(net541),
    .Y(_0967_));
 sg13g2_nand2b_1 _3416_ (.Y(_0968_),
    .B(_0967_),
    .A_N(_0966_));
 sg13g2_o21ai_1 _3417_ (.B1(_0965_),
    .Y(_0158_),
    .A1(_0964_),
    .A2(_0968_));
 sg13g2_nand2_1 _3418_ (.Y(_0969_),
    .A(net268),
    .B(net292));
 sg13g2_or2_1 _3419_ (.X(_0970_),
    .B(_0967_),
    .A(_1185_));
 sg13g2_xnor2_1 _3420_ (.Y(_0971_),
    .A(_1185_),
    .B(net542));
 sg13g2_o21ai_1 _3421_ (.B1(_0969_),
    .Y(_0159_),
    .A1(_0964_),
    .A2(_0971_));
 sg13g2_nand2_1 _3422_ (.Y(_0972_),
    .A(net246),
    .B(net292));
 sg13g2_xnor2_1 _3423_ (.Y(_0973_),
    .A(_0054_),
    .B(_0970_));
 sg13g2_o21ai_1 _3424_ (.B1(_0972_),
    .Y(_0160_),
    .A1(_0964_),
    .A2(_0973_));
 sg13g2_nand3b_1 _3425_ (.B(\clock_sec_d[1] ),
    .C(\clock_sec_d[2] ),
    .Y(_0974_),
    .A_N(\clock_sec_d[0] ));
 sg13g2_nand2_2 _3426_ (.Y(_0975_),
    .A(_0891_),
    .B(_0974_));
 sg13g2_inv_1 _3427_ (.Y(_0976_),
    .A(_0975_));
 sg13g2_o21ai_1 _3428_ (.B1(net363),
    .Y(_0977_),
    .A1(\clock_color_offset[0] ),
    .A2(_0975_));
 sg13g2_a21oi_1 _3429_ (.A1(_1184_),
    .A2(_0975_),
    .Y(_0161_),
    .B1(_0977_));
 sg13g2_a21oi_1 _3430_ (.A1(\clock_color_offset[0] ),
    .A2(_0975_),
    .Y(_0978_),
    .B1(net403));
 sg13g2_and3_1 _3431_ (.X(_0979_),
    .A(net403),
    .B(\clock_color_offset[0] ),
    .C(_0975_));
 sg13g2_nor3_1 _3432_ (.A(net352),
    .B(net404),
    .C(_0979_),
    .Y(_0162_));
 sg13g2_o21ai_1 _3433_ (.B1(net363),
    .Y(_0980_),
    .A1(net372),
    .A2(_0979_));
 sg13g2_a21oi_1 _3434_ (.A1(net372),
    .A2(_0979_),
    .Y(_0163_),
    .B1(_0980_));
 sg13g2_nor2_1 _3435_ (.A(net444),
    .B(\clock_hrs_u[0] ),
    .Y(_0981_));
 sg13g2_nand3_1 _3436_ (.B(\clock_hrs_d[1] ),
    .C(_0981_),
    .A(\clock_hrs_u[2] ),
    .Y(_0982_));
 sg13g2_nor3_1 _3437_ (.A(\clock_hrs_u[3] ),
    .B(\clock_hrs_d[0] ),
    .C(_0982_),
    .Y(_0983_));
 sg13g2_nand2b_1 _3438_ (.Y(_0984_),
    .B(net358),
    .A_N(_0983_));
 sg13g2_nand2_1 _3439_ (.Y(_0985_),
    .A(\clock_hrs_u[3] ),
    .B(\clock_hrs_u[1] ));
 sg13g2_nor3_2 _3440_ (.A(\clock_hrs_u[2] ),
    .B(\clock_hrs_u[0] ),
    .C(_0985_),
    .Y(_0986_));
 sg13g2_nand2b_1 _3441_ (.Y(_0987_),
    .B(\clock_hrs_d[0] ),
    .A_N(_0986_));
 sg13g2_nand2_1 _3442_ (.Y(_0988_),
    .A(net225),
    .B(_0986_));
 sg13g2_a21oi_1 _3443_ (.A1(_0987_),
    .A2(net226),
    .Y(_0164_),
    .B1(_0984_));
 sg13g2_nand2_1 _3444_ (.Y(_0989_),
    .A(\clock_hrs_d[0] ),
    .B(_0986_));
 sg13g2_xor2_1 _3445_ (.B(_0989_),
    .A(net409),
    .X(_0990_));
 sg13g2_nor2_1 _3446_ (.A(_0984_),
    .B(net410),
    .Y(_0165_));
 sg13g2_nand3_1 _3447_ (.B(\clock_min_d[1] ),
    .C(_1182_),
    .A(\clock_min_d[2] ),
    .Y(_0991_));
 sg13g2_nor2_1 _3448_ (.A(_0983_),
    .B(_0986_),
    .Y(_0992_));
 sg13g2_nand3_1 _3449_ (.B(_0991_),
    .C(_0992_),
    .A(_0862_),
    .Y(_0993_));
 sg13g2_nor4_1 _3450_ (.A(\clock_hrs_u[0] ),
    .B(_0861_),
    .C(_0983_),
    .D(_0986_),
    .Y(_0994_));
 sg13g2_a21oi_1 _3451_ (.A1(net378),
    .A2(_0861_),
    .Y(_0995_),
    .B1(_0994_));
 sg13g2_o21ai_1 _3452_ (.B1(net358),
    .Y(_0996_),
    .A1(_0993_),
    .A2(_0995_));
 sg13g2_a21oi_1 _3453_ (.A1(_0993_),
    .A2(net379),
    .Y(_0166_),
    .B1(_0996_));
 sg13g2_nand2_1 _3454_ (.Y(_0997_),
    .A(net444),
    .B(\clock_hrs_u[0] ));
 sg13g2_a21oi_1 _3455_ (.A1(_0862_),
    .A2(_0986_),
    .Y(_0998_),
    .B1(_0981_));
 sg13g2_nand2_1 _3456_ (.Y(_0999_),
    .A(_0997_),
    .B(_0998_));
 sg13g2_o21ai_1 _3457_ (.B1(net358),
    .Y(_1000_),
    .A1(net444),
    .A2(_0993_));
 sg13g2_a21oi_1 _3458_ (.A1(_0993_),
    .A2(_0999_),
    .Y(_0167_),
    .B1(_1000_));
 sg13g2_nor2_1 _3459_ (.A(_0861_),
    .B(_0992_),
    .Y(_1001_));
 sg13g2_nor2_1 _3460_ (.A(_0036_),
    .B(_0997_),
    .Y(_1002_));
 sg13g2_xnor2_1 _3461_ (.Y(_1003_),
    .A(_0036_),
    .B(_0997_));
 sg13g2_o21ai_1 _3462_ (.B1(_0993_),
    .Y(_1004_),
    .A1(_1001_),
    .A2(_1003_));
 sg13g2_o21ai_1 _3463_ (.B1(net358),
    .Y(_1005_),
    .A1(net458),
    .A2(_0993_));
 sg13g2_nor2b_1 _3464_ (.A(_1005_),
    .B_N(_1004_),
    .Y(_0168_));
 sg13g2_xor2_1 _3465_ (.B(_1002_),
    .A(_0033_),
    .X(_1006_));
 sg13g2_o21ai_1 _3466_ (.B1(_0993_),
    .Y(_1007_),
    .A1(_1001_),
    .A2(_1006_));
 sg13g2_o21ai_1 _3467_ (.B1(_1007_),
    .Y(_1008_),
    .A1(net449),
    .A2(_0993_));
 sg13g2_nor2_1 _3468_ (.A(net350),
    .B(net450),
    .Y(_0169_));
 sg13g2_nor4_1 _3469_ (.A(_1180_),
    .B(net248),
    .C(_1181_),
    .D(\clock_min_u[0] ),
    .Y(_1009_));
 sg13g2_nor2_1 _3470_ (.A(\clock_min_d[0] ),
    .B(net303),
    .Y(_1010_));
 sg13g2_nand2_1 _3471_ (.Y(_1011_),
    .A(net357),
    .B(_0991_));
 sg13g2_nor2b_1 _3472_ (.A(net223),
    .B_N(net303),
    .Y(_1012_));
 sg13g2_nor3_1 _3473_ (.A(_1010_),
    .B(_1011_),
    .C(_1012_),
    .Y(_0170_));
 sg13g2_nand3_1 _3474_ (.B(net494),
    .C(net303),
    .A(\clock_min_d[1] ),
    .Y(_1013_));
 sg13g2_a21oi_1 _3475_ (.A1(net494),
    .A2(net303),
    .Y(_1014_),
    .B1(\clock_min_d[1] ));
 sg13g2_nor2_1 _3476_ (.A(_1011_),
    .B(net495),
    .Y(_1015_));
 sg13g2_and2_1 _3477_ (.A(_1013_),
    .B(_1015_),
    .X(_0171_));
 sg13g2_xor2_1 _3478_ (.B(_1013_),
    .A(net400),
    .X(_1016_));
 sg13g2_nor2_1 _3479_ (.A(_1011_),
    .B(net401),
    .Y(_0172_));
 sg13g2_nor2_1 _3480_ (.A(_0975_),
    .B(_1009_),
    .Y(_1017_));
 sg13g2_or2_1 _3481_ (.X(_1018_),
    .B(net303),
    .A(_0975_));
 sg13g2_nor2_1 _3482_ (.A(\clock_min_u[0] ),
    .B(net303),
    .Y(_1019_));
 sg13g2_mux2_1 _3483_ (.A0(net386),
    .A1(_1019_),
    .S(_0891_),
    .X(_1020_));
 sg13g2_o21ai_1 _3484_ (.B1(net357),
    .Y(_1021_),
    .A1(_1017_),
    .A2(_1020_));
 sg13g2_a21oi_1 _3485_ (.A1(_1017_),
    .A2(_1020_),
    .Y(_0173_),
    .B1(_1021_));
 sg13g2_nand2_1 _3486_ (.Y(_1022_),
    .A(\clock_min_u[0] ),
    .B(_0975_));
 sg13g2_a21o_1 _3487_ (.A2(net303),
    .A1(_0891_),
    .B1(net350),
    .X(_1023_));
 sg13g2_nand2_1 _3488_ (.Y(_1024_),
    .A(\clock_min_u[1] ),
    .B(\clock_min_u[0] ));
 sg13g2_xnor2_1 _3489_ (.Y(_1025_),
    .A(_1181_),
    .B(_1022_));
 sg13g2_nor2_1 _3490_ (.A(_1023_),
    .B(net498),
    .Y(_0174_));
 sg13g2_nor2_1 _3491_ (.A(_0038_),
    .B(_1024_),
    .Y(_1026_));
 sg13g2_a22oi_1 _3492_ (.Y(_1027_),
    .B1(_1024_),
    .B2(_0038_),
    .A2(net303),
    .A1(_0891_));
 sg13g2_nor2b_1 _3493_ (.A(_1026_),
    .B_N(_1027_),
    .Y(_1028_));
 sg13g2_a22oi_1 _3494_ (.Y(_1029_),
    .B1(_1018_),
    .B2(_1028_),
    .A2(_0976_),
    .A1(net248));
 sg13g2_nor2_1 _3495_ (.A(net350),
    .B(net249),
    .Y(_0175_));
 sg13g2_xor2_1 _3496_ (.B(_1026_),
    .A(_0034_),
    .X(_1030_));
 sg13g2_a221oi_1 _3497_ (.B2(_1030_),
    .C1(_1023_),
    .B1(_1018_),
    .A1(_1180_),
    .Y(_0176_),
    .A2(_0976_));
 sg13g2_nand2_1 _3498_ (.Y(_1031_),
    .A(net265),
    .B(\clock_sec_u[1] ));
 sg13g2_nor3_2 _3499_ (.A(net273),
    .B(\clock_sec_u[0] ),
    .C(_1031_),
    .Y(_1032_));
 sg13g2_nor2b_1 _3500_ (.A(_0062_),
    .B_N(_1032_),
    .Y(_1033_));
 sg13g2_nand2_1 _3501_ (.Y(_1034_),
    .A(net357),
    .B(_0974_));
 sg13g2_nor2_1 _3502_ (.A(net390),
    .B(_1032_),
    .Y(_1035_));
 sg13g2_nor3_1 _3503_ (.A(_1033_),
    .B(_1034_),
    .C(net391),
    .Y(_0177_));
 sg13g2_nand3_1 _3504_ (.B(net390),
    .C(_1032_),
    .A(net513),
    .Y(_1036_));
 sg13g2_a21oi_1 _3505_ (.A1(net390),
    .A2(_1032_),
    .Y(_1037_),
    .B1(net513));
 sg13g2_nor2_1 _3506_ (.A(_1034_),
    .B(_1037_),
    .Y(_1038_));
 sg13g2_and2_1 _3507_ (.A(_1036_),
    .B(_1038_),
    .X(_0178_));
 sg13g2_xor2_1 _3508_ (.B(_1036_),
    .A(net407),
    .X(_1039_));
 sg13g2_nor2_1 _3509_ (.A(_1034_),
    .B(net408),
    .Y(_0179_));
 sg13g2_and3_1 _3510_ (.X(_1040_),
    .A(net232),
    .B(\matt_venn_clock.sec_counter[1] ),
    .C(\matt_venn_clock.sec_counter[0] ));
 sg13g2_and2_1 _3511_ (.A(net263),
    .B(_1040_),
    .X(_1041_));
 sg13g2_and2_1 _3512_ (.A(net267),
    .B(_1041_),
    .X(_1042_));
 sg13g2_and2_1 _3513_ (.A(net244),
    .B(_1042_),
    .X(_1043_));
 sg13g2_and2_1 _3514_ (.A(net374),
    .B(_1043_),
    .X(_1044_));
 sg13g2_and2_1 _3515_ (.A(net275),
    .B(_1044_),
    .X(_1045_));
 sg13g2_nand3_1 _3516_ (.B(net457),
    .C(_1045_),
    .A(net479),
    .Y(_1046_));
 sg13g2_nor2_1 _3517_ (.A(_1212_),
    .B(_1046_),
    .Y(_1047_));
 sg13g2_and2_1 _3518_ (.A(\matt_venn_clock.sec_counter[11] ),
    .B(_1047_),
    .X(_1048_));
 sg13g2_and3_1 _3519_ (.X(_1049_),
    .A(\matt_venn_clock.sec_counter[12] ),
    .B(net416),
    .C(_1048_));
 sg13g2_and2_1 _3520_ (.A(net540),
    .B(_1049_),
    .X(_1050_));
 sg13g2_and2_1 _3521_ (.A(net388),
    .B(_1050_),
    .X(_1051_));
 sg13g2_and2_1 _3522_ (.A(net543),
    .B(_1051_),
    .X(_1052_));
 sg13g2_and2_1 _3523_ (.A(net370),
    .B(_1052_),
    .X(_1053_));
 sg13g2_and3_1 _3524_ (.X(_1054_),
    .A(\matt_venn_clock.sec_counter[19] ),
    .B(\matt_venn_clock.sec_counter[18] ),
    .C(_1053_));
 sg13g2_and3_1 _3525_ (.X(_1055_),
    .A(net238),
    .B(net539),
    .C(_1054_));
 sg13g2_xnor2_1 _3526_ (.Y(_1056_),
    .A(net491),
    .B(_1055_));
 sg13g2_nand2b_1 _3527_ (.Y(_1057_),
    .B(_1053_),
    .A_N(net398));
 sg13g2_xor2_1 _3528_ (.B(_1057_),
    .A(net486),
    .X(_1058_));
 sg13g2_xnor2_1 _3529_ (.Y(_1059_),
    .A(net454),
    .B(_1051_));
 sg13g2_xnor2_1 _3530_ (.Y(_1060_),
    .A(net431),
    .B(_1049_));
 sg13g2_nor2b_1 _3531_ (.A(net412),
    .B_N(_1048_),
    .Y(_1061_));
 sg13g2_xnor2_1 _3532_ (.Y(_1062_),
    .A(net416),
    .B(_1061_));
 sg13g2_xnor2_1 _3533_ (.Y(_1063_),
    .A(net434),
    .B(_1047_));
 sg13g2_xnor2_1 _3534_ (.Y(_1064_),
    .A(_1212_),
    .B(_1046_));
 sg13g2_a21o_1 _3535_ (.A2(_1045_),
    .A1(net457),
    .B1(net479),
    .X(_1065_));
 sg13g2_nand2_1 _3536_ (.Y(_1066_),
    .A(_1046_),
    .B(_1065_));
 sg13g2_xnor2_1 _3537_ (.Y(_1067_),
    .A(net457),
    .B(_1045_));
 sg13g2_nand2b_1 _3538_ (.Y(_1068_),
    .B(\matt_venn_clock.sec_counter[24] ),
    .A_N(\matt_venn_clock.sec_counter[17] ));
 sg13g2_nor4_1 _3539_ (.A(\matt_venn_clock.sec_counter[6] ),
    .B(\matt_venn_clock.sec_counter[7] ),
    .C(_0048_),
    .D(\matt_venn_clock.sec_counter[23] ),
    .Y(_1069_));
 sg13g2_nand3_1 _3540_ (.B(\matt_venn_clock.sec_counter[20] ),
    .C(_1069_),
    .A(\matt_venn_clock.sec_counter[21] ),
    .Y(_1070_));
 sg13g2_nor4_1 _3541_ (.A(\matt_venn_clock.sec_counter[15] ),
    .B(_0049_),
    .C(_1068_),
    .D(_1070_),
    .Y(_1071_));
 sg13g2_and2_1 _3542_ (.A(_1043_),
    .B(_1071_),
    .X(_1072_));
 sg13g2_nand4_1 _3543_ (.B(_1066_),
    .C(_1067_),
    .A(_1064_),
    .Y(_1073_),
    .D(_1072_));
 sg13g2_or4_1 _3544_ (.A(_1060_),
    .B(_1062_),
    .C(_1063_),
    .D(_1073_),
    .X(_1074_));
 sg13g2_nor4_2 _3545_ (.A(_1056_),
    .B(_1058_),
    .C(_1059_),
    .Y(_1075_),
    .D(_1074_));
 sg13g2_inv_2 _3546_ (.Y(_1076_),
    .A(_1075_));
 sg13g2_nor3_1 _3547_ (.A(\clock_sec_u[0] ),
    .B(_0946_),
    .C(_1076_),
    .Y(_1077_));
 sg13g2_or2_2 _3548_ (.X(_1078_),
    .B(_1075_),
    .A(_0946_));
 sg13g2_inv_1 _3549_ (.Y(_1079_),
    .A(_1078_));
 sg13g2_a221oi_1 _3550_ (.B2(\clock_sec_u[0] ),
    .C1(_1077_),
    .B1(_1079_),
    .A1(net438),
    .Y(_1080_),
    .A2(_0946_));
 sg13g2_nor2_1 _3551_ (.A(net350),
    .B(net439),
    .Y(_0180_));
 sg13g2_nor2_1 _3552_ (.A(_1032_),
    .B(_1078_),
    .Y(_1081_));
 sg13g2_nand2_1 _3553_ (.Y(_1082_),
    .A(\clock_sec_u[1] ),
    .B(\clock_sec_u[0] ));
 sg13g2_xor2_1 _3554_ (.B(\clock_sec_u[0] ),
    .A(net460),
    .X(_1083_));
 sg13g2_a22oi_1 _3555_ (.Y(_1084_),
    .B1(_1083_),
    .B2(_1078_),
    .A2(_1081_),
    .A1(net460));
 sg13g2_nor2_1 _3556_ (.A(net350),
    .B(net461),
    .Y(_0181_));
 sg13g2_nor2_1 _3557_ (.A(_0040_),
    .B(_1082_),
    .Y(_1085_));
 sg13g2_xor2_1 _3558_ (.B(_1082_),
    .A(_0040_),
    .X(_1086_));
 sg13g2_nor2_1 _3559_ (.A(net273),
    .B(_1078_),
    .Y(_1087_));
 sg13g2_nor2_1 _3560_ (.A(_1079_),
    .B(_1086_),
    .Y(_1088_));
 sg13g2_nor3_1 _3561_ (.A(net350),
    .B(_1087_),
    .C(_1088_),
    .Y(_0182_));
 sg13g2_xnor2_1 _3562_ (.Y(_1089_),
    .A(_0035_),
    .B(_1085_));
 sg13g2_a22oi_1 _3563_ (.Y(_1090_),
    .B1(_1089_),
    .B2(_1078_),
    .A2(_1081_),
    .A1(net265));
 sg13g2_nor2_1 _3564_ (.A(net350),
    .B(net266),
    .Y(_0183_));
 sg13g2_nand2b_1 _3565_ (.Y(_1091_),
    .B(_0568_),
    .A_N(_0565_));
 sg13g2_nor2b_1 _3566_ (.A(_0571_),
    .B_N(_1091_),
    .Y(_0184_));
 sg13g2_a21oi_1 _3567_ (.A1(_0567_),
    .A2(_1091_),
    .Y(_0185_),
    .B1(_0572_));
 sg13g2_and2_1 _3568_ (.A(_0567_),
    .B(_0571_),
    .X(_0186_));
 sg13g2_nor4_1 _3569_ (.A(\matt_venn_vga.x_block_q[5] ),
    .B(\matt_venn_vga.y_block_q[4] ),
    .C(net240),
    .D(\matt_venn_vga.y_block_q[5] ),
    .Y(_1092_));
 sg13g2_nor3_1 _3570_ (.A(\matt_venn_vga.font_0.dout[3] ),
    .B(\matt_venn_vga.col_index_q[0] ),
    .C(\matt_venn_vga.col_index_q[1] ),
    .Y(_1093_));
 sg13g2_o21ai_1 _3571_ (.B1(\matt_venn_vga.y_block_q[2] ),
    .Y(_1094_),
    .A1(\matt_venn_vga.y_block_q[1] ),
    .A2(\matt_venn_vga.y_block_q[0] ));
 sg13g2_o21ai_1 _3572_ (.B1(\matt_venn_vga.col_index_q[0] ),
    .Y(_1095_),
    .A1(_1232_),
    .A2(\matt_venn_vga.col_index_q[1] ));
 sg13g2_nand2_1 _3573_ (.Y(_1096_),
    .A(_1094_),
    .B(_1095_));
 sg13g2_o21ai_1 _3574_ (.B1(net241),
    .Y(_1097_),
    .A1(\matt_venn_vga.font_0.dout[1] ),
    .A2(_1233_));
 sg13g2_nor3_1 _3575_ (.A(_1093_),
    .B(_1096_),
    .C(net242),
    .Y(_0187_));
 sg13g2_nand2_1 _3576_ (.Y(_1098_),
    .A(net365),
    .B(_1076_));
 sg13g2_and3_1 _3577_ (.X(_0188_),
    .A(net366),
    .B(net219),
    .C(_1076_));
 sg13g2_xnor2_1 _3578_ (.Y(_1099_),
    .A(net380),
    .B(\matt_venn_clock.sec_counter[0] ));
 sg13g2_nor2_1 _3579_ (.A(net278),
    .B(net381),
    .Y(_0189_));
 sg13g2_a21oi_1 _3580_ (.A1(\matt_venn_clock.sec_counter[1] ),
    .A2(\matt_venn_clock.sec_counter[0] ),
    .Y(_1100_),
    .B1(net232));
 sg13g2_nor3_1 _3581_ (.A(_1040_),
    .B(net278),
    .C(net233),
    .Y(_0190_));
 sg13g2_nor2_1 _3582_ (.A(net263),
    .B(_1040_),
    .Y(_1101_));
 sg13g2_nor3_1 _3583_ (.A(_1041_),
    .B(net278),
    .C(net264),
    .Y(_0191_));
 sg13g2_nor2_1 _3584_ (.A(net267),
    .B(_1041_),
    .Y(_1102_));
 sg13g2_nor3_1 _3585_ (.A(_1042_),
    .B(net278),
    .C(_1102_),
    .Y(_0192_));
 sg13g2_nor2_1 _3586_ (.A(net244),
    .B(_1042_),
    .Y(_1103_));
 sg13g2_nor3_1 _3587_ (.A(_1043_),
    .B(net278),
    .C(net245),
    .Y(_0193_));
 sg13g2_nor2_1 _3588_ (.A(net374),
    .B(_1043_),
    .Y(_1104_));
 sg13g2_nor3_1 _3589_ (.A(_1044_),
    .B(_1098_),
    .C(_1104_),
    .Y(_0194_));
 sg13g2_nor2_1 _3590_ (.A(net275),
    .B(_1044_),
    .Y(_1105_));
 sg13g2_nor3_1 _3591_ (.A(_1045_),
    .B(net278),
    .C(net368),
    .Y(_0195_));
 sg13g2_nor2_1 _3592_ (.A(_1067_),
    .B(net277),
    .Y(_0196_));
 sg13g2_nor2_1 _3593_ (.A(_1066_),
    .B(net277),
    .Y(_0197_));
 sg13g2_nor2_1 _3594_ (.A(net477),
    .B(net277),
    .Y(_0198_));
 sg13g2_nor2_1 _3595_ (.A(net435),
    .B(net276),
    .Y(_0199_));
 sg13g2_nor2b_1 _3596_ (.A(_1048_),
    .B_N(net412),
    .Y(_1106_));
 sg13g2_nor3_1 _3597_ (.A(_1061_),
    .B(net276),
    .C(net413),
    .Y(_0200_));
 sg13g2_nor2_1 _3598_ (.A(_1062_),
    .B(net276),
    .Y(_0201_));
 sg13g2_nor2_1 _3599_ (.A(net432),
    .B(net276),
    .Y(_0202_));
 sg13g2_nor2_1 _3600_ (.A(net388),
    .B(_1050_),
    .Y(_1107_));
 sg13g2_nor3_1 _3601_ (.A(_1051_),
    .B(net276),
    .C(net389),
    .Y(_0203_));
 sg13g2_nor2_1 _3602_ (.A(_1059_),
    .B(net276),
    .Y(_0204_));
 sg13g2_nor2_1 _3603_ (.A(net370),
    .B(_1052_),
    .Y(_1108_));
 sg13g2_nor3_1 _3604_ (.A(_1053_),
    .B(net276),
    .C(net371),
    .Y(_0205_));
 sg13g2_nand2b_1 _3605_ (.Y(_1109_),
    .B(net398),
    .A_N(_1053_));
 sg13g2_and4_1 _3606_ (.A(net365),
    .B(_1057_),
    .C(_1076_),
    .D(_1109_),
    .X(_0206_));
 sg13g2_nor2_1 _3607_ (.A(_1058_),
    .B(net276),
    .Y(_0207_));
 sg13g2_a21oi_1 _3608_ (.A1(net466),
    .A2(_1054_),
    .Y(_1110_),
    .B1(net277));
 sg13g2_o21ai_1 _3609_ (.B1(_1110_),
    .Y(_1111_),
    .A1(net466),
    .A2(_1054_));
 sg13g2_inv_1 _3610_ (.Y(_0208_),
    .A(net467));
 sg13g2_a21oi_1 _3611_ (.A1(\matt_venn_clock.sec_counter[20] ),
    .A2(_1054_),
    .Y(_1112_),
    .B1(net238));
 sg13g2_nor3_1 _3612_ (.A(_1055_),
    .B(net277),
    .C(net239),
    .Y(_0209_));
 sg13g2_nor2_1 _3613_ (.A(_1056_),
    .B(net277),
    .Y(_0210_));
 sg13g2_a21oi_1 _3614_ (.A1(\matt_venn_clock.sec_counter[22] ),
    .A2(_1055_),
    .Y(_1113_),
    .B1(net260));
 sg13g2_and3_1 _3615_ (.X(_1114_),
    .A(net260),
    .B(\matt_venn_clock.sec_counter[22] ),
    .C(_1055_));
 sg13g2_nor3_1 _3616_ (.A(net277),
    .B(net261),
    .C(_1114_),
    .Y(_0211_));
 sg13g2_xnor2_1 _3617_ (.Y(_1115_),
    .A(net271),
    .B(_1114_));
 sg13g2_nor2_1 _3618_ (.A(net277),
    .B(net272),
    .Y(_0212_));
 sg13g2_and2_1 _3619_ (.A(net362),
    .B(_0306_),
    .X(_0213_));
 sg13g2_a21oi_1 _3620_ (.A1(_1271_),
    .A2(net526),
    .Y(_0214_),
    .B1(net352));
 sg13g2_and2_1 _3621_ (.A(net362),
    .B(_0417_),
    .X(_0215_));
 sg13g2_and2_1 _3622_ (.A(net362),
    .B(_0416_),
    .X(_0216_));
 sg13g2_and2_1 _3623_ (.A(net362),
    .B(_0415_),
    .X(_0217_));
 sg13g2_and2_1 _3624_ (.A(net362),
    .B(_0429_),
    .X(_0218_));
 sg13g2_and2_1 _3625_ (.A(net362),
    .B(_0445_),
    .X(_0219_));
 sg13g2_nand2b_1 _3626_ (.Y(_1116_),
    .B(net337),
    .A_N(_0768_));
 sg13g2_and2_1 _3627_ (.A(_0773_),
    .B(_1116_),
    .X(_1117_));
 sg13g2_and2_1 _3628_ (.A(_0574_),
    .B(_1117_),
    .X(_1118_));
 sg13g2_and3_2 _3629_ (.X(_1119_),
    .A(_0580_),
    .B(_0773_),
    .C(_1116_));
 sg13g2_nand2_1 _3630_ (.Y(_1120_),
    .A(net296),
    .B(_1117_));
 sg13g2_o21ai_1 _3631_ (.B1(net359),
    .Y(_1121_),
    .A1(\product_comp[1] ),
    .A2(net284));
 sg13g2_a21oi_1 _3632_ (.A1(_1179_),
    .A2(net284),
    .Y(_0220_),
    .B1(_1121_));
 sg13g2_nor2b_1 _3633_ (.A(net338),
    .B_N(\product_comp[2] ),
    .Y(_1122_));
 sg13g2_nand2b_1 _3634_ (.Y(_1123_),
    .B(net338),
    .A_N(\product_comp[2] ));
 sg13g2_nor2b_1 _3635_ (.A(_1122_),
    .B_N(_1123_),
    .Y(_1124_));
 sg13g2_xnor2_1 _3636_ (.Y(_1125_),
    .A(_1179_),
    .B(_1124_));
 sg13g2_o21ai_1 _3637_ (.B1(net359),
    .Y(_1126_),
    .A1(net427),
    .A2(net284));
 sg13g2_a21oi_1 _3638_ (.A1(_1119_),
    .A2(_1125_),
    .Y(_0221_),
    .B1(_1126_));
 sg13g2_nand2_1 _3639_ (.Y(_1127_),
    .A(net455),
    .B(_1120_));
 sg13g2_xnor2_1 _3640_ (.Y(_1128_),
    .A(\product_comp[3] ),
    .B(net338));
 sg13g2_o21ai_1 _3641_ (.B1(_1123_),
    .Y(_1129_),
    .A1(\product_comp[1] ),
    .A2(_1122_));
 sg13g2_nor2_1 _3642_ (.A(_1128_),
    .B(_1129_),
    .Y(_1130_));
 sg13g2_nand2_1 _3643_ (.Y(_1131_),
    .A(_1128_),
    .B(_1129_));
 sg13g2_nand3b_1 _3644_ (.B(_1131_),
    .C(net284),
    .Y(_1132_),
    .A_N(_1130_));
 sg13g2_nand3_1 _3645_ (.B(_1127_),
    .C(_1132_),
    .A(net359),
    .Y(_0222_));
 sg13g2_nand2_1 _3646_ (.Y(_1133_),
    .A(\product_comp[4] ),
    .B(_1202_));
 sg13g2_xor2_1 _3647_ (.B(net338),
    .A(\product_comp[4] ),
    .X(_1134_));
 sg13g2_a21oi_1 _3648_ (.A1(net455),
    .A2(net338),
    .Y(_1135_),
    .B1(_1130_));
 sg13g2_xnor2_1 _3649_ (.Y(_1136_),
    .A(_1134_),
    .B(_1135_));
 sg13g2_o21ai_1 _3650_ (.B1(net359),
    .Y(_1137_),
    .A1(net485),
    .A2(net284));
 sg13g2_a21oi_1 _3651_ (.A1(net284),
    .A2(_1136_),
    .Y(_0223_),
    .B1(_1137_));
 sg13g2_nor2b_1 _3652_ (.A(net338),
    .B_N(\product_comp[5] ),
    .Y(_1138_));
 sg13g2_xnor2_1 _3653_ (.Y(_1139_),
    .A(\product_comp[5] ),
    .B(net338));
 sg13g2_o21ai_1 _3654_ (.B1(_1133_),
    .Y(_1140_),
    .A1(_1134_),
    .A2(_1135_));
 sg13g2_xnor2_1 _3655_ (.Y(_1141_),
    .A(_1139_),
    .B(_1140_));
 sg13g2_o21ai_1 _3656_ (.B1(net360),
    .Y(_1142_),
    .A1(net520),
    .A2(_1118_));
 sg13g2_a21oi_1 _3657_ (.A1(_1118_),
    .A2(_1141_),
    .Y(_0224_),
    .B1(_1142_));
 sg13g2_o21ai_1 _3658_ (.B1(net359),
    .Y(_1143_),
    .A1(net515),
    .A2(net284));
 sg13g2_xnor2_1 _3659_ (.Y(_1144_),
    .A(\product_comp[6] ),
    .B(net337));
 sg13g2_a21o_1 _3660_ (.A2(_1140_),
    .A1(_1139_),
    .B1(_1138_),
    .X(_1145_));
 sg13g2_xnor2_1 _3661_ (.Y(_1146_),
    .A(_1144_),
    .B(_1145_));
 sg13g2_a21oi_1 _3662_ (.A1(_1119_),
    .A2(_1146_),
    .Y(_0225_),
    .B1(_1143_));
 sg13g2_xor2_1 _3663_ (.B(net337),
    .A(\product_comp[7] ),
    .X(_1147_));
 sg13g2_nand3_1 _3664_ (.B(_1140_),
    .C(_1144_),
    .A(_1139_),
    .Y(_1148_));
 sg13g2_o21ai_1 _3665_ (.B1(_1202_),
    .Y(_1149_),
    .A1(\product_comp[6] ),
    .A2(\product_comp[5] ));
 sg13g2_and3_1 _3666_ (.X(_1150_),
    .A(_1147_),
    .B(_1148_),
    .C(_1149_));
 sg13g2_a21oi_1 _3667_ (.A1(_1148_),
    .A2(_1149_),
    .Y(_1151_),
    .B1(_1147_));
 sg13g2_nand2b_1 _3668_ (.Y(_1152_),
    .B(_1120_),
    .A_N(net516));
 sg13g2_o21ai_1 _3669_ (.B1(_1119_),
    .Y(_1153_),
    .A1(_1150_),
    .A2(_1151_));
 sg13g2_and3_1 _3670_ (.X(_0226_),
    .A(net359),
    .B(_1152_),
    .C(_1153_));
 sg13g2_o21ai_1 _3671_ (.B1(net359),
    .Y(_1154_),
    .A1(net499),
    .A2(net284));
 sg13g2_xnor2_1 _3672_ (.Y(_1155_),
    .A(\product_comp[8] ),
    .B(net337));
 sg13g2_a21oi_1 _3673_ (.A1(net548),
    .A2(_1202_),
    .Y(_1156_),
    .B1(_1151_));
 sg13g2_xor2_1 _3674_ (.B(_1156_),
    .A(_1155_),
    .X(_1157_));
 sg13g2_a21oi_1 _3675_ (.A1(_1119_),
    .A2(_1157_),
    .Y(_0227_),
    .B1(_1154_));
 sg13g2_nand2b_1 _3676_ (.Y(_1158_),
    .B(_1155_),
    .A_N(_1147_));
 sg13g2_nor2_1 _3677_ (.A(_1148_),
    .B(_1158_),
    .Y(_1159_));
 sg13g2_o21ai_1 _3678_ (.B1(_1202_),
    .Y(_1160_),
    .A1(\product_comp[8] ),
    .A2(\product_comp[7] ));
 sg13g2_nand2_1 _3679_ (.Y(_1161_),
    .A(_1149_),
    .B(_1160_));
 sg13g2_nor2_1 _3680_ (.A(_1159_),
    .B(_1161_),
    .Y(_1162_));
 sg13g2_xnor2_1 _3681_ (.Y(_1163_),
    .A(_1202_),
    .B(_1162_));
 sg13g2_and2_1 _3682_ (.A(_1119_),
    .B(_1163_),
    .X(_1164_));
 sg13g2_o21ai_1 _3683_ (.B1(net360),
    .Y(_1165_),
    .A1(net411),
    .A2(_1164_));
 sg13g2_a21oi_1 _3684_ (.A1(net411),
    .A2(_1164_),
    .Y(_0228_),
    .B1(_1165_));
 sg13g2_nor4_1 _3685_ (.A(\product_comp[9] ),
    .B(_1202_),
    .C(_1159_),
    .D(_1161_),
    .Y(_1166_));
 sg13g2_a21oi_1 _3686_ (.A1(_1177_),
    .A2(_1162_),
    .Y(_1167_),
    .B1(net337));
 sg13g2_nor3_1 _3687_ (.A(_1120_),
    .B(_1166_),
    .C(_1167_),
    .Y(_1168_));
 sg13g2_o21ai_1 _3688_ (.B1(net359),
    .Y(_1169_),
    .A1(net387),
    .A2(_1168_));
 sg13g2_a21oi_1 _3689_ (.A1(net387),
    .A2(_1168_),
    .Y(_0229_),
    .B1(_1169_));
 sg13g2_nor4_1 _3690_ (.A(\matt_venn_vga_shadow.x_block_q[5] ),
    .B(\matt_venn_vga_shadow.y_block_q[4] ),
    .C(\matt_venn_vga_shadow.y_block_q[3] ),
    .D(net256),
    .Y(_1170_));
 sg13g2_nor3_1 _3691_ (.A(\matt_venn_vga_shadow.font_0.dout[3] ),
    .B(\matt_venn_vga_shadow.col_index_q[0] ),
    .C(\matt_venn_vga_shadow.col_index_q[1] ),
    .Y(_1171_));
 sg13g2_o21ai_1 _3692_ (.B1(\matt_venn_vga_shadow.y_block_q[2] ),
    .Y(_1172_),
    .A1(\matt_venn_vga_shadow.y_block_q[1] ),
    .A2(\matt_venn_vga_shadow.y_block_q[0] ));
 sg13g2_o21ai_1 _3693_ (.B1(\matt_venn_vga_shadow.col_index_q[0] ),
    .Y(_1173_),
    .A1(_1234_),
    .A2(\matt_venn_vga_shadow.col_index_q[1] ));
 sg13g2_nand2_1 _3694_ (.Y(_1174_),
    .A(_1172_),
    .B(_1173_));
 sg13g2_o21ai_1 _3695_ (.B1(net257),
    .Y(_1175_),
    .A1(\matt_venn_vga_shadow.font_0.dout[1] ),
    .A2(_1235_));
 sg13g2_nor3_1 _3696_ (.A(_1171_),
    .B(_1174_),
    .C(net258),
    .Y(_0230_));
 sg13g2_or2_1 _3697_ (.X(_0231_),
    .B(net301),
    .A(net314));
 sg13g2_or2_1 _3698_ (.X(_0232_),
    .B(net301),
    .A(net311));
 sg13g2_nor2_1 _3699_ (.A(net352),
    .B(_0364_),
    .Y(_0233_));
 sg13g2_and2_1 _3700_ (.A(net363),
    .B(_0486_),
    .X(_0234_));
 sg13g2_and2_1 _3701_ (.A(net363),
    .B(_0484_),
    .X(_0235_));
 sg13g2_and2_1 _3702_ (.A(net362),
    .B(_0492_),
    .X(_0236_));
 sg13g2_and2_1 _3703_ (.A(net362),
    .B(_0498_),
    .X(_0237_));
 sg13g2_nor2_1 _3704_ (.A(net352),
    .B(_0504_),
    .Y(_0238_));
 sg13g2_and2_1 _3705_ (.A(net363),
    .B(_0510_),
    .X(_0239_));
 sg13g2_dfrbp_1 _3706_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net14),
    .D(_0000_),
    .Q_N(_1821_),
    .Q(\matt_venn_vga.digit_0.digit_index[0] ));
 sg13g2_dfrbp_1 _3707_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net15),
    .D(_0001_),
    .Q_N(_1822_),
    .Q(\matt_venn_vga.digit_0.digit_index[1] ));
 sg13g2_dfrbp_1 _3708_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net16),
    .D(_0002_),
    .Q_N(_1823_),
    .Q(\matt_venn_vga.digit_0.digit_index[2] ));
 sg13g2_dfrbp_1 _3709_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net17),
    .D(_0003_),
    .Q_N(_1824_),
    .Q(\matt_venn_vga.digit_0.digit_index[3] ));
 sg13g2_dfrbp_1 _3710_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net18),
    .D(_0004_),
    .Q_N(_1825_),
    .Q(\matt_venn_vga.digit_0.digit_index[4] ));
 sg13g2_dfrbp_1 _3711_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net19),
    .D(_0005_),
    .Q_N(_1826_),
    .Q(\matt_venn_vga.digit_0.digit_index[5] ));
 sg13g2_dfrbp_1 _3712_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net20),
    .D(_0011_),
    .Q_N(_1827_),
    .Q(\matt_venn_vga_shadow.digit_0.digit_index[0] ));
 sg13g2_dfrbp_1 _3713_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net21),
    .D(_0012_),
    .Q_N(_1828_),
    .Q(\matt_venn_vga_shadow.digit_0.digit_index[1] ));
 sg13g2_dfrbp_1 _3714_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net22),
    .D(_0013_),
    .Q_N(_1829_),
    .Q(\matt_venn_vga_shadow.digit_0.digit_index[2] ));
 sg13g2_dfrbp_1 _3715_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net23),
    .D(_0014_),
    .Q_N(_1830_),
    .Q(\matt_venn_vga_shadow.digit_0.digit_index[3] ));
 sg13g2_dfrbp_1 _3716_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net24),
    .D(_0015_),
    .Q_N(_1831_),
    .Q(\matt_venn_vga_shadow.digit_0.digit_index[4] ));
 sg13g2_dfrbp_1 _3717_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net25),
    .D(_0016_),
    .Q_N(_1832_),
    .Q(\matt_venn_vga_shadow.digit_0.digit_index[5] ));
 sg13g2_dfrbp_1 _3718_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net26),
    .D(_0017_),
    .Q_N(_1833_),
    .Q(\matt_venn_vga_shadow.color[4] ));
 sg13g2_dfrbp_1 _3719_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net27),
    .D(_0018_),
    .Q_N(_1834_),
    .Q(\matt_venn_vga_shadow.color[5] ));
 sg13g2_dfrbp_1 _3720_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net28),
    .D(_0006_),
    .Q_N(_1835_),
    .Q(\matt_venn_vga.color[4] ));
 sg13g2_dfrbp_1 _3721_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net29),
    .D(_0007_),
    .Q_N(_1836_),
    .Q(\matt_venn_vga.color[5] ));
 sg13g2_dfrbp_1 _3722_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net30),
    .D(_0008_),
    .Q_N(_1837_),
    .Q(\matt_venn_vga.font_0.dout[1] ));
 sg13g2_dfrbp_1 _3723_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net66),
    .D(_0009_),
    .Q_N(_1838_),
    .Q(\matt_venn_vga.font_0.dout[2] ));
 sg13g2_dfrbp_1 _3724_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net13),
    .D(_0010_),
    .Q_N(_1820_),
    .Q(\matt_venn_vga.font_0.dout[3] ));
 sg13g2_dfrbp_1 _3725_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net35),
    .D(_0068_),
    .Q_N(_1819_),
    .Q(\matt_venn_vga_shadow.color[3] ));
 sg13g2_dfrbp_1 _3726_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net34),
    .D(_0069_),
    .Q_N(_1818_),
    .Q(\matt_venn_vga_shadow.color[0] ));
 sg13g2_dfrbp_1 _3727_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net33),
    .D(_0070_),
    .Q_N(_1817_),
    .Q(\matt_venn_vga_shadow.color[1] ));
 sg13g2_dfrbp_1 _3728_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net32),
    .D(net236),
    .Q_N(_0044_),
    .Q(\ydelta[0] ));
 sg13g2_dfrbp_1 _3729_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net12),
    .D(_0072_),
    .Q_N(_1816_),
    .Q(\ydelta[1] ));
 sg13g2_dfrbp_1 _3730_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net208),
    .D(_0073_),
    .Q_N(_1815_),
    .Q(\ydelta[2] ));
 sg13g2_dfrbp_1 _3731_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net206),
    .D(_0074_),
    .Q_N(_1814_),
    .Q(\ydelta[3] ));
 sg13g2_dfrbp_1 _3732_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net204),
    .D(_0075_),
    .Q_N(_1813_),
    .Q(\ydelta[4] ));
 sg13g2_dfrbp_1 _3733_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net202),
    .D(_0076_),
    .Q_N(_1812_),
    .Q(\ydelta[5] ));
 sg13g2_dfrbp_1 _3734_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net200),
    .D(_0077_),
    .Q_N(_1811_),
    .Q(\ydelta[6] ));
 sg13g2_dfrbp_1 _3735_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net198),
    .D(net394),
    .Q_N(_0043_),
    .Q(\ydelta[7] ));
 sg13g2_dfrbp_1 _3736_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net194),
    .D(_0079_),
    .Q_N(_0067_),
    .Q(\pxm[0] ));
 sg13g2_dfrbp_1 _3737_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net192),
    .D(_0080_),
    .Q_N(_1810_),
    .Q(\pxm[1] ));
 sg13g2_dfrbp_1 _3738_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net190),
    .D(_0081_),
    .Q_N(_0045_),
    .Q(\px[0] ));
 sg13g2_dfrbp_1 _3739_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net188),
    .D(_0082_),
    .Q_N(_1809_),
    .Q(\px[1] ));
 sg13g2_dfrbp_1 _3740_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net186),
    .D(_0083_),
    .Q_N(_1808_),
    .Q(\px[2] ));
 sg13g2_dfrbp_1 _3741_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net184),
    .D(_0084_),
    .Q_N(_1807_),
    .Q(\px[3] ));
 sg13g2_dfrbp_1 _3742_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net182),
    .D(_0085_),
    .Q_N(_1806_),
    .Q(\px[4] ));
 sg13g2_dfrbp_1 _3743_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net180),
    .D(_0086_),
    .Q_N(_1805_),
    .Q(\px[5] ));
 sg13g2_dfrbp_1 _3744_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net178),
    .D(_0087_),
    .Q_N(_1804_),
    .Q(\px[6] ));
 sg13g2_dfrbp_1 _3745_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net176),
    .D(_0088_),
    .Q_N(_0059_),
    .Q(\px[7] ));
 sg13g2_dfrbp_1 _3746_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net174),
    .D(_0089_),
    .Q_N(_1803_),
    .Q(\px[8] ));
 sg13g2_dfrbp_1 _3747_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net172),
    .D(_0090_),
    .Q_N(_1802_),
    .Q(\px[9] ));
 sg13g2_dfrbp_1 _3748_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net168),
    .D(net523),
    .Q_N(_1801_),
    .Q(\py[0] ));
 sg13g2_dfrbp_1 _3749_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net166),
    .D(_0092_),
    .Q_N(_1800_),
    .Q(\py[1] ));
 sg13g2_dfrbp_1 _3750_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net164),
    .D(_0093_),
    .Q_N(_1799_),
    .Q(\py[2] ));
 sg13g2_dfrbp_1 _3751_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net162),
    .D(_0094_),
    .Q_N(_1798_),
    .Q(\py[3] ));
 sg13g2_dfrbp_1 _3752_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net160),
    .D(_0095_),
    .Q_N(_1797_),
    .Q(\py[4] ));
 sg13g2_dfrbp_1 _3753_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net158),
    .D(_0096_),
    .Q_N(_1796_),
    .Q(\py[5] ));
 sg13g2_dfrbp_1 _3754_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net157),
    .D(_0097_),
    .Q_N(_1795_),
    .Q(\py[6] ));
 sg13g2_dfrbp_1 _3755_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net155),
    .D(_0098_),
    .Q_N(_0022_),
    .Q(\py[7] ));
 sg13g2_dfrbp_1 _3756_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net154),
    .D(_0099_),
    .Q_N(_1794_),
    .Q(\py[8] ));
 sg13g2_dfrbp_1 _3757_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net152),
    .D(_0100_),
    .Q_N(_1793_),
    .Q(\py[9] ));
 sg13g2_dfrbp_1 _3758_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net151),
    .D(_0101_),
    .Q_N(_1792_),
    .Q(\pym[10] ));
 sg13g2_dfrbp_1 _3759_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net149),
    .D(_0102_),
    .Q_N(_1791_),
    .Q(\pym[11] ));
 sg13g2_dfrbp_1 _3760_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net147),
    .D(_0103_),
    .Q_N(_1790_),
    .Q(product_comp_dir));
 sg13g2_dfrbp_1 _3761_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net67),
    .D(_0104_),
    .Q_N(_1839_),
    .Q(dx));
 sg13g2_dfrbp_1 _3762_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net68),
    .D(_0019_),
    .Q_N(_1840_),
    .Q(\matt_venn_vga_shadow.font_0.dout[1] ));
 sg13g2_dfrbp_1 _3763_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net169),
    .D(_0020_),
    .Q_N(_1841_),
    .Q(\matt_venn_vga_shadow.font_0.dout[2] ));
 sg13g2_dfrbp_1 _3764_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net145),
    .D(_0021_),
    .Q_N(_1789_),
    .Q(\matt_venn_vga_shadow.font_0.dout[3] ));
 sg13g2_dfrbp_1 _3765_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net143),
    .D(_0105_),
    .Q_N(_1788_),
    .Q(\matt_venn_vga.color[2] ));
 sg13g2_dfrbp_1 _3766_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net142),
    .D(_0106_),
    .Q_N(_0058_),
    .Q(\vga_sync.hsync ));
 sg13g2_dfrbp_1 _3767_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net141),
    .D(_0107_),
    .Q_N(_1787_),
    .Q(\matt_venn_vga.y_px[0] ));
 sg13g2_dfrbp_1 _3768_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net139),
    .D(_0108_),
    .Q_N(_1786_),
    .Q(\matt_venn_vga.y_px[1] ));
 sg13g2_dfrbp_1 _3769_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net137),
    .D(_0109_),
    .Q_N(_0026_),
    .Q(\matt_venn_vga.y_px[2] ));
 sg13g2_dfrbp_1 _3770_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net135),
    .D(net406),
    .Q_N(_0027_),
    .Q(\matt_venn_vga.y_px[3] ));
 sg13g2_dfrbp_1 _3771_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net133),
    .D(_0111_),
    .Q_N(_0025_),
    .Q(\matt_venn_vga.y_px[4] ));
 sg13g2_dfrbp_1 _3772_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net131),
    .D(net502),
    .Q_N(_0057_),
    .Q(\matt_venn_vga.y_px[5] ));
 sg13g2_dfrbp_1 _3773_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net129),
    .D(_0113_),
    .Q_N(_0024_),
    .Q(\matt_venn_vga.y_px[6] ));
 sg13g2_dfrbp_1 _3774_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net127),
    .D(_0114_),
    .Q_N(_0031_),
    .Q(\matt_venn_vga.y_px[7] ));
 sg13g2_dfrbp_1 _3775_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net125),
    .D(_0115_),
    .Q_N(_0023_),
    .Q(\matt_venn_vga.y_px[8] ));
 sg13g2_dfrbp_1 _3776_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net123),
    .D(net490),
    .Q_N(_0052_),
    .Q(\matt_venn_vga.y_px[9] ));
 sg13g2_dfrbp_1 _3777_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net121),
    .D(_0117_),
    .Q_N(_1785_),
    .Q(\vga_sync.vsync ));
 sg13g2_dfrbp_1 _3778_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net120),
    .D(_0118_),
    .Q_N(_1784_),
    .Q(\matt_venn_vga_shadow.col_index[0] ));
 sg13g2_dfrbp_1 _3779_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net119),
    .D(_0119_),
    .Q_N(_1783_),
    .Q(\matt_venn_vga_shadow.col_index[1] ));
 sg13g2_dfrbp_1 _3780_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net118),
    .D(_0120_),
    .Q_N(_1782_),
    .Q(\matt_venn_vga_shadow.color[2] ));
 sg13g2_dfrbp_1 _3781_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net117),
    .D(_0121_),
    .Q_N(_0066_),
    .Q(\h[0] ));
 sg13g2_dfrbp_1 _3782_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net116),
    .D(net506),
    .Q_N(_1781_),
    .Q(\h[1] ));
 sg13g2_dfrbp_1 _3783_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net115),
    .D(_0123_),
    .Q_N(_1780_),
    .Q(\h[2] ));
 sg13g2_dfrbp_1 _3784_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net114),
    .D(_0124_),
    .Q_N(_1779_),
    .Q(\h[3] ));
 sg13g2_dfrbp_1 _3785_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net113),
    .D(_0125_),
    .Q_N(_1778_),
    .Q(\h[4] ));
 sg13g2_dfrbp_1 _3786_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net112),
    .D(_0126_),
    .Q_N(_1777_),
    .Q(\h[5] ));
 sg13g2_dfrbp_1 _3787_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net111),
    .D(_0127_),
    .Q_N(\matt_venn_vga.digit_0.char[0] ),
    .Q(\h[6] ));
 sg13g2_dfrbp_1 _3788_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net110),
    .D(_0128_),
    .Q_N(_1776_),
    .Q(\h[7] ));
 sg13g2_dfrbp_1 _3789_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net109),
    .D(_0129_),
    .Q_N(_0050_),
    .Q(\h[8] ));
 sg13g2_dfrbp_1 _3790_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net108),
    .D(_0130_),
    .Q_N(_1775_),
    .Q(\h[9] ));
 sg13g2_dfrbp_1 _3791_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net107),
    .D(_0131_),
    .Q_N(_1774_),
    .Q(\matt_venn_clock.pulse_hrs.comp[0] ));
 sg13g2_dfrbp_1 _3792_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net105),
    .D(_0132_),
    .Q_N(_1773_),
    .Q(\matt_venn_clock.pulse_hrs.comp[1] ));
 sg13g2_dfrbp_1 _3793_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net103),
    .D(net465),
    .Q_N(_1772_),
    .Q(\matt_venn_clock.pulse_hrs.comp[2] ));
 sg13g2_dfrbp_1 _3794_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net101),
    .D(_0134_),
    .Q_N(_1771_),
    .Q(\matt_venn_clock.pulse_hrs.comp[3] ));
 sg13g2_dfrbp_1 _3795_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net99),
    .D(_0135_),
    .Q_N(_1770_),
    .Q(\matt_venn_clock.pulse_hrs.comp[4] ));
 sg13g2_dfrbp_1 _3796_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net97),
    .D(_0136_),
    .Q_N(_1769_),
    .Q(\matt_venn_clock.pulse_hrs.count[0] ));
 sg13g2_dfrbp_1 _3797_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net95),
    .D(net437),
    .Q_N(_1768_),
    .Q(\matt_venn_clock.pulse_hrs.count[1] ));
 sg13g2_dfrbp_1 _3798_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net93),
    .D(net396),
    .Q_N(_1767_),
    .Q(\matt_venn_clock.pulse_hrs.count[2] ));
 sg13g2_dfrbp_1 _3799_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net91),
    .D(net270),
    .Q_N(_1766_),
    .Q(\matt_venn_clock.pulse_hrs.count[3] ));
 sg13g2_dfrbp_1 _3800_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net89),
    .D(net255),
    .Q_N(_0056_),
    .Q(\matt_venn_clock.pulse_hrs.count[4] ));
 sg13g2_dfrbp_1 _3801_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net87),
    .D(_0141_),
    .Q_N(_1765_),
    .Q(\matt_venn_clock.pulse_min.comp[0] ));
 sg13g2_dfrbp_1 _3802_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net85),
    .D(_0142_),
    .Q_N(_1764_),
    .Q(\matt_venn_clock.pulse_min.comp[1] ));
 sg13g2_dfrbp_1 _3803_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net83),
    .D(_0143_),
    .Q_N(_1763_),
    .Q(\matt_venn_clock.pulse_min.comp[2] ));
 sg13g2_dfrbp_1 _3804_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net81),
    .D(_0144_),
    .Q_N(_1762_),
    .Q(\matt_venn_clock.pulse_min.comp[3] ));
 sg13g2_dfrbp_1 _3805_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net79),
    .D(net415),
    .Q_N(_1761_),
    .Q(\matt_venn_clock.pulse_min.comp[4] ));
 sg13g2_dfrbp_1 _3806_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net77),
    .D(_0146_),
    .Q_N(_1760_),
    .Q(\matt_venn_clock.pulse_min.count[0] ));
 sg13g2_dfrbp_1 _3807_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net76),
    .D(net448),
    .Q_N(_1759_),
    .Q(\matt_venn_clock.pulse_min.count[1] ));
 sg13g2_dfrbp_1 _3808_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net75),
    .D(net423),
    .Q_N(_1758_),
    .Q(\matt_venn_clock.pulse_min.count[2] ));
 sg13g2_dfrbp_1 _3809_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net74),
    .D(net426),
    .Q_N(_1757_),
    .Q(\matt_venn_clock.pulse_min.count[3] ));
 sg13g2_dfrbp_1 _3810_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net73),
    .D(net252),
    .Q_N(_0055_),
    .Q(\matt_venn_clock.pulse_min.count[4] ));
 sg13g2_dfrbp_1 _3811_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net72),
    .D(_0151_),
    .Q_N(_1756_),
    .Q(\matt_venn_clock.pulse_sec.comp[0] ));
 sg13g2_dfrbp_1 _3812_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net70),
    .D(_0152_),
    .Q_N(_1755_),
    .Q(\matt_venn_clock.pulse_sec.comp[1] ));
 sg13g2_dfrbp_1 _3813_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net65),
    .D(net442),
    .Q_N(_1754_),
    .Q(\matt_venn_clock.pulse_sec.comp[2] ));
 sg13g2_dfrbp_1 _3814_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net63),
    .D(_0154_),
    .Q_N(_1753_),
    .Q(\matt_venn_clock.pulse_sec.comp[3] ));
 sg13g2_dfrbp_1 _3815_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net61),
    .D(net385),
    .Q_N(_1752_),
    .Q(\matt_venn_clock.pulse_sec.comp[4] ));
 sg13g2_dfrbp_1 _3816_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net59),
    .D(net488),
    .Q_N(_1751_),
    .Q(\matt_venn_clock.pulse_sec.count[0] ));
 sg13g2_dfrbp_1 _3817_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net57),
    .D(net446),
    .Q_N(_1750_),
    .Q(\matt_venn_clock.pulse_sec.count[1] ));
 sg13g2_dfrbp_1 _3818_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net55),
    .D(net430),
    .Q_N(_1749_),
    .Q(\matt_venn_clock.pulse_sec.count[2] ));
 sg13g2_dfrbp_1 _3819_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net53),
    .D(_0159_),
    .Q_N(_1748_),
    .Q(\matt_venn_clock.pulse_sec.count[3] ));
 sg13g2_dfrbp_1 _3820_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net52),
    .D(net247),
    .Q_N(_0054_),
    .Q(\matt_venn_clock.pulse_sec.count[4] ));
 sg13g2_dfrbp_1 _3821_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net50),
    .D(net222),
    .Q_N(_0065_),
    .Q(\clock_color_offset[0] ));
 sg13g2_dfrbp_1 _3822_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net49),
    .D(_0162_),
    .Q_N(_0051_),
    .Q(\clock_color_offset[1] ));
 sg13g2_dfrbp_1 _3823_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net47),
    .D(net373),
    .Q_N(_1747_),
    .Q(\clock_color_offset[2] ));
 sg13g2_dfrbp_1 _3824_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net45),
    .D(net227),
    .Q_N(_0064_),
    .Q(\clock_hrs_d[0] ));
 sg13g2_dfrbp_1 _3825_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net43),
    .D(_0165_),
    .Q_N(_0041_),
    .Q(\clock_hrs_d[1] ));
 sg13g2_dfrbp_1 _3826_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net41),
    .D(_0166_),
    .Q_N(_0047_),
    .Q(\clock_hrs_u[0] ));
 sg13g2_dfrbp_1 _3827_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net39),
    .D(_0167_),
    .Q_N(_0042_),
    .Q(\clock_hrs_u[1] ));
 sg13g2_dfrbp_1 _3828_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net37),
    .D(net459),
    .Q_N(_0036_),
    .Q(\clock_hrs_u[2] ));
 sg13g2_dfrbp_1 _3829_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net31),
    .D(_0169_),
    .Q_N(_0033_),
    .Q(\clock_hrs_u[3] ));
 sg13g2_dfrbp_1 _3830_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net207),
    .D(net224),
    .Q_N(_0063_),
    .Q(\clock_min_d[0] ));
 sg13g2_dfrbp_1 _3831_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net203),
    .D(net496),
    .Q_N(_1746_),
    .Q(\clock_min_d[1] ));
 sg13g2_dfrbp_1 _3832_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net199),
    .D(net402),
    .Q_N(_0037_),
    .Q(\clock_min_d[2] ));
 sg13g2_dfrbp_1 _3833_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net193),
    .D(_0173_),
    .Q_N(_0046_),
    .Q(\clock_min_u[0] ));
 sg13g2_dfrbp_1 _3834_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net189),
    .D(_0174_),
    .Q_N(_1745_),
    .Q(\clock_min_u[1] ));
 sg13g2_dfrbp_1 _3835_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net185),
    .D(_0175_),
    .Q_N(_0038_),
    .Q(\clock_min_u[2] ));
 sg13g2_dfrbp_1 _3836_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net181),
    .D(net376),
    .Q_N(_0034_),
    .Q(\clock_min_u[3] ));
 sg13g2_dfrbp_1 _3837_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net177),
    .D(net392),
    .Q_N(_0062_),
    .Q(\clock_sec_d[0] ));
 sg13g2_dfrbp_1 _3838_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net173),
    .D(_0178_),
    .Q_N(_1744_),
    .Q(\clock_sec_d[1] ));
 sg13g2_dfrbp_1 _3839_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net167),
    .D(_0179_),
    .Q_N(_0039_),
    .Q(\clock_sec_d[2] ));
 sg13g2_dfrbp_1 _3840_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net163),
    .D(_0180_),
    .Q_N(_0032_),
    .Q(\clock_sec_u[0] ));
 sg13g2_dfrbp_1 _3841_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net159),
    .D(_0181_),
    .Q_N(_1743_),
    .Q(\clock_sec_u[1] ));
 sg13g2_dfrbp_1 _3842_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net156),
    .D(net274),
    .Q_N(_0040_),
    .Q(\clock_sec_u[2] ));
 sg13g2_dfrbp_1 _3843_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net153),
    .D(_0183_),
    .Q_N(_0035_),
    .Q(\clock_sec_u[3] ));
 sg13g2_dfrbp_1 _3844_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net150),
    .D(_0184_),
    .Q_N(_1742_),
    .Q(\matt_venn_vga.color[3] ));
 sg13g2_dfrbp_1 _3845_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net148),
    .D(_0185_),
    .Q_N(_1741_),
    .Q(\matt_venn_vga.color[0] ));
 sg13g2_dfrbp_1 _3846_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net146),
    .D(_0186_),
    .Q_N(_1740_),
    .Q(\matt_venn_vga.color[1] ));
 sg13g2_dfrbp_1 _3847_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net144),
    .D(net243),
    .Q_N(_1739_),
    .Q(\matt_venn_vga.draw ));
 sg13g2_dfrbp_1 _3848_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net140),
    .D(_0188_),
    .Q_N(_0061_),
    .Q(\matt_venn_clock.sec_counter[0] ));
 sg13g2_dfrbp_1 _3849_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net138),
    .D(_0189_),
    .Q_N(_1738_),
    .Q(\matt_venn_clock.sec_counter[1] ));
 sg13g2_dfrbp_1 _3850_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net136),
    .D(net234),
    .Q_N(_1737_),
    .Q(\matt_venn_clock.sec_counter[2] ));
 sg13g2_dfrbp_1 _3851_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net134),
    .D(_0191_),
    .Q_N(_1736_),
    .Q(\matt_venn_clock.sec_counter[3] ));
 sg13g2_dfrbp_1 _3852_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net132),
    .D(_0192_),
    .Q_N(_1735_),
    .Q(\matt_venn_clock.sec_counter[4] ));
 sg13g2_dfrbp_1 _3853_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net130),
    .D(_0193_),
    .Q_N(_1734_),
    .Q(\matt_venn_clock.sec_counter[5] ));
 sg13g2_dfrbp_1 _3854_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net128),
    .D(_0194_),
    .Q_N(_1733_),
    .Q(\matt_venn_clock.sec_counter[6] ));
 sg13g2_dfrbp_1 _3855_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net126),
    .D(_0195_),
    .Q_N(_1732_),
    .Q(\matt_venn_clock.sec_counter[7] ));
 sg13g2_dfrbp_1 _3856_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net124),
    .D(_0196_),
    .Q_N(_1731_),
    .Q(\matt_venn_clock.sec_counter[8] ));
 sg13g2_dfrbp_1 _3857_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net122),
    .D(_0197_),
    .Q_N(_1730_),
    .Q(\matt_venn_clock.sec_counter[9] ));
 sg13g2_dfrbp_1 _3858_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net106),
    .D(_0198_),
    .Q_N(_1729_),
    .Q(\matt_venn_clock.sec_counter[10] ));
 sg13g2_dfrbp_1 _3859_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net104),
    .D(_0199_),
    .Q_N(_1728_),
    .Q(\matt_venn_clock.sec_counter[11] ));
 sg13g2_dfrbp_1 _3860_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net102),
    .D(_0200_),
    .Q_N(_0048_),
    .Q(\matt_venn_clock.sec_counter[12] ));
 sg13g2_dfrbp_1 _3861_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net100),
    .D(_0201_),
    .Q_N(_1727_),
    .Q(\matt_venn_clock.sec_counter[13] ));
 sg13g2_dfrbp_1 _3862_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net98),
    .D(_0202_),
    .Q_N(_1726_),
    .Q(\matt_venn_clock.sec_counter[14] ));
 sg13g2_dfrbp_1 _3863_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net96),
    .D(_0203_),
    .Q_N(_1725_),
    .Q(\matt_venn_clock.sec_counter[15] ));
 sg13g2_dfrbp_1 _3864_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net94),
    .D(_0204_),
    .Q_N(_1724_),
    .Q(\matt_venn_clock.sec_counter[16] ));
 sg13g2_dfrbp_1 _3865_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net92),
    .D(_0205_),
    .Q_N(_1723_),
    .Q(\matt_venn_clock.sec_counter[17] ));
 sg13g2_dfrbp_1 _3866_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net90),
    .D(_0206_),
    .Q_N(_0049_),
    .Q(\matt_venn_clock.sec_counter[18] ));
 sg13g2_dfrbp_1 _3867_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net88),
    .D(_0207_),
    .Q_N(_1722_),
    .Q(\matt_venn_clock.sec_counter[19] ));
 sg13g2_dfrbp_1 _3868_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net86),
    .D(_0208_),
    .Q_N(_1721_),
    .Q(\matt_venn_clock.sec_counter[20] ));
 sg13g2_dfrbp_1 _3869_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net84),
    .D(_0209_),
    .Q_N(_1720_),
    .Q(\matt_venn_clock.sec_counter[21] ));
 sg13g2_dfrbp_1 _3870_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net82),
    .D(_0210_),
    .Q_N(_1719_),
    .Q(\matt_venn_clock.sec_counter[22] ));
 sg13g2_dfrbp_1 _3871_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net80),
    .D(net262),
    .Q_N(_1718_),
    .Q(\matt_venn_clock.sec_counter[23] ));
 sg13g2_dfrbp_1 _3872_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net170),
    .D(_0212_),
    .Q_N(_1842_),
    .Q(\matt_venn_clock.sec_counter[24] ));
 sg13g2_dfrbp_1 _3873_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net196),
    .D(net218),
    .Q_N(_1843_),
    .Q(\matt_venn_vga.col_index_q[0] ));
 sg13g2_dfrbp_1 _3874_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net78),
    .D(net217),
    .Q_N(_1717_),
    .Q(\matt_venn_vga.col_index_q[1] ));
 sg13g2_dfrbp_1 _3875_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net71),
    .D(_0213_),
    .Q_N(_1716_),
    .Q(\matt_venn_vga.x_block_q[5] ));
 sg13g2_dfrbp_1 _3876_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net69),
    .D(_0214_),
    .Q_N(_1715_),
    .Q(\matt_venn_vga.y_block_q[0] ));
 sg13g2_dfrbp_1 _3877_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net64),
    .D(_0215_),
    .Q_N(_1714_),
    .Q(\matt_venn_vga.y_block_q[1] ));
 sg13g2_dfrbp_1 _3878_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net62),
    .D(_0216_),
    .Q_N(_1713_),
    .Q(\matt_venn_vga.y_block_q[2] ));
 sg13g2_dfrbp_1 _3879_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net60),
    .D(_0217_),
    .Q_N(_1712_),
    .Q(\matt_venn_vga.y_block_q[3] ));
 sg13g2_dfrbp_1 _3880_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net58),
    .D(_0218_),
    .Q_N(_1711_),
    .Q(\matt_venn_vga.y_block_q[4] ));
 sg13g2_dfrbp_1 _3881_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net56),
    .D(_0219_),
    .Q_N(_1710_),
    .Q(\matt_venn_vga.y_block_q[5] ));
 sg13g2_dfrbp_1 _3882_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net54),
    .D(net231),
    .Q_N(_0060_),
    .Q(\product_comp[1] ));
 sg13g2_dfrbp_1 _3883_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net51),
    .D(net428),
    .Q_N(_1709_),
    .Q(\product_comp[2] ));
 sg13g2_dfrbp_1 _3884_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net48),
    .D(_0222_),
    .Q_N(_0030_),
    .Q(\product_comp[3] ));
 sg13g2_dfrbp_1 _3885_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net44),
    .D(_0223_),
    .Q_N(_1708_),
    .Q(\product_comp[4] ));
 sg13g2_dfrbp_1 _3886_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net40),
    .D(_0224_),
    .Q_N(_1707_),
    .Q(\product_comp[5] ));
 sg13g2_dfrbp_1 _3887_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net36),
    .D(_0225_),
    .Q_N(_1706_),
    .Q(\product_comp[6] ));
 sg13g2_dfrbp_1 _3888_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net205),
    .D(_0226_),
    .Q_N(_0029_),
    .Q(\product_comp[7] ));
 sg13g2_dfrbp_1 _3889_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net195),
    .D(_0227_),
    .Q_N(_1705_),
    .Q(\product_comp[8] ));
 sg13g2_dfrbp_1 _3890_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net187),
    .D(_0228_),
    .Q_N(_0028_),
    .Q(\product_comp[9] ));
 sg13g2_dfrbp_1 _3891_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net179),
    .D(_0229_),
    .Q_N(_0053_),
    .Q(\product_comp[10] ));
 sg13g2_dfrbp_1 _3892_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net171),
    .D(net259),
    .Q_N(_1704_),
    .Q(\matt_venn_vga_shadow.draw ));
 sg13g2_dfrbp_1 _3893_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net165),
    .D(_0231_),
    .Q_N(_1703_),
    .Q(\matt_venn_vga.col_index[0] ));
 sg13g2_dfrbp_1 _3894_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net197),
    .D(_0232_),
    .Q_N(_1844_),
    .Q(\matt_venn_vga.col_index[1] ));
 sg13g2_dfrbp_1 _3895_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net175),
    .D(net216),
    .Q_N(_1845_),
    .Q(\matt_venn_vga_shadow.col_index_q[0] ));
 sg13g2_dfrbp_1 _3896_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net161),
    .D(net215),
    .Q_N(_1702_),
    .Q(\matt_venn_vga_shadow.col_index_q[1] ));
 sg13g2_dfrbp_1 _3897_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net46),
    .D(_0233_),
    .Q_N(_1701_),
    .Q(\matt_venn_vga_shadow.x_block_q[5] ));
 sg13g2_dfrbp_1 _3898_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net42),
    .D(_0234_),
    .Q_N(_1700_),
    .Q(\matt_venn_vga_shadow.y_block_q[0] ));
 sg13g2_dfrbp_1 _3899_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net38),
    .D(_0235_),
    .Q_N(_1699_),
    .Q(\matt_venn_vga_shadow.y_block_q[1] ));
 sg13g2_dfrbp_1 _3900_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net209),
    .D(_0236_),
    .Q_N(_1698_),
    .Q(\matt_venn_vga_shadow.y_block_q[2] ));
 sg13g2_dfrbp_1 _3901_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net201),
    .D(_0237_),
    .Q_N(_1697_),
    .Q(\matt_venn_vga_shadow.y_block_q[3] ));
 sg13g2_dfrbp_1 _3902_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net191),
    .D(_0238_),
    .Q_N(_1696_),
    .Q(\matt_venn_vga_shadow.y_block_q[4] ));
 sg13g2_dfrbp_1 _3903_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net183),
    .D(_0239_),
    .Q_N(_1695_),
    .Q(\matt_venn_vga_shadow.y_block_q[5] ));
 sg13g2_tiehi _3724__13 (.L_HI(net13));
 sg13g2_tiehi _3706__14 (.L_HI(net14));
 sg13g2_tiehi _3707__15 (.L_HI(net15));
 sg13g2_tiehi _3708__16 (.L_HI(net16));
 sg13g2_tiehi _3709__17 (.L_HI(net17));
 sg13g2_tiehi _3710__18 (.L_HI(net18));
 sg13g2_tiehi _3711__19 (.L_HI(net19));
 sg13g2_tiehi _3712__20 (.L_HI(net20));
 sg13g2_tiehi _3713__21 (.L_HI(net21));
 sg13g2_tiehi _3714__22 (.L_HI(net22));
 sg13g2_tiehi _3715__23 (.L_HI(net23));
 sg13g2_tiehi _3716__24 (.L_HI(net24));
 sg13g2_tiehi _3717__25 (.L_HI(net25));
 sg13g2_tiehi _3718__26 (.L_HI(net26));
 sg13g2_tiehi _3719__27 (.L_HI(net27));
 sg13g2_tiehi _3720__28 (.L_HI(net28));
 sg13g2_tiehi _3721__29 (.L_HI(net29));
 sg13g2_tiehi _3722__30 (.L_HI(net30));
 sg13g2_tiehi _3829__31 (.L_HI(net31));
 sg13g2_tiehi _3728__32 (.L_HI(net32));
 sg13g2_tiehi _3727__33 (.L_HI(net33));
 sg13g2_tiehi _3726__34 (.L_HI(net34));
 sg13g2_tiehi _3725__35 (.L_HI(net35));
 sg13g2_tiehi _3887__36 (.L_HI(net36));
 sg13g2_tiehi _3828__37 (.L_HI(net37));
 sg13g2_tiehi _3899__38 (.L_HI(net38));
 sg13g2_tiehi _3827__39 (.L_HI(net39));
 sg13g2_tiehi _3886__40 (.L_HI(net40));
 sg13g2_tiehi _3826__41 (.L_HI(net41));
 sg13g2_tiehi _3898__42 (.L_HI(net42));
 sg13g2_tiehi _3825__43 (.L_HI(net43));
 sg13g2_tiehi _3885__44 (.L_HI(net44));
 sg13g2_tiehi _3824__45 (.L_HI(net45));
 sg13g2_tiehi _3897__46 (.L_HI(net46));
 sg13g2_tiehi _3823__47 (.L_HI(net47));
 sg13g2_tiehi _3884__48 (.L_HI(net48));
 sg13g2_tiehi _3822__49 (.L_HI(net49));
 sg13g2_tiehi _3821__50 (.L_HI(net50));
 sg13g2_tiehi _3883__51 (.L_HI(net51));
 sg13g2_tiehi _3820__52 (.L_HI(net52));
 sg13g2_tiehi _3819__53 (.L_HI(net53));
 sg13g2_tiehi _3882__54 (.L_HI(net54));
 sg13g2_tiehi _3818__55 (.L_HI(net55));
 sg13g2_tiehi _3881__56 (.L_HI(net56));
 sg13g2_tiehi _3817__57 (.L_HI(net57));
 sg13g2_tiehi _3880__58 (.L_HI(net58));
 sg13g2_tiehi _3816__59 (.L_HI(net59));
 sg13g2_tiehi _3879__60 (.L_HI(net60));
 sg13g2_tiehi _3815__61 (.L_HI(net61));
 sg13g2_tiehi _3878__62 (.L_HI(net62));
 sg13g2_tiehi _3814__63 (.L_HI(net63));
 sg13g2_tiehi _3877__64 (.L_HI(net64));
 sg13g2_tiehi _3813__65 (.L_HI(net65));
 sg13g2_tiehi _3723__66 (.L_HI(net66));
 sg13g2_tiehi _3761__67 (.L_HI(net67));
 sg13g2_tiehi _3762__68 (.L_HI(net68));
 sg13g2_tiehi _3876__69 (.L_HI(net69));
 sg13g2_tiehi _3812__70 (.L_HI(net70));
 sg13g2_tiehi _3875__71 (.L_HI(net71));
 sg13g2_tiehi _3811__72 (.L_HI(net72));
 sg13g2_tiehi _3810__73 (.L_HI(net73));
 sg13g2_tiehi _3809__74 (.L_HI(net74));
 sg13g2_tiehi _3808__75 (.L_HI(net75));
 sg13g2_tiehi _3807__76 (.L_HI(net76));
 sg13g2_tiehi _3806__77 (.L_HI(net77));
 sg13g2_tiehi _3874__78 (.L_HI(net78));
 sg13g2_tiehi _3805__79 (.L_HI(net79));
 sg13g2_tiehi _3871__80 (.L_HI(net80));
 sg13g2_tiehi _3804__81 (.L_HI(net81));
 sg13g2_tiehi _3870__82 (.L_HI(net82));
 sg13g2_tiehi _3803__83 (.L_HI(net83));
 sg13g2_tiehi _3869__84 (.L_HI(net84));
 sg13g2_tiehi _3802__85 (.L_HI(net85));
 sg13g2_tiehi _3868__86 (.L_HI(net86));
 sg13g2_tiehi _3801__87 (.L_HI(net87));
 sg13g2_tiehi _3867__88 (.L_HI(net88));
 sg13g2_tiehi _3800__89 (.L_HI(net89));
 sg13g2_tiehi _3866__90 (.L_HI(net90));
 sg13g2_tiehi _3799__91 (.L_HI(net91));
 sg13g2_tiehi _3865__92 (.L_HI(net92));
 sg13g2_tiehi _3798__93 (.L_HI(net93));
 sg13g2_tiehi _3864__94 (.L_HI(net94));
 sg13g2_tiehi _3797__95 (.L_HI(net95));
 sg13g2_tiehi _3863__96 (.L_HI(net96));
 sg13g2_tiehi _3796__97 (.L_HI(net97));
 sg13g2_tiehi _3862__98 (.L_HI(net98));
 sg13g2_tiehi _3795__99 (.L_HI(net99));
 sg13g2_tiehi _3861__100 (.L_HI(net100));
 sg13g2_tiehi _3794__101 (.L_HI(net101));
 sg13g2_tiehi _3860__102 (.L_HI(net102));
 sg13g2_tiehi _3793__103 (.L_HI(net103));
 sg13g2_tiehi _3859__104 (.L_HI(net104));
 sg13g2_tiehi _3792__105 (.L_HI(net105));
 sg13g2_tiehi _3858__106 (.L_HI(net106));
 sg13g2_tiehi _3791__107 (.L_HI(net107));
 sg13g2_tiehi _3790__108 (.L_HI(net108));
 sg13g2_tiehi _3789__109 (.L_HI(net109));
 sg13g2_tiehi _3788__110 (.L_HI(net110));
 sg13g2_tiehi _3787__111 (.L_HI(net111));
 sg13g2_tiehi _3786__112 (.L_HI(net112));
 sg13g2_tiehi _3785__113 (.L_HI(net113));
 sg13g2_tiehi _3784__114 (.L_HI(net114));
 sg13g2_tiehi _3783__115 (.L_HI(net115));
 sg13g2_tiehi _3782__116 (.L_HI(net116));
 sg13g2_tiehi _3781__117 (.L_HI(net117));
 sg13g2_tiehi _3780__118 (.L_HI(net118));
 sg13g2_tiehi _3779__119 (.L_HI(net119));
 sg13g2_tiehi _3778__120 (.L_HI(net120));
 sg13g2_tiehi _3777__121 (.L_HI(net121));
 sg13g2_tiehi _3857__122 (.L_HI(net122));
 sg13g2_tiehi _3776__123 (.L_HI(net123));
 sg13g2_tiehi _3856__124 (.L_HI(net124));
 sg13g2_tiehi _3775__125 (.L_HI(net125));
 sg13g2_tiehi _3855__126 (.L_HI(net126));
 sg13g2_tiehi _3774__127 (.L_HI(net127));
 sg13g2_tiehi _3854__128 (.L_HI(net128));
 sg13g2_tiehi _3773__129 (.L_HI(net129));
 sg13g2_tiehi _3853__130 (.L_HI(net130));
 sg13g2_tiehi _3772__131 (.L_HI(net131));
 sg13g2_tiehi _3852__132 (.L_HI(net132));
 sg13g2_tiehi _3771__133 (.L_HI(net133));
 sg13g2_tiehi _3851__134 (.L_HI(net134));
 sg13g2_tiehi _3770__135 (.L_HI(net135));
 sg13g2_tiehi _3850__136 (.L_HI(net136));
 sg13g2_tiehi _3769__137 (.L_HI(net137));
 sg13g2_tiehi _3849__138 (.L_HI(net138));
 sg13g2_tiehi _3768__139 (.L_HI(net139));
 sg13g2_tiehi _3848__140 (.L_HI(net140));
 sg13g2_tiehi _3767__141 (.L_HI(net141));
 sg13g2_tiehi _3766__142 (.L_HI(net142));
 sg13g2_tiehi _3765__143 (.L_HI(net143));
 sg13g2_tiehi _3847__144 (.L_HI(net144));
 sg13g2_tiehi _3764__145 (.L_HI(net145));
 sg13g2_tiehi _3846__146 (.L_HI(net146));
 sg13g2_tiehi _3760__147 (.L_HI(net147));
 sg13g2_tiehi _3845__148 (.L_HI(net148));
 sg13g2_tiehi _3759__149 (.L_HI(net149));
 sg13g2_tiehi _3844__150 (.L_HI(net150));
 sg13g2_tiehi _3758__151 (.L_HI(net151));
 sg13g2_tiehi _3757__152 (.L_HI(net152));
 sg13g2_tiehi _3843__153 (.L_HI(net153));
 sg13g2_tiehi _3756__154 (.L_HI(net154));
 sg13g2_tiehi _3755__155 (.L_HI(net155));
 sg13g2_tiehi _3842__156 (.L_HI(net156));
 sg13g2_tiehi _3754__157 (.L_HI(net157));
 sg13g2_tiehi _3753__158 (.L_HI(net158));
 sg13g2_tiehi _3841__159 (.L_HI(net159));
 sg13g2_tiehi _3752__160 (.L_HI(net160));
 sg13g2_tiehi _3896__161 (.L_HI(net161));
 sg13g2_tiehi _3751__162 (.L_HI(net162));
 sg13g2_tiehi _3840__163 (.L_HI(net163));
 sg13g2_tiehi _3750__164 (.L_HI(net164));
 sg13g2_tiehi _3893__165 (.L_HI(net165));
 sg13g2_tiehi _3749__166 (.L_HI(net166));
 sg13g2_tiehi _3839__167 (.L_HI(net167));
 sg13g2_tiehi _3748__168 (.L_HI(net168));
 sg13g2_tiehi _3763__169 (.L_HI(net169));
 sg13g2_tiehi _3872__170 (.L_HI(net170));
 sg13g2_tiehi _3892__171 (.L_HI(net171));
 sg13g2_tiehi _3747__172 (.L_HI(net172));
 sg13g2_tiehi _3838__173 (.L_HI(net173));
 sg13g2_tiehi _3746__174 (.L_HI(net174));
 sg13g2_tiehi _3895__175 (.L_HI(net175));
 sg13g2_tiehi _3745__176 (.L_HI(net176));
 sg13g2_tiehi _3837__177 (.L_HI(net177));
 sg13g2_tiehi _3744__178 (.L_HI(net178));
 sg13g2_tiehi _3891__179 (.L_HI(net179));
 sg13g2_tiehi _3743__180 (.L_HI(net180));
 sg13g2_tiehi _3836__181 (.L_HI(net181));
 sg13g2_tiehi _3742__182 (.L_HI(net182));
 sg13g2_tiehi _3903__183 (.L_HI(net183));
 sg13g2_tiehi _3741__184 (.L_HI(net184));
 sg13g2_tiehi _3835__185 (.L_HI(net185));
 sg13g2_tiehi _3740__186 (.L_HI(net186));
 sg13g2_tiehi _3890__187 (.L_HI(net187));
 sg13g2_tiehi _3739__188 (.L_HI(net188));
 sg13g2_tiehi _3834__189 (.L_HI(net189));
 sg13g2_tiehi _3738__190 (.L_HI(net190));
 sg13g2_tiehi _3902__191 (.L_HI(net191));
 sg13g2_tiehi _3737__192 (.L_HI(net192));
 sg13g2_tiehi _3833__193 (.L_HI(net193));
 sg13g2_tiehi _3736__194 (.L_HI(net194));
 sg13g2_tiehi _3889__195 (.L_HI(net195));
 sg13g2_tiehi _3873__196 (.L_HI(net196));
 sg13g2_tiehi _3894__197 (.L_HI(net197));
 sg13g2_tiehi _3735__198 (.L_HI(net198));
 sg13g2_tiehi _3832__199 (.L_HI(net199));
 sg13g2_tiehi _3734__200 (.L_HI(net200));
 sg13g2_tiehi _3901__201 (.L_HI(net201));
 sg13g2_tiehi _3733__202 (.L_HI(net202));
 sg13g2_tiehi _3831__203 (.L_HI(net203));
 sg13g2_tiehi _3732__204 (.L_HI(net204));
 sg13g2_tiehi _3888__205 (.L_HI(net205));
 sg13g2_tiehi _3731__206 (.L_HI(net206));
 sg13g2_tiehi _3830__207 (.L_HI(net207));
 sg13g2_tiehi _3730__208 (.L_HI(net208));
 sg13g2_tiehi _3900__209 (.L_HI(net209));
 sg13g2_tiehi tt_um_algofoogle_vga_210 (.L_HI(net210));
 sg13g2_tiehi tt_um_algofoogle_vga_211 (.L_HI(net211));
 sg13g2_tiehi tt_um_algofoogle_vga_212 (.L_HI(net212));
 sg13g2_tiehi tt_um_algofoogle_vga_213 (.L_HI(net213));
 sg13g2_tiehi tt_um_algofoogle_vga_214 (.L_HI(net214));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_algofoogle_vga_7 (.L_LO(net7));
 sg13g2_tielo tt_um_algofoogle_vga_8 (.L_LO(net8));
 sg13g2_tielo tt_um_algofoogle_vga_9 (.L_LO(net9));
 sg13g2_tielo tt_um_algofoogle_vga_10 (.L_LO(net10));
 sg13g2_tielo tt_um_algofoogle_vga_11 (.L_LO(net11));
 sg13g2_tiehi _3729__12 (.L_HI(net12));
 sg13g2_buf_2 _4113_ (.A(hmax),
    .X(uio_out[0]));
 sg13g2_buf_2 _4114_ (.A(\vga_sync.o_vmax ),
    .X(uio_out[1]));
 sg13g2_buf_2 _4115_ (.A(hblank),
    .X(uio_out[2]));
 sg13g2_buf_2 _4116_ (.A(vblank),
    .X(uio_out[3]));
 sg13g2_buf_2 _4117_ (.A(\matt_venn_vga.activevideo ),
    .X(uio_out[4]));
 sg13g2_buf_2 fanout276 (.A(net278),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(net278),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_1098_),
    .X(net278));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(net280));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(_0641_));
 sg13g2_buf_2 fanout281 (.A(_0513_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_0432_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_0501_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_1118_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(net286),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_0435_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(net288),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(net293),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(net293),
    .X(net290));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(net293));
 sg13g2_buf_4 fanout292 (.X(net292),
    .A(net293));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(_0635_));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(_0575_));
 sg13g2_buf_2 fanout295 (.A(_0496_),
    .X(net295));
 sg13g2_buf_4 fanout296 (.X(net296),
    .A(_0581_));
 sg13g2_buf_2 fanout297 (.A(_0433_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_1445_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_1438_),
    .X(net299));
 sg13g2_buf_1 fanout300 (.A(_1438_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_0306_),
    .X(net301));
 sg13g2_buf_4 fanout302 (.X(net302),
    .A(_1455_));
 sg13g2_buf_2 fanout303 (.A(_1009_),
    .X(net303));
 sg13g2_buf_4 fanout304 (.X(net304),
    .A(_1410_));
 sg13g2_buf_2 fanout305 (.A(\h[9] ),
    .X(net305));
 sg13g2_buf_4 fanout306 (.X(net306),
    .A(net308));
 sg13g2_buf_2 fanout307 (.A(net308),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(\h[7] ),
    .X(net308));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(net310));
 sg13g2_buf_2 fanout310 (.A(\h[6] ),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(net312),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(net511),
    .X(net312));
 sg13g2_buf_4 fanout313 (.X(net313),
    .A(net478));
 sg13g2_buf_2 fanout314 (.A(net478),
    .X(net314));
 sg13g2_buf_4 fanout315 (.X(net315),
    .A(net519));
 sg13g2_buf_4 fanout316 (.X(net316),
    .A(net505));
 sg13g2_buf_2 fanout317 (.A(net318),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(net489),
    .X(net318));
 sg13g2_buf_4 fanout319 (.X(net319),
    .A(net528));
 sg13g2_buf_2 fanout320 (.A(net321),
    .X(net320));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(\matt_venn_vga.y_px[7] ));
 sg13g2_buf_2 fanout322 (.A(net323),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(net512),
    .X(net323));
 sg13g2_buf_4 fanout324 (.X(net324),
    .A(net501));
 sg13g2_buf_2 fanout325 (.A(\matt_venn_vga.y_px[5] ),
    .X(net325));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(net532));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(net525));
 sg13g2_buf_2 fanout328 (.A(\matt_venn_vga.y_px[3] ),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(net509),
    .X(net329));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(\matt_venn_vga.y_px[2] ));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(net531));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(net518));
 sg13g2_buf_1 fanout333 (.A(\matt_venn_vga.y_px[0] ),
    .X(net333));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(net336));
 sg13g2_buf_2 fanout335 (.A(net336),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(dx),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(net338),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(product_comp_dir),
    .X(net338));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(net529));
 sg13g2_buf_2 fanout340 (.A(\py[1] ),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(net522),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(net534),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(net538),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(net517),
    .X(net344));
 sg13g2_buf_4 fanout345 (.X(net345),
    .A(net484));
 sg13g2_buf_1 fanout346 (.A(\px[1] ),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(\px[0] ),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(net349),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(\ydelta[7] ),
    .X(net349));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(net353));
 sg13g2_buf_2 fanout351 (.A(net353),
    .X(net351));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(net353));
 sg13g2_buf_2 fanout353 (.A(_1219_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(net355),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(ui_in[7]),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(net4),
    .X(net356));
 sg13g2_buf_4 fanout357 (.X(net357),
    .A(net361));
 sg13g2_buf_1 fanout358 (.A(net361),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(net360),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(net361),
    .X(net360));
 sg13g2_buf_4 fanout361 (.X(net361),
    .A(net367));
 sg13g2_buf_2 fanout362 (.A(net367),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(net367),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(net366),
    .X(net364));
 sg13g2_buf_4 fanout365 (.X(net365),
    .A(net366));
 sg13g2_buf_2 fanout366 (.A(net367),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(rst_n),
    .X(net367));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_tielo tt_um_algofoogle_vga_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_25__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\matt_venn_vga_shadow.col_index[1] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold2 (.A(\matt_venn_vga_shadow.col_index[0] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold3 (.A(\matt_venn_vga.col_index[1] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold4 (.A(\matt_venn_vga.col_index[0] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0061_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0066_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0065_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0161_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0063_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0170_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0064_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0988_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0164_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0067_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0656_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0060_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0220_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold18 (.A(\matt_venn_clock.sec_counter[2] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold19 (.A(_1100_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0190_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0045_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0071_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold23 (.A(\py[1] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold24 (.A(\matt_venn_clock.sec_counter[21] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold25 (.A(_1112_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold26 (.A(\matt_venn_vga.y_block_q[3] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold27 (.A(_1092_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold28 (.A(_1097_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0187_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold30 (.A(\matt_venn_clock.sec_counter[5] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold31 (.A(_1103_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold32 (.A(\matt_venn_clock.pulse_sec.count[4] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0160_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold34 (.A(\clock_min_u[2] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold35 (.A(_1029_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold36 (.A(\pxm[1] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold37 (.A(\matt_venn_clock.pulse_min.count[4] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0150_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold39 (.A(\vga_sync.vsync ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold40 (.A(\matt_venn_clock.pulse_hrs.count[4] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0140_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold42 (.A(\matt_venn_vga_shadow.y_block_q[5] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold43 (.A(_1170_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold44 (.A(_1175_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0230_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold46 (.A(\matt_venn_clock.sec_counter[23] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold47 (.A(_1113_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0211_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold49 (.A(\matt_venn_clock.sec_counter[3] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold50 (.A(_1101_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold51 (.A(\clock_sec_u[3] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold52 (.A(_1090_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold53 (.A(\matt_venn_clock.sec_counter[4] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold54 (.A(\matt_venn_clock.pulse_sec.count[3] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold55 (.A(\matt_venn_clock.pulse_hrs.count[3] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0139_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold57 (.A(\matt_venn_clock.sec_counter[24] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold58 (.A(_1115_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold59 (.A(\clock_sec_u[2] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0182_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold61 (.A(\matt_venn_clock.sec_counter[7] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold62 (.A(_1105_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold63 (.A(\pym[11] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold64 (.A(\matt_venn_clock.sec_counter[17] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold65 (.A(_1108_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold66 (.A(\clock_color_offset[2] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0163_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold68 (.A(\matt_venn_clock.sec_counter[6] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold69 (.A(\clock_min_u[3] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0176_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold71 (.A(\px[9] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0047_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0995_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold74 (.A(\matt_venn_clock.sec_counter[1] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold75 (.A(_1099_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold76 (.A(\pym[10] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold77 (.A(\matt_venn_clock.pulse_sec.comp[4] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0950_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0155_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0046_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold81 (.A(\product_comp[10] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold82 (.A(\matt_venn_clock.sec_counter[15] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold83 (.A(_1107_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold84 (.A(\clock_sec_d[0] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold85 (.A(_1035_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0177_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0043_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0078_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold89 (.A(\matt_venn_clock.pulse_hrs.count[2] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0138_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold91 (.A(\matt_venn_clock.pulse_min.comp[1] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0049_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold93 (.A(\ydelta[5] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold94 (.A(\clock_min_d[2] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold95 (.A(_1016_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0172_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold97 (.A(\clock_color_offset[1] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0978_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0026_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0110_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold101 (.A(\clock_sec_d[2] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold102 (.A(_1039_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold103 (.A(\clock_hrs_d[1] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0990_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold105 (.A(\product_comp[9] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0048_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold107 (.A(_1106_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold108 (.A(\matt_venn_clock.pulse_min.comp[4] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0145_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold110 (.A(\matt_venn_clock.sec_counter[13] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold111 (.A(\px[3] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold112 (.A(\matt_venn_clock.pulse_hrs.comp[4] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0866_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold114 (.A(\vga_sync.hsync ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0790_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold116 (.A(\matt_venn_clock.pulse_min.count[2] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0148_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold118 (.A(\ydelta[6] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold119 (.A(\matt_venn_clock.pulse_min.count[3] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0149_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold121 (.A(\product_comp[2] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0221_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold123 (.A(\matt_venn_clock.pulse_sec.count[2] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0158_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold125 (.A(\matt_venn_clock.sec_counter[14] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold126 (.A(_1060_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold127 (.A(\ydelta[3] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold128 (.A(\matt_venn_clock.sec_counter[11] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold129 (.A(_1063_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold130 (.A(\matt_venn_clock.pulse_hrs.count[1] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0137_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0032_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold133 (.A(_1080_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold134 (.A(\matt_venn_clock.pulse_min.comp[0] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold135 (.A(\matt_venn_clock.pulse_sec.comp[2] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0153_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold137 (.A(\matt_venn_clock.pulse_hrs.count[0] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold138 (.A(\clock_hrs_u[1] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold139 (.A(\matt_venn_clock.pulse_sec.count[1] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0157_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold141 (.A(\matt_venn_clock.pulse_min.count[1] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0147_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold143 (.A(\clock_hrs_u[3] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold144 (.A(_1008_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold145 (.A(\matt_venn_clock.pulse_sec.comp[1] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold146 (.A(\matt_venn_clock.pulse_min.comp[3] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0053_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold148 (.A(\matt_venn_clock.sec_counter[16] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold149 (.A(\product_comp[3] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold150 (.A(\matt_venn_clock.pulse_hrs.comp[1] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold151 (.A(\matt_venn_clock.sec_counter[8] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold152 (.A(\clock_hrs_u[2] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0168_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold154 (.A(\clock_sec_u[1] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold155 (.A(_1084_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold156 (.A(\matt_venn_clock.pulse_min.comp[2] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold157 (.A(\py[7] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold158 (.A(\matt_venn_clock.pulse_hrs.comp[2] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0133_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold160 (.A(\matt_venn_clock.sec_counter[20] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold161 (.A(_1111_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold162 (.A(\ydelta[4] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold163 (.A(\py[8] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold164 (.A(\matt_venn_clock.pulse_sec.comp[3] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0949_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold166 (.A(\ydelta[2] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold167 (.A(\ydelta[1] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold168 (.A(\px[2] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold169 (.A(\matt_venn_clock.pulse_hrs.comp[0] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold170 (.A(\matt_venn_clock.sec_counter[10] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold171 (.A(_1064_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold172 (.A(\h[4] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold173 (.A(\matt_venn_clock.sec_counter[9] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0024_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold175 (.A(\matt_venn_vga.digit_0.char[0] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0840_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold177 (.A(\py[9] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold178 (.A(\px[1] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold179 (.A(\product_comp[4] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold180 (.A(\matt_venn_clock.sec_counter[19] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold181 (.A(\matt_venn_clock.pulse_sec.count[0] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0156_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold183 (.A(\matt_venn_vga.y_px[9] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0116_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold185 (.A(\matt_venn_clock.sec_counter[22] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold186 (.A(\py[2] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold187 (.A(\matt_venn_clock.pulse_min.count[0] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold188 (.A(\clock_min_d[0] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold189 (.A(_1014_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0171_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold191 (.A(\clock_min_u[1] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold192 (.A(_1025_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold193 (.A(\product_comp[8] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold194 (.A(\py[5] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold195 (.A(\matt_venn_vga.y_px[5] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0112_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold197 (.A(\px[4] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold198 (.A(\py[6] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold199 (.A(\h[1] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0122_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold201 (.A(\px[8] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold202 (.A(\h[3] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold203 (.A(\matt_venn_vga.y_px[2] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0799_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold205 (.A(\h[5] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold206 (.A(\matt_venn_vga.y_px[6] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold207 (.A(\clock_sec_d[1] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold208 (.A(\py[3] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold209 (.A(\product_comp[6] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold210 (.A(\product_comp[7] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold211 (.A(\px[5] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold212 (.A(\matt_venn_vga.y_px[0] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold213 (.A(\h[2] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold214 (.A(\product_comp[5] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold215 (.A(\h[8] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold216 (.A(\py[0] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0091_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold218 (.A(\matt_venn_clock.pulse_hrs.comp[3] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold219 (.A(\matt_venn_vga.y_px[3] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold220 (.A(_1281_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0041_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold222 (.A(\matt_venn_vga.y_px[8] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold223 (.A(\py[4] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold224 (.A(\matt_venn_clock.pulse_sec.comp[0] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold225 (.A(\matt_venn_vga.y_px[1] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold226 (.A(\matt_venn_vga.y_px[4] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0031_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold228 (.A(\px[7] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0033_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0050_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0033_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold232 (.A(\px[6] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold233 (.A(\matt_venn_clock.sec_counter[20] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold234 (.A(\matt_venn_clock.sec_counter[14] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold235 (.A(\matt_venn_clock.pulse_sec.count[2] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0967_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold237 (.A(\matt_venn_clock.sec_counter[16] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold238 (.A(\clock_color_offset[1] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold239 (.A(\matt_venn_clock.pulse_min.comp[3] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold240 (.A(\pym[10] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0041_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold242 (.A(\product_comp[7] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold243 (.A(\clock_color_offset[1] ),
    .X(net549));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_fill_1 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_202 ();
 sg13g2_decap_8 FILLER_5_209 ();
 sg13g2_decap_8 FILLER_5_216 ();
 sg13g2_decap_8 FILLER_5_223 ();
 sg13g2_decap_8 FILLER_5_230 ();
 sg13g2_decap_8 FILLER_5_237 ();
 sg13g2_decap_8 FILLER_5_244 ();
 sg13g2_decap_8 FILLER_5_251 ();
 sg13g2_decap_8 FILLER_5_258 ();
 sg13g2_decap_8 FILLER_5_265 ();
 sg13g2_decap_8 FILLER_5_272 ();
 sg13g2_decap_8 FILLER_5_279 ();
 sg13g2_decap_8 FILLER_5_286 ();
 sg13g2_decap_8 FILLER_5_293 ();
 sg13g2_decap_8 FILLER_5_300 ();
 sg13g2_decap_8 FILLER_5_307 ();
 sg13g2_decap_8 FILLER_5_314 ();
 sg13g2_decap_8 FILLER_5_321 ();
 sg13g2_decap_8 FILLER_5_328 ();
 sg13g2_decap_8 FILLER_5_335 ();
 sg13g2_decap_8 FILLER_5_342 ();
 sg13g2_decap_8 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_356 ();
 sg13g2_decap_8 FILLER_5_363 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_fill_2 FILLER_6_168 ();
 sg13g2_fill_1 FILLER_6_170 ();
 sg13g2_decap_8 FILLER_6_213 ();
 sg13g2_decap_8 FILLER_6_220 ();
 sg13g2_decap_8 FILLER_6_227 ();
 sg13g2_decap_8 FILLER_6_234 ();
 sg13g2_decap_8 FILLER_6_241 ();
 sg13g2_decap_8 FILLER_6_248 ();
 sg13g2_decap_8 FILLER_6_255 ();
 sg13g2_decap_8 FILLER_6_262 ();
 sg13g2_decap_8 FILLER_6_269 ();
 sg13g2_decap_8 FILLER_6_276 ();
 sg13g2_decap_8 FILLER_6_283 ();
 sg13g2_decap_8 FILLER_6_290 ();
 sg13g2_decap_8 FILLER_6_297 ();
 sg13g2_decap_8 FILLER_6_304 ();
 sg13g2_decap_8 FILLER_6_311 ();
 sg13g2_decap_8 FILLER_6_318 ();
 sg13g2_decap_8 FILLER_6_325 ();
 sg13g2_decap_8 FILLER_6_332 ();
 sg13g2_decap_8 FILLER_6_339 ();
 sg13g2_decap_8 FILLER_6_346 ();
 sg13g2_decap_8 FILLER_6_353 ();
 sg13g2_decap_8 FILLER_6_360 ();
 sg13g2_decap_8 FILLER_6_367 ();
 sg13g2_decap_8 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_381 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_decap_8 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_4 FILLER_7_168 ();
 sg13g2_fill_1 FILLER_7_202 ();
 sg13g2_decap_8 FILLER_7_233 ();
 sg13g2_decap_8 FILLER_7_240 ();
 sg13g2_decap_8 FILLER_7_247 ();
 sg13g2_decap_8 FILLER_7_254 ();
 sg13g2_decap_8 FILLER_7_261 ();
 sg13g2_decap_8 FILLER_7_268 ();
 sg13g2_decap_8 FILLER_7_275 ();
 sg13g2_decap_8 FILLER_7_282 ();
 sg13g2_decap_8 FILLER_7_289 ();
 sg13g2_decap_8 FILLER_7_296 ();
 sg13g2_decap_8 FILLER_7_303 ();
 sg13g2_decap_8 FILLER_7_310 ();
 sg13g2_decap_8 FILLER_7_317 ();
 sg13g2_decap_8 FILLER_7_324 ();
 sg13g2_decap_8 FILLER_7_331 ();
 sg13g2_decap_8 FILLER_7_338 ();
 sg13g2_decap_8 FILLER_7_345 ();
 sg13g2_decap_8 FILLER_7_352 ();
 sg13g2_decap_8 FILLER_7_359 ();
 sg13g2_decap_8 FILLER_7_366 ();
 sg13g2_decap_8 FILLER_7_373 ();
 sg13g2_decap_8 FILLER_7_380 ();
 sg13g2_decap_8 FILLER_7_387 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_4 FILLER_9_182 ();
 sg13g2_fill_2 FILLER_9_204 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_fill_2 FILLER_9_287 ();
 sg13g2_fill_1 FILLER_9_289 ();
 sg13g2_fill_2 FILLER_9_302 ();
 sg13g2_fill_1 FILLER_9_304 ();
 sg13g2_decap_8 FILLER_9_318 ();
 sg13g2_decap_8 FILLER_9_325 ();
 sg13g2_decap_8 FILLER_9_332 ();
 sg13g2_decap_8 FILLER_9_339 ();
 sg13g2_decap_8 FILLER_9_346 ();
 sg13g2_decap_8 FILLER_9_353 ();
 sg13g2_decap_8 FILLER_9_360 ();
 sg13g2_decap_8 FILLER_9_367 ();
 sg13g2_decap_8 FILLER_9_374 ();
 sg13g2_decap_8 FILLER_9_381 ();
 sg13g2_decap_8 FILLER_9_388 ();
 sg13g2_decap_8 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_4 FILLER_10_168 ();
 sg13g2_fill_2 FILLER_10_172 ();
 sg13g2_decap_8 FILLER_10_192 ();
 sg13g2_fill_1 FILLER_10_199 ();
 sg13g2_decap_4 FILLER_10_204 ();
 sg13g2_fill_2 FILLER_10_208 ();
 sg13g2_fill_2 FILLER_10_231 ();
 sg13g2_fill_1 FILLER_10_233 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_decap_8 FILLER_10_271 ();
 sg13g2_fill_2 FILLER_10_278 ();
 sg13g2_fill_1 FILLER_10_280 ();
 sg13g2_fill_2 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_328 ();
 sg13g2_decap_8 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_4 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_226 ();
 sg13g2_fill_1 FILLER_11_237 ();
 sg13g2_fill_2 FILLER_11_246 ();
 sg13g2_fill_1 FILLER_11_248 ();
 sg13g2_decap_4 FILLER_11_275 ();
 sg13g2_decap_4 FILLER_11_289 ();
 sg13g2_fill_1 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_fill_2 FILLER_12_154 ();
 sg13g2_fill_1 FILLER_12_156 ();
 sg13g2_fill_1 FILLER_12_174 ();
 sg13g2_fill_2 FILLER_12_189 ();
 sg13g2_fill_1 FILLER_12_191 ();
 sg13g2_fill_2 FILLER_12_212 ();
 sg13g2_fill_1 FILLER_12_241 ();
 sg13g2_fill_2 FILLER_12_250 ();
 sg13g2_fill_1 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_257 ();
 sg13g2_fill_2 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_295 ();
 sg13g2_decap_4 FILLER_12_302 ();
 sg13g2_fill_2 FILLER_12_311 ();
 sg13g2_decap_4 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_4 FILLER_13_161 ();
 sg13g2_fill_1 FILLER_13_178 ();
 sg13g2_fill_1 FILLER_13_184 ();
 sg13g2_decap_8 FILLER_13_192 ();
 sg13g2_fill_1 FILLER_13_199 ();
 sg13g2_fill_1 FILLER_13_216 ();
 sg13g2_fill_1 FILLER_13_232 ();
 sg13g2_decap_8 FILLER_13_257 ();
 sg13g2_decap_4 FILLER_13_264 ();
 sg13g2_fill_2 FILLER_13_282 ();
 sg13g2_fill_2 FILLER_13_302 ();
 sg13g2_fill_2 FILLER_13_317 ();
 sg13g2_fill_1 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_4 FILLER_14_154 ();
 sg13g2_fill_1 FILLER_14_158 ();
 sg13g2_fill_1 FILLER_14_246 ();
 sg13g2_fill_2 FILLER_14_300 ();
 sg13g2_fill_1 FILLER_14_302 ();
 sg13g2_fill_2 FILLER_14_319 ();
 sg13g2_fill_1 FILLER_14_321 ();
 sg13g2_decap_8 FILLER_14_339 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_decap_8 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_decap_8 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_4 FILLER_15_126 ();
 sg13g2_fill_1 FILLER_15_130 ();
 sg13g2_decap_8 FILLER_15_157 ();
 sg13g2_decap_4 FILLER_15_164 ();
 sg13g2_fill_1 FILLER_15_168 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_fill_1 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_222 ();
 sg13g2_fill_1 FILLER_15_277 ();
 sg13g2_fill_2 FILLER_15_300 ();
 sg13g2_fill_2 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_decap_8 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_decap_8 FILLER_15_369 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_4 FILLER_16_126 ();
 sg13g2_fill_1 FILLER_16_130 ();
 sg13g2_decap_4 FILLER_16_168 ();
 sg13g2_fill_1 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_decap_4 FILLER_16_230 ();
 sg13g2_decap_8 FILLER_16_255 ();
 sg13g2_fill_2 FILLER_16_262 ();
 sg13g2_fill_1 FILLER_16_264 ();
 sg13g2_decap_8 FILLER_16_290 ();
 sg13g2_decap_8 FILLER_16_297 ();
 sg13g2_decap_8 FILLER_16_304 ();
 sg13g2_decap_8 FILLER_16_311 ();
 sg13g2_decap_8 FILLER_16_318 ();
 sg13g2_decap_8 FILLER_16_325 ();
 sg13g2_decap_8 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_4 FILLER_17_126 ();
 sg13g2_fill_1 FILLER_17_130 ();
 sg13g2_fill_1 FILLER_17_153 ();
 sg13g2_fill_1 FILLER_17_182 ();
 sg13g2_decap_4 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_200 ();
 sg13g2_decap_8 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_214 ();
 sg13g2_fill_1 FILLER_17_216 ();
 sg13g2_decap_8 FILLER_17_221 ();
 sg13g2_fill_2 FILLER_17_228 ();
 sg13g2_decap_8 FILLER_17_239 ();
 sg13g2_decap_4 FILLER_17_246 ();
 sg13g2_fill_1 FILLER_17_250 ();
 sg13g2_decap_8 FILLER_17_256 ();
 sg13g2_fill_2 FILLER_17_288 ();
 sg13g2_decap_4 FILLER_17_299 ();
 sg13g2_fill_1 FILLER_17_303 ();
 sg13g2_fill_2 FILLER_17_327 ();
 sg13g2_decap_8 FILLER_17_338 ();
 sg13g2_decap_8 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_fill_2 FILLER_18_140 ();
 sg13g2_fill_1 FILLER_18_142 ();
 sg13g2_decap_4 FILLER_18_159 ();
 sg13g2_fill_2 FILLER_18_171 ();
 sg13g2_fill_1 FILLER_18_173 ();
 sg13g2_decap_4 FILLER_18_183 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_2 FILLER_18_214 ();
 sg13g2_fill_1 FILLER_18_216 ();
 sg13g2_fill_2 FILLER_18_222 ();
 sg13g2_decap_8 FILLER_18_236 ();
 sg13g2_decap_4 FILLER_18_243 ();
 sg13g2_fill_1 FILLER_18_247 ();
 sg13g2_fill_1 FILLER_18_278 ();
 sg13g2_fill_2 FILLER_18_286 ();
 sg13g2_fill_2 FILLER_18_304 ();
 sg13g2_decap_4 FILLER_18_311 ();
 sg13g2_decap_8 FILLER_18_344 ();
 sg13g2_decap_8 FILLER_18_351 ();
 sg13g2_decap_8 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_365 ();
 sg13g2_decap_8 FILLER_18_372 ();
 sg13g2_decap_8 FILLER_18_379 ();
 sg13g2_decap_8 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_fill_2 FILLER_19_133 ();
 sg13g2_fill_1 FILLER_19_135 ();
 sg13g2_decap_8 FILLER_19_141 ();
 sg13g2_decap_4 FILLER_19_148 ();
 sg13g2_fill_1 FILLER_19_152 ();
 sg13g2_fill_2 FILLER_19_182 ();
 sg13g2_fill_1 FILLER_19_184 ();
 sg13g2_fill_2 FILLER_19_270 ();
 sg13g2_fill_1 FILLER_19_285 ();
 sg13g2_fill_1 FILLER_19_294 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_341 ();
 sg13g2_decap_8 FILLER_19_348 ();
 sg13g2_decap_8 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_362 ();
 sg13g2_decap_8 FILLER_19_369 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_fill_2 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_decap_4 FILLER_20_234 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_260 ();
 sg13g2_fill_2 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_271 ();
 sg13g2_decap_4 FILLER_20_294 ();
 sg13g2_decap_4 FILLER_20_312 ();
 sg13g2_fill_2 FILLER_20_316 ();
 sg13g2_fill_2 FILLER_20_323 ();
 sg13g2_decap_8 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_342 ();
 sg13g2_decap_8 FILLER_20_349 ();
 sg13g2_decap_8 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_4 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_123 ();
 sg13g2_fill_2 FILLER_21_128 ();
 sg13g2_fill_2 FILLER_21_159 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_decap_8 FILLER_21_229 ();
 sg13g2_decap_8 FILLER_21_236 ();
 sg13g2_fill_2 FILLER_21_247 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_fill_2 FILLER_21_283 ();
 sg13g2_fill_1 FILLER_21_285 ();
 sg13g2_decap_8 FILLER_21_309 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_fill_2 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_135 ();
 sg13g2_fill_1 FILLER_22_155 ();
 sg13g2_decap_8 FILLER_22_160 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_fill_2 FILLER_22_176 ();
 sg13g2_fill_1 FILLER_22_178 ();
 sg13g2_decap_8 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_216 ();
 sg13g2_fill_2 FILLER_22_223 ();
 sg13g2_fill_1 FILLER_22_236 ();
 sg13g2_fill_2 FILLER_22_249 ();
 sg13g2_fill_1 FILLER_22_251 ();
 sg13g2_fill_2 FILLER_22_261 ();
 sg13g2_fill_1 FILLER_22_263 ();
 sg13g2_fill_1 FILLER_22_290 ();
 sg13g2_decap_4 FILLER_22_324 ();
 sg13g2_fill_1 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_decap_8 FILLER_22_341 ();
 sg13g2_decap_8 FILLER_22_348 ();
 sg13g2_decap_8 FILLER_22_355 ();
 sg13g2_decap_8 FILLER_22_362 ();
 sg13g2_decap_8 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_fill_1 FILLER_23_133 ();
 sg13g2_fill_1 FILLER_23_139 ();
 sg13g2_fill_2 FILLER_23_162 ();
 sg13g2_fill_1 FILLER_23_180 ();
 sg13g2_fill_2 FILLER_23_194 ();
 sg13g2_fill_2 FILLER_23_210 ();
 sg13g2_decap_4 FILLER_23_294 ();
 sg13g2_fill_2 FILLER_23_298 ();
 sg13g2_fill_2 FILLER_23_304 ();
 sg13g2_decap_8 FILLER_23_344 ();
 sg13g2_decap_8 FILLER_23_351 ();
 sg13g2_decap_8 FILLER_23_358 ();
 sg13g2_decap_8 FILLER_23_365 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_4 FILLER_24_105 ();
 sg13g2_decap_4 FILLER_24_135 ();
 sg13g2_fill_2 FILLER_24_151 ();
 sg13g2_fill_2 FILLER_24_160 ();
 sg13g2_fill_1 FILLER_24_167 ();
 sg13g2_decap_4 FILLER_24_178 ();
 sg13g2_fill_1 FILLER_24_201 ();
 sg13g2_fill_2 FILLER_24_234 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_fill_2 FILLER_24_273 ();
 sg13g2_fill_2 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_295 ();
 sg13g2_decap_4 FILLER_24_307 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_178 ();
 sg13g2_fill_2 FILLER_25_189 ();
 sg13g2_fill_1 FILLER_25_228 ();
 sg13g2_decap_8 FILLER_25_237 ();
 sg13g2_fill_2 FILLER_25_285 ();
 sg13g2_decap_8 FILLER_25_304 ();
 sg13g2_fill_2 FILLER_25_311 ();
 sg13g2_fill_1 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_324 ();
 sg13g2_fill_2 FILLER_25_330 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_decap_8 FILLER_25_341 ();
 sg13g2_decap_8 FILLER_25_348 ();
 sg13g2_decap_8 FILLER_25_355 ();
 sg13g2_decap_8 FILLER_25_362 ();
 sg13g2_decap_8 FILLER_25_369 ();
 sg13g2_decap_8 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_119 ();
 sg13g2_decap_4 FILLER_26_128 ();
 sg13g2_fill_1 FILLER_26_132 ();
 sg13g2_fill_2 FILLER_26_138 ();
 sg13g2_fill_1 FILLER_26_140 ();
 sg13g2_fill_2 FILLER_26_150 ();
 sg13g2_fill_1 FILLER_26_162 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_223 ();
 sg13g2_decap_8 FILLER_26_229 ();
 sg13g2_decap_8 FILLER_26_236 ();
 sg13g2_decap_8 FILLER_26_243 ();
 sg13g2_decap_4 FILLER_26_250 ();
 sg13g2_decap_4 FILLER_26_265 ();
 sg13g2_fill_1 FILLER_26_269 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_298 ();
 sg13g2_decap_8 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_decap_8 FILLER_26_319 ();
 sg13g2_decap_4 FILLER_26_326 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_decap_8 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_4 FILLER_27_126 ();
 sg13g2_decap_4 FILLER_27_135 ();
 sg13g2_fill_2 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_155 ();
 sg13g2_fill_1 FILLER_27_162 ();
 sg13g2_fill_2 FILLER_27_195 ();
 sg13g2_decap_8 FILLER_27_201 ();
 sg13g2_decap_4 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_217 ();
 sg13g2_fill_1 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_decap_4 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_fill_2 FILLER_27_316 ();
 sg13g2_fill_2 FILLER_27_328 ();
 sg13g2_decap_8 FILLER_27_338 ();
 sg13g2_decap_8 FILLER_27_345 ();
 sg13g2_decap_8 FILLER_27_352 ();
 sg13g2_decap_8 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_fill_2 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_104 ();
 sg13g2_decap_4 FILLER_28_109 ();
 sg13g2_fill_2 FILLER_28_113 ();
 sg13g2_fill_2 FILLER_28_141 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_fill_2 FILLER_28_149 ();
 sg13g2_fill_2 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_177 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_fill_2 FILLER_28_225 ();
 sg13g2_fill_1 FILLER_28_227 ();
 sg13g2_fill_2 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_287 ();
 sg13g2_fill_2 FILLER_28_330 ();
 sg13g2_decap_8 FILLER_28_345 ();
 sg13g2_decap_8 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_28_359 ();
 sg13g2_decap_8 FILLER_28_366 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_4 FILLER_29_77 ();
 sg13g2_fill_1 FILLER_29_81 ();
 sg13g2_fill_1 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_162 ();
 sg13g2_decap_8 FILLER_29_177 ();
 sg13g2_decap_8 FILLER_29_184 ();
 sg13g2_decap_4 FILLER_29_191 ();
 sg13g2_fill_1 FILLER_29_218 ();
 sg13g2_fill_2 FILLER_29_245 ();
 sg13g2_fill_2 FILLER_29_286 ();
 sg13g2_fill_1 FILLER_29_294 ();
 sg13g2_fill_2 FILLER_29_330 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_decap_8 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_decap_8 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_29_370 ();
 sg13g2_decap_8 FILLER_29_377 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_fill_1 FILLER_30_106 ();
 sg13g2_fill_1 FILLER_30_163 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_fill_2 FILLER_30_197 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_269 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_fill_2 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_353 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_367 ();
 sg13g2_decap_8 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_65 ();
 sg13g2_fill_2 FILLER_31_92 ();
 sg13g2_fill_2 FILLER_31_128 ();
 sg13g2_fill_2 FILLER_31_135 ();
 sg13g2_fill_1 FILLER_31_137 ();
 sg13g2_decap_8 FILLER_31_142 ();
 sg13g2_fill_2 FILLER_31_208 ();
 sg13g2_decap_4 FILLER_31_225 ();
 sg13g2_decap_4 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_decap_4 FILLER_31_260 ();
 sg13g2_fill_2 FILLER_31_272 ();
 sg13g2_fill_1 FILLER_31_274 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_fill_1 FILLER_31_307 ();
 sg13g2_decap_8 FILLER_31_313 ();
 sg13g2_fill_1 FILLER_31_320 ();
 sg13g2_fill_2 FILLER_31_325 ();
 sg13g2_fill_1 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_353 ();
 sg13g2_decap_8 FILLER_31_360 ();
 sg13g2_decap_8 FILLER_31_367 ();
 sg13g2_decap_8 FILLER_31_374 ();
 sg13g2_decap_8 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_fill_2 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_144 ();
 sg13g2_fill_1 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_166 ();
 sg13g2_decap_8 FILLER_32_173 ();
 sg13g2_fill_1 FILLER_32_180 ();
 sg13g2_fill_2 FILLER_32_191 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_decap_8 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_226 ();
 sg13g2_decap_4 FILLER_32_233 ();
 sg13g2_fill_1 FILLER_32_237 ();
 sg13g2_decap_4 FILLER_32_272 ();
 sg13g2_fill_2 FILLER_32_276 ();
 sg13g2_fill_2 FILLER_32_314 ();
 sg13g2_fill_2 FILLER_32_324 ();
 sg13g2_decap_8 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_fill_2 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_fill_2 FILLER_33_147 ();
 sg13g2_fill_1 FILLER_33_149 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_fill_1 FILLER_33_182 ();
 sg13g2_fill_1 FILLER_33_213 ();
 sg13g2_fill_1 FILLER_33_226 ();
 sg13g2_fill_2 FILLER_33_287 ();
 sg13g2_fill_1 FILLER_33_289 ();
 sg13g2_fill_2 FILLER_33_310 ();
 sg13g2_fill_1 FILLER_33_312 ();
 sg13g2_decap_4 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_346 ();
 sg13g2_decap_8 FILLER_33_353 ();
 sg13g2_decap_8 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_33_367 ();
 sg13g2_decap_8 FILLER_33_374 ();
 sg13g2_decap_8 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_33_388 ();
 sg13g2_decap_8 FILLER_33_395 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_fill_2 FILLER_34_89 ();
 sg13g2_fill_2 FILLER_34_115 ();
 sg13g2_fill_1 FILLER_34_117 ();
 sg13g2_fill_1 FILLER_34_156 ();
 sg13g2_fill_1 FILLER_34_162 ();
 sg13g2_fill_2 FILLER_34_198 ();
 sg13g2_fill_1 FILLER_34_200 ();
 sg13g2_decap_4 FILLER_34_222 ();
 sg13g2_fill_1 FILLER_34_226 ();
 sg13g2_decap_4 FILLER_34_235 ();
 sg13g2_decap_8 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_fill_2 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_298 ();
 sg13g2_decap_8 FILLER_34_305 ();
 sg13g2_fill_1 FILLER_34_312 ();
 sg13g2_decap_4 FILLER_34_317 ();
 sg13g2_fill_1 FILLER_34_321 ();
 sg13g2_decap_8 FILLER_34_338 ();
 sg13g2_decap_8 FILLER_34_345 ();
 sg13g2_decap_8 FILLER_34_352 ();
 sg13g2_decap_8 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_34_366 ();
 sg13g2_decap_8 FILLER_34_373 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_4 FILLER_35_42 ();
 sg13g2_fill_1 FILLER_35_121 ();
 sg13g2_fill_1 FILLER_35_146 ();
 sg13g2_fill_2 FILLER_35_178 ();
 sg13g2_fill_1 FILLER_35_180 ();
 sg13g2_decap_4 FILLER_35_190 ();
 sg13g2_fill_1 FILLER_35_206 ();
 sg13g2_fill_2 FILLER_35_215 ();
 sg13g2_decap_8 FILLER_35_222 ();
 sg13g2_decap_4 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_233 ();
 sg13g2_decap_8 FILLER_35_249 ();
 sg13g2_decap_4 FILLER_35_266 ();
 sg13g2_fill_1 FILLER_35_270 ();
 sg13g2_fill_2 FILLER_35_276 ();
 sg13g2_fill_1 FILLER_35_278 ();
 sg13g2_fill_2 FILLER_35_295 ();
 sg13g2_decap_8 FILLER_35_325 ();
 sg13g2_decap_8 FILLER_35_332 ();
 sg13g2_decap_8 FILLER_35_339 ();
 sg13g2_decap_8 FILLER_35_346 ();
 sg13g2_decap_8 FILLER_35_353 ();
 sg13g2_decap_8 FILLER_35_360 ();
 sg13g2_decap_8 FILLER_35_367 ();
 sg13g2_decap_8 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_49 ();
 sg13g2_fill_1 FILLER_36_55 ();
 sg13g2_decap_8 FILLER_36_122 ();
 sg13g2_decap_4 FILLER_36_129 ();
 sg13g2_fill_2 FILLER_36_146 ();
 sg13g2_fill_2 FILLER_36_153 ();
 sg13g2_decap_4 FILLER_36_159 ();
 sg13g2_fill_2 FILLER_36_163 ();
 sg13g2_decap_8 FILLER_36_219 ();
 sg13g2_decap_4 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_230 ();
 sg13g2_decap_4 FILLER_36_236 ();
 sg13g2_fill_1 FILLER_36_240 ();
 sg13g2_decap_8 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_fill_2 FILLER_36_271 ();
 sg13g2_decap_4 FILLER_36_291 ();
 sg13g2_fill_2 FILLER_36_316 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_fill_2 FILLER_36_334 ();
 sg13g2_decap_8 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_fill_2 FILLER_37_63 ();
 sg13g2_fill_1 FILLER_37_69 ();
 sg13g2_fill_2 FILLER_37_86 ();
 sg13g2_fill_1 FILLER_37_92 ();
 sg13g2_fill_1 FILLER_37_111 ();
 sg13g2_fill_1 FILLER_37_122 ();
 sg13g2_decap_4 FILLER_37_131 ();
 sg13g2_fill_2 FILLER_37_135 ();
 sg13g2_decap_8 FILLER_37_145 ();
 sg13g2_decap_8 FILLER_37_152 ();
 sg13g2_decap_8 FILLER_37_159 ();
 sg13g2_decap_8 FILLER_37_166 ();
 sg13g2_fill_2 FILLER_37_173 ();
 sg13g2_fill_1 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_180 ();
 sg13g2_decap_8 FILLER_37_187 ();
 sg13g2_decap_4 FILLER_37_194 ();
 sg13g2_fill_1 FILLER_37_198 ();
 sg13g2_fill_1 FILLER_37_207 ();
 sg13g2_fill_2 FILLER_37_216 ();
 sg13g2_fill_2 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_241 ();
 sg13g2_fill_2 FILLER_37_250 ();
 sg13g2_fill_1 FILLER_37_252 ();
 sg13g2_fill_2 FILLER_37_266 ();
 sg13g2_fill_1 FILLER_37_268 ();
 sg13g2_fill_1 FILLER_37_321 ();
 sg13g2_decap_8 FILLER_37_339 ();
 sg13g2_decap_8 FILLER_37_346 ();
 sg13g2_decap_8 FILLER_37_353 ();
 sg13g2_decap_8 FILLER_37_360 ();
 sg13g2_decap_8 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_374 ();
 sg13g2_decap_8 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_4 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_32 ();
 sg13g2_fill_2 FILLER_38_107 ();
 sg13g2_fill_1 FILLER_38_113 ();
 sg13g2_fill_1 FILLER_38_145 ();
 sg13g2_decap_8 FILLER_38_177 ();
 sg13g2_decap_8 FILLER_38_184 ();
 sg13g2_decap_8 FILLER_38_191 ();
 sg13g2_decap_8 FILLER_38_198 ();
 sg13g2_fill_2 FILLER_38_205 ();
 sg13g2_fill_2 FILLER_38_239 ();
 sg13g2_fill_1 FILLER_38_241 ();
 sg13g2_fill_2 FILLER_38_250 ();
 sg13g2_fill_1 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_289 ();
 sg13g2_fill_2 FILLER_38_296 ();
 sg13g2_fill_2 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_373 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_4 FILLER_39_28 ();
 sg13g2_fill_2 FILLER_39_32 ();
 sg13g2_fill_2 FILLER_39_65 ();
 sg13g2_fill_1 FILLER_39_67 ();
 sg13g2_fill_1 FILLER_39_90 ();
 sg13g2_fill_2 FILLER_39_111 ();
 sg13g2_fill_1 FILLER_39_139 ();
 sg13g2_fill_1 FILLER_39_159 ();
 sg13g2_decap_8 FILLER_39_188 ();
 sg13g2_fill_1 FILLER_39_195 ();
 sg13g2_decap_8 FILLER_39_200 ();
 sg13g2_fill_2 FILLER_39_211 ();
 sg13g2_fill_1 FILLER_39_213 ();
 sg13g2_fill_2 FILLER_39_220 ();
 sg13g2_decap_4 FILLER_39_242 ();
 sg13g2_fill_2 FILLER_39_246 ();
 sg13g2_decap_8 FILLER_39_279 ();
 sg13g2_decap_8 FILLER_39_286 ();
 sg13g2_decap_8 FILLER_39_293 ();
 sg13g2_fill_2 FILLER_39_300 ();
 sg13g2_fill_1 FILLER_39_302 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_fill_2 FILLER_39_322 ();
 sg13g2_fill_1 FILLER_39_324 ();
 sg13g2_decap_4 FILLER_39_342 ();
 sg13g2_fill_1 FILLER_39_346 ();
 sg13g2_decap_8 FILLER_39_373 ();
 sg13g2_decap_8 FILLER_39_380 ();
 sg13g2_decap_8 FILLER_39_387 ();
 sg13g2_decap_8 FILLER_39_394 ();
 sg13g2_decap_8 FILLER_39_401 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_fill_1 FILLER_40_28 ();
 sg13g2_fill_1 FILLER_40_78 ();
 sg13g2_fill_1 FILLER_40_84 ();
 sg13g2_fill_2 FILLER_40_94 ();
 sg13g2_fill_1 FILLER_40_96 ();
 sg13g2_fill_1 FILLER_40_144 ();
 sg13g2_fill_2 FILLER_40_158 ();
 sg13g2_fill_1 FILLER_40_160 ();
 sg13g2_decap_4 FILLER_40_241 ();
 sg13g2_fill_2 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_260 ();
 sg13g2_decap_8 FILLER_40_267 ();
 sg13g2_decap_8 FILLER_40_274 ();
 sg13g2_decap_4 FILLER_40_281 ();
 sg13g2_decap_8 FILLER_40_303 ();
 sg13g2_decap_8 FILLER_40_310 ();
 sg13g2_decap_8 FILLER_40_317 ();
 sg13g2_decap_4 FILLER_40_324 ();
 sg13g2_fill_2 FILLER_40_339 ();
 sg13g2_fill_1 FILLER_40_341 ();
 sg13g2_decap_8 FILLER_40_379 ();
 sg13g2_decap_8 FILLER_40_386 ();
 sg13g2_decap_8 FILLER_40_393 ();
 sg13g2_decap_8 FILLER_40_400 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_fill_2 FILLER_41_35 ();
 sg13g2_fill_1 FILLER_41_37 ();
 sg13g2_fill_1 FILLER_41_56 ();
 sg13g2_fill_1 FILLER_41_74 ();
 sg13g2_fill_2 FILLER_41_167 ();
 sg13g2_decap_4 FILLER_41_211 ();
 sg13g2_fill_2 FILLER_41_215 ();
 sg13g2_fill_2 FILLER_41_220 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_fill_2 FILLER_41_266 ();
 sg13g2_fill_2 FILLER_41_284 ();
 sg13g2_fill_2 FILLER_41_312 ();
 sg13g2_fill_1 FILLER_41_314 ();
 sg13g2_fill_1 FILLER_41_341 ();
 sg13g2_fill_1 FILLER_41_352 ();
 sg13g2_decap_8 FILLER_41_379 ();
 sg13g2_decap_8 FILLER_41_386 ();
 sg13g2_decap_8 FILLER_41_393 ();
 sg13g2_decap_8 FILLER_41_400 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_4 FILLER_42_28 ();
 sg13g2_fill_1 FILLER_42_32 ();
 sg13g2_decap_4 FILLER_42_61 ();
 sg13g2_fill_1 FILLER_42_98 ();
 sg13g2_fill_1 FILLER_42_190 ();
 sg13g2_decap_8 FILLER_42_195 ();
 sg13g2_decap_4 FILLER_42_202 ();
 sg13g2_fill_1 FILLER_42_235 ();
 sg13g2_decap_4 FILLER_42_267 ();
 sg13g2_decap_4 FILLER_42_279 ();
 sg13g2_fill_1 FILLER_42_283 ();
 sg13g2_fill_1 FILLER_42_304 ();
 sg13g2_fill_2 FILLER_42_336 ();
 sg13g2_fill_1 FILLER_42_338 ();
 sg13g2_fill_2 FILLER_42_368 ();
 sg13g2_decap_8 FILLER_42_379 ();
 sg13g2_decap_8 FILLER_42_386 ();
 sg13g2_decap_8 FILLER_42_393 ();
 sg13g2_decap_8 FILLER_42_400 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_fill_2 FILLER_43_21 ();
 sg13g2_fill_1 FILLER_43_23 ();
 sg13g2_fill_1 FILLER_43_64 ();
 sg13g2_decap_8 FILLER_43_74 ();
 sg13g2_decap_4 FILLER_43_81 ();
 sg13g2_decap_4 FILLER_43_151 ();
 sg13g2_fill_1 FILLER_43_155 ();
 sg13g2_fill_1 FILLER_43_174 ();
 sg13g2_fill_2 FILLER_43_215 ();
 sg13g2_decap_8 FILLER_43_299 ();
 sg13g2_decap_4 FILLER_43_310 ();
 sg13g2_fill_2 FILLER_43_314 ();
 sg13g2_fill_1 FILLER_43_329 ();
 sg13g2_fill_2 FILLER_43_339 ();
 sg13g2_fill_1 FILLER_43_341 ();
 sg13g2_decap_4 FILLER_43_355 ();
 sg13g2_decap_8 FILLER_43_368 ();
 sg13g2_decap_8 FILLER_43_375 ();
 sg13g2_decap_8 FILLER_43_382 ();
 sg13g2_decap_8 FILLER_43_389 ();
 sg13g2_decap_8 FILLER_43_396 ();
 sg13g2_decap_4 FILLER_43_403 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_fill_1 FILLER_44_62 ();
 sg13g2_fill_2 FILLER_44_88 ();
 sg13g2_fill_1 FILLER_44_90 ();
 sg13g2_decap_8 FILLER_44_94 ();
 sg13g2_decap_8 FILLER_44_114 ();
 sg13g2_fill_1 FILLER_44_121 ();
 sg13g2_decap_8 FILLER_44_151 ();
 sg13g2_decap_8 FILLER_44_158 ();
 sg13g2_decap_4 FILLER_44_165 ();
 sg13g2_decap_4 FILLER_44_179 ();
 sg13g2_fill_1 FILLER_44_183 ();
 sg13g2_fill_2 FILLER_44_206 ();
 sg13g2_fill_1 FILLER_44_286 ();
 sg13g2_decap_8 FILLER_44_377 ();
 sg13g2_decap_8 FILLER_44_384 ();
 sg13g2_decap_8 FILLER_44_391 ();
 sg13g2_decap_8 FILLER_44_398 ();
 sg13g2_decap_4 FILLER_44_405 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_14 ();
 sg13g2_fill_1 FILLER_45_16 ();
 sg13g2_fill_2 FILLER_45_31 ();
 sg13g2_fill_2 FILLER_45_42 ();
 sg13g2_fill_1 FILLER_45_44 ();
 sg13g2_fill_2 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_108 ();
 sg13g2_decap_8 FILLER_45_115 ();
 sg13g2_decap_4 FILLER_45_122 ();
 sg13g2_fill_2 FILLER_45_126 ();
 sg13g2_fill_2 FILLER_45_184 ();
 sg13g2_fill_2 FILLER_45_207 ();
 sg13g2_fill_2 FILLER_45_246 ();
 sg13g2_fill_1 FILLER_45_248 ();
 sg13g2_fill_2 FILLER_45_275 ();
 sg13g2_fill_1 FILLER_45_308 ();
 sg13g2_fill_2 FILLER_45_332 ();
 sg13g2_fill_1 FILLER_45_351 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_fill_2 FILLER_45_406 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_4 FILLER_46_14 ();
 sg13g2_fill_1 FILLER_46_18 ();
 sg13g2_decap_4 FILLER_46_127 ();
 sg13g2_fill_1 FILLER_46_179 ();
 sg13g2_fill_1 FILLER_46_202 ();
 sg13g2_fill_1 FILLER_46_218 ();
 sg13g2_fill_2 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_274 ();
 sg13g2_decap_4 FILLER_46_281 ();
 sg13g2_fill_2 FILLER_46_285 ();
 sg13g2_fill_2 FILLER_46_291 ();
 sg13g2_fill_2 FILLER_46_311 ();
 sg13g2_fill_1 FILLER_46_325 ();
 sg13g2_fill_1 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_377 ();
 sg13g2_decap_8 FILLER_46_384 ();
 sg13g2_decap_8 FILLER_46_391 ();
 sg13g2_decap_8 FILLER_46_398 ();
 sg13g2_decap_4 FILLER_46_405 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_fill_2 FILLER_47_21 ();
 sg13g2_fill_1 FILLER_47_23 ();
 sg13g2_fill_1 FILLER_47_99 ();
 sg13g2_fill_2 FILLER_47_156 ();
 sg13g2_fill_1 FILLER_47_180 ();
 sg13g2_fill_1 FILLER_47_191 ();
 sg13g2_fill_2 FILLER_47_205 ();
 sg13g2_fill_1 FILLER_47_224 ();
 sg13g2_fill_2 FILLER_47_242 ();
 sg13g2_fill_1 FILLER_47_244 ();
 sg13g2_decap_8 FILLER_47_271 ();
 sg13g2_decap_4 FILLER_47_278 ();
 sg13g2_fill_1 FILLER_47_282 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_fill_1 FILLER_47_301 ();
 sg13g2_fill_2 FILLER_47_310 ();
 sg13g2_decap_8 FILLER_47_368 ();
 sg13g2_decap_8 FILLER_47_375 ();
 sg13g2_decap_8 FILLER_47_382 ();
 sg13g2_decap_8 FILLER_47_389 ();
 sg13g2_decap_8 FILLER_47_396 ();
 sg13g2_decap_4 FILLER_47_403 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_4 FILLER_48_21 ();
 sg13g2_fill_1 FILLER_48_25 ();
 sg13g2_fill_1 FILLER_48_83 ();
 sg13g2_fill_2 FILLER_48_97 ();
 sg13g2_fill_1 FILLER_48_104 ();
 sg13g2_fill_1 FILLER_48_120 ();
 sg13g2_decap_4 FILLER_48_141 ();
 sg13g2_decap_4 FILLER_48_161 ();
 sg13g2_fill_1 FILLER_48_165 ();
 sg13g2_fill_2 FILLER_48_170 ();
 sg13g2_decap_4 FILLER_48_177 ();
 sg13g2_decap_4 FILLER_48_211 ();
 sg13g2_fill_2 FILLER_48_215 ();
 sg13g2_decap_8 FILLER_48_227 ();
 sg13g2_fill_1 FILLER_48_234 ();
 sg13g2_fill_1 FILLER_48_249 ();
 sg13g2_decap_8 FILLER_48_302 ();
 sg13g2_fill_1 FILLER_48_309 ();
 sg13g2_fill_1 FILLER_48_319 ();
 sg13g2_fill_2 FILLER_48_329 ();
 sg13g2_fill_1 FILLER_48_331 ();
 sg13g2_decap_8 FILLER_48_356 ();
 sg13g2_decap_8 FILLER_48_363 ();
 sg13g2_decap_8 FILLER_48_370 ();
 sg13g2_decap_8 FILLER_48_377 ();
 sg13g2_decap_8 FILLER_48_384 ();
 sg13g2_decap_8 FILLER_48_391 ();
 sg13g2_decap_8 FILLER_48_398 ();
 sg13g2_decap_4 FILLER_48_405 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_fill_2 FILLER_49_35 ();
 sg13g2_fill_1 FILLER_49_37 ();
 sg13g2_fill_1 FILLER_49_55 ();
 sg13g2_fill_1 FILLER_49_66 ();
 sg13g2_fill_2 FILLER_49_75 ();
 sg13g2_fill_2 FILLER_49_89 ();
 sg13g2_decap_8 FILLER_49_104 ();
 sg13g2_fill_2 FILLER_49_111 ();
 sg13g2_fill_1 FILLER_49_113 ();
 sg13g2_decap_4 FILLER_49_151 ();
 sg13g2_fill_2 FILLER_49_155 ();
 sg13g2_decap_8 FILLER_49_176 ();
 sg13g2_decap_8 FILLER_49_183 ();
 sg13g2_fill_2 FILLER_49_190 ();
 sg13g2_fill_1 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_223 ();
 sg13g2_fill_1 FILLER_49_230 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_fill_1 FILLER_49_242 ();
 sg13g2_fill_2 FILLER_49_253 ();
 sg13g2_fill_1 FILLER_49_255 ();
 sg13g2_fill_1 FILLER_49_264 ();
 sg13g2_fill_2 FILLER_49_300 ();
 sg13g2_fill_2 FILLER_49_328 ();
 sg13g2_fill_1 FILLER_49_330 ();
 sg13g2_decap_8 FILLER_49_367 ();
 sg13g2_decap_8 FILLER_49_374 ();
 sg13g2_decap_8 FILLER_49_381 ();
 sg13g2_decap_8 FILLER_49_388 ();
 sg13g2_decap_8 FILLER_49_395 ();
 sg13g2_decap_8 FILLER_49_402 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_fill_2 FILLER_50_28 ();
 sg13g2_fill_1 FILLER_50_30 ();
 sg13g2_fill_1 FILLER_50_51 ();
 sg13g2_fill_1 FILLER_50_66 ();
 sg13g2_fill_2 FILLER_50_93 ();
 sg13g2_fill_1 FILLER_50_113 ();
 sg13g2_fill_2 FILLER_50_134 ();
 sg13g2_fill_1 FILLER_50_154 ();
 sg13g2_fill_2 FILLER_50_189 ();
 sg13g2_fill_1 FILLER_50_191 ();
 sg13g2_fill_2 FILLER_50_202 ();
 sg13g2_fill_1 FILLER_50_204 ();
 sg13g2_fill_2 FILLER_50_218 ();
 sg13g2_fill_1 FILLER_50_220 ();
 sg13g2_fill_2 FILLER_50_251 ();
 sg13g2_fill_1 FILLER_50_253 ();
 sg13g2_decap_4 FILLER_50_306 ();
 sg13g2_fill_2 FILLER_50_330 ();
 sg13g2_fill_1 FILLER_50_332 ();
 sg13g2_decap_8 FILLER_50_374 ();
 sg13g2_decap_8 FILLER_50_381 ();
 sg13g2_decap_8 FILLER_50_388 ();
 sg13g2_decap_8 FILLER_50_395 ();
 sg13g2_decap_8 FILLER_50_402 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_4 FILLER_51_21 ();
 sg13g2_fill_1 FILLER_51_30 ();
 sg13g2_fill_1 FILLER_51_58 ();
 sg13g2_decap_4 FILLER_51_67 ();
 sg13g2_fill_1 FILLER_51_71 ();
 sg13g2_fill_2 FILLER_51_80 ();
 sg13g2_fill_1 FILLER_51_108 ();
 sg13g2_decap_8 FILLER_51_120 ();
 sg13g2_decap_8 FILLER_51_127 ();
 sg13g2_decap_8 FILLER_51_134 ();
 sg13g2_decap_4 FILLER_51_141 ();
 sg13g2_fill_2 FILLER_51_180 ();
 sg13g2_decap_8 FILLER_51_190 ();
 sg13g2_decap_4 FILLER_51_197 ();
 sg13g2_fill_1 FILLER_51_201 ();
 sg13g2_fill_1 FILLER_51_212 ();
 sg13g2_fill_1 FILLER_51_221 ();
 sg13g2_fill_2 FILLER_51_244 ();
 sg13g2_fill_1 FILLER_51_246 ();
 sg13g2_decap_4 FILLER_51_315 ();
 sg13g2_fill_1 FILLER_51_324 ();
 sg13g2_decap_4 FILLER_51_330 ();
 sg13g2_fill_1 FILLER_51_334 ();
 sg13g2_decap_8 FILLER_51_365 ();
 sg13g2_decap_8 FILLER_51_372 ();
 sg13g2_decap_8 FILLER_51_379 ();
 sg13g2_decap_8 FILLER_51_386 ();
 sg13g2_decap_8 FILLER_51_393 ();
 sg13g2_decap_8 FILLER_51_400 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_4 FILLER_52_7 ();
 sg13g2_fill_1 FILLER_52_11 ();
 sg13g2_fill_2 FILLER_52_37 ();
 sg13g2_fill_2 FILLER_52_49 ();
 sg13g2_fill_1 FILLER_52_51 ();
 sg13g2_decap_8 FILLER_52_65 ();
 sg13g2_decap_4 FILLER_52_72 ();
 sg13g2_fill_2 FILLER_52_106 ();
 sg13g2_fill_1 FILLER_52_108 ();
 sg13g2_decap_4 FILLER_52_114 ();
 sg13g2_fill_2 FILLER_52_118 ();
 sg13g2_decap_8 FILLER_52_130 ();
 sg13g2_decap_8 FILLER_52_137 ();
 sg13g2_decap_8 FILLER_52_144 ();
 sg13g2_fill_2 FILLER_52_151 ();
 sg13g2_fill_2 FILLER_52_159 ();
 sg13g2_fill_2 FILLER_52_183 ();
 sg13g2_decap_4 FILLER_52_194 ();
 sg13g2_fill_1 FILLER_52_211 ();
 sg13g2_fill_1 FILLER_52_225 ();
 sg13g2_fill_2 FILLER_52_237 ();
 sg13g2_decap_4 FILLER_52_256 ();
 sg13g2_fill_2 FILLER_52_260 ();
 sg13g2_fill_2 FILLER_52_291 ();
 sg13g2_fill_2 FILLER_52_302 ();
 sg13g2_fill_1 FILLER_52_304 ();
 sg13g2_fill_2 FILLER_52_319 ();
 sg13g2_decap_8 FILLER_52_352 ();
 sg13g2_decap_8 FILLER_52_359 ();
 sg13g2_decap_8 FILLER_52_366 ();
 sg13g2_decap_8 FILLER_52_373 ();
 sg13g2_decap_8 FILLER_52_380 ();
 sg13g2_decap_8 FILLER_52_387 ();
 sg13g2_decap_8 FILLER_52_394 ();
 sg13g2_decap_8 FILLER_52_401 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_fill_1 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_27 ();
 sg13g2_decap_8 FILLER_53_34 ();
 sg13g2_fill_1 FILLER_53_41 ();
 sg13g2_decap_8 FILLER_53_71 ();
 sg13g2_decap_8 FILLER_53_78 ();
 sg13g2_fill_2 FILLER_53_85 ();
 sg13g2_fill_1 FILLER_53_87 ();
 sg13g2_decap_4 FILLER_53_108 ();
 sg13g2_fill_2 FILLER_53_112 ();
 sg13g2_decap_4 FILLER_53_154 ();
 sg13g2_fill_1 FILLER_53_158 ();
 sg13g2_fill_1 FILLER_53_170 ();
 sg13g2_fill_1 FILLER_53_217 ();
 sg13g2_fill_1 FILLER_53_229 ();
 sg13g2_decap_4 FILLER_53_240 ();
 sg13g2_fill_1 FILLER_53_244 ();
 sg13g2_fill_2 FILLER_53_261 ();
 sg13g2_fill_1 FILLER_53_263 ();
 sg13g2_decap_4 FILLER_53_326 ();
 sg13g2_fill_2 FILLER_53_330 ();
 sg13g2_decap_8 FILLER_53_336 ();
 sg13g2_fill_2 FILLER_53_343 ();
 sg13g2_fill_1 FILLER_53_345 ();
 sg13g2_decap_8 FILLER_53_351 ();
 sg13g2_decap_4 FILLER_53_358 ();
 sg13g2_fill_2 FILLER_53_362 ();
 sg13g2_decap_8 FILLER_53_369 ();
 sg13g2_decap_8 FILLER_53_376 ();
 sg13g2_decap_8 FILLER_53_383 ();
 sg13g2_decap_8 FILLER_53_390 ();
 sg13g2_decap_8 FILLER_53_397 ();
 sg13g2_decap_4 FILLER_53_404 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_4 FILLER_54_35 ();
 sg13g2_fill_1 FILLER_54_39 ();
 sg13g2_decap_8 FILLER_54_78 ();
 sg13g2_decap_8 FILLER_54_85 ();
 sg13g2_decap_4 FILLER_54_92 ();
 sg13g2_fill_2 FILLER_54_96 ();
 sg13g2_decap_8 FILLER_54_102 ();
 sg13g2_fill_2 FILLER_54_109 ();
 sg13g2_fill_1 FILLER_54_111 ();
 sg13g2_decap_4 FILLER_54_164 ();
 sg13g2_fill_2 FILLER_54_168 ();
 sg13g2_decap_4 FILLER_54_190 ();
 sg13g2_fill_1 FILLER_54_194 ();
 sg13g2_decap_4 FILLER_54_215 ();
 sg13g2_fill_1 FILLER_54_219 ();
 sg13g2_fill_2 FILLER_54_244 ();
 sg13g2_fill_1 FILLER_54_246 ();
 sg13g2_decap_8 FILLER_54_261 ();
 sg13g2_fill_1 FILLER_54_268 ();
 sg13g2_fill_1 FILLER_54_293 ();
 sg13g2_fill_1 FILLER_54_324 ();
 sg13g2_decap_8 FILLER_54_351 ();
 sg13g2_decap_8 FILLER_54_358 ();
 sg13g2_decap_8 FILLER_54_365 ();
 sg13g2_decap_8 FILLER_54_372 ();
 sg13g2_decap_8 FILLER_54_379 ();
 sg13g2_decap_8 FILLER_54_386 ();
 sg13g2_decap_8 FILLER_54_393 ();
 sg13g2_decap_8 FILLER_54_400 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_fill_1 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_59 ();
 sg13g2_fill_1 FILLER_55_66 ();
 sg13g2_fill_2 FILLER_55_75 ();
 sg13g2_fill_1 FILLER_55_77 ();
 sg13g2_fill_1 FILLER_55_82 ();
 sg13g2_fill_1 FILLER_55_87 ();
 sg13g2_decap_8 FILLER_55_113 ();
 sg13g2_decap_4 FILLER_55_120 ();
 sg13g2_fill_2 FILLER_55_124 ();
 sg13g2_fill_2 FILLER_55_134 ();
 sg13g2_decap_8 FILLER_55_166 ();
 sg13g2_decap_8 FILLER_55_173 ();
 sg13g2_fill_2 FILLER_55_180 ();
 sg13g2_decap_4 FILLER_55_190 ();
 sg13g2_fill_2 FILLER_55_202 ();
 sg13g2_decap_8 FILLER_55_213 ();
 sg13g2_fill_1 FILLER_55_220 ();
 sg13g2_fill_1 FILLER_55_243 ();
 sg13g2_fill_1 FILLER_55_267 ();
 sg13g2_fill_1 FILLER_55_325 ();
 sg13g2_decap_8 FILLER_55_343 ();
 sg13g2_decap_8 FILLER_55_350 ();
 sg13g2_decap_8 FILLER_55_357 ();
 sg13g2_decap_8 FILLER_55_364 ();
 sg13g2_decap_8 FILLER_55_371 ();
 sg13g2_decap_8 FILLER_55_378 ();
 sg13g2_decap_8 FILLER_55_385 ();
 sg13g2_decap_8 FILLER_55_392 ();
 sg13g2_decap_8 FILLER_55_399 ();
 sg13g2_fill_2 FILLER_55_406 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_48 ();
 sg13g2_fill_1 FILLER_56_55 ();
 sg13g2_fill_1 FILLER_56_65 ();
 sg13g2_decap_4 FILLER_56_132 ();
 sg13g2_fill_1 FILLER_56_136 ();
 sg13g2_fill_2 FILLER_56_146 ();
 sg13g2_fill_1 FILLER_56_148 ();
 sg13g2_fill_2 FILLER_56_153 ();
 sg13g2_fill_2 FILLER_56_181 ();
 sg13g2_fill_1 FILLER_56_191 ();
 sg13g2_fill_1 FILLER_56_205 ();
 sg13g2_fill_1 FILLER_56_239 ();
 sg13g2_fill_1 FILLER_56_251 ();
 sg13g2_fill_2 FILLER_56_262 ();
 sg13g2_fill_1 FILLER_56_264 ();
 sg13g2_fill_1 FILLER_56_315 ();
 sg13g2_decap_8 FILLER_56_342 ();
 sg13g2_decap_8 FILLER_56_349 ();
 sg13g2_decap_8 FILLER_56_356 ();
 sg13g2_decap_8 FILLER_56_363 ();
 sg13g2_fill_2 FILLER_56_370 ();
 sg13g2_decap_8 FILLER_56_376 ();
 sg13g2_decap_8 FILLER_56_383 ();
 sg13g2_decap_8 FILLER_56_390 ();
 sg13g2_decap_8 FILLER_56_397 ();
 sg13g2_decap_4 FILLER_56_404 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_21 ();
 sg13g2_fill_1 FILLER_57_48 ();
 sg13g2_decap_8 FILLER_57_180 ();
 sg13g2_decap_4 FILLER_57_187 ();
 sg13g2_fill_2 FILLER_57_191 ();
 sg13g2_decap_8 FILLER_57_207 ();
 sg13g2_decap_8 FILLER_57_214 ();
 sg13g2_decap_4 FILLER_57_221 ();
 sg13g2_fill_1 FILLER_57_234 ();
 sg13g2_fill_1 FILLER_57_245 ();
 sg13g2_fill_2 FILLER_57_250 ();
 sg13g2_fill_1 FILLER_57_252 ();
 sg13g2_decap_4 FILLER_57_261 ();
 sg13g2_decap_4 FILLER_57_270 ();
 sg13g2_fill_1 FILLER_57_274 ();
 sg13g2_fill_2 FILLER_57_280 ();
 sg13g2_fill_1 FILLER_57_285 ();
 sg13g2_fill_1 FILLER_57_300 ();
 sg13g2_fill_2 FILLER_57_343 ();
 sg13g2_fill_2 FILLER_57_349 ();
 sg13g2_fill_1 FILLER_57_351 ();
 sg13g2_fill_1 FILLER_57_357 ();
 sg13g2_decap_8 FILLER_57_393 ();
 sg13g2_decap_8 FILLER_57_400 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_fill_1 FILLER_58_28 ();
 sg13g2_fill_1 FILLER_58_66 ();
 sg13g2_fill_1 FILLER_58_115 ();
 sg13g2_decap_8 FILLER_58_156 ();
 sg13g2_fill_2 FILLER_58_163 ();
 sg13g2_fill_2 FILLER_58_173 ();
 sg13g2_fill_1 FILLER_58_175 ();
 sg13g2_fill_2 FILLER_58_260 ();
 sg13g2_decap_8 FILLER_58_267 ();
 sg13g2_fill_1 FILLER_58_274 ();
 sg13g2_fill_2 FILLER_58_283 ();
 sg13g2_fill_1 FILLER_58_285 ();
 sg13g2_fill_1 FILLER_58_329 ();
 sg13g2_decap_4 FILLER_58_404 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_4 FILLER_59_21 ();
 sg13g2_fill_1 FILLER_59_25 ();
 sg13g2_fill_1 FILLER_59_30 ();
 sg13g2_fill_2 FILLER_59_44 ();
 sg13g2_fill_1 FILLER_59_46 ();
 sg13g2_fill_2 FILLER_59_67 ();
 sg13g2_fill_1 FILLER_59_146 ();
 sg13g2_decap_4 FILLER_59_162 ();
 sg13g2_fill_1 FILLER_59_166 ();
 sg13g2_fill_1 FILLER_59_201 ();
 sg13g2_decap_8 FILLER_59_220 ();
 sg13g2_decap_4 FILLER_59_227 ();
 sg13g2_fill_1 FILLER_59_231 ();
 sg13g2_fill_2 FILLER_59_241 ();
 sg13g2_fill_1 FILLER_59_243 ();
 sg13g2_fill_2 FILLER_59_266 ();
 sg13g2_fill_1 FILLER_59_311 ();
 sg13g2_fill_2 FILLER_59_338 ();
 sg13g2_fill_1 FILLER_59_340 ();
 sg13g2_fill_2 FILLER_59_384 ();
 sg13g2_decap_4 FILLER_59_404 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_4 FILLER_60_70 ();
 sg13g2_fill_2 FILLER_60_109 ();
 sg13g2_decap_8 FILLER_60_168 ();
 sg13g2_fill_2 FILLER_60_184 ();
 sg13g2_fill_1 FILLER_60_186 ();
 sg13g2_decap_8 FILLER_60_195 ();
 sg13g2_decap_4 FILLER_60_202 ();
 sg13g2_decap_8 FILLER_60_218 ();
 sg13g2_fill_2 FILLER_60_230 ();
 sg13g2_fill_1 FILLER_60_232 ();
 sg13g2_fill_2 FILLER_60_248 ();
 sg13g2_fill_2 FILLER_60_302 ();
 sg13g2_fill_1 FILLER_60_304 ();
 sg13g2_fill_2 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_fill_2 FILLER_61_35 ();
 sg13g2_decap_4 FILLER_61_41 ();
 sg13g2_fill_2 FILLER_61_45 ();
 sg13g2_fill_2 FILLER_61_62 ();
 sg13g2_fill_2 FILLER_61_74 ();
 sg13g2_decap_4 FILLER_61_135 ();
 sg13g2_fill_2 FILLER_61_153 ();
 sg13g2_fill_1 FILLER_61_155 ();
 sg13g2_decap_8 FILLER_61_178 ();
 sg13g2_decap_8 FILLER_61_185 ();
 sg13g2_decap_8 FILLER_61_192 ();
 sg13g2_decap_8 FILLER_61_203 ();
 sg13g2_decap_8 FILLER_61_210 ();
 sg13g2_decap_8 FILLER_61_217 ();
 sg13g2_fill_2 FILLER_61_224 ();
 sg13g2_decap_8 FILLER_61_238 ();
 sg13g2_decap_4 FILLER_61_245 ();
 sg13g2_fill_1 FILLER_61_249 ();
 sg13g2_decap_8 FILLER_61_270 ();
 sg13g2_fill_2 FILLER_61_277 ();
 sg13g2_fill_2 FILLER_61_283 ();
 sg13g2_fill_1 FILLER_61_333 ();
 sg13g2_fill_1 FILLER_61_361 ();
 sg13g2_fill_2 FILLER_61_372 ();
 sg13g2_fill_1 FILLER_61_374 ();
 sg13g2_fill_2 FILLER_61_390 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_fill_1 FILLER_62_42 ();
 sg13g2_fill_2 FILLER_62_52 ();
 sg13g2_decap_4 FILLER_62_73 ();
 sg13g2_decap_8 FILLER_62_134 ();
 sg13g2_fill_1 FILLER_62_146 ();
 sg13g2_fill_1 FILLER_62_187 ();
 sg13g2_fill_2 FILLER_62_219 ();
 sg13g2_fill_1 FILLER_62_221 ();
 sg13g2_decap_8 FILLER_62_251 ();
 sg13g2_fill_1 FILLER_62_258 ();
 sg13g2_decap_8 FILLER_62_272 ();
 sg13g2_decap_8 FILLER_62_279 ();
 sg13g2_decap_8 FILLER_62_286 ();
 sg13g2_fill_2 FILLER_62_293 ();
 sg13g2_fill_2 FILLER_62_303 ();
 sg13g2_fill_1 FILLER_62_305 ();
 sg13g2_fill_2 FILLER_62_309 ();
 sg13g2_fill_2 FILLER_62_316 ();
 sg13g2_fill_2 FILLER_62_344 ();
 sg13g2_fill_2 FILLER_62_358 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_4 FILLER_63_28 ();
 sg13g2_fill_2 FILLER_63_57 ();
 sg13g2_fill_1 FILLER_63_59 ();
 sg13g2_decap_8 FILLER_63_68 ();
 sg13g2_decap_8 FILLER_63_75 ();
 sg13g2_decap_4 FILLER_63_82 ();
 sg13g2_fill_1 FILLER_63_86 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_fill_1 FILLER_63_112 ();
 sg13g2_fill_1 FILLER_63_126 ();
 sg13g2_fill_2 FILLER_63_143 ();
 sg13g2_fill_1 FILLER_63_163 ();
 sg13g2_fill_2 FILLER_63_169 ();
 sg13g2_fill_1 FILLER_63_171 ();
 sg13g2_decap_8 FILLER_63_198 ();
 sg13g2_decap_8 FILLER_63_257 ();
 sg13g2_decap_4 FILLER_63_264 ();
 sg13g2_decap_8 FILLER_63_272 ();
 sg13g2_fill_1 FILLER_63_279 ();
 sg13g2_fill_2 FILLER_63_288 ();
 sg13g2_fill_2 FILLER_63_324 ();
 sg13g2_fill_1 FILLER_63_326 ();
 sg13g2_fill_2 FILLER_63_339 ();
 sg13g2_fill_2 FILLER_63_381 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_fill_1 FILLER_64_21 ();
 sg13g2_decap_4 FILLER_64_72 ();
 sg13g2_decap_8 FILLER_64_102 ();
 sg13g2_fill_1 FILLER_64_109 ();
 sg13g2_decap_8 FILLER_64_203 ();
 sg13g2_fill_2 FILLER_64_210 ();
 sg13g2_fill_1 FILLER_64_212 ();
 sg13g2_fill_1 FILLER_64_235 ();
 sg13g2_fill_2 FILLER_64_254 ();
 sg13g2_fill_1 FILLER_64_256 ();
 sg13g2_fill_1 FILLER_64_323 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_4 FILLER_65_28 ();
 sg13g2_fill_2 FILLER_65_45 ();
 sg13g2_fill_1 FILLER_65_128 ();
 sg13g2_fill_1 FILLER_65_136 ();
 sg13g2_fill_1 FILLER_65_145 ();
 sg13g2_fill_1 FILLER_65_180 ();
 sg13g2_decap_8 FILLER_65_207 ();
 sg13g2_decap_4 FILLER_65_214 ();
 sg13g2_decap_8 FILLER_65_252 ();
 sg13g2_fill_2 FILLER_65_259 ();
 sg13g2_fill_2 FILLER_65_287 ();
 sg13g2_fill_1 FILLER_65_289 ();
 sg13g2_fill_1 FILLER_65_347 ();
 sg13g2_fill_1 FILLER_65_362 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_fill_1 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_4 FILLER_66_84 ();
 sg13g2_fill_1 FILLER_66_88 ();
 sg13g2_decap_8 FILLER_66_97 ();
 sg13g2_fill_1 FILLER_66_104 ();
 sg13g2_fill_2 FILLER_66_222 ();
 sg13g2_fill_1 FILLER_66_224 ();
 sg13g2_fill_2 FILLER_66_235 ();
 sg13g2_fill_1 FILLER_66_262 ();
 sg13g2_fill_1 FILLER_66_272 ();
 sg13g2_fill_1 FILLER_66_327 ();
 sg13g2_fill_2 FILLER_66_381 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_4 FILLER_67_42 ();
 sg13g2_fill_2 FILLER_67_54 ();
 sg13g2_decap_8 FILLER_67_60 ();
 sg13g2_decap_8 FILLER_67_67 ();
 sg13g2_decap_8 FILLER_67_74 ();
 sg13g2_decap_8 FILLER_67_81 ();
 sg13g2_decap_4 FILLER_67_88 ();
 sg13g2_fill_2 FILLER_67_92 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_fill_1 FILLER_67_112 ();
 sg13g2_fill_1 FILLER_67_121 ();
 sg13g2_fill_1 FILLER_67_127 ();
 sg13g2_fill_2 FILLER_67_206 ();
 sg13g2_fill_2 FILLER_67_212 ();
 sg13g2_fill_1 FILLER_67_214 ();
 sg13g2_decap_4 FILLER_67_240 ();
 sg13g2_fill_2 FILLER_67_244 ();
 sg13g2_fill_2 FILLER_67_255 ();
 sg13g2_fill_1 FILLER_67_257 ();
 sg13g2_fill_1 FILLER_67_305 ();
 sg13g2_fill_2 FILLER_67_389 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_4 FILLER_68_56 ();
 sg13g2_fill_2 FILLER_68_60 ();
 sg13g2_fill_2 FILLER_68_71 ();
 sg13g2_fill_1 FILLER_68_73 ();
 sg13g2_decap_8 FILLER_68_78 ();
 sg13g2_decap_4 FILLER_68_111 ();
 sg13g2_decap_4 FILLER_68_130 ();
 sg13g2_fill_1 FILLER_68_134 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_fill_2 FILLER_68_158 ();
 sg13g2_fill_1 FILLER_68_160 ();
 sg13g2_fill_2 FILLER_68_177 ();
 sg13g2_fill_1 FILLER_68_179 ();
 sg13g2_decap_8 FILLER_68_210 ();
 sg13g2_decap_8 FILLER_68_217 ();
 sg13g2_fill_1 FILLER_68_224 ();
 sg13g2_decap_4 FILLER_68_235 ();
 sg13g2_fill_2 FILLER_68_239 ();
 sg13g2_fill_2 FILLER_68_257 ();
 sg13g2_fill_2 FILLER_68_297 ();
 sg13g2_fill_1 FILLER_68_312 ();
 sg13g2_fill_1 FILLER_68_339 ();
 sg13g2_fill_2 FILLER_68_381 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_4 FILLER_69_49 ();
 sg13g2_fill_1 FILLER_69_82 ();
 sg13g2_fill_1 FILLER_69_109 ();
 sg13g2_decap_8 FILLER_69_136 ();
 sg13g2_fill_2 FILLER_69_143 ();
 sg13g2_decap_4 FILLER_69_150 ();
 sg13g2_fill_2 FILLER_69_154 ();
 sg13g2_decap_8 FILLER_69_169 ();
 sg13g2_decap_8 FILLER_69_176 ();
 sg13g2_decap_4 FILLER_69_187 ();
 sg13g2_decap_8 FILLER_69_195 ();
 sg13g2_decap_8 FILLER_69_202 ();
 sg13g2_decap_8 FILLER_69_209 ();
 sg13g2_decap_8 FILLER_69_216 ();
 sg13g2_decap_8 FILLER_69_223 ();
 sg13g2_decap_4 FILLER_69_236 ();
 sg13g2_fill_1 FILLER_69_252 ();
 sg13g2_fill_1 FILLER_69_299 ();
 sg13g2_fill_2 FILLER_69_310 ();
 sg13g2_fill_2 FILLER_69_326 ();
 sg13g2_fill_1 FILLER_69_361 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_4 FILLER_70_49 ();
 sg13g2_fill_2 FILLER_70_53 ();
 sg13g2_fill_1 FILLER_70_119 ();
 sg13g2_fill_1 FILLER_70_163 ();
 sg13g2_fill_1 FILLER_70_172 ();
 sg13g2_decap_4 FILLER_70_181 ();
 sg13g2_decap_4 FILLER_70_189 ();
 sg13g2_fill_2 FILLER_70_193 ();
 sg13g2_fill_2 FILLER_70_200 ();
 sg13g2_fill_1 FILLER_70_282 ();
 sg13g2_fill_2 FILLER_70_300 ();
 sg13g2_fill_2 FILLER_70_384 ();
 sg13g2_fill_1 FILLER_70_386 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_fill_2 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_74 ();
 sg13g2_fill_1 FILLER_71_81 ();
 sg13g2_fill_1 FILLER_71_86 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_fill_1 FILLER_71_98 ();
 sg13g2_fill_1 FILLER_71_112 ();
 sg13g2_fill_2 FILLER_71_121 ();
 sg13g2_fill_2 FILLER_71_180 ();
 sg13g2_decap_4 FILLER_71_197 ();
 sg13g2_fill_2 FILLER_71_235 ();
 sg13g2_decap_8 FILLER_71_241 ();
 sg13g2_decap_8 FILLER_71_248 ();
 sg13g2_decap_4 FILLER_71_255 ();
 sg13g2_fill_2 FILLER_71_259 ();
 sg13g2_fill_2 FILLER_71_347 ();
 sg13g2_fill_1 FILLER_71_354 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_fill_1 FILLER_72_70 ();
 sg13g2_fill_2 FILLER_72_106 ();
 sg13g2_decap_8 FILLER_72_118 ();
 sg13g2_fill_1 FILLER_72_125 ();
 sg13g2_decap_4 FILLER_72_230 ();
 sg13g2_fill_1 FILLER_72_234 ();
 sg13g2_fill_2 FILLER_72_248 ();
 sg13g2_fill_2 FILLER_72_268 ();
 sg13g2_fill_1 FILLER_72_299 ();
 sg13g2_fill_2 FILLER_72_327 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_fill_1 FILLER_73_63 ();
 sg13g2_fill_2 FILLER_73_90 ();
 sg13g2_fill_1 FILLER_73_92 ();
 sg13g2_fill_1 FILLER_73_101 ();
 sg13g2_decap_8 FILLER_73_118 ();
 sg13g2_decap_8 FILLER_73_125 ();
 sg13g2_decap_8 FILLER_73_132 ();
 sg13g2_decap_4 FILLER_73_139 ();
 sg13g2_fill_2 FILLER_73_155 ();
 sg13g2_fill_1 FILLER_73_157 ();
 sg13g2_decap_4 FILLER_73_203 ();
 sg13g2_fill_1 FILLER_73_207 ();
 sg13g2_decap_8 FILLER_73_217 ();
 sg13g2_decap_4 FILLER_73_224 ();
 sg13g2_fill_1 FILLER_73_228 ();
 sg13g2_fill_2 FILLER_73_241 ();
 sg13g2_fill_1 FILLER_73_256 ();
 sg13g2_fill_2 FILLER_73_279 ();
 sg13g2_fill_1 FILLER_73_378 ();
 sg13g2_fill_1 FILLER_73_396 ();
 sg13g2_fill_2 FILLER_73_406 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_fill_1 FILLER_74_63 ();
 sg13g2_decap_4 FILLER_74_90 ();
 sg13g2_fill_1 FILLER_74_94 ();
 sg13g2_decap_8 FILLER_74_107 ();
 sg13g2_decap_8 FILLER_74_114 ();
 sg13g2_fill_1 FILLER_74_121 ();
 sg13g2_decap_8 FILLER_74_138 ();
 sg13g2_decap_8 FILLER_74_145 ();
 sg13g2_decap_8 FILLER_74_152 ();
 sg13g2_decap_8 FILLER_74_159 ();
 sg13g2_decap_8 FILLER_74_166 ();
 sg13g2_decap_4 FILLER_74_173 ();
 sg13g2_fill_1 FILLER_74_177 ();
 sg13g2_fill_1 FILLER_74_182 ();
 sg13g2_fill_1 FILLER_74_195 ();
 sg13g2_fill_2 FILLER_74_265 ();
 sg13g2_fill_2 FILLER_74_282 ();
 sg13g2_fill_1 FILLER_74_284 ();
 sg13g2_fill_2 FILLER_74_309 ();
 sg13g2_fill_2 FILLER_74_360 ();
 sg13g2_fill_2 FILLER_74_367 ();
 sg13g2_fill_1 FILLER_74_369 ();
 sg13g2_fill_2 FILLER_74_388 ();
 sg13g2_fill_2 FILLER_74_397 ();
 sg13g2_fill_1 FILLER_74_399 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_4 FILLER_75_70 ();
 sg13g2_fill_1 FILLER_75_74 ();
 sg13g2_decap_8 FILLER_75_83 ();
 sg13g2_fill_2 FILLER_75_90 ();
 sg13g2_fill_1 FILLER_75_92 ();
 sg13g2_fill_2 FILLER_75_110 ();
 sg13g2_fill_2 FILLER_75_122 ();
 sg13g2_fill_2 FILLER_75_151 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_fill_2 FILLER_75_168 ();
 sg13g2_fill_1 FILLER_75_170 ();
 sg13g2_fill_2 FILLER_75_176 ();
 sg13g2_decap_8 FILLER_75_183 ();
 sg13g2_fill_1 FILLER_75_190 ();
 sg13g2_fill_1 FILLER_75_196 ();
 sg13g2_decap_8 FILLER_75_202 ();
 sg13g2_decap_8 FILLER_75_213 ();
 sg13g2_decap_4 FILLER_75_220 ();
 sg13g2_fill_1 FILLER_75_224 ();
 sg13g2_decap_8 FILLER_75_270 ();
 sg13g2_decap_8 FILLER_75_277 ();
 sg13g2_fill_2 FILLER_75_307 ();
 sg13g2_fill_2 FILLER_75_339 ();
 sg13g2_fill_1 FILLER_75_370 ();
 sg13g2_fill_2 FILLER_75_406 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_4 FILLER_76_201 ();
 sg13g2_fill_1 FILLER_76_253 ();
 sg13g2_decap_8 FILLER_76_272 ();
 sg13g2_fill_2 FILLER_76_288 ();
 sg13g2_fill_1 FILLER_76_290 ();
 sg13g2_fill_2 FILLER_76_331 ();
 sg13g2_fill_2 FILLER_76_346 ();
 sg13g2_fill_1 FILLER_76_348 ();
 sg13g2_fill_2 FILLER_76_358 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_fill_1 FILLER_77_128 ();
 sg13g2_fill_1 FILLER_77_185 ();
 sg13g2_fill_2 FILLER_77_225 ();
 sg13g2_fill_1 FILLER_77_227 ();
 sg13g2_fill_2 FILLER_77_254 ();
 sg13g2_fill_2 FILLER_77_325 ();
 sg13g2_fill_2 FILLER_77_353 ();
 sg13g2_fill_2 FILLER_77_360 ();
 sg13g2_fill_1 FILLER_77_362 ();
 sg13g2_fill_1 FILLER_77_401 ();
 sg13g2_fill_2 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_4 FILLER_78_84 ();
 sg13g2_fill_2 FILLER_78_88 ();
 sg13g2_fill_2 FILLER_78_123 ();
 sg13g2_decap_4 FILLER_78_136 ();
 sg13g2_fill_2 FILLER_78_166 ();
 sg13g2_fill_1 FILLER_78_220 ();
 sg13g2_decap_4 FILLER_78_321 ();
 sg13g2_fill_2 FILLER_78_325 ();
 sg13g2_fill_1 FILLER_78_379 ();
 sg13g2_decap_8 FILLER_78_402 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_fill_2 FILLER_79_98 ();
 sg13g2_fill_1 FILLER_79_100 ();
 sg13g2_fill_1 FILLER_79_110 ();
 sg13g2_fill_1 FILLER_79_121 ();
 sg13g2_decap_8 FILLER_79_132 ();
 sg13g2_decap_8 FILLER_79_139 ();
 sg13g2_fill_2 FILLER_79_146 ();
 sg13g2_fill_2 FILLER_79_204 ();
 sg13g2_fill_1 FILLER_79_232 ();
 sg13g2_fill_2 FILLER_79_255 ();
 sg13g2_fill_2 FILLER_79_271 ();
 sg13g2_fill_2 FILLER_79_290 ();
 sg13g2_fill_1 FILLER_79_292 ();
 sg13g2_fill_2 FILLER_79_328 ();
 sg13g2_fill_1 FILLER_79_330 ();
 sg13g2_fill_1 FILLER_79_344 ();
 sg13g2_fill_2 FILLER_79_366 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_fill_1 FILLER_80_111 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_8 FILLER_80_140 ();
 sg13g2_decap_8 FILLER_80_147 ();
 sg13g2_decap_8 FILLER_80_154 ();
 sg13g2_decap_8 FILLER_80_161 ();
 sg13g2_fill_2 FILLER_80_175 ();
 sg13g2_fill_1 FILLER_80_177 ();
 sg13g2_fill_2 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_193 ();
 sg13g2_decap_8 FILLER_80_200 ();
 sg13g2_decap_8 FILLER_80_207 ();
 sg13g2_fill_2 FILLER_80_214 ();
 sg13g2_fill_1 FILLER_80_216 ();
 sg13g2_decap_8 FILLER_80_221 ();
 sg13g2_decap_4 FILLER_80_228 ();
 sg13g2_decap_4 FILLER_80_239 ();
 sg13g2_fill_1 FILLER_80_243 ();
 sg13g2_fill_1 FILLER_80_263 ();
 sg13g2_fill_2 FILLER_80_268 ();
 sg13g2_fill_1 FILLER_80_270 ();
 sg13g2_fill_1 FILLER_80_288 ();
 sg13g2_fill_1 FILLER_80_293 ();
 sg13g2_decap_8 FILLER_80_320 ();
 sg13g2_decap_8 FILLER_80_327 ();
 sg13g2_fill_1 FILLER_80_334 ();
 sg13g2_fill_2 FILLER_80_345 ();
 sg13g2_decap_8 FILLER_80_385 ();
 sg13g2_decap_8 FILLER_80_392 ();
 sg13g2_decap_8 FILLER_80_399 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net210;
 assign uio_oe[1] = net211;
 assign uio_oe[2] = net212;
 assign uio_oe[3] = net213;
 assign uio_oe[4] = net214;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[5] = net9;
 assign uio_out[6] = net10;
 assign uio_out[7] = net11;
endmodule

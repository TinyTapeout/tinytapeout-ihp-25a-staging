module tt_um_strau0106_simple_viii (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire clknet_leaf_0_clk;
 wire \cpu_instance.addr_reg_op[0] ;
 wire \cpu_instance.addr_reg_op[1] ;
 wire \cpu_instance.addr_reg_op[2] ;
 wire \cpu_instance.addr_sel ;
 wire \cpu_instance.alu_instance.op[0] ;
 wire \cpu_instance.alu_instance.op[1] ;
 wire \cpu_instance.alu_instance.op[2] ;
 wire \cpu_instance.alu_instance.op[3] ;
 wire \cpu_instance.ctrl_instance.flag_carry ;
 wire \cpu_instance.ctrl_instance.flag_zero ;
 wire \cpu_instance.ctrl_instance.jmp_op_addr_sel ;
 wire \cpu_instance.ctrl_instance.mem_ctrl_op[0] ;
 wire \cpu_instance.ctrl_instance.mem_ctrl_op[1] ;
 wire \cpu_instance.ctrl_instance.mem_ctrl_op[2] ;
 wire \cpu_instance.ctrl_instance.mem_op_done ;
 wire \cpu_instance.ctrl_instance.mux_sel[0] ;
 wire \cpu_instance.ctrl_instance.mux_sel[1] ;
 wire \cpu_instance.ctrl_instance.mux_sel[2] ;
 wire \cpu_instance.ctrl_instance.reg_op ;
 wire \cpu_instance.ctrl_instance.reg_sel_1[0] ;
 wire \cpu_instance.ctrl_instance.reg_sel_1[1] ;
 wire \cpu_instance.ctrl_instance.reg_sel_2[0] ;
 wire \cpu_instance.ctrl_instance.reg_sel_2[1] ;
 wire \cpu_instance.ctrl_instance.reg_sel_in[0] ;
 wire \cpu_instance.ctrl_instance.reg_sel_in[1] ;
 wire \cpu_instance.ctrl_instance.state[0] ;
 wire \cpu_instance.ctrl_instance.state[1] ;
 wire \cpu_instance.ctrl_instance.state[2] ;
 wire \cpu_instance.ctrl_instance.state[3] ;
 wire \cpu_instance.ctrl_instance.state[4] ;
 wire \cpu_instance.ctrl_instance.state[5] ;
 wire \cpu_instance.ctrl_instance.state[6] ;
 wire \cpu_instance.ctrl_instance.state[7] ;
 wire \cpu_instance.ctrl_instance.use_register_bank_in ;
 wire \cpu_instance.ctrl_instance.use_register_bank_out_1 ;
 wire \cpu_instance.mem_instance.addr[24] ;
 wire \cpu_instance.mem_instance.bus_data_out[0] ;
 wire \cpu_instance.mem_instance.bus_data_out[1] ;
 wire \cpu_instance.mem_instance.bus_data_out[2] ;
 wire \cpu_instance.mem_instance.bus_data_out[3] ;
 wire \cpu_instance.mem_instance.bus_data_out[4] ;
 wire \cpu_instance.mem_instance.bus_data_out[5] ;
 wire \cpu_instance.mem_instance.bus_data_out[6] ;
 wire \cpu_instance.mem_instance.bus_data_out[7] ;
 wire \cpu_instance.mem_instance.data_qi_mo[0] ;
 wire \cpu_instance.mem_instance.data_qi_mo[1] ;
 wire \cpu_instance.mem_instance.data_qi_mo[2] ;
 wire \cpu_instance.mem_instance.data_qi_mo[3] ;
 wire \cpu_instance.mem_instance.data_qi_mo[4] ;
 wire \cpu_instance.mem_instance.data_qi_mo[5] ;
 wire \cpu_instance.mem_instance.data_qi_mo[6] ;
 wire \cpu_instance.mem_instance.data_qi_mo[7] ;
 wire \cpu_instance.mem_instance.data_qo_mi[0] ;
 wire \cpu_instance.mem_instance.data_qo_mi[1] ;
 wire \cpu_instance.mem_instance.data_qo_mi[2] ;
 wire \cpu_instance.mem_instance.data_qo_mi[3] ;
 wire \cpu_instance.mem_instance.data_qo_mi[4] ;
 wire \cpu_instance.mem_instance.data_qo_mi[5] ;
 wire \cpu_instance.mem_instance.data_qo_mi[6] ;
 wire \cpu_instance.mem_instance.data_qo_mi[7] ;
 wire \cpu_instance.mem_instance.data_ready ;
 wire \cpu_instance.mem_instance.data_req ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][0] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][10] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][11] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][12] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][13] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][14] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][15] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][1] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][2] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][3] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][4] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][5] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][6] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][7] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][8] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][9] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][0] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][10] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][11] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][12] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][13] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][14] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][15] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][1] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][2] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][3] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][4] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][5] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][6] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][7] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][8] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][9] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[0] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[10] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[11] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[12] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[13] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[14] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[15] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[16] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[17] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[18] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[19] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[1] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[20] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[21] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[22] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[23] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[24] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[25] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[26] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[27] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[28] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[29] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[2] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[30] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[31] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[32] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[33] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[34] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[35] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[36] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[37] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[38] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[39] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[3] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[40] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[41] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[42] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[43] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[44] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[45] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[46] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[47] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[48] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[49] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[4] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[50] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[51] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[52] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[53] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[54] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[55] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[56] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[57] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[58] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[59] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[5] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[60] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[61] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[62] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[63] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[6] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[7] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[8] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[9] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.stall_txn ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.start_read ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.start_write ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.state[0] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.state[1] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.state[2] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.state[3] ;
 wire \cpu_instance.mem_instance.mem_ctrl_instance.stop_txn ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[10] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[11] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[12] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[13] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[14] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[15] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[16] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[17] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[18] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[19] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[1] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[20] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[21] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[22] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[23] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[2] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[3] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[4] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[5] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[6] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[7] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[8] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.addr[9] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[1] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[1] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[2] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.is_writing ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.last_ram_a_sel ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[1] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[2] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_clk_out ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_data_oe[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[0] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[1] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[2] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[3] ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.spi_ram_a_select ;
 wire \cpu_instance.mem_instance.qspi_ctrl_instance.stop_txn_reg ;
 wire \cpu_instance.registers_instance.register_bank[10][0] ;
 wire \cpu_instance.registers_instance.register_bank[10][1] ;
 wire \cpu_instance.registers_instance.register_bank[10][2] ;
 wire \cpu_instance.registers_instance.register_bank[10][3] ;
 wire \cpu_instance.registers_instance.register_bank[10][4] ;
 wire \cpu_instance.registers_instance.register_bank[10][5] ;
 wire \cpu_instance.registers_instance.register_bank[10][6] ;
 wire \cpu_instance.registers_instance.register_bank[10][7] ;
 wire \cpu_instance.registers_instance.register_bank[11][0] ;
 wire \cpu_instance.registers_instance.register_bank[11][1] ;
 wire \cpu_instance.registers_instance.register_bank[11][2] ;
 wire \cpu_instance.registers_instance.register_bank[11][3] ;
 wire \cpu_instance.registers_instance.register_bank[11][4] ;
 wire \cpu_instance.registers_instance.register_bank[11][5] ;
 wire \cpu_instance.registers_instance.register_bank[11][6] ;
 wire \cpu_instance.registers_instance.register_bank[11][7] ;
 wire \cpu_instance.registers_instance.register_bank[12][0] ;
 wire \cpu_instance.registers_instance.register_bank[12][1] ;
 wire \cpu_instance.registers_instance.register_bank[12][2] ;
 wire \cpu_instance.registers_instance.register_bank[12][3] ;
 wire \cpu_instance.registers_instance.register_bank[12][4] ;
 wire \cpu_instance.registers_instance.register_bank[12][5] ;
 wire \cpu_instance.registers_instance.register_bank[12][6] ;
 wire \cpu_instance.registers_instance.register_bank[12][7] ;
 wire \cpu_instance.registers_instance.register_bank[13][0] ;
 wire \cpu_instance.registers_instance.register_bank[13][1] ;
 wire \cpu_instance.registers_instance.register_bank[13][2] ;
 wire \cpu_instance.registers_instance.register_bank[13][3] ;
 wire \cpu_instance.registers_instance.register_bank[13][4] ;
 wire \cpu_instance.registers_instance.register_bank[13][5] ;
 wire \cpu_instance.registers_instance.register_bank[13][6] ;
 wire \cpu_instance.registers_instance.register_bank[13][7] ;
 wire \cpu_instance.registers_instance.register_bank[14][0] ;
 wire \cpu_instance.registers_instance.register_bank[14][1] ;
 wire \cpu_instance.registers_instance.register_bank[14][2] ;
 wire \cpu_instance.registers_instance.register_bank[14][3] ;
 wire \cpu_instance.registers_instance.register_bank[14][4] ;
 wire \cpu_instance.registers_instance.register_bank[14][5] ;
 wire \cpu_instance.registers_instance.register_bank[14][6] ;
 wire \cpu_instance.registers_instance.register_bank[14][7] ;
 wire \cpu_instance.registers_instance.register_bank[15][0] ;
 wire \cpu_instance.registers_instance.register_bank[15][1] ;
 wire \cpu_instance.registers_instance.register_bank[15][2] ;
 wire \cpu_instance.registers_instance.register_bank[15][3] ;
 wire \cpu_instance.registers_instance.register_bank[15][4] ;
 wire \cpu_instance.registers_instance.register_bank[15][5] ;
 wire \cpu_instance.registers_instance.register_bank[15][6] ;
 wire \cpu_instance.registers_instance.register_bank[15][7] ;
 wire \cpu_instance.registers_instance.register_bank[8][0] ;
 wire \cpu_instance.registers_instance.register_bank[8][1] ;
 wire \cpu_instance.registers_instance.register_bank[8][2] ;
 wire \cpu_instance.registers_instance.register_bank[8][3] ;
 wire \cpu_instance.registers_instance.register_bank[8][4] ;
 wire \cpu_instance.registers_instance.register_bank[8][5] ;
 wire \cpu_instance.registers_instance.register_bank[8][6] ;
 wire \cpu_instance.registers_instance.register_bank[8][7] ;
 wire \cpu_instance.registers_instance.register_bank[9][0] ;
 wire \cpu_instance.registers_instance.register_bank[9][1] ;
 wire \cpu_instance.registers_instance.register_bank[9][2] ;
 wire \cpu_instance.registers_instance.register_bank[9][3] ;
 wire \cpu_instance.registers_instance.register_bank[9][4] ;
 wire \cpu_instance.registers_instance.register_bank[9][5] ;
 wire \cpu_instance.registers_instance.register_bank[9][6] ;
 wire \cpu_instance.registers_instance.register_bank[9][7] ;
 wire \cpu_instance.registers_instance.registers[0][0] ;
 wire \cpu_instance.registers_instance.registers[0][1] ;
 wire \cpu_instance.registers_instance.registers[0][2] ;
 wire \cpu_instance.registers_instance.registers[0][3] ;
 wire \cpu_instance.registers_instance.registers[0][4] ;
 wire \cpu_instance.registers_instance.registers[0][5] ;
 wire \cpu_instance.registers_instance.registers[0][6] ;
 wire \cpu_instance.registers_instance.registers[0][7] ;
 wire \cpu_instance.registers_instance.registers[1][0] ;
 wire \cpu_instance.registers_instance.registers[1][1] ;
 wire \cpu_instance.registers_instance.registers[1][2] ;
 wire \cpu_instance.registers_instance.registers[1][3] ;
 wire \cpu_instance.registers_instance.registers[1][4] ;
 wire \cpu_instance.registers_instance.registers[1][5] ;
 wire \cpu_instance.registers_instance.registers[1][6] ;
 wire \cpu_instance.registers_instance.registers[1][7] ;
 wire \cpu_instance.registers_instance.registers[2][0] ;
 wire \cpu_instance.registers_instance.registers[2][1] ;
 wire \cpu_instance.registers_instance.registers[2][2] ;
 wire \cpu_instance.registers_instance.registers[2][3] ;
 wire \cpu_instance.registers_instance.registers[2][4] ;
 wire \cpu_instance.registers_instance.registers[2][5] ;
 wire \cpu_instance.registers_instance.registers[2][6] ;
 wire \cpu_instance.registers_instance.registers[2][7] ;
 wire net12;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;

 sg13g2_inv_1 _2202_ (.Y(_1276_),
    .A(uo_out[2]));
 sg13g2_inv_1 _2203_ (.Y(_1277_),
    .A(\cpu_instance.registers_instance.registers[2][4] ));
 sg13g2_inv_1 _2204_ (.Y(_1278_),
    .A(\cpu_instance.registers_instance.registers[2][2] ));
 sg13g2_inv_1 _2205_ (.Y(_1279_),
    .A(\cpu_instance.registers_instance.registers[1][4] ));
 sg13g2_inv_1 _2206_ (.Y(_1280_),
    .A(\cpu_instance.registers_instance.registers[1][2] ));
 sg13g2_inv_1 _2207_ (.Y(_1281_),
    .A(\cpu_instance.registers_instance.registers[0][7] ));
 sg13g2_inv_1 _2208_ (.Y(_1282_),
    .A(\cpu_instance.registers_instance.registers[0][2] ));
 sg13g2_inv_1 _2209_ (.Y(_1283_),
    .A(net392));
 sg13g2_inv_4 _2210_ (.A(net721),
    .Y(_1284_));
 sg13g2_inv_4 _2211_ (.A(net725),
    .Y(_1285_));
 sg13g2_inv_1 _2212_ (.Y(_1286_),
    .A(\cpu_instance.alu_instance.op[3] ));
 sg13g2_inv_2 _2213_ (.Y(_1287_),
    .A(\cpu_instance.ctrl_instance.reg_sel_in[1] ));
 sg13g2_inv_2 _2214_ (.Y(_1288_),
    .A(\cpu_instance.ctrl_instance.reg_sel_in[0] ));
 sg13g2_inv_1 _2215_ (.Y(_1289_),
    .A(net728));
 sg13g2_inv_2 _2216_ (.Y(_1290_),
    .A(net733));
 sg13g2_inv_1 _2217_ (.Y(_1291_),
    .A(net400));
 sg13g2_inv_1 _2218_ (.Y(_1292_),
    .A(_0032_));
 sg13g2_inv_1 _2219_ (.Y(_1293_),
    .A(_0031_));
 sg13g2_inv_1 _2220_ (.Y(_1294_),
    .A(_0034_));
 sg13g2_inv_1 _2221_ (.Y(_1295_),
    .A(_0036_));
 sg13g2_inv_1 _2222_ (.Y(_1296_),
    .A(_0035_));
 sg13g2_inv_4 _2223_ (.A(\cpu_instance.ctrl_instance.reg_sel_2[1] ),
    .Y(_1297_));
 sg13g2_inv_1 _2224_ (.Y(_1298_),
    .A(_0037_));
 sg13g2_inv_1 _2225_ (.Y(_1299_),
    .A(_0044_));
 sg13g2_inv_1 _2226_ (.Y(_1300_),
    .A(\cpu_instance.ctrl_instance.mux_sel[0] ));
 sg13g2_inv_1 _2227_ (.Y(_1301_),
    .A(_0020_));
 sg13g2_inv_1 _2228_ (.Y(_1302_),
    .A(net359));
 sg13g2_inv_1 _2229_ (.Y(_1303_),
    .A(net771));
 sg13g2_inv_1 _2230_ (.Y(_1304_),
    .A(net395));
 sg13g2_inv_1 _2231_ (.Y(_1305_),
    .A(net816));
 sg13g2_inv_1 _2232_ (.Y(_1306_),
    .A(net804));
 sg13g2_inv_1 _2233_ (.Y(_1307_),
    .A(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ));
 sg13g2_inv_1 _2234_ (.Y(_1308_),
    .A(net364));
 sg13g2_inv_1 _2235_ (.Y(_1309_),
    .A(net367));
 sg13g2_inv_1 _2236_ (.Y(_1310_),
    .A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[7] ));
 sg13g2_inv_1 _2237_ (.Y(_1311_),
    .A(net340));
 sg13g2_inv_1 _2238_ (.Y(_1312_),
    .A(net343));
 sg13g2_inv_1 _2239_ (.Y(_1313_),
    .A(net333));
 sg13g2_inv_1 _2240_ (.Y(_1314_),
    .A(net387));
 sg13g2_inv_1 _2241_ (.Y(_1315_),
    .A(net461));
 sg13g2_or2_1 _2242_ (.X(_1316_),
    .B(net356),
    .A(net445));
 sg13g2_o21ai_1 _2243_ (.B1(net769),
    .Y(_1317_),
    .A1(net505),
    .A2(net715));
 sg13g2_and2_2 _2244_ (.A(net719),
    .B(net773),
    .X(_1318_));
 sg13g2_nor2_2 _2245_ (.A(net718),
    .B(net741),
    .Y(_1319_));
 sg13g2_nand2_2 _2246_ (.Y(_1320_),
    .A(net585),
    .B(net769));
 sg13g2_a22oi_1 _2247_ (.Y(_1321_),
    .B1(_1319_),
    .B2(net570),
    .A2(_1318_),
    .A1(net583));
 sg13g2_nand3_1 _2248_ (.B(_1320_),
    .C(_1321_),
    .A(_1317_),
    .Y(_0002_));
 sg13g2_nor2b_1 _2249_ (.A(\cpu_instance.alu_instance.op[0] ),
    .B_N(\cpu_instance.alu_instance.op[1] ),
    .Y(_1322_));
 sg13g2_nand2b_2 _2250_ (.Y(_1323_),
    .B(\cpu_instance.alu_instance.op[1] ),
    .A_N(\cpu_instance.alu_instance.op[0] ));
 sg13g2_nor2_2 _2251_ (.A(\cpu_instance.alu_instance.op[3] ),
    .B(\cpu_instance.alu_instance.op[2] ),
    .Y(_1324_));
 sg13g2_and2_2 _2252_ (.A(_1322_),
    .B(_1324_),
    .X(_1325_));
 sg13g2_nand2_1 _2253_ (.Y(_1326_),
    .A(_1322_),
    .B(_1324_));
 sg13g2_nand3b_1 _2254_ (.B(net729),
    .C(\cpu_instance.registers_instance.registers[2][2] ),
    .Y(_1327_),
    .A_N(net733));
 sg13g2_nor2_1 _2255_ (.A(net729),
    .B(_1290_),
    .Y(_1328_));
 sg13g2_nor2_2 _2256_ (.A(net716),
    .B(_1290_),
    .Y(_1329_));
 sg13g2_nand3_1 _2257_ (.B(net729),
    .C(net733),
    .A(uo_out[2]),
    .Y(_1330_));
 sg13g2_nor2_2 _2258_ (.A(net729),
    .B(net733),
    .Y(_1331_));
 sg13g2_or2_1 _2259_ (.X(_1332_),
    .B(net733),
    .A(net729));
 sg13g2_nand2b_1 _2260_ (.Y(_1333_),
    .B(\cpu_instance.registers_instance.registers[1][2] ),
    .A_N(net729));
 sg13g2_nand4_1 _2261_ (.B(_1330_),
    .C(_1332_),
    .A(_1327_),
    .Y(_1334_),
    .D(_1333_));
 sg13g2_nor3_1 _2262_ (.A(\cpu_instance.registers_instance.registers[0][2] ),
    .B(net728),
    .C(net732),
    .Y(_1335_));
 sg13g2_mux4_1 _2263_ (.S0(\cpu_instance.ctrl_instance.reg_sel_1[0] ),
    .A0(\cpu_instance.registers_instance.registers[0][2] ),
    .A1(\cpu_instance.registers_instance.registers[1][2] ),
    .A2(\cpu_instance.registers_instance.registers[2][2] ),
    .A3(uo_out[2]),
    .S1(\cpu_instance.ctrl_instance.reg_sel_1[1] ),
    .X(_1336_));
 sg13g2_mux4_1 _2264_ (.S0(_1290_),
    .A0(_1276_),
    .A1(_1278_),
    .A2(_1280_),
    .A3(_1282_),
    .S1(_1289_),
    .X(_1337_));
 sg13g2_nand3b_1 _2265_ (.B(net726),
    .C(\cpu_instance.registers_instance.registers[2][3] ),
    .Y(_1338_),
    .A_N(net730));
 sg13g2_nand3b_1 _2266_ (.B(net730),
    .C(net726),
    .Y(_1339_),
    .A_N(_0036_));
 sg13g2_nand3b_1 _2267_ (.B(net731),
    .C(\cpu_instance.registers_instance.registers[1][3] ),
    .Y(_1340_),
    .A_N(net727));
 sg13g2_nand3_1 _2268_ (.B(_1339_),
    .C(_1340_),
    .A(_1338_),
    .Y(_1341_));
 sg13g2_or3_1 _2269_ (.A(net726),
    .B(net730),
    .C(_0035_),
    .X(_1342_));
 sg13g2_and4_1 _2270_ (.A(_1338_),
    .B(_1339_),
    .C(_1340_),
    .D(_1342_),
    .X(_1343_));
 sg13g2_nand4_1 _2271_ (.B(_1339_),
    .C(_1340_),
    .A(_1338_),
    .Y(_1344_),
    .D(_1342_));
 sg13g2_nand3b_1 _2272_ (.B(net730),
    .C(\cpu_instance.registers_instance.registers[1][0] ),
    .Y(_1345_),
    .A_N(net726));
 sg13g2_nand3b_1 _2273_ (.B(net730),
    .C(net726),
    .Y(_1346_),
    .A_N(_0032_));
 sg13g2_nand3b_1 _2274_ (.B(net726),
    .C(\cpu_instance.registers_instance.registers[2][0] ),
    .Y(_1347_),
    .A_N(net730));
 sg13g2_nand3_1 _2275_ (.B(_1346_),
    .C(_1347_),
    .A(_1345_),
    .Y(_1348_));
 sg13g2_mux4_1 _2276_ (.S0(net716),
    .A0(\cpu_instance.registers_instance.registers[2][0] ),
    .A1(\cpu_instance.registers_instance.registers[0][0] ),
    .A2(_1292_),
    .A3(\cpu_instance.registers_instance.registers[1][0] ),
    .S1(net730),
    .X(_1349_));
 sg13g2_nand3b_1 _2277_ (.B(net730),
    .C(\cpu_instance.registers_instance.registers[1][1] ),
    .Y(_1350_),
    .A_N(net727));
 sg13g2_nand3b_1 _2278_ (.B(net731),
    .C(net726),
    .Y(_1351_),
    .A_N(_0034_));
 sg13g2_nand3b_1 _2279_ (.B(net726),
    .C(\cpu_instance.registers_instance.registers[2][1] ),
    .Y(_1352_),
    .A_N(net731));
 sg13g2_nand3_1 _2280_ (.B(_1351_),
    .C(_1352_),
    .A(_1350_),
    .Y(_1353_));
 sg13g2_mux4_1 _2281_ (.S0(net716),
    .A0(\cpu_instance.registers_instance.registers[2][1] ),
    .A1(\cpu_instance.registers_instance.registers[0][1] ),
    .A2(_1294_),
    .A3(\cpu_instance.registers_instance.registers[1][1] ),
    .S1(net732),
    .X(_1354_));
 sg13g2_nor4_2 _2282_ (.A(_1336_),
    .B(net706),
    .C(_1349_),
    .Y(_1355_),
    .D(_1354_));
 sg13g2_nor4_2 _2283_ (.A(_1337_),
    .B(net706),
    .C(_1349_),
    .Y(_1356_),
    .D(_1354_));
 sg13g2_or3_1 _2284_ (.A(net727),
    .B(net731),
    .C(_0031_),
    .X(_1357_));
 sg13g2_and4_1 _2285_ (.A(_1345_),
    .B(_1346_),
    .C(_1347_),
    .D(_1357_),
    .X(_1358_));
 sg13g2_nor4_2 _2286_ (.A(_1336_),
    .B(net706),
    .C(_1354_),
    .Y(_1359_),
    .D(net705));
 sg13g2_or3_1 _2287_ (.A(net727),
    .B(net731),
    .C(_0033_),
    .X(_1360_));
 sg13g2_and4_2 _2288_ (.A(_1350_),
    .B(_1351_),
    .C(_1352_),
    .D(_1360_),
    .X(_1361_));
 sg13g2_nor4_2 _2289_ (.A(_1337_),
    .B(net706),
    .C(_1349_),
    .Y(_1362_),
    .D(net704));
 sg13g2_nor2_1 _2290_ (.A(_1334_),
    .B(_1341_),
    .Y(_1363_));
 sg13g2_nor2_1 _2291_ (.A(_1348_),
    .B(_1353_),
    .Y(_1364_));
 sg13g2_nor4_2 _2292_ (.A(_1334_),
    .B(_1341_),
    .C(_1348_),
    .Y(_1365_),
    .D(_1353_));
 sg13g2_nand3_1 _2293_ (.B(_0033_),
    .C(_1331_),
    .A(\cpu_instance.registers_instance.registers[0][1] ),
    .Y(_1366_));
 sg13g2_and2_1 _2294_ (.A(_0033_),
    .B(_0035_),
    .X(_1367_));
 sg13g2_a22oi_1 _2295_ (.Y(_1368_),
    .B1(_1335_),
    .B2(_1367_),
    .A2(_1331_),
    .A1(\cpu_instance.registers_instance.registers[0][0] ));
 sg13g2_o21ai_1 _2296_ (.B1(_1366_),
    .Y(_1369_),
    .A1(_1293_),
    .A2(_1368_));
 sg13g2_nor2_2 _2297_ (.A(_1365_),
    .B(_1369_),
    .Y(_1370_));
 sg13g2_or2_2 _2298_ (.X(_1371_),
    .B(_1369_),
    .A(_1365_));
 sg13g2_nor4_2 _2299_ (.A(_1336_),
    .B(net706),
    .C(_1349_),
    .Y(_1372_),
    .D(net704));
 sg13g2_nor4_2 _2300_ (.A(_1337_),
    .B(_1344_),
    .C(_1354_),
    .Y(_1373_),
    .D(net705));
 sg13g2_nor4_2 _2301_ (.A(_1336_),
    .B(_1344_),
    .C(_1354_),
    .Y(_1374_),
    .D(net705));
 sg13g2_nor4_2 _2302_ (.A(_1336_),
    .B(_1344_),
    .C(_1349_),
    .Y(_1375_),
    .D(net704));
 sg13g2_nor4_2 _2303_ (.A(_1337_),
    .B(net706),
    .C(_1354_),
    .Y(_1376_),
    .D(net705));
 sg13g2_nand2_1 _2304_ (.Y(_1377_),
    .A(\cpu_instance.registers_instance.register_bank[13][5] ),
    .B(_1376_));
 sg13g2_nor4_2 _2305_ (.A(_1337_),
    .B(_1344_),
    .C(_1349_),
    .Y(_1378_),
    .D(net704));
 sg13g2_nor4_2 _2306_ (.A(_1337_),
    .B(net706),
    .C(net705),
    .Y(_1379_),
    .D(net704));
 sg13g2_nor4_2 _2307_ (.A(_1336_),
    .B(net706),
    .C(net705),
    .Y(_1380_),
    .D(net704));
 sg13g2_nor4_2 _2308_ (.A(_1336_),
    .B(_1344_),
    .C(net705),
    .Y(_1381_),
    .D(net704));
 sg13g2_nor4_2 _2309_ (.A(_1337_),
    .B(_1344_),
    .C(net705),
    .Y(_1382_),
    .D(_1361_));
 sg13g2_nor4_2 _2310_ (.A(_1337_),
    .B(_1344_),
    .C(_1349_),
    .Y(_1383_),
    .D(_1354_));
 sg13g2_a22oi_1 _2311_ (.Y(_1384_),
    .B1(_1373_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[45] ),
    .A2(_1372_),
    .A1(\cpu_instance.registers_instance.register_bank[10][5] ));
 sg13g2_a22oi_1 _2312_ (.Y(_1385_),
    .B1(_1379_),
    .B2(\cpu_instance.registers_instance.register_bank[15][5] ),
    .A2(_1362_),
    .A1(\cpu_instance.registers_instance.register_bank[14][5] ));
 sg13g2_a22oi_1 _2313_ (.Y(_1386_),
    .B1(_1359_),
    .B2(\cpu_instance.registers_instance.register_bank[9][5] ),
    .A2(_1355_),
    .A1(\cpu_instance.registers_instance.register_bank[8][5] ));
 sg13g2_a22oi_1 _2314_ (.Y(_1387_),
    .B1(_1382_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[61] ),
    .A2(_1378_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[53] ));
 sg13g2_a22oi_1 _2315_ (.Y(_1388_),
    .B1(_1383_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[37] ),
    .A2(_1380_),
    .A1(\cpu_instance.registers_instance.register_bank[11][5] ));
 sg13g2_nand4_1 _2316_ (.B(_1386_),
    .C(_1387_),
    .A(_1384_),
    .Y(_1389_),
    .D(_1388_));
 sg13g2_a22oi_1 _2317_ (.Y(_1390_),
    .B1(_1381_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[29] ),
    .A2(_1374_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[13] ));
 sg13g2_a22oi_1 _2318_ (.Y(_1391_),
    .B1(_1375_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[21] ),
    .A2(_1356_),
    .A1(\cpu_instance.registers_instance.register_bank[12][5] ));
 sg13g2_nand4_1 _2319_ (.B(_1385_),
    .C(_1390_),
    .A(_1377_),
    .Y(_1392_),
    .D(_1391_));
 sg13g2_nor3_2 _2320_ (.A(_1371_),
    .B(_1389_),
    .C(_1392_),
    .Y(_1393_));
 sg13g2_o21ai_1 _2321_ (.B1(\cpu_instance.ctrl_instance.use_register_bank_out_1 ),
    .Y(_1394_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[5] ),
    .A2(_1370_));
 sg13g2_o21ai_1 _2322_ (.B1(_1290_),
    .Y(_1395_),
    .A1(\cpu_instance.registers_instance.registers[2][5] ),
    .A2(net716));
 sg13g2_a22oi_1 _2323_ (.Y(_1396_),
    .B1(_1329_),
    .B2(uo_out[5]),
    .A2(net716),
    .A1(\cpu_instance.registers_instance.registers[1][5] ));
 sg13g2_o21ai_1 _2324_ (.B1(_1285_),
    .Y(_1397_),
    .A1(\cpu_instance.registers_instance.registers[0][5] ),
    .A2(_1332_));
 sg13g2_a21o_1 _2325_ (.A2(_1396_),
    .A1(_1395_),
    .B1(_1397_),
    .X(_1398_));
 sg13g2_o21ai_1 _2326_ (.B1(_1398_),
    .Y(_1399_),
    .A1(_1393_),
    .A2(_1394_));
 sg13g2_inv_1 _2327_ (.Y(_1400_),
    .A(_1399_));
 sg13g2_nor2b_2 _2328_ (.A(\cpu_instance.ctrl_instance.reg_sel_2[1] ),
    .B_N(\cpu_instance.ctrl_instance.reg_sel_2[0] ),
    .Y(_1401_));
 sg13g2_nand2_1 _2329_ (.Y(_1402_),
    .A(\cpu_instance.ctrl_instance.reg_sel_2[0] ),
    .B(\cpu_instance.ctrl_instance.reg_sel_2[1] ));
 sg13g2_inv_1 _2330_ (.Y(_1403_),
    .A(_1402_));
 sg13g2_nor2_1 _2331_ (.A(\cpu_instance.ctrl_instance.reg_sel_2[0] ),
    .B(\cpu_instance.ctrl_instance.reg_sel_2[1] ),
    .Y(_1404_));
 sg13g2_nor2_2 _2332_ (.A(\cpu_instance.ctrl_instance.reg_sel_2[0] ),
    .B(_1297_),
    .Y(_1405_));
 sg13g2_a21oi_1 _2333_ (.A1(uo_out[5]),
    .A2(_1403_),
    .Y(_1406_),
    .B1(net714));
 sg13g2_a22oi_1 _2334_ (.Y(_1407_),
    .B1(_1405_),
    .B2(\cpu_instance.registers_instance.registers[2][5] ),
    .A2(_1401_),
    .A1(\cpu_instance.registers_instance.registers[1][5] ));
 sg13g2_a22oi_1 _2335_ (.Y(_1408_),
    .B1(_1406_),
    .B2(_1407_),
    .A2(net714),
    .A1(_0038_));
 sg13g2_inv_1 _2336_ (.Y(_1409_),
    .A(_1408_));
 sg13g2_nand2_1 _2337_ (.Y(_1410_),
    .A(_1400_),
    .B(_1408_));
 sg13g2_nor2_1 _2338_ (.A(_1400_),
    .B(_1408_),
    .Y(_1411_));
 sg13g2_xnor2_1 _2339_ (.Y(_1412_),
    .A(_1399_),
    .B(_1409_));
 sg13g2_a22oi_1 _2340_ (.Y(_1413_),
    .B1(_1379_),
    .B2(\cpu_instance.registers_instance.register_bank[15][4] ),
    .A2(_1372_),
    .A1(\cpu_instance.registers_instance.register_bank[10][4] ));
 sg13g2_nand2_1 _2341_ (.Y(_1414_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[20] ),
    .B(_1375_));
 sg13g2_a22oi_1 _2342_ (.Y(_1415_),
    .B1(_1382_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[60] ),
    .A2(_1362_),
    .A1(\cpu_instance.registers_instance.register_bank[14][4] ));
 sg13g2_a22oi_1 _2343_ (.Y(_1416_),
    .B1(_1374_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[12] ),
    .A2(_1359_),
    .A1(\cpu_instance.registers_instance.register_bank[9][4] ));
 sg13g2_a22oi_1 _2344_ (.Y(_1417_),
    .B1(_1373_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[44] ),
    .A2(_1355_),
    .A1(\cpu_instance.registers_instance.register_bank[8][4] ));
 sg13g2_a22oi_1 _2345_ (.Y(_1418_),
    .B1(_1376_),
    .B2(\cpu_instance.registers_instance.register_bank[13][4] ),
    .A2(_1356_),
    .A1(\cpu_instance.registers_instance.register_bank[12][4] ));
 sg13g2_a22oi_1 _2346_ (.Y(_1419_),
    .B1(_1383_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[36] ),
    .A2(_1380_),
    .A1(\cpu_instance.registers_instance.register_bank[11][4] ));
 sg13g2_o21ai_1 _2347_ (.B1(net725),
    .Y(_1420_),
    .A1(_0041_),
    .A2(_1370_));
 sg13g2_a22oi_1 _2348_ (.Y(_1421_),
    .B1(_1381_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[28] ),
    .A2(_1378_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[52] ));
 sg13g2_nand4_1 _2349_ (.B(_1418_),
    .C(_1419_),
    .A(_1417_),
    .Y(_1422_),
    .D(_1421_));
 sg13g2_nand4_1 _2350_ (.B(_1414_),
    .C(_1415_),
    .A(_1413_),
    .Y(_1423_),
    .D(_1416_));
 sg13g2_nor3_2 _2351_ (.A(_1420_),
    .B(_1422_),
    .C(_1423_),
    .Y(_1424_));
 sg13g2_mux4_1 _2352_ (.S0(net733),
    .A0(_1277_),
    .A1(_0040_),
    .A2(_0039_),
    .A3(_1279_),
    .S1(net716),
    .X(_1425_));
 sg13g2_a21oi_2 _2353_ (.B1(_1424_),
    .Y(_1426_),
    .A2(_1425_),
    .A1(_1285_));
 sg13g2_inv_1 _2354_ (.Y(_1427_),
    .A(_1426_));
 sg13g2_mux4_1 _2355_ (.S0(\cpu_instance.ctrl_instance.reg_sel_2[0] ),
    .A0(_1277_),
    .A1(_0040_),
    .A2(_0039_),
    .A3(_1279_),
    .S1(_1297_),
    .X(_1428_));
 sg13g2_nor2_1 _2356_ (.A(_1427_),
    .B(_1428_),
    .Y(_1429_));
 sg13g2_xnor2_1 _2357_ (.Y(_1430_),
    .A(_1426_),
    .B(_1428_));
 sg13g2_inv_1 _2358_ (.Y(_1431_),
    .A(_1430_));
 sg13g2_nand2_1 _2359_ (.Y(_1432_),
    .A(\cpu_instance.registers_instance.register_bank[12][3] ),
    .B(_1356_));
 sg13g2_a22oi_1 _2360_ (.Y(_1433_),
    .B1(_1380_),
    .B2(\cpu_instance.registers_instance.register_bank[11][3] ),
    .A2(_1374_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[11] ));
 sg13g2_a22oi_1 _2361_ (.Y(_1434_),
    .B1(_1382_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[59] ),
    .A2(_1376_),
    .A1(\cpu_instance.registers_instance.register_bank[13][3] ));
 sg13g2_a22oi_1 _2362_ (.Y(_1435_),
    .B1(_1375_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[19] ),
    .A2(_1362_),
    .A1(\cpu_instance.registers_instance.register_bank[14][3] ));
 sg13g2_a22oi_1 _2363_ (.Y(_1436_),
    .B1(_1381_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[27] ),
    .A2(_1378_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[51] ));
 sg13g2_a22oi_1 _2364_ (.Y(_1437_),
    .B1(_1379_),
    .B2(\cpu_instance.registers_instance.register_bank[15][3] ),
    .A2(_1359_),
    .A1(\cpu_instance.registers_instance.register_bank[9][3] ));
 sg13g2_nand4_1 _2365_ (.B(_1435_),
    .C(_1436_),
    .A(_1432_),
    .Y(_1438_),
    .D(_1437_));
 sg13g2_a22oi_1 _2366_ (.Y(_1439_),
    .B1(_1383_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[35] ),
    .A2(_1373_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[43] ));
 sg13g2_o21ai_1 _2367_ (.B1(net725),
    .Y(_1440_),
    .A1(_0042_),
    .A2(_1370_));
 sg13g2_a22oi_1 _2368_ (.Y(_1441_),
    .B1(_1372_),
    .B2(\cpu_instance.registers_instance.register_bank[10][3] ),
    .A2(_1355_),
    .A1(\cpu_instance.registers_instance.register_bank[8][3] ));
 sg13g2_nand4_1 _2369_ (.B(_1434_),
    .C(_1439_),
    .A(_1433_),
    .Y(_1442_),
    .D(_1441_));
 sg13g2_nor3_2 _2370_ (.A(_1438_),
    .B(_1440_),
    .C(_1442_),
    .Y(_1443_));
 sg13g2_a21oi_2 _2371_ (.B1(_1443_),
    .Y(_1444_),
    .A2(_1343_),
    .A1(_1285_));
 sg13g2_a21oi_1 _2372_ (.A1(_1295_),
    .A2(_1403_),
    .Y(_1445_),
    .B1(net714));
 sg13g2_a22oi_1 _2373_ (.Y(_1446_),
    .B1(_1405_),
    .B2(\cpu_instance.registers_instance.registers[2][3] ),
    .A2(_1401_),
    .A1(\cpu_instance.registers_instance.registers[1][3] ));
 sg13g2_a22oi_1 _2374_ (.Y(_1447_),
    .B1(_1445_),
    .B2(_1446_),
    .A2(net714),
    .A1(_0035_));
 sg13g2_nor2b_1 _2375_ (.A(_1447_),
    .B_N(_1444_),
    .Y(_1448_));
 sg13g2_nor2b_1 _2376_ (.A(_1444_),
    .B_N(_1447_),
    .Y(_1449_));
 sg13g2_nor2_1 _2377_ (.A(net725),
    .B(_1336_),
    .Y(_1450_));
 sg13g2_nand2_1 _2378_ (.Y(_1451_),
    .A(\cpu_instance.registers_instance.register_bank[14][2] ),
    .B(_1362_));
 sg13g2_a22oi_1 _2379_ (.Y(_1452_),
    .B1(_1381_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[26] ),
    .A2(_1374_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[10] ));
 sg13g2_a22oi_1 _2380_ (.Y(_1453_),
    .B1(_1380_),
    .B2(\cpu_instance.registers_instance.register_bank[11][2] ),
    .A2(_1356_),
    .A1(\cpu_instance.registers_instance.register_bank[12][2] ));
 sg13g2_a22oi_1 _2381_ (.Y(_1454_),
    .B1(_1379_),
    .B2(\cpu_instance.registers_instance.register_bank[15][2] ),
    .A2(_1375_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[18] ));
 sg13g2_a22oi_1 _2382_ (.Y(_1455_),
    .B1(_1383_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[34] ),
    .A2(_1373_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[42] ));
 sg13g2_a22oi_1 _2383_ (.Y(_1456_),
    .B1(_1376_),
    .B2(\cpu_instance.registers_instance.register_bank[13][2] ),
    .A2(_1355_),
    .A1(\cpu_instance.registers_instance.register_bank[8][2] ));
 sg13g2_nand4_1 _2384_ (.B(_1454_),
    .C(_1455_),
    .A(_1451_),
    .Y(_1457_),
    .D(_1456_));
 sg13g2_a22oi_1 _2385_ (.Y(_1458_),
    .B1(_1382_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[58] ),
    .A2(_1359_),
    .A1(\cpu_instance.registers_instance.register_bank[9][2] ));
 sg13g2_o21ai_1 _2386_ (.B1(net725),
    .Y(_1459_),
    .A1(_0043_),
    .A2(_1370_));
 sg13g2_a22oi_1 _2387_ (.Y(_1460_),
    .B1(_1378_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[50] ),
    .A2(_1372_),
    .A1(\cpu_instance.registers_instance.register_bank[10][2] ));
 sg13g2_nand4_1 _2388_ (.B(_1453_),
    .C(_1458_),
    .A(_1452_),
    .Y(_1461_),
    .D(_1460_));
 sg13g2_nor3_2 _2389_ (.A(_1457_),
    .B(_1459_),
    .C(_1461_),
    .Y(_1462_));
 sg13g2_nor2_2 _2390_ (.A(_1450_),
    .B(_1462_),
    .Y(_1463_));
 sg13g2_a21oi_1 _2391_ (.A1(_1278_),
    .A2(\cpu_instance.ctrl_instance.reg_sel_2[1] ),
    .Y(_1464_),
    .B1(\cpu_instance.ctrl_instance.reg_sel_2[0] ));
 sg13g2_a221oi_1 _2392_ (.B2(uo_out[2]),
    .C1(_1464_),
    .B1(_1403_),
    .A1(\cpu_instance.registers_instance.registers[1][2] ),
    .Y(_1465_),
    .A2(_1297_));
 sg13g2_a21oi_2 _2393_ (.B1(_1465_),
    .Y(_1466_),
    .A2(_1404_),
    .A1(_0044_));
 sg13g2_nor3_2 _2394_ (.A(_1450_),
    .B(_1462_),
    .C(_1466_),
    .Y(_1467_));
 sg13g2_and2_1 _2395_ (.A(_1463_),
    .B(_1466_),
    .X(_1468_));
 sg13g2_xor2_1 _2396_ (.B(_1466_),
    .A(_1463_),
    .X(_1469_));
 sg13g2_and2_1 _2397_ (.A(_1285_),
    .B(net704),
    .X(_1470_));
 sg13g2_nand2_1 _2398_ (.Y(_1471_),
    .A(_1285_),
    .B(_1361_));
 sg13g2_a22oi_1 _2399_ (.Y(_1472_),
    .B1(_1375_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[17] ),
    .A2(_1356_),
    .A1(\cpu_instance.registers_instance.register_bank[12][1] ));
 sg13g2_nand2_1 _2400_ (.Y(_1473_),
    .A(\cpu_instance.registers_instance.register_bank[8][1] ),
    .B(_1355_));
 sg13g2_a22oi_1 _2401_ (.Y(_1474_),
    .B1(_1379_),
    .B2(\cpu_instance.registers_instance.register_bank[15][1] ),
    .A2(_1378_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[49] ));
 sg13g2_a22oi_1 _2402_ (.Y(_1475_),
    .B1(_1383_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[33] ),
    .A2(_1382_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[57] ));
 sg13g2_a22oi_1 _2403_ (.Y(_1476_),
    .B1(_1374_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[9] ),
    .A2(_1362_),
    .A1(\cpu_instance.registers_instance.register_bank[14][1] ));
 sg13g2_a22oi_1 _2404_ (.Y(_1477_),
    .B1(_1381_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[25] ),
    .A2(_1373_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[41] ));
 sg13g2_nand4_1 _2405_ (.B(_1475_),
    .C(_1476_),
    .A(_1474_),
    .Y(_1478_),
    .D(_1477_));
 sg13g2_a22oi_1 _2406_ (.Y(_1479_),
    .B1(_1372_),
    .B2(\cpu_instance.registers_instance.register_bank[10][1] ),
    .A2(_1359_),
    .A1(\cpu_instance.registers_instance.register_bank[9][1] ));
 sg13g2_a22oi_1 _2407_ (.Y(_1480_),
    .B1(_1380_),
    .B2(\cpu_instance.registers_instance.register_bank[11][1] ),
    .A2(_1376_),
    .A1(\cpu_instance.registers_instance.register_bank[13][1] ));
 sg13g2_nand4_1 _2408_ (.B(_1473_),
    .C(_1479_),
    .A(_1472_),
    .Y(_1481_),
    .D(_1480_));
 sg13g2_o21ai_1 _2409_ (.B1(net725),
    .Y(_1482_),
    .A1(_0045_),
    .A2(_1370_));
 sg13g2_nor3_2 _2410_ (.A(_1478_),
    .B(_1481_),
    .C(_1482_),
    .Y(_1483_));
 sg13g2_or3_1 _2411_ (.A(_1478_),
    .B(_1481_),
    .C(_1482_),
    .X(_1484_));
 sg13g2_nor2_2 _2412_ (.A(_1470_),
    .B(_1483_),
    .Y(_1485_));
 sg13g2_nand2_1 _2413_ (.Y(_1486_),
    .A(_0033_),
    .B(net714));
 sg13g2_a221oi_1 _2414_ (.B2(\cpu_instance.registers_instance.registers[2][1] ),
    .C1(net714),
    .B1(_1405_),
    .A1(\cpu_instance.registers_instance.registers[1][1] ),
    .Y(_1487_),
    .A2(_1297_));
 sg13g2_o21ai_1 _2415_ (.B1(_1487_),
    .Y(_1488_),
    .A1(_0034_),
    .A2(_1402_));
 sg13g2_nand2_2 _2416_ (.Y(_1489_),
    .A(_1486_),
    .B(_1488_));
 sg13g2_inv_1 _2417_ (.Y(_1490_),
    .A(_1489_));
 sg13g2_nor3_2 _2418_ (.A(_1470_),
    .B(_1483_),
    .C(_1489_),
    .Y(_1491_));
 sg13g2_nand3_1 _2419_ (.B(_1484_),
    .C(_1490_),
    .A(_1471_),
    .Y(_1492_));
 sg13g2_a21oi_2 _2420_ (.B1(_1490_),
    .Y(_1493_),
    .A2(_1484_),
    .A1(_1471_));
 sg13g2_o21ai_1 _2421_ (.B1(_1489_),
    .Y(_1494_),
    .A1(_1470_),
    .A2(_1483_));
 sg13g2_a22oi_1 _2422_ (.Y(_1495_),
    .B1(_1375_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[16] ),
    .A2(_1356_),
    .A1(\cpu_instance.registers_instance.register_bank[12][0] ));
 sg13g2_a22oi_1 _2423_ (.Y(_1496_),
    .B1(_1378_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[48] ),
    .A2(_1376_),
    .A1(\cpu_instance.registers_instance.register_bank[13][0] ));
 sg13g2_a22oi_1 _2424_ (.Y(_1497_),
    .B1(_1374_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[8] ),
    .A2(_1362_),
    .A1(\cpu_instance.registers_instance.register_bank[14][0] ));
 sg13g2_a22oi_1 _2425_ (.Y(_1498_),
    .B1(_1372_),
    .B2(\cpu_instance.registers_instance.register_bank[10][0] ),
    .A2(_1355_),
    .A1(\cpu_instance.registers_instance.register_bank[8][0] ));
 sg13g2_a22oi_1 _2426_ (.Y(_1499_),
    .B1(_1381_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[24] ),
    .A2(_1380_),
    .A1(\cpu_instance.registers_instance.register_bank[11][0] ));
 sg13g2_a22oi_1 _2427_ (.Y(_1500_),
    .B1(_1379_),
    .B2(\cpu_instance.registers_instance.register_bank[15][0] ),
    .A2(_1373_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[40] ));
 sg13g2_a221oi_1 _2428_ (.B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[56] ),
    .C1(_1369_),
    .B1(_1382_),
    .A1(_1363_),
    .Y(_1501_),
    .A2(_1364_));
 sg13g2_a22oi_1 _2429_ (.Y(_1502_),
    .B1(_1383_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[32] ),
    .A2(_1359_),
    .A1(\cpu_instance.registers_instance.register_bank[9][0] ));
 sg13g2_nand4_1 _2430_ (.B(_1497_),
    .C(_1499_),
    .A(_1495_),
    .Y(_1503_),
    .D(_1501_));
 sg13g2_nand4_1 _2431_ (.B(_1498_),
    .C(_1500_),
    .A(_1496_),
    .Y(_1504_),
    .D(_1502_));
 sg13g2_a21oi_1 _2432_ (.A1(_0046_),
    .A2(_1371_),
    .Y(_1505_),
    .B1(_1285_));
 sg13g2_o21ai_1 _2433_ (.B1(_1505_),
    .Y(_1506_),
    .A1(_1503_),
    .A2(_1504_));
 sg13g2_or2_2 _2434_ (.X(_1507_),
    .B(_1358_),
    .A(net725));
 sg13g2_and2_1 _2435_ (.A(_1506_),
    .B(_1507_),
    .X(_1508_));
 sg13g2_nand2_2 _2436_ (.Y(_1509_),
    .A(_1506_),
    .B(_1507_));
 sg13g2_a21oi_1 _2437_ (.A1(_1292_),
    .A2(_1403_),
    .Y(_1510_),
    .B1(net714));
 sg13g2_a22oi_1 _2438_ (.Y(_1511_),
    .B1(_1405_),
    .B2(\cpu_instance.registers_instance.registers[2][0] ),
    .A2(_1401_),
    .A1(\cpu_instance.registers_instance.registers[1][0] ));
 sg13g2_a22oi_1 _2439_ (.Y(_1512_),
    .B1(_1510_),
    .B2(_1511_),
    .A2(net714),
    .A1(_0031_));
 sg13g2_inv_1 _2440_ (.Y(_1513_),
    .A(_1512_));
 sg13g2_nand3_1 _2441_ (.B(_1507_),
    .C(_1512_),
    .A(_1506_),
    .Y(_1514_));
 sg13g2_o21ai_1 _2442_ (.B1(_1514_),
    .Y(_1515_),
    .A1(_1491_),
    .A2(_1493_));
 sg13g2_nand2_1 _2443_ (.Y(_1516_),
    .A(_1485_),
    .B(_1489_));
 sg13g2_a21oi_2 _2444_ (.B1(_1469_),
    .Y(_1517_),
    .A2(_1516_),
    .A1(_1515_));
 sg13g2_nor3_1 _2445_ (.A(_1448_),
    .B(_1467_),
    .C(_1517_),
    .Y(_1518_));
 sg13g2_nor3_2 _2446_ (.A(_1430_),
    .B(_1449_),
    .C(_1518_),
    .Y(_1519_));
 sg13g2_and2_1 _2447_ (.A(_1426_),
    .B(_1428_),
    .X(_1520_));
 sg13g2_nor2_1 _2448_ (.A(_1519_),
    .B(_1520_),
    .Y(_1521_));
 sg13g2_xor2_1 _2449_ (.B(_1521_),
    .A(_1412_),
    .X(_1522_));
 sg13g2_nor2b_1 _2450_ (.A(\cpu_instance.alu_instance.op[1] ),
    .B_N(\cpu_instance.alu_instance.op[0] ),
    .Y(_1523_));
 sg13g2_nand2b_2 _2451_ (.Y(_1524_),
    .B(\cpu_instance.alu_instance.op[0] ),
    .A_N(\cpu_instance.alu_instance.op[1] ));
 sg13g2_nand2b_2 _2452_ (.Y(_1525_),
    .B(\cpu_instance.alu_instance.op[3] ),
    .A_N(\cpu_instance.alu_instance.op[2] ));
 sg13g2_nor2_2 _2453_ (.A(_1524_),
    .B(_1525_),
    .Y(_1526_));
 sg13g2_nor2_1 _2454_ (.A(\cpu_instance.alu_instance.op[1] ),
    .B(\cpu_instance.alu_instance.op[0] ),
    .Y(_1527_));
 sg13g2_nor3_2 _2455_ (.A(\cpu_instance.alu_instance.op[2] ),
    .B(\cpu_instance.alu_instance.op[1] ),
    .C(\cpu_instance.alu_instance.op[0] ),
    .Y(_1528_));
 sg13g2_and2_2 _2456_ (.A(\cpu_instance.alu_instance.op[3] ),
    .B(_1528_),
    .X(_1529_));
 sg13g2_inv_1 _2457_ (.Y(_1530_),
    .A(_1529_));
 sg13g2_nor2_1 _2458_ (.A(_1400_),
    .B(_1409_),
    .Y(_1531_));
 sg13g2_inv_1 _2459_ (.Y(_1532_),
    .A(_1531_));
 sg13g2_nor2b_1 _2460_ (.A(\cpu_instance.alu_instance.op[3] ),
    .B_N(\cpu_instance.alu_instance.op[2] ),
    .Y(_1533_));
 sg13g2_nand2_2 _2461_ (.Y(_1534_),
    .A(_1286_),
    .B(\cpu_instance.alu_instance.op[2] ));
 sg13g2_nand2_1 _2462_ (.Y(_1535_),
    .A(\cpu_instance.alu_instance.op[1] ),
    .B(\cpu_instance.alu_instance.op[0] ));
 sg13g2_nor2_2 _2463_ (.A(_1534_),
    .B(_1535_),
    .Y(_1536_));
 sg13g2_nor2_2 _2464_ (.A(_1323_),
    .B(_1525_),
    .Y(_1537_));
 sg13g2_nor2_1 _2465_ (.A(_1524_),
    .B(_1534_),
    .Y(_1538_));
 sg13g2_a21oi_2 _2466_ (.B1(_1534_),
    .Y(_1539_),
    .A2(_1524_),
    .A1(_1323_));
 sg13g2_nand2_1 _2467_ (.Y(_1540_),
    .A(\cpu_instance.registers_instance.register_bank[12][6] ),
    .B(_1356_));
 sg13g2_a22oi_1 _2468_ (.Y(_1541_),
    .B1(_1382_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[62] ),
    .A2(_1375_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[22] ));
 sg13g2_a22oi_1 _2469_ (.Y(_1542_),
    .B1(_1381_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[30] ),
    .A2(_1378_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[54] ));
 sg13g2_a22oi_1 _2470_ (.Y(_1543_),
    .B1(_1383_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[38] ),
    .A2(_1379_),
    .A1(\cpu_instance.registers_instance.register_bank[15][6] ));
 sg13g2_a22oi_1 _2471_ (.Y(_1544_),
    .B1(_1374_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[14] ),
    .A2(_1373_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[46] ));
 sg13g2_nand4_1 _2472_ (.B(_1542_),
    .C(_1543_),
    .A(_1541_),
    .Y(_1545_),
    .D(_1544_));
 sg13g2_a22oi_1 _2473_ (.Y(_1546_),
    .B1(_1380_),
    .B2(\cpu_instance.registers_instance.register_bank[11][6] ),
    .A2(_1372_),
    .A1(\cpu_instance.registers_instance.register_bank[10][6] ));
 sg13g2_a22oi_1 _2474_ (.Y(_1547_),
    .B1(_1359_),
    .B2(\cpu_instance.registers_instance.register_bank[9][6] ),
    .A2(_1355_),
    .A1(\cpu_instance.registers_instance.register_bank[8][6] ));
 sg13g2_a22oi_1 _2475_ (.Y(_1548_),
    .B1(_1376_),
    .B2(\cpu_instance.registers_instance.register_bank[13][6] ),
    .A2(_1362_),
    .A1(\cpu_instance.registers_instance.register_bank[14][6] ));
 sg13g2_nand4_1 _2476_ (.B(_1546_),
    .C(_1547_),
    .A(_1540_),
    .Y(_1549_),
    .D(_1548_));
 sg13g2_nor3_2 _2477_ (.A(_1371_),
    .B(_1545_),
    .C(_1549_),
    .Y(_1550_));
 sg13g2_o21ai_1 _2478_ (.B1(\cpu_instance.ctrl_instance.use_register_bank_out_1 ),
    .Y(_1551_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[6] ),
    .A2(_1370_));
 sg13g2_o21ai_1 _2479_ (.B1(_1290_),
    .Y(_1552_),
    .A1(\cpu_instance.registers_instance.registers[2][6] ),
    .A2(net716));
 sg13g2_a22oi_1 _2480_ (.Y(_1553_),
    .B1(_1329_),
    .B2(uo_out[6]),
    .A2(_1328_),
    .A1(\cpu_instance.registers_instance.registers[1][6] ));
 sg13g2_o21ai_1 _2481_ (.B1(_1285_),
    .Y(_1554_),
    .A1(\cpu_instance.registers_instance.registers[0][6] ),
    .A2(_1332_));
 sg13g2_a21o_1 _2482_ (.A2(_1553_),
    .A1(_1552_),
    .B1(_1554_),
    .X(_1555_));
 sg13g2_o21ai_1 _2483_ (.B1(_1555_),
    .Y(_1556_),
    .A1(_1550_),
    .A2(_1551_));
 sg13g2_inv_1 _2484_ (.Y(_1557_),
    .A(_1556_));
 sg13g2_and2_1 _2485_ (.A(_1527_),
    .B(_1533_),
    .X(_1558_));
 sg13g2_nor3_1 _2486_ (.A(\cpu_instance.alu_instance.op[3] ),
    .B(\cpu_instance.alu_instance.op[2] ),
    .C(_1535_),
    .Y(_1559_));
 sg13g2_or2_2 _2487_ (.X(_1560_),
    .B(_1559_),
    .A(_1558_));
 sg13g2_a22oi_1 _2488_ (.Y(_1561_),
    .B1(_1539_),
    .B2(_1556_),
    .A2(_1528_),
    .A1(_1399_));
 sg13g2_a22oi_1 _2489_ (.Y(_1562_),
    .B1(_1560_),
    .B2(_1426_),
    .A2(_1537_),
    .A1(_1400_));
 sg13g2_nor2_1 _2490_ (.A(_1410_),
    .B(_1530_),
    .Y(_1563_));
 sg13g2_a221oi_1 _2491_ (.B2(_1536_),
    .C1(_1563_),
    .B1(_1531_),
    .A1(_1412_),
    .Y(_1564_),
    .A2(_1526_));
 sg13g2_or2_1 _2492_ (.X(_1565_),
    .B(_1447_),
    .A(_1444_));
 sg13g2_inv_1 _2493_ (.Y(_1566_),
    .A(_1565_));
 sg13g2_and2_1 _2494_ (.A(_1444_),
    .B(_1447_),
    .X(_1567_));
 sg13g2_a21oi_2 _2495_ (.B1(_1513_),
    .Y(_1568_),
    .A2(_1507_),
    .A1(_1506_));
 sg13g2_nand3_1 _2496_ (.B(_1494_),
    .C(_1568_),
    .A(_1492_),
    .Y(_1569_));
 sg13g2_a21o_1 _2497_ (.A2(_1568_),
    .A1(_1494_),
    .B1(_1491_),
    .X(_1570_));
 sg13g2_a21o_1 _2498_ (.A2(_1570_),
    .A1(_1469_),
    .B1(_1468_),
    .X(_1571_));
 sg13g2_a221oi_1 _2499_ (.B2(_1570_),
    .C1(_1468_),
    .B1(_1469_),
    .A1(_1444_),
    .Y(_1572_),
    .A2(_1447_));
 sg13g2_nor3_2 _2500_ (.A(_1431_),
    .B(_1566_),
    .C(_1572_),
    .Y(_1573_));
 sg13g2_o21ai_1 _2501_ (.B1(_1412_),
    .Y(_1574_),
    .A1(_1429_),
    .A2(_1573_));
 sg13g2_and2_2 _2502_ (.A(_1324_),
    .B(_1523_),
    .X(_1575_));
 sg13g2_nand2_2 _2503_ (.Y(_1576_),
    .A(_1324_),
    .B(_1523_));
 sg13g2_or3_1 _2504_ (.A(_1412_),
    .B(_1429_),
    .C(_1573_),
    .X(_1577_));
 sg13g2_nand3_1 _2505_ (.B(_1575_),
    .C(_1577_),
    .A(_1574_),
    .Y(_1578_));
 sg13g2_nand4_1 _2506_ (.B(_1562_),
    .C(_1564_),
    .A(_1561_),
    .Y(_1579_),
    .D(_1578_));
 sg13g2_a21o_1 _2507_ (.A2(_1522_),
    .A1(_1325_),
    .B1(_1579_),
    .X(_1580_));
 sg13g2_and2_1 _2508_ (.A(\cpu_instance.ctrl_instance.mux_sel[1] ),
    .B(net4),
    .X(_1581_));
 sg13g2_a221oi_1 _2509_ (.B2(_1580_),
    .C1(_1581_),
    .B1(\cpu_instance.ctrl_instance.mux_sel[0] ),
    .A1(\cpu_instance.mem_instance.bus_data_out[5] ),
    .Y(_1582_),
    .A2(\cpu_instance.ctrl_instance.mux_sel[2] ));
 sg13g2_inv_1 _2510_ (.Y(_1583_),
    .A(net608));
 sg13g2_o21ai_1 _2511_ (.B1(_1431_),
    .Y(_1584_),
    .A1(_1566_),
    .A2(_1572_));
 sg13g2_nor2_1 _2512_ (.A(_1573_),
    .B(_1576_),
    .Y(_1585_));
 sg13g2_nand2_1 _2513_ (.Y(_1586_),
    .A(_1430_),
    .B(_1526_));
 sg13g2_nand2_1 _2514_ (.Y(_1587_),
    .A(_1427_),
    .B(_1537_));
 sg13g2_a22oi_1 _2515_ (.Y(_1588_),
    .B1(_1560_),
    .B2(_1444_),
    .A2(_1539_),
    .A1(_1399_));
 sg13g2_o21ai_1 _2516_ (.B1(_1427_),
    .Y(_1589_),
    .A1(_1286_),
    .A2(_1428_));
 sg13g2_a22oi_1 _2517_ (.Y(_1590_),
    .B1(_1589_),
    .B2(_1528_),
    .A2(_1536_),
    .A1(_1429_));
 sg13g2_and2_1 _2518_ (.A(_1286_),
    .B(_1528_),
    .X(_1591_));
 sg13g2_nand4_1 _2519_ (.B(_1587_),
    .C(_1588_),
    .A(_1586_),
    .Y(_1592_),
    .D(_1590_));
 sg13g2_o21ai_1 _2520_ (.B1(_1430_),
    .Y(_1593_),
    .A1(_1449_),
    .A2(_1518_));
 sg13g2_nor2b_1 _2521_ (.A(_1519_),
    .B_N(_1593_),
    .Y(_1594_));
 sg13g2_a221oi_1 _2522_ (.B2(_1325_),
    .C1(_1592_),
    .B1(_1594_),
    .A1(_1584_),
    .Y(_1595_),
    .A2(_1585_));
 sg13g2_nor2_1 _2523_ (.A(_1300_),
    .B(_1595_),
    .Y(_1596_));
 sg13g2_a22oi_1 _2524_ (.Y(_1597_),
    .B1(net3),
    .B2(\cpu_instance.ctrl_instance.mux_sel[1] ),
    .A2(\cpu_instance.ctrl_instance.mux_sel[2] ),
    .A1(\cpu_instance.mem_instance.bus_data_out[4] ));
 sg13g2_nor2b_1 _2525_ (.A(_1596_),
    .B_N(_1597_),
    .Y(_1598_));
 sg13g2_o21ai_1 _2526_ (.B1(_1597_),
    .Y(_1599_),
    .A1(_1300_),
    .A2(_1595_));
 sg13g2_nor2_1 _2527_ (.A(_1583_),
    .B(_1599_),
    .Y(_1600_));
 sg13g2_nand2_2 _2528_ (.Y(_1601_),
    .A(net612),
    .B(_1598_));
 sg13g2_nand2_1 _2529_ (.Y(_1602_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[63] ),
    .B(_1382_));
 sg13g2_a22oi_1 _2530_ (.Y(_1603_),
    .B1(_1376_),
    .B2(\cpu_instance.registers_instance.register_bank[13][7] ),
    .A2(_1372_),
    .A1(\cpu_instance.registers_instance.register_bank[10][7] ));
 sg13g2_a22oi_1 _2531_ (.Y(_1604_),
    .B1(_1381_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[31] ),
    .A2(_1374_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[15] ));
 sg13g2_a22oi_1 _2532_ (.Y(_1605_),
    .B1(_1359_),
    .B2(\cpu_instance.registers_instance.register_bank[9][7] ),
    .A2(_1355_),
    .A1(\cpu_instance.registers_instance.register_bank[8][7] ));
 sg13g2_a22oi_1 _2533_ (.Y(_1606_),
    .B1(_1380_),
    .B2(\cpu_instance.registers_instance.register_bank[11][7] ),
    .A2(_1362_),
    .A1(\cpu_instance.registers_instance.register_bank[14][7] ));
 sg13g2_a22oi_1 _2534_ (.Y(_1607_),
    .B1(_1379_),
    .B2(\cpu_instance.registers_instance.register_bank[15][7] ),
    .A2(_1356_),
    .A1(\cpu_instance.registers_instance.register_bank[12][7] ));
 sg13g2_nand4_1 _2535_ (.B(_1605_),
    .C(_1606_),
    .A(_1603_),
    .Y(_1608_),
    .D(_1607_));
 sg13g2_a22oi_1 _2536_ (.Y(_1609_),
    .B1(_1383_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[39] ),
    .A2(_1375_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[23] ));
 sg13g2_a22oi_1 _2537_ (.Y(_1610_),
    .B1(_1378_),
    .B2(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[55] ),
    .A2(_1373_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[47] ));
 sg13g2_nand4_1 _2538_ (.B(_1604_),
    .C(_1609_),
    .A(_1602_),
    .Y(_1611_),
    .D(_1610_));
 sg13g2_nor3_2 _2539_ (.A(_1371_),
    .B(_1608_),
    .C(_1611_),
    .Y(_1612_));
 sg13g2_o21ai_1 _2540_ (.B1(net725),
    .Y(_1613_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[7] ),
    .A2(_1370_));
 sg13g2_o21ai_1 _2541_ (.B1(_1290_),
    .Y(_0337_),
    .A1(\cpu_instance.registers_instance.registers[2][7] ),
    .A2(net716));
 sg13g2_a22oi_1 _2542_ (.Y(_0338_),
    .B1(_1329_),
    .B2(uo_out[7]),
    .A2(_1328_),
    .A1(\cpu_instance.registers_instance.registers[1][7] ));
 sg13g2_a22oi_1 _2543_ (.Y(_0339_),
    .B1(_0337_),
    .B2(_0338_),
    .A2(_1331_),
    .A1(_1281_));
 sg13g2_nand2_1 _2544_ (.Y(_0340_),
    .A(_1285_),
    .B(_0339_));
 sg13g2_o21ai_1 _2545_ (.B1(_0340_),
    .Y(_0341_),
    .A1(_1612_),
    .A2(_1613_));
 sg13g2_mux4_1 _2546_ (.S0(_1297_),
    .A0(\cpu_instance.registers_instance.registers[2][7] ),
    .A1(_1301_),
    .A2(uo_out[7]),
    .A3(\cpu_instance.registers_instance.registers[1][7] ),
    .S1(\cpu_instance.ctrl_instance.reg_sel_2[0] ),
    .X(_0342_));
 sg13g2_inv_1 _2547_ (.Y(_0343_),
    .A(_0342_));
 sg13g2_nand2_1 _2548_ (.Y(_0344_),
    .A(_0341_),
    .B(_0343_));
 sg13g2_nand2_1 _2549_ (.Y(_0345_),
    .A(net629),
    .B(_0342_));
 sg13g2_xnor2_1 _2550_ (.Y(_0346_),
    .A(net629),
    .B(_0342_));
 sg13g2_inv_1 _2551_ (.Y(_0347_),
    .A(_0346_));
 sg13g2_mux4_1 _2552_ (.S0(_1297_),
    .A0(\cpu_instance.registers_instance.registers[2][6] ),
    .A1(_1298_),
    .A2(uo_out[6]),
    .A3(\cpu_instance.registers_instance.registers[1][6] ),
    .S1(\cpu_instance.ctrl_instance.reg_sel_2[0] ),
    .X(_0348_));
 sg13g2_nor2_1 _2553_ (.A(_1557_),
    .B(_0348_),
    .Y(_0349_));
 sg13g2_nand2_1 _2554_ (.Y(_0350_),
    .A(_1556_),
    .B(_0348_));
 sg13g2_inv_1 _2555_ (.Y(_0351_),
    .A(_0350_));
 sg13g2_xnor2_1 _2556_ (.Y(_0352_),
    .A(_1556_),
    .B(_0348_));
 sg13g2_or3_1 _2557_ (.A(_1411_),
    .B(_1519_),
    .C(_1520_),
    .X(_0353_));
 sg13g2_and3_1 _2558_ (.X(_0354_),
    .A(_1410_),
    .B(_0352_),
    .C(_0353_));
 sg13g2_or3_1 _2559_ (.A(_0346_),
    .B(_0349_),
    .C(_0354_),
    .X(_0355_));
 sg13g2_o21ai_1 _2560_ (.B1(_0346_),
    .Y(_0356_),
    .A1(_0349_),
    .A2(_0354_));
 sg13g2_and3_1 _2561_ (.X(_0357_),
    .A(_1325_),
    .B(_0355_),
    .C(_0356_));
 sg13g2_nand3_1 _2562_ (.B(_1509_),
    .C(_1533_),
    .A(_1322_),
    .Y(_0358_));
 sg13g2_nor3_1 _2563_ (.A(_1323_),
    .B(_1525_),
    .C(net629),
    .Y(_0359_));
 sg13g2_nand3_1 _2564_ (.B(net629),
    .C(_0342_),
    .A(_1536_),
    .Y(_0360_));
 sg13g2_a21o_1 _2565_ (.A2(_0342_),
    .A1(\cpu_instance.alu_instance.op[3] ),
    .B1(net629),
    .X(_0361_));
 sg13g2_a221oi_1 _2566_ (.B2(_1528_),
    .C1(_0359_),
    .B1(_0361_),
    .A1(_1556_),
    .Y(_0362_),
    .A2(_1560_));
 sg13g2_nand3_1 _2567_ (.B(_0360_),
    .C(_0362_),
    .A(_0358_),
    .Y(_0363_));
 sg13g2_a21oi_1 _2568_ (.A1(_1526_),
    .A2(_0347_),
    .Y(_0364_),
    .B1(_0363_));
 sg13g2_a21oi_1 _2569_ (.A1(_1532_),
    .A2(_1574_),
    .Y(_0365_),
    .B1(_0352_));
 sg13g2_nor3_1 _2570_ (.A(_0347_),
    .B(_0351_),
    .C(_0365_),
    .Y(_0366_));
 sg13g2_o21ai_1 _2571_ (.B1(_0347_),
    .Y(_0367_),
    .A1(_0351_),
    .A2(_0365_));
 sg13g2_nand2_1 _2572_ (.Y(_0368_),
    .A(_1575_),
    .B(_0367_));
 sg13g2_o21ai_1 _2573_ (.B1(_0364_),
    .Y(_0369_),
    .A1(_0366_),
    .A2(_0368_));
 sg13g2_o21ai_1 _2574_ (.B1(\cpu_instance.ctrl_instance.mux_sel[0] ),
    .Y(_0370_),
    .A1(_0357_),
    .A2(_0369_));
 sg13g2_a22oi_1 _2575_ (.Y(_0371_),
    .B1(net6),
    .B2(\cpu_instance.ctrl_instance.mux_sel[1] ),
    .A2(\cpu_instance.ctrl_instance.mux_sel[2] ),
    .A1(net429));
 sg13g2_and2_1 _2576_ (.A(_0370_),
    .B(_0371_),
    .X(_0372_));
 sg13g2_nand2_1 _2577_ (.Y(_0373_),
    .A(_0370_),
    .B(_0371_));
 sg13g2_a21oi_1 _2578_ (.A1(_1410_),
    .A2(_0353_),
    .Y(_0374_),
    .B1(_0352_));
 sg13g2_nor3_1 _2579_ (.A(_1326_),
    .B(_0354_),
    .C(_0374_),
    .Y(_0375_));
 sg13g2_and3_1 _2580_ (.X(_0376_),
    .A(_1532_),
    .B(_1574_),
    .C(_0352_));
 sg13g2_nor3_1 _2581_ (.A(_1576_),
    .B(_0365_),
    .C(_0376_),
    .Y(_0377_));
 sg13g2_nand2b_1 _2582_ (.Y(_0378_),
    .B(_1526_),
    .A_N(_0352_));
 sg13g2_a22oi_1 _2583_ (.Y(_0379_),
    .B1(_1560_),
    .B2(_1399_),
    .A2(_1557_),
    .A1(_1537_));
 sg13g2_a22oi_1 _2584_ (.Y(_0380_),
    .B1(_0348_),
    .B2(_1529_),
    .A2(net629),
    .A1(_1539_));
 sg13g2_a22oi_1 _2585_ (.Y(_0381_),
    .B1(_0351_),
    .B2(_1536_),
    .A2(_1556_),
    .A1(_1528_));
 sg13g2_nand4_1 _2586_ (.B(_0379_),
    .C(_0380_),
    .A(_0378_),
    .Y(_0382_),
    .D(_0381_));
 sg13g2_or3_2 _2587_ (.A(_0375_),
    .B(_0377_),
    .C(_0382_),
    .X(_0383_));
 sg13g2_and2_1 _2588_ (.A(\cpu_instance.mem_instance.bus_data_out[6] ),
    .B(\cpu_instance.ctrl_instance.mux_sel[2] ),
    .X(_0384_));
 sg13g2_a221oi_1 _2589_ (.B2(_0383_),
    .C1(_0384_),
    .B1(\cpu_instance.ctrl_instance.mux_sel[0] ),
    .A1(net5),
    .Y(_0385_),
    .A2(\cpu_instance.ctrl_instance.mux_sel[1] ));
 sg13g2_inv_4 _2590_ (.A(net599),
    .Y(_0386_));
 sg13g2_nor2_2 _2591_ (.A(net595),
    .B(_0386_),
    .Y(_0387_));
 sg13g2_and2_1 _2592_ (.A(net717),
    .B(net775),
    .X(_0388_));
 sg13g2_nand2_1 _2593_ (.Y(_0389_),
    .A(net717),
    .B(net773));
 sg13g2_nand3_1 _2594_ (.B(_0387_),
    .C(_0388_),
    .A(net570),
    .Y(_0390_));
 sg13g2_or2_1 _2595_ (.X(_0391_),
    .B(_0390_),
    .A(_1601_));
 sg13g2_nor2_1 _2596_ (.A(net719),
    .B(\cpu_instance.ctrl_instance.state[5] ),
    .Y(_0392_));
 sg13g2_nand2b_1 _2597_ (.Y(_0393_),
    .B(_0392_),
    .A_N(\cpu_instance.ctrl_instance.state[7] ));
 sg13g2_or3_1 _2598_ (.A(net847),
    .B(net715),
    .C(_0393_),
    .X(_0394_));
 sg13g2_nand2_1 _2599_ (.Y(_0395_),
    .A(net832),
    .B(net717));
 sg13g2_a21oi_2 _2600_ (.B1(net741),
    .Y(_0396_),
    .A2(net717),
    .A1(net838));
 sg13g2_nand4_1 _2601_ (.B(_0394_),
    .C(_0395_),
    .A(_0391_),
    .Y(_0003_),
    .D(_0396_));
 sg13g2_o21ai_1 _2602_ (.B1(_0391_),
    .Y(_0001_),
    .A1(net741),
    .A2(_1304_));
 sg13g2_nand2b_1 _2603_ (.Y(_0397_),
    .B(_1601_),
    .A_N(_0390_));
 sg13g2_nor2b_2 _2604_ (.A(net583),
    .B_N(net822),
    .Y(_0398_));
 sg13g2_inv_1 _2605_ (.Y(_0399_),
    .A(_0398_));
 sg13g2_nand2_2 _2606_ (.Y(_0400_),
    .A(net770),
    .B(_0398_));
 sg13g2_or2_1 _2607_ (.X(_0401_),
    .B(_0400_),
    .A(_0387_));
 sg13g2_nand2b_1 _2608_ (.Y(_0402_),
    .B(_1304_),
    .A_N(_0394_));
 sg13g2_nand4_1 _2609_ (.B(_0397_),
    .C(_0401_),
    .A(_0396_),
    .Y(_0000_),
    .D(_0402_));
 sg13g2_nand2_1 _2610_ (.Y(_0403_),
    .A(net596),
    .B(_0386_));
 sg13g2_or2_1 _2611_ (.X(_0404_),
    .B(_0400_),
    .A(net600));
 sg13g2_nand2b_1 _2612_ (.Y(_0405_),
    .B(_1318_),
    .A_N(net717));
 sg13g2_o21ai_1 _2613_ (.B1(_0405_),
    .Y(_0009_),
    .A1(_0373_),
    .A2(_0404_));
 sg13g2_nand2_1 _2614_ (.Y(_0406_),
    .A(net395),
    .B(_1319_));
 sg13g2_nand3_1 _2615_ (.B(_0387_),
    .C(_0398_),
    .A(net769),
    .Y(_0407_));
 sg13g2_nand2_1 _2616_ (.Y(_0408_),
    .A(_1600_),
    .B(_0387_));
 sg13g2_o21ai_1 _2617_ (.B1(_0406_),
    .Y(_0010_),
    .A1(_1601_),
    .A2(_0407_));
 sg13g2_a22oi_1 _2618_ (.Y(_0409_),
    .B1(_1319_),
    .B2(\cpu_instance.ctrl_instance.state[5] ),
    .A2(net505),
    .A1(net769));
 sg13g2_inv_1 _2619_ (.Y(_0011_),
    .A(net506));
 sg13g2_nor3_1 _2620_ (.A(net611),
    .B(net616),
    .C(_0407_),
    .Y(_0410_));
 sg13g2_a21o_1 _2621_ (.A2(_1319_),
    .A1(net356),
    .B1(_0410_),
    .X(_0012_));
 sg13g2_xnor2_1 _2622_ (.Y(_0411_),
    .A(\cpu_instance.ctrl_instance.flag_zero ),
    .B(net616));
 sg13g2_a21oi_1 _2623_ (.A1(\cpu_instance.ctrl_instance.flag_carry ),
    .A2(net602),
    .Y(_0412_),
    .B1(_0411_));
 sg13g2_o21ai_1 _2624_ (.B1(_0412_),
    .Y(_0413_),
    .A1(\cpu_instance.ctrl_instance.flag_carry ),
    .A2(net602));
 sg13g2_nand3_1 _2625_ (.B(_0386_),
    .C(_0413_),
    .A(net591),
    .Y(_0414_));
 sg13g2_nand2_1 _2626_ (.Y(_0415_),
    .A(net585),
    .B(_1319_));
 sg13g2_o21ai_1 _2627_ (.B1(_0415_),
    .Y(_0013_),
    .A1(_0400_),
    .A2(_0414_));
 sg13g2_nor2_2 _2628_ (.A(\cpu_instance.ctrl_instance.mem_ctrl_op[0] ),
    .B(net798),
    .Y(_0416_));
 sg13g2_or2_1 _2629_ (.X(_0417_),
    .B(net798),
    .A(\cpu_instance.ctrl_instance.mem_ctrl_op[0] ));
 sg13g2_nor2b_1 _2630_ (.A(net827),
    .B_N(\cpu_instance.mem_instance.mem_ctrl_instance.state[2] ),
    .Y(_0418_));
 sg13g2_o21ai_1 _2631_ (.B1(_0417_),
    .Y(_0419_),
    .A1(net819),
    .A2(_0418_));
 sg13g2_nor3_2 _2632_ (.A(\cpu_instance.ctrl_instance.mem_ctrl_op[0] ),
    .B(net816),
    .C(\cpu_instance.ctrl_instance.mem_ctrl_op[2] ),
    .Y(_0420_));
 sg13g2_nand2b_1 _2633_ (.Y(_0421_),
    .B(net557),
    .A_N(_0420_));
 sg13g2_nor2_1 _2634_ (.A(net798),
    .B(\cpu_instance.ctrl_instance.mem_ctrl_op[2] ),
    .Y(_0422_));
 sg13g2_a21oi_1 _2635_ (.A1(net369),
    .A2(_0422_),
    .Y(_0423_),
    .B1(net738));
 sg13g2_nand3_1 _2636_ (.B(net558),
    .C(_0423_),
    .A(_0419_),
    .Y(_0014_));
 sg13g2_a22oi_1 _2637_ (.Y(_0424_),
    .B1(net799),
    .B2(_0418_),
    .A2(net369),
    .A1(\cpu_instance.ctrl_instance.mem_ctrl_op[2] ));
 sg13g2_nor2_1 _2638_ (.A(net738),
    .B(net800),
    .Y(_0016_));
 sg13g2_nor2b_1 _2639_ (.A(\cpu_instance.ctrl_instance.mem_ctrl_op[2] ),
    .B_N(net798),
    .Y(_0425_));
 sg13g2_nand2_1 _2640_ (.Y(_0426_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.state[3] ),
    .B(_0420_));
 sg13g2_a22oi_1 _2641_ (.Y(_0427_),
    .B1(_0425_),
    .B2(net369),
    .A2(_0420_),
    .A1(net557));
 sg13g2_nor2_1 _2642_ (.A(net738),
    .B(_0427_),
    .Y(_0017_));
 sg13g2_a21oi_1 _2643_ (.A1(net800),
    .A2(_0427_),
    .Y(_0018_),
    .B1(net738));
 sg13g2_nand2_1 _2644_ (.Y(_0428_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.state[2] ),
    .B(net827));
 sg13g2_a22oi_1 _2645_ (.Y(_0429_),
    .B1(net799),
    .B2(net819),
    .A2(\cpu_instance.mem_instance.data_ready ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.state[2] ));
 sg13g2_nor2_1 _2646_ (.A(net738),
    .B(net820),
    .Y(_0015_));
 sg13g2_a21oi_1 _2647_ (.A1(_0427_),
    .A2(net820),
    .Y(_0019_),
    .B1(net738));
 sg13g2_nor3_1 _2648_ (.A(net602),
    .B(net605),
    .C(_0407_),
    .Y(_0430_));
 sg13g2_a21o_1 _2649_ (.A2(_1319_),
    .A1(net445),
    .B1(_0430_),
    .X(_0008_));
 sg13g2_nor2_2 _2650_ (.A(net591),
    .B(_0386_),
    .Y(_0431_));
 sg13g2_nand3_1 _2651_ (.B(_0371_),
    .C(net601),
    .A(_0370_),
    .Y(_0432_));
 sg13g2_nor3_1 _2652_ (.A(net595),
    .B(net600),
    .C(_0413_),
    .Y(_0433_));
 sg13g2_nor2_1 _2653_ (.A(_0431_),
    .B(_0433_),
    .Y(_0434_));
 sg13g2_nand2_2 _2654_ (.Y(_0435_),
    .A(net602),
    .B(_1599_));
 sg13g2_nor2_2 _2655_ (.A(net585),
    .B(net395),
    .Y(_0436_));
 sg13g2_nand2b_2 _2656_ (.Y(_0437_),
    .B(_0436_),
    .A_N(net719));
 sg13g2_o21ai_1 _2657_ (.B1(_0388_),
    .Y(_0438_),
    .A1(net715),
    .A2(_0437_));
 sg13g2_o21ai_1 _2658_ (.B1(_0438_),
    .Y(_0439_),
    .A1(_0390_),
    .A2(_0435_));
 sg13g2_inv_1 _2659_ (.Y(_0440_),
    .A(_0439_));
 sg13g2_o21ai_1 _2660_ (.B1(_0440_),
    .Y(_0007_),
    .A1(_0400_),
    .A2(_0434_));
 sg13g2_nand2b_1 _2661_ (.Y(_0006_),
    .B(net769),
    .A_N(net327));
 sg13g2_nor3_2 _2662_ (.A(net509),
    .B(_0389_),
    .C(_0432_),
    .Y(_0441_));
 sg13g2_a22oi_1 _2663_ (.Y(_0442_),
    .B1(_0441_),
    .B2(net611),
    .A2(_0393_),
    .A1(_1319_));
 sg13g2_nand4_1 _2664_ (.B(_0397_),
    .C(_0404_),
    .A(_1317_),
    .Y(_0005_),
    .D(_0442_));
 sg13g2_and2_1 _2665_ (.A(net602),
    .B(_0441_),
    .X(_0004_));
 sg13g2_and2_1 _2666_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_data_oe[0] ),
    .B(net772),
    .X(uio_oe[5]));
 sg13g2_nor2b_1 _2667_ (.A(net723),
    .B_N(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[0] ),
    .Y(_0443_));
 sg13g2_nand2_2 _2668_ (.Y(_0444_),
    .A(_0023_),
    .B(_0443_));
 sg13g2_and2_1 _2669_ (.A(net722),
    .B(net724),
    .X(_0445_));
 sg13g2_nor2b_2 _2670_ (.A(net723),
    .B_N(net712),
    .Y(_0446_));
 sg13g2_nand2b_1 _2671_ (.Y(_0447_),
    .B(net712),
    .A_N(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[1] ));
 sg13g2_nor2b_2 _2672_ (.A(net724),
    .B_N(net723),
    .Y(_0448_));
 sg13g2_nand2b_1 _2673_ (.Y(_0449_),
    .B(_0448_),
    .A_N(net722));
 sg13g2_nand3_1 _2674_ (.B(_0447_),
    .C(_0449_),
    .A(_0444_),
    .Y(_0450_));
 sg13g2_inv_1 _2675_ (.Y(_0451_),
    .A(_0450_));
 sg13g2_nor2_1 _2676_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[0] ),
    .B(_0444_),
    .Y(_0452_));
 sg13g2_nor3_1 _2677_ (.A(net720),
    .B(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[0] ),
    .C(_0444_),
    .Y(_0453_));
 sg13g2_nand2_1 _2678_ (.Y(_0454_),
    .A(net723),
    .B(_0023_));
 sg13g2_nor2_2 _2679_ (.A(net724),
    .B(_0454_),
    .Y(_0455_));
 sg13g2_nand2_1 _2680_ (.Y(_0456_),
    .A(_0023_),
    .B(_0448_));
 sg13g2_a221oi_1 _2681_ (.B2(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[20] ),
    .C1(_0453_),
    .B1(_0455_),
    .A1(\cpu_instance.mem_instance.data_qo_mi[4] ),
    .Y(_0457_),
    .A2(_0446_));
 sg13g2_nor2_2 _2682_ (.A(_0451_),
    .B(_0457_),
    .Y(uio_out[1]));
 sg13g2_a221oi_1 _2683_ (.B2(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[21] ),
    .C1(_0452_),
    .B1(_0455_),
    .A1(\cpu_instance.mem_instance.data_qo_mi[5] ),
    .Y(_0458_),
    .A2(_0446_));
 sg13g2_nand2_2 _2684_ (.Y(uio_out[2]),
    .A(_0450_),
    .B(_0458_));
 sg13g2_nand3_1 _2685_ (.B(_0450_),
    .C(_0455_),
    .A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[22] ),
    .Y(_0459_));
 sg13g2_o21ai_1 _2686_ (.B1(_0459_),
    .Y(uio_out[4]),
    .A1(_1315_),
    .A2(_0447_));
 sg13g2_nand2_1 _2687_ (.Y(_0460_),
    .A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[23] ),
    .B(_0455_));
 sg13g2_a21oi_1 _2688_ (.A1(\cpu_instance.mem_instance.data_qo_mi[7] ),
    .A2(_0446_),
    .Y(_0461_),
    .B1(_0453_));
 sg13g2_nand3_1 _2689_ (.B(_0460_),
    .C(_0461_),
    .A(_0450_),
    .Y(uio_out[5]));
 sg13g2_nor2_2 _2690_ (.A(net854),
    .B(\cpu_instance.mem_instance.mem_ctrl_instance.state[2] ),
    .Y(_0462_));
 sg13g2_o21ai_1 _2691_ (.B1(_0421_),
    .Y(_0463_),
    .A1(_0416_),
    .A2(_0462_));
 sg13g2_a21oi_1 _2692_ (.A1(net359),
    .A2(_0462_),
    .Y(_0464_),
    .B1(net738));
 sg13g2_and2_1 _2693_ (.A(_0463_),
    .B(_0464_),
    .X(_0047_));
 sg13g2_nand2_1 _2694_ (.Y(_0465_),
    .A(net600),
    .B(_0398_));
 sg13g2_nand4_1 _2695_ (.B(net595),
    .C(net600),
    .A(net602),
    .Y(_0466_),
    .D(_0398_));
 sg13g2_o21ai_1 _2696_ (.B1(net717),
    .Y(_0467_),
    .A1(net719),
    .A2(net715));
 sg13g2_a21oi_1 _2697_ (.A1(_0466_),
    .A2(_0467_),
    .Y(_0048_),
    .B1(net741));
 sg13g2_o21ai_1 _2698_ (.B1(_0387_),
    .Y(_0468_),
    .A1(net609),
    .A2(net616));
 sg13g2_nand3_1 _2699_ (.B(_0434_),
    .C(_0468_),
    .A(_0398_),
    .Y(_0469_));
 sg13g2_nor2_1 _2700_ (.A(net595),
    .B(_0395_),
    .Y(_0470_));
 sg13g2_nor2_1 _2701_ (.A(net327),
    .B(_0470_),
    .Y(_0471_));
 sg13g2_o21ai_1 _2702_ (.B1(net769),
    .Y(_0472_),
    .A1(net570),
    .A2(net327));
 sg13g2_a22oi_1 _2703_ (.Y(_0049_),
    .B1(_0472_),
    .B2(_1320_),
    .A2(_0471_),
    .A1(_0469_));
 sg13g2_nor3_1 _2704_ (.A(net583),
    .B(_1320_),
    .C(net600),
    .Y(_0050_));
 sg13g2_nor3_1 _2705_ (.A(net583),
    .B(_1320_),
    .C(net609),
    .Y(_0051_));
 sg13g2_o21ai_1 _2706_ (.B1(net320),
    .Y(_0473_),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_clk_out ),
    .A2(_1284_));
 sg13g2_nand2_1 _2707_ (.Y(_0474_),
    .A(net771),
    .B(_0473_));
 sg13g2_nor2_2 _2708_ (.A(net390),
    .B(_0474_),
    .Y(_0475_));
 sg13g2_or2_2 _2709_ (.X(_0476_),
    .B(_0474_),
    .A(net390));
 sg13g2_and2_1 _2710_ (.A(net320),
    .B(_0475_),
    .X(_0052_));
 sg13g2_nor2_2 _2711_ (.A(_0024_),
    .B(_0456_),
    .Y(_0477_));
 sg13g2_nand2b_2 _2712_ (.Y(_0478_),
    .B(_0455_),
    .A_N(_0024_));
 sg13g2_nor2_1 _2713_ (.A(net723),
    .B(net724),
    .Y(_0479_));
 sg13g2_and2_2 _2714_ (.A(_0023_),
    .B(_0479_),
    .X(_0480_));
 sg13g2_nand2_2 _2715_ (.Y(_0481_),
    .A(_0023_),
    .B(_0479_));
 sg13g2_nor2_1 _2716_ (.A(\cpu_instance.mem_instance.mem_ctrl_instance.start_write ),
    .B(\cpu_instance.mem_instance.mem_ctrl_instance.start_read ),
    .Y(_0482_));
 sg13g2_nor2_1 _2717_ (.A(_0481_),
    .B(_0482_),
    .Y(_0483_));
 sg13g2_nand2b_2 _2718_ (.Y(_0484_),
    .B(_0480_),
    .A_N(_0482_));
 sg13g2_nor2_2 _2719_ (.A(net691),
    .B(net688),
    .Y(_0485_));
 sg13g2_nand2_2 _2720_ (.Y(_0486_),
    .A(net689),
    .B(_0484_));
 sg13g2_a22oi_1 _2721_ (.Y(_0487_),
    .B1(_0485_),
    .B2(net328),
    .A2(net690),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[12] ));
 sg13g2_inv_1 _2722_ (.Y(_0053_),
    .A(net329));
 sg13g2_a22oi_1 _2723_ (.Y(_0488_),
    .B1(_0485_),
    .B2(net335),
    .A2(net691),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[13] ));
 sg13g2_inv_1 _2724_ (.Y(_0054_),
    .A(net336));
 sg13g2_a22oi_1 _2725_ (.Y(_0489_),
    .B1(_0485_),
    .B2(net330),
    .A2(net691),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[14] ));
 sg13g2_inv_1 _2726_ (.Y(_0055_),
    .A(net331));
 sg13g2_a22oi_1 _2727_ (.Y(_0490_),
    .B1(net685),
    .B2(net324),
    .A2(net691),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[15] ));
 sg13g2_inv_1 _2728_ (.Y(_0056_),
    .A(net325));
 sg13g2_a22oi_1 _2729_ (.Y(_0491_),
    .B1(net685),
    .B2(net355),
    .A2(net691),
    .A1(net328));
 sg13g2_inv_1 _2730_ (.Y(_0057_),
    .A(_0491_));
 sg13g2_a22oi_1 _2731_ (.Y(_0492_),
    .B1(net685),
    .B2(net376),
    .A2(net690),
    .A1(net335));
 sg13g2_inv_1 _2732_ (.Y(_0058_),
    .A(_0492_));
 sg13g2_a22oi_1 _2733_ (.Y(_0493_),
    .B1(net685),
    .B2(net389),
    .A2(net690),
    .A1(net330));
 sg13g2_inv_1 _2734_ (.Y(_0059_),
    .A(_0493_));
 sg13g2_a21o_1 _2735_ (.A2(_1494_),
    .A1(_1492_),
    .B1(_1568_),
    .X(_0494_));
 sg13g2_nand3_1 _2736_ (.B(_1575_),
    .C(_0494_),
    .A(_1569_),
    .Y(_0495_));
 sg13g2_nand4_1 _2737_ (.B(_1494_),
    .C(_1508_),
    .A(_1492_),
    .Y(_0496_),
    .D(_1512_));
 sg13g2_nand3_1 _2738_ (.B(_1515_),
    .C(_0496_),
    .A(_1325_),
    .Y(_0497_));
 sg13g2_nor4_1 _2739_ (.A(_1491_),
    .B(_1493_),
    .C(_1524_),
    .D(_1525_),
    .Y(_0498_));
 sg13g2_mux2_1 _2740_ (.A0(_1537_),
    .A1(_1591_),
    .S(_1485_),
    .X(_0499_));
 sg13g2_a221oi_1 _2741_ (.B2(_1509_),
    .C1(_0498_),
    .B1(_1560_),
    .A1(_1463_),
    .Y(_0500_),
    .A2(_1539_));
 sg13g2_a221oi_1 _2742_ (.B2(_1491_),
    .C1(_0499_),
    .B1(_1536_),
    .A1(_1494_),
    .Y(_0501_),
    .A2(_1529_));
 sg13g2_nand4_1 _2743_ (.B(_0497_),
    .C(_0500_),
    .A(_0495_),
    .Y(_0502_),
    .D(_0501_));
 sg13g2_and2_1 _2744_ (.A(net782),
    .B(\cpu_instance.ctrl_instance.mux_sel[2] ),
    .X(_0503_));
 sg13g2_a21oi_2 _2745_ (.B1(_0503_),
    .Y(_0504_),
    .A2(_0502_),
    .A1(\cpu_instance.ctrl_instance.mux_sel[0] ));
 sg13g2_a21o_2 _2746_ (.A2(_0502_),
    .A1(\cpu_instance.ctrl_instance.mux_sel[0] ),
    .B1(_0503_),
    .X(_0505_));
 sg13g2_or4_1 _2747_ (.A(\cpu_instance.ctrl_instance.state[7] ),
    .B(_0400_),
    .C(_0414_),
    .D(_0504_),
    .X(_0506_));
 sg13g2_o21ai_1 _2748_ (.B1(_0506_),
    .Y(_0060_),
    .A1(_1291_),
    .A2(_1320_));
 sg13g2_nand3_1 _2749_ (.B(net609),
    .C(_0387_),
    .A(net717),
    .Y(_0507_));
 sg13g2_nand3b_1 _2750_ (.B(net509),
    .C(_0436_),
    .Y(_0508_),
    .A_N(net445));
 sg13g2_nand2_1 _2751_ (.Y(_0509_),
    .A(_1291_),
    .B(net717));
 sg13g2_a22oi_1 _2752_ (.Y(_0510_),
    .B1(_0509_),
    .B2(net585),
    .A2(_0507_),
    .A1(net570));
 sg13g2_a21oi_1 _2753_ (.A1(_0508_),
    .A2(_0510_),
    .Y(_0061_),
    .B1(net741));
 sg13g2_a21oi_1 _2754_ (.A1(_1469_),
    .A2(_1570_),
    .Y(_0511_),
    .B1(_1576_));
 sg13g2_o21ai_1 _2755_ (.B1(_0511_),
    .Y(_0512_),
    .A1(_1469_),
    .A2(_1570_));
 sg13g2_nand3_1 _2756_ (.B(_1515_),
    .C(_1516_),
    .A(_1469_),
    .Y(_0513_));
 sg13g2_nand3b_1 _2757_ (.B(_0513_),
    .C(_1325_),
    .Y(_0514_),
    .A_N(_1517_));
 sg13g2_nand2_1 _2758_ (.Y(_0515_),
    .A(_1469_),
    .B(_1526_));
 sg13g2_nor2b_1 _2759_ (.A(_1463_),
    .B_N(_1537_),
    .Y(_0516_));
 sg13g2_o21ai_1 _2760_ (.B1(_1529_),
    .Y(_0517_),
    .A1(_1463_),
    .A2(_1466_));
 sg13g2_a22oi_1 _2761_ (.Y(_0518_),
    .B1(_1560_),
    .B2(_1485_),
    .A2(_1536_),
    .A1(_1468_));
 sg13g2_a221oi_1 _2762_ (.B2(_1463_),
    .C1(_0516_),
    .B1(_1591_),
    .A1(_1444_),
    .Y(_0519_),
    .A2(_1539_));
 sg13g2_nand4_1 _2763_ (.B(_0517_),
    .C(_0518_),
    .A(_0515_),
    .Y(_0520_),
    .D(_0519_));
 sg13g2_nand3b_1 _2764_ (.B(_0514_),
    .C(_0512_),
    .Y(_0521_),
    .A_N(_0520_));
 sg13g2_and2_1 _2765_ (.A(\cpu_instance.ctrl_instance.mux_sel[1] ),
    .B(net1),
    .X(_0522_));
 sg13g2_a221oi_1 _2766_ (.B2(_0521_),
    .C1(_0522_),
    .B1(\cpu_instance.ctrl_instance.mux_sel[0] ),
    .A1(\cpu_instance.mem_instance.bus_data_out[2] ),
    .Y(_0523_),
    .A2(\cpu_instance.ctrl_instance.mux_sel[2] ));
 sg13g2_inv_1 _2767_ (.Y(_0524_),
    .A(_0523_));
 sg13g2_nand2_1 _2768_ (.Y(_0525_),
    .A(_0408_),
    .B(_0414_));
 sg13g2_nand2_1 _2769_ (.Y(_0526_),
    .A(_0524_),
    .B(_0525_));
 sg13g2_nor2b_1 _2770_ (.A(_1527_),
    .B_N(_1324_),
    .Y(_0527_));
 sg13g2_a21oi_1 _2771_ (.A1(_1535_),
    .A2(_0527_),
    .Y(_0528_),
    .B1(_1526_));
 sg13g2_o21ai_1 _2772_ (.B1(_1530_),
    .Y(_0529_),
    .A1(_1568_),
    .A2(_0528_));
 sg13g2_nand2_1 _2773_ (.Y(_0530_),
    .A(_1508_),
    .B(_1513_));
 sg13g2_a22oi_1 _2774_ (.Y(_0531_),
    .B1(_1558_),
    .B2(net629),
    .A2(_1537_),
    .A1(_1508_));
 sg13g2_a21oi_1 _2775_ (.A1(_1512_),
    .A2(_1536_),
    .Y(_0532_),
    .B1(_1591_));
 sg13g2_nor2_1 _2776_ (.A(_1508_),
    .B(_0532_),
    .Y(_0533_));
 sg13g2_a221oi_1 _2777_ (.B2(_0530_),
    .C1(_0533_),
    .B1(_0529_),
    .A1(_1485_),
    .Y(_0534_),
    .A2(_1539_));
 sg13g2_nand2_1 _2778_ (.Y(_0535_),
    .A(_0531_),
    .B(_0534_));
 sg13g2_a21oi_2 _2779_ (.B1(_1300_),
    .Y(_0536_),
    .A2(_0534_),
    .A1(_0531_));
 sg13g2_and2_1 _2780_ (.A(\cpu_instance.mem_instance.bus_data_out[0] ),
    .B(\cpu_instance.ctrl_instance.mux_sel[2] ),
    .X(_0537_));
 sg13g2_nor2_1 _2781_ (.A(_0536_),
    .B(_0537_),
    .Y(_0538_));
 sg13g2_inv_1 _2782_ (.Y(_0539_),
    .A(net624));
 sg13g2_o21ai_1 _2783_ (.B1(_0526_),
    .Y(_0540_),
    .A1(_0403_),
    .A2(net623));
 sg13g2_nor3_2 _2784_ (.A(_0399_),
    .B(_0431_),
    .C(_0437_),
    .Y(_0541_));
 sg13g2_a22oi_1 _2785_ (.Y(_0542_),
    .B1(_0540_),
    .B2(_0541_),
    .A2(_0437_),
    .A1(net733));
 sg13g2_nor2_1 _2786_ (.A(net742),
    .B(_0542_),
    .Y(_0062_));
 sg13g2_nor2_1 _2787_ (.A(_1566_),
    .B(_1567_),
    .Y(_0543_));
 sg13g2_nand2b_1 _2788_ (.Y(_0544_),
    .B(_1575_),
    .A_N(_1571_));
 sg13g2_o21ai_1 _2789_ (.B1(_1325_),
    .Y(_0545_),
    .A1(_1467_),
    .A2(_1517_));
 sg13g2_nand3b_1 _2790_ (.B(_0544_),
    .C(_0545_),
    .Y(_0546_),
    .A_N(_1526_));
 sg13g2_and2_1 _2791_ (.A(_0543_),
    .B(_0546_),
    .X(_0547_));
 sg13g2_or3_1 _2792_ (.A(_1326_),
    .B(_1467_),
    .C(_1517_),
    .X(_0548_));
 sg13g2_nand2_1 _2793_ (.Y(_0549_),
    .A(_1571_),
    .B(_1575_));
 sg13g2_a21oi_1 _2794_ (.A1(_0548_),
    .A2(_0549_),
    .Y(_0550_),
    .B1(_0543_));
 sg13g2_mux2_1 _2795_ (.A0(_1537_),
    .A1(_1591_),
    .S(_1444_),
    .X(_0551_));
 sg13g2_a221oi_1 _2796_ (.B2(_1463_),
    .C1(_0551_),
    .B1(_1560_),
    .A1(_1426_),
    .Y(_0552_),
    .A2(_1539_));
 sg13g2_a22oi_1 _2797_ (.Y(_0553_),
    .B1(_1567_),
    .B2(_1536_),
    .A2(_1565_),
    .A1(_1529_));
 sg13g2_nand3b_1 _2798_ (.B(_0552_),
    .C(_0553_),
    .Y(_0554_),
    .A_N(_0550_));
 sg13g2_o21ai_1 _2799_ (.B1(\cpu_instance.ctrl_instance.mux_sel[0] ),
    .Y(_0555_),
    .A1(_0547_),
    .A2(_0554_));
 sg13g2_and2_1 _2800_ (.A(\cpu_instance.mem_instance.bus_data_out[3] ),
    .B(\cpu_instance.ctrl_instance.mux_sel[2] ),
    .X(_0556_));
 sg13g2_a21o_1 _2801_ (.A2(net2),
    .A1(\cpu_instance.ctrl_instance.mux_sel[1] ),
    .B1(_0556_),
    .X(_0557_));
 sg13g2_nor2b_2 _2802_ (.A(_0557_),
    .B_N(_0555_),
    .Y(_0558_));
 sg13g2_inv_4 _2803_ (.A(net613),
    .Y(_0559_));
 sg13g2_nand2_1 _2804_ (.Y(_0560_),
    .A(_0525_),
    .B(_0559_));
 sg13g2_o21ai_1 _2805_ (.B1(_0560_),
    .Y(_0561_),
    .A1(_0403_),
    .A2(_0504_));
 sg13g2_a22oi_1 _2806_ (.Y(_0562_),
    .B1(_0541_),
    .B2(_0561_),
    .A2(_0437_),
    .A1(net729));
 sg13g2_nor2_1 _2807_ (.A(net742),
    .B(_0562_),
    .Y(_0063_));
 sg13g2_nor2_1 _2808_ (.A(net715),
    .B(_0392_),
    .Y(_0563_));
 sg13g2_o21ai_1 _2809_ (.B1(_0431_),
    .Y(_0564_),
    .A1(net608),
    .A2(_0558_));
 sg13g2_nand3_1 _2810_ (.B(_0435_),
    .C(_0524_),
    .A(_1601_),
    .Y(_0565_));
 sg13g2_a21oi_1 _2811_ (.A1(net591),
    .A2(_0565_),
    .Y(_0566_),
    .B1(_0465_));
 sg13g2_nand2_1 _2812_ (.Y(_0567_),
    .A(_0564_),
    .B(_0566_));
 sg13g2_nand2_1 _2813_ (.Y(_0568_),
    .A(net718),
    .B(_1599_));
 sg13g2_o21ai_1 _2814_ (.B1(_0567_),
    .Y(_0569_),
    .A1(net526),
    .A2(_0568_));
 sg13g2_a22oi_1 _2815_ (.Y(_0570_),
    .B1(_0563_),
    .B2(net527),
    .A2(_1316_),
    .A1(\cpu_instance.ctrl_instance.reg_sel_in[0] ));
 sg13g2_nor2_1 _2816_ (.A(net741),
    .B(net528),
    .Y(_0064_));
 sg13g2_nand2_1 _2817_ (.Y(_0571_),
    .A(net809),
    .B(net715));
 sg13g2_nand3_1 _2818_ (.B(_0435_),
    .C(_0559_),
    .A(_1601_),
    .Y(_0572_));
 sg13g2_a221oi_1 _2819_ (.B2(net591),
    .C1(_0465_),
    .B1(_0572_),
    .A1(_0431_),
    .Y(_0573_),
    .A2(_0435_));
 sg13g2_nor3_1 _2820_ (.A(net583),
    .B(net526),
    .C(net609),
    .Y(_0574_));
 sg13g2_o21ai_1 _2821_ (.B1(_0563_),
    .Y(_0575_),
    .A1(_0573_),
    .A2(_0574_));
 sg13g2_a21oi_1 _2822_ (.A1(_0571_),
    .A2(_0575_),
    .Y(_0065_),
    .B1(net741));
 sg13g2_nand2_2 _2823_ (.Y(_0576_),
    .A(net718),
    .B(_1318_));
 sg13g2_or4_1 _2824_ (.A(_0502_),
    .B(_0521_),
    .C(_0535_),
    .D(_0576_),
    .X(_0577_));
 sg13g2_nor3_1 _2825_ (.A(_0547_),
    .B(_0554_),
    .C(_0577_),
    .Y(_0578_));
 sg13g2_nand3b_1 _2826_ (.B(_1595_),
    .C(_0578_),
    .Y(_0579_),
    .A_N(_1580_));
 sg13g2_nor4_2 _2827_ (.A(_0357_),
    .B(_0369_),
    .C(_0383_),
    .Y(_0580_),
    .D(_0579_));
 sg13g2_a21o_1 _2828_ (.A2(_0396_),
    .A1(net384),
    .B1(_0580_),
    .X(_0066_));
 sg13g2_nand3_1 _2829_ (.B(_0344_),
    .C(_0356_),
    .A(_1325_),
    .Y(_0581_));
 sg13g2_a21oi_1 _2830_ (.A1(_0345_),
    .A2(_0367_),
    .Y(_0582_),
    .B1(_1576_));
 sg13g2_a221oi_1 _2831_ (.B2(net629),
    .C1(_0582_),
    .B1(_1559_),
    .A1(_1509_),
    .Y(_0583_),
    .A2(_1538_));
 sg13g2_a21oi_1 _2832_ (.A1(_0581_),
    .A2(_0583_),
    .Y(_0584_),
    .B1(_0576_));
 sg13g2_a21o_1 _2833_ (.A2(_0396_),
    .A1(net419),
    .B1(_0584_),
    .X(_0067_));
 sg13g2_nand2_1 _2834_ (.Y(_0585_),
    .A(net790),
    .B(_1318_));
 sg13g2_or3_2 _2835_ (.A(\cpu_instance.ctrl_instance.state[3] ),
    .B(net591),
    .C(_0404_),
    .X(_0586_));
 sg13g2_o21ai_1 _2836_ (.B1(_0585_),
    .Y(_0068_),
    .A1(net620),
    .A2(_0586_));
 sg13g2_nand2_1 _2837_ (.Y(_0587_),
    .A(net793),
    .B(_1318_));
 sg13g2_o21ai_1 _2838_ (.B1(_0587_),
    .Y(_0069_),
    .A1(net615),
    .A2(_0586_));
 sg13g2_nand2_1 _2839_ (.Y(_0588_),
    .A(net813),
    .B(_1318_));
 sg13g2_o21ai_1 _2840_ (.B1(_0588_),
    .Y(_0070_),
    .A1(net605),
    .A2(_0586_));
 sg13g2_nand2_1 _2841_ (.Y(_0589_),
    .A(net807),
    .B(_1318_));
 sg13g2_o21ai_1 _2842_ (.B1(_0589_),
    .Y(_0071_),
    .A1(net611),
    .A2(_0586_));
 sg13g2_nand3_1 _2843_ (.B(_0387_),
    .C(_0505_),
    .A(_1600_),
    .Y(_0590_));
 sg13g2_o21ai_1 _2844_ (.B1(_0590_),
    .Y(_0591_),
    .A1(_0414_),
    .A2(net624));
 sg13g2_or2_1 _2845_ (.X(_0592_),
    .B(_0392_),
    .A(net853));
 sg13g2_a21oi_1 _2846_ (.A1(net719),
    .A2(net620),
    .Y(_0593_),
    .B1(_0592_));
 sg13g2_o21ai_1 _2847_ (.B1(_0593_),
    .Y(_0594_),
    .A1(net719),
    .A2(_0591_));
 sg13g2_o21ai_1 _2848_ (.B1(net773),
    .Y(_0595_),
    .A1(net796),
    .A2(_0436_));
 sg13g2_a21oi_1 _2849_ (.A1(_0436_),
    .A2(_0594_),
    .Y(_0072_),
    .B1(_0595_));
 sg13g2_and4_1 _2850_ (.A(_1601_),
    .B(_0387_),
    .C(_0435_),
    .D(_0505_),
    .X(_0596_));
 sg13g2_nor3_1 _2851_ (.A(net609),
    .B(_0432_),
    .C(net620),
    .Y(_0597_));
 sg13g2_nor3_1 _2852_ (.A(net719),
    .B(_0596_),
    .C(_0597_),
    .Y(_0598_));
 sg13g2_nand2_1 _2853_ (.Y(_0599_),
    .A(net719),
    .B(_0558_));
 sg13g2_nor3_1 _2854_ (.A(net715),
    .B(_0592_),
    .C(_0598_),
    .Y(_0600_));
 sg13g2_a22oi_1 _2855_ (.Y(_0601_),
    .B1(_0599_),
    .B2(_0600_),
    .A2(net715),
    .A1(net393));
 sg13g2_nor2_1 _2856_ (.A(net741),
    .B(_0601_),
    .Y(_0073_));
 sg13g2_nand2_1 _2857_ (.Y(_0602_),
    .A(\cpu_instance.addr_reg_op[1] ),
    .B(\cpu_instance.addr_reg_op[0] ));
 sg13g2_nor2_1 _2858_ (.A(\cpu_instance.addr_reg_op[1] ),
    .B(\cpu_instance.addr_reg_op[0] ),
    .Y(_0603_));
 sg13g2_or2_1 _2859_ (.X(_0604_),
    .B(\cpu_instance.addr_reg_op[0] ),
    .A(\cpu_instance.addr_reg_op[1] ));
 sg13g2_nand3_1 _2860_ (.B(_0602_),
    .C(_0604_),
    .A(_0026_),
    .Y(_0605_));
 sg13g2_nor2_2 _2861_ (.A(\cpu_instance.addr_reg_op[2] ),
    .B(_0602_),
    .Y(_0606_));
 sg13g2_or2_2 _2862_ (.X(_0607_),
    .B(_0602_),
    .A(\cpu_instance.addr_reg_op[2] ));
 sg13g2_and2_1 _2863_ (.A(\cpu_instance.addr_reg_op[2] ),
    .B(_0603_),
    .X(_0608_));
 sg13g2_nand2_1 _2864_ (.Y(_0609_),
    .A(\cpu_instance.addr_reg_op[2] ),
    .B(_0603_));
 sg13g2_nor2_1 _2865_ (.A(_0606_),
    .B(_0608_),
    .Y(_0610_));
 sg13g2_nor2_1 _2866_ (.A(\cpu_instance.mem_instance.addr[24] ),
    .B(_0605_),
    .Y(_0611_));
 sg13g2_o21ai_1 _2867_ (.B1(_0607_),
    .Y(_0612_),
    .A1(_0026_),
    .A2(_0604_));
 sg13g2_a221oi_1 _2868_ (.B2(net736),
    .C1(_0611_),
    .B1(_0612_),
    .A1(_0605_),
    .Y(_0613_),
    .A2(_0610_));
 sg13g2_nand3b_1 _2869_ (.B(_0026_),
    .C(\cpu_instance.addr_reg_op[1] ),
    .Y(_0614_),
    .A_N(\cpu_instance.addr_reg_op[0] ));
 sg13g2_nor2b_1 _2870_ (.A(_0612_),
    .B_N(_0614_),
    .Y(_0615_));
 sg13g2_nand2b_1 _2871_ (.Y(_0616_),
    .B(_0614_),
    .A_N(_0612_));
 sg13g2_mux2_1 _2872_ (.A0(_0026_),
    .A1(net622),
    .S(net702),
    .X(_0617_));
 sg13g2_mux2_1 _2873_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][0] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][0] ),
    .S(net735),
    .X(_0618_));
 sg13g2_nand2b_1 _2874_ (.Y(_0619_),
    .B(net711),
    .A_N(_0617_));
 sg13g2_xnor2_1 _2875_ (.Y(_0620_),
    .A(_0617_),
    .B(net711));
 sg13g2_nand2_1 _2876_ (.Y(_0621_),
    .A(net622),
    .B(net677));
 sg13g2_o21ai_1 _2877_ (.B1(_0621_),
    .Y(_0622_),
    .A1(net677),
    .A2(_0620_));
 sg13g2_o21ai_1 _2878_ (.B1(net745),
    .Y(_0623_),
    .A1(net440),
    .A2(net681));
 sg13g2_a21oi_1 _2879_ (.A1(net681),
    .A2(_0622_),
    .Y(_0074_),
    .B1(_0623_));
 sg13g2_o21ai_1 _2880_ (.B1(_0607_),
    .Y(_0624_),
    .A1(_0536_),
    .A2(_0537_));
 sg13g2_xnor2_1 _2881_ (.Y(_0625_),
    .A(_0505_),
    .B(_0624_));
 sg13g2_mux2_1 _2882_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][1] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][1] ),
    .S(net735),
    .X(_0626_));
 sg13g2_nand3_1 _2883_ (.B(_0625_),
    .C(_0626_),
    .A(net702),
    .Y(_0627_));
 sg13g2_a21oi_1 _2884_ (.A1(net701),
    .A2(_0625_),
    .Y(_0628_),
    .B1(_0626_));
 sg13g2_a21o_1 _2885_ (.A2(_0625_),
    .A1(net701),
    .B1(net707),
    .X(_0629_));
 sg13g2_nand2_1 _2886_ (.Y(_0630_),
    .A(_0627_),
    .B(_0629_));
 sg13g2_a21oi_1 _2887_ (.A1(_0619_),
    .A2(_0630_),
    .Y(_0631_),
    .B1(net677));
 sg13g2_o21ai_1 _2888_ (.B1(_0631_),
    .Y(_0632_),
    .A1(_0619_),
    .A2(_0630_));
 sg13g2_o21ai_1 _2889_ (.B1(_0632_),
    .Y(_0633_),
    .A1(net626),
    .A2(net676));
 sg13g2_inv_1 _2890_ (.Y(_0634_),
    .A(_0633_));
 sg13g2_o21ai_1 _2891_ (.B1(net745),
    .Y(_0635_),
    .A1(net566),
    .A2(net681));
 sg13g2_a21oi_1 _2892_ (.A1(net681),
    .A2(_0634_),
    .Y(_0075_),
    .B1(_0635_));
 sg13g2_nor2_1 _2893_ (.A(net619),
    .B(net676),
    .Y(_0636_));
 sg13g2_a21oi_1 _2894_ (.A1(net625),
    .A2(net622),
    .Y(_0637_),
    .B1(_0606_));
 sg13g2_xnor2_1 _2895_ (.Y(_0638_),
    .A(net619),
    .B(_0637_));
 sg13g2_mux2_2 _2896_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][2] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][2] ),
    .S(net735),
    .X(_0639_));
 sg13g2_a21o_1 _2897_ (.A2(_0638_),
    .A1(net702),
    .B1(_0639_),
    .X(_0640_));
 sg13g2_nand3_1 _2898_ (.B(_0638_),
    .C(_0639_),
    .A(net702),
    .Y(_0641_));
 sg13g2_nand2_1 _2899_ (.Y(_0642_),
    .A(_0640_),
    .B(_0641_));
 sg13g2_o21ai_1 _2900_ (.B1(_0627_),
    .Y(_0643_),
    .A1(_0619_),
    .A2(_0628_));
 sg13g2_nand3_1 _2901_ (.B(_0641_),
    .C(_0643_),
    .A(_0640_),
    .Y(_0644_));
 sg13g2_xnor2_1 _2902_ (.Y(_0645_),
    .A(_0642_),
    .B(_0643_));
 sg13g2_a21oi_1 _2903_ (.A1(net676),
    .A2(_0645_),
    .Y(_0646_),
    .B1(_0636_));
 sg13g2_o21ai_1 _2904_ (.B1(net745),
    .Y(_0647_),
    .A1(net405),
    .A2(net681));
 sg13g2_a21oi_1 _2905_ (.A1(net681),
    .A2(_0646_),
    .Y(_0076_),
    .B1(_0647_));
 sg13g2_and2_1 _2906_ (.A(_0641_),
    .B(_0644_),
    .X(_0648_));
 sg13g2_and3_2 _2907_ (.X(_0649_),
    .A(net627),
    .B(net620),
    .C(net622));
 sg13g2_nor2_1 _2908_ (.A(_0606_),
    .B(_0649_),
    .Y(_0650_));
 sg13g2_xnor2_1 _2909_ (.Y(_0651_),
    .A(net613),
    .B(_0650_));
 sg13g2_mux2_2 _2910_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][3] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][3] ),
    .S(net735),
    .X(_0652_));
 sg13g2_nand3_1 _2911_ (.B(_0651_),
    .C(_0652_),
    .A(net701),
    .Y(_0653_));
 sg13g2_a21oi_1 _2912_ (.A1(net701),
    .A2(_0651_),
    .Y(_0654_),
    .B1(_0652_));
 sg13g2_a21o_1 _2913_ (.A2(_0651_),
    .A1(net701),
    .B1(_0652_),
    .X(_0655_));
 sg13g2_nand2_1 _2914_ (.Y(_0656_),
    .A(_0653_),
    .B(_0655_));
 sg13g2_xnor2_1 _2915_ (.Y(_0657_),
    .A(_0648_),
    .B(_0656_));
 sg13g2_nand2_1 _2916_ (.Y(_0658_),
    .A(net676),
    .B(_0657_));
 sg13g2_o21ai_1 _2917_ (.B1(_0658_),
    .Y(_0659_),
    .A1(_0559_),
    .A2(net676));
 sg13g2_o21ai_1 _2918_ (.B1(net746),
    .Y(_0660_),
    .A1(net361),
    .A2(net681));
 sg13g2_a21oi_1 _2919_ (.A1(net681),
    .A2(_0659_),
    .Y(_0077_),
    .B1(_0660_));
 sg13g2_o21ai_1 _2920_ (.B1(_0653_),
    .Y(_0661_),
    .A1(_0648_),
    .A2(_0654_));
 sg13g2_nand3b_1 _2921_ (.B(_0649_),
    .C(_0555_),
    .Y(_0662_),
    .A_N(_0557_));
 sg13g2_nand3_1 _2922_ (.B(_0607_),
    .C(_0662_),
    .A(net616),
    .Y(_0663_));
 sg13g2_a21o_1 _2923_ (.A2(_0662_),
    .A1(_0607_),
    .B1(net616),
    .X(_0664_));
 sg13g2_nand3_1 _2924_ (.B(_0663_),
    .C(_0664_),
    .A(net703),
    .Y(_0665_));
 sg13g2_mux2_2 _2925_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][4] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][4] ),
    .S(net736),
    .X(_0666_));
 sg13g2_inv_1 _2926_ (.Y(_0667_),
    .A(_0666_));
 sg13g2_nor2_1 _2927_ (.A(_0665_),
    .B(_0667_),
    .Y(_0668_));
 sg13g2_xnor2_1 _2928_ (.Y(_0669_),
    .A(_0665_),
    .B(_0666_));
 sg13g2_o21ai_1 _2929_ (.B1(net675),
    .Y(_0670_),
    .A1(_0661_),
    .A2(_0669_));
 sg13g2_a21oi_1 _2930_ (.A1(_0661_),
    .A2(_0669_),
    .Y(_0671_),
    .B1(_0670_));
 sg13g2_a21oi_1 _2931_ (.A1(net616),
    .A2(net677),
    .Y(_0672_),
    .B1(_0671_));
 sg13g2_o21ai_1 _2932_ (.B1(net769),
    .Y(_0673_),
    .A1(net421),
    .A2(net683));
 sg13g2_a21oi_1 _2933_ (.A1(net683),
    .A2(_0672_),
    .Y(_0078_),
    .B1(_0673_));
 sg13g2_a21oi_1 _2934_ (.A1(_0661_),
    .A2(_0669_),
    .Y(_0674_),
    .B1(_0668_));
 sg13g2_nor2_2 _2935_ (.A(net616),
    .B(_0662_),
    .Y(_0675_));
 sg13g2_o21ai_1 _2936_ (.B1(net608),
    .Y(_0676_),
    .A1(_0606_),
    .A2(_0675_));
 sg13g2_or3_1 _2937_ (.A(net608),
    .B(_0606_),
    .C(_0675_),
    .X(_0677_));
 sg13g2_and3_1 _2938_ (.X(_0678_),
    .A(net703),
    .B(_0676_),
    .C(_0677_));
 sg13g2_mux2_2 _2939_ (.A0(net380),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][5] ),
    .S(net735),
    .X(_0679_));
 sg13g2_inv_1 _2940_ (.Y(_0680_),
    .A(_0679_));
 sg13g2_nor2_1 _2941_ (.A(_0678_),
    .B(_0679_),
    .Y(_0681_));
 sg13g2_xnor2_1 _2942_ (.Y(_0682_),
    .A(_0678_),
    .B(_0679_));
 sg13g2_xnor2_1 _2943_ (.Y(_0683_),
    .A(_0674_),
    .B(_0682_));
 sg13g2_nor2_1 _2944_ (.A(net678),
    .B(_0683_),
    .Y(_0684_));
 sg13g2_a21oi_2 _2945_ (.B1(_0684_),
    .Y(_0685_),
    .A2(net677),
    .A1(net602));
 sg13g2_o21ai_1 _2946_ (.B1(net746),
    .Y(_0686_),
    .A1(net380),
    .A2(net683));
 sg13g2_a21oi_1 _2947_ (.A1(net683),
    .A2(_0685_),
    .Y(_0079_),
    .B1(_0686_));
 sg13g2_and2_1 _2948_ (.A(net608),
    .B(_0675_),
    .X(_0687_));
 sg13g2_nand2_1 _2949_ (.Y(_0688_),
    .A(net608),
    .B(_0675_));
 sg13g2_a21oi_1 _2950_ (.A1(net608),
    .A2(_0675_),
    .Y(_0689_),
    .B1(_0606_));
 sg13g2_xnor2_1 _2951_ (.Y(_0690_),
    .A(net599),
    .B(_0689_));
 sg13g2_mux2_2 _2952_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][6] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][6] ),
    .S(net735),
    .X(_0691_));
 sg13g2_and3_1 _2953_ (.X(_0692_),
    .A(net701),
    .B(_0690_),
    .C(_0691_));
 sg13g2_nand3_1 _2954_ (.B(_0690_),
    .C(_0691_),
    .A(net701),
    .Y(_0693_));
 sg13g2_a21oi_1 _2955_ (.A1(net701),
    .A2(_0690_),
    .Y(_0694_),
    .B1(_0691_));
 sg13g2_or2_1 _2956_ (.X(_0695_),
    .B(_0694_),
    .A(_0692_));
 sg13g2_a221oi_1 _2957_ (.B2(_0679_),
    .C1(_0668_),
    .B1(_0678_),
    .A1(_0661_),
    .Y(_0696_),
    .A2(_0669_));
 sg13g2_or2_1 _2958_ (.X(_0697_),
    .B(_0696_),
    .A(_0681_));
 sg13g2_or4_1 _2959_ (.A(_0681_),
    .B(_0692_),
    .C(_0694_),
    .D(_0696_),
    .X(_0698_));
 sg13g2_a21oi_1 _2960_ (.A1(_0695_),
    .A2(_0697_),
    .Y(_0699_),
    .B1(net677));
 sg13g2_a22oi_1 _2961_ (.Y(_0700_),
    .B1(_0698_),
    .B2(_0699_),
    .A2(net677),
    .A1(_0386_));
 sg13g2_o21ai_1 _2962_ (.B1(net745),
    .Y(_0701_),
    .A1(net394),
    .A2(net682));
 sg13g2_a21oi_1 _2963_ (.A1(net682),
    .A2(_0700_),
    .Y(_0080_),
    .B1(_0701_));
 sg13g2_a21oi_1 _2964_ (.A1(net599),
    .A2(_0687_),
    .Y(_0702_),
    .B1(_0606_));
 sg13g2_nand2b_1 _2965_ (.Y(_0703_),
    .B(net594),
    .A_N(_0702_));
 sg13g2_a21oi_1 _2966_ (.A1(net591),
    .A2(_0702_),
    .Y(_0704_),
    .B1(_0608_));
 sg13g2_mux2_2 _2967_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][7] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][7] ),
    .S(net734),
    .X(_0705_));
 sg13g2_inv_1 _2968_ (.Y(_0706_),
    .A(_0705_));
 sg13g2_and3_1 _2969_ (.X(_0707_),
    .A(_0703_),
    .B(_0704_),
    .C(_0705_));
 sg13g2_a21o_1 _2970_ (.A2(_0704_),
    .A1(_0703_),
    .B1(_0706_),
    .X(_0708_));
 sg13g2_nand3_1 _2971_ (.B(_0704_),
    .C(_0706_),
    .A(_0703_),
    .Y(_0709_));
 sg13g2_nand4_1 _2972_ (.B(_0698_),
    .C(_0708_),
    .A(_0693_),
    .Y(_0710_),
    .D(_0709_));
 sg13g2_a22oi_1 _2973_ (.Y(_0711_),
    .B1(_0708_),
    .B2(_0709_),
    .A2(_0698_),
    .A1(_0693_));
 sg13g2_nor2_1 _2974_ (.A(net678),
    .B(_0711_),
    .Y(_0712_));
 sg13g2_a22oi_1 _2975_ (.Y(_0713_),
    .B1(_0710_),
    .B2(_0712_),
    .A2(net677),
    .A1(net591));
 sg13g2_o21ai_1 _2976_ (.B1(net746),
    .Y(_0714_),
    .A1(net787),
    .A2(net682));
 sg13g2_a21oi_1 _2977_ (.A1(net682),
    .A2(_0713_),
    .Y(_0081_),
    .B1(_0714_));
 sg13g2_a221oi_1 _2978_ (.B2(_0431_),
    .C1(_0606_),
    .B1(_0687_),
    .A1(\cpu_instance.addr_reg_op[2] ),
    .Y(_0715_),
    .A2(_0603_));
 sg13g2_o21ai_1 _2979_ (.B1(_0610_),
    .Y(_0716_),
    .A1(_0432_),
    .A2(_0688_));
 sg13g2_mux2_2 _2980_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][8] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][8] ),
    .S(net734),
    .X(_0717_));
 sg13g2_inv_2 _2981_ (.Y(_0718_),
    .A(_0717_));
 sg13g2_nand2_1 _2982_ (.Y(_0719_),
    .A(_0715_),
    .B(_0717_));
 sg13g2_xnor2_1 _2983_ (.Y(_0720_),
    .A(net589),
    .B(_0717_));
 sg13g2_xnor2_1 _2984_ (.Y(_0721_),
    .A(net589),
    .B(_0718_));
 sg13g2_or3_1 _2985_ (.A(_0707_),
    .B(_0711_),
    .C(_0720_),
    .X(_0722_));
 sg13g2_o21ai_1 _2986_ (.B1(_0720_),
    .Y(_0723_),
    .A1(_0707_),
    .A2(_0711_));
 sg13g2_nand3_1 _2987_ (.B(_0722_),
    .C(_0723_),
    .A(net675),
    .Y(_0724_));
 sg13g2_o21ai_1 _2988_ (.B1(net743),
    .Y(_0725_),
    .A1(net379),
    .A2(net679));
 sg13g2_a21oi_1 _2989_ (.A1(net679),
    .A2(_0724_),
    .Y(_0082_),
    .B1(_0725_));
 sg13g2_nor2_1 _2990_ (.A(net734),
    .B(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][9] ),
    .Y(_0726_));
 sg13g2_nand2b_1 _2991_ (.Y(_0727_),
    .B(net734),
    .A_N(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][9] ));
 sg13g2_nor2b_2 _2992_ (.A(_0726_),
    .B_N(_0727_),
    .Y(_0728_));
 sg13g2_nand2b_1 _2993_ (.Y(_0729_),
    .B(_0727_),
    .A_N(_0726_));
 sg13g2_nor2_1 _2994_ (.A(_0715_),
    .B(_0728_),
    .Y(_0730_));
 sg13g2_xnor2_1 _2995_ (.Y(_0731_),
    .A(net589),
    .B(_0729_));
 sg13g2_a21o_1 _2996_ (.A2(_0723_),
    .A1(_0719_),
    .B1(_0731_),
    .X(_0732_));
 sg13g2_nand3_1 _2997_ (.B(_0723_),
    .C(_0731_),
    .A(_0719_),
    .Y(_0733_));
 sg13g2_nand3_1 _2998_ (.B(_0732_),
    .C(_0733_),
    .A(net675),
    .Y(_0734_));
 sg13g2_o21ai_1 _2999_ (.B1(net743),
    .Y(_0735_),
    .A1(net548),
    .A2(net680));
 sg13g2_a21oi_1 _3000_ (.A1(net680),
    .A2(_0734_),
    .Y(_0083_),
    .B1(_0735_));
 sg13g2_mux2_2 _3001_ (.A0(net381),
    .A1(net855),
    .S(net734),
    .X(_0736_));
 sg13g2_nor2b_1 _3002_ (.A(net589),
    .B_N(_0736_),
    .Y(_0737_));
 sg13g2_xor2_1 _3003_ (.B(_0736_),
    .A(net589),
    .X(_0738_));
 sg13g2_o21ai_1 _3004_ (.B1(_0715_),
    .Y(_0739_),
    .A1(_0717_),
    .A2(_0728_));
 sg13g2_a21oi_1 _3005_ (.A1(_0718_),
    .A2(_0729_),
    .Y(_0740_),
    .B1(net589));
 sg13g2_a21o_1 _3006_ (.A2(_0739_),
    .A1(_0723_),
    .B1(_0730_),
    .X(_0741_));
 sg13g2_nor2_1 _3007_ (.A(_0738_),
    .B(_0741_),
    .Y(_0742_));
 sg13g2_a21oi_1 _3008_ (.A1(_0738_),
    .A2(_0741_),
    .Y(_0743_),
    .B1(net678));
 sg13g2_nand2b_1 _3009_ (.Y(_0744_),
    .B(_0743_),
    .A_N(_0742_));
 sg13g2_o21ai_1 _3010_ (.B1(net743),
    .Y(_0745_),
    .A1(net381),
    .A2(net679));
 sg13g2_a21oi_1 _3011_ (.A1(net679),
    .A2(_0744_),
    .Y(_0084_),
    .B1(_0745_));
 sg13g2_mux2_2 _3012_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][11] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][11] ),
    .S(net734),
    .X(_0746_));
 sg13g2_inv_1 _3013_ (.Y(_0747_),
    .A(_0746_));
 sg13g2_xnor2_1 _3014_ (.Y(_0748_),
    .A(net589),
    .B(_0746_));
 sg13g2_xnor2_1 _3015_ (.Y(_0749_),
    .A(net590),
    .B(_0747_));
 sg13g2_o21ai_1 _3016_ (.B1(_0748_),
    .Y(_0750_),
    .A1(_0737_),
    .A2(_0742_));
 sg13g2_or3_1 _3017_ (.A(_0737_),
    .B(_0742_),
    .C(_0748_),
    .X(_0751_));
 sg13g2_nand3_1 _3018_ (.B(_0750_),
    .C(_0751_),
    .A(net675),
    .Y(_0752_));
 sg13g2_o21ai_1 _3019_ (.B1(net743),
    .Y(_0753_),
    .A1(net508),
    .A2(net679));
 sg13g2_a21oi_1 _3020_ (.A1(net679),
    .A2(_0752_),
    .Y(_0085_),
    .B1(_0753_));
 sg13g2_nor2_1 _3021_ (.A(_0738_),
    .B(_0749_),
    .Y(_0754_));
 sg13g2_nor4_1 _3022_ (.A(_0721_),
    .B(_0731_),
    .C(_0738_),
    .D(_0749_),
    .Y(_0755_));
 sg13g2_o21ai_1 _3023_ (.B1(_0755_),
    .Y(_0756_),
    .A1(_0707_),
    .A2(_0711_));
 sg13g2_a221oi_1 _3024_ (.B2(_0740_),
    .C1(_0737_),
    .B1(_0754_),
    .A1(_0715_),
    .Y(_0757_),
    .A2(_0746_));
 sg13g2_mux2_2 _3025_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][12] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][12] ),
    .S(net734),
    .X(_0758_));
 sg13g2_nand2_1 _3026_ (.Y(_0759_),
    .A(_0715_),
    .B(_0758_));
 sg13g2_xor2_1 _3027_ (.B(_0758_),
    .A(net589),
    .X(_0760_));
 sg13g2_nand3_1 _3028_ (.B(_0757_),
    .C(_0760_),
    .A(_0756_),
    .Y(_0761_));
 sg13g2_a21o_1 _3029_ (.A2(_0757_),
    .A1(_0756_),
    .B1(_0760_),
    .X(_0762_));
 sg13g2_nand3_1 _3030_ (.B(_0761_),
    .C(_0762_),
    .A(net675),
    .Y(_0763_));
 sg13g2_o21ai_1 _3031_ (.B1(net744),
    .Y(_0764_),
    .A1(net563),
    .A2(net679));
 sg13g2_a21oi_1 _3032_ (.A1(net679),
    .A2(_0763_),
    .Y(_0086_),
    .B1(_0764_));
 sg13g2_mux2_2 _3033_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][13] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][13] ),
    .S(net736),
    .X(_0765_));
 sg13g2_nand2_1 _3034_ (.Y(_0766_),
    .A(_0715_),
    .B(_0765_));
 sg13g2_xnor2_1 _3035_ (.Y(_0767_),
    .A(net590),
    .B(_0765_));
 sg13g2_nand2_1 _3036_ (.Y(_0768_),
    .A(_0759_),
    .B(_0762_));
 sg13g2_o21ai_1 _3037_ (.B1(net675),
    .Y(_0769_),
    .A1(_0767_),
    .A2(_0768_));
 sg13g2_a21o_1 _3038_ (.A2(_0768_),
    .A1(_0767_),
    .B1(_0769_),
    .X(_0770_));
 sg13g2_o21ai_1 _3039_ (.B1(net744),
    .Y(_0771_),
    .A1(net463),
    .A2(net680));
 sg13g2_a21oi_1 _3040_ (.A1(net680),
    .A2(_0770_),
    .Y(_0087_),
    .B1(_0771_));
 sg13g2_nand2b_1 _3041_ (.Y(_0772_),
    .B(_0767_),
    .A_N(_0760_));
 sg13g2_a21o_1 _3042_ (.A2(_0757_),
    .A1(_0756_),
    .B1(_0772_),
    .X(_0773_));
 sg13g2_nand2_1 _3043_ (.Y(_0774_),
    .A(_0759_),
    .B(_0766_));
 sg13g2_inv_1 _3044_ (.Y(_0775_),
    .A(_0774_));
 sg13g2_mux2_2 _3045_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][14] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][14] ),
    .S(net734),
    .X(_0776_));
 sg13g2_nand2_1 _3046_ (.Y(_0777_),
    .A(_0715_),
    .B(_0776_));
 sg13g2_xnor2_1 _3047_ (.Y(_0778_),
    .A(net590),
    .B(_0776_));
 sg13g2_inv_1 _3048_ (.Y(_0779_),
    .A(_0778_));
 sg13g2_nand3_1 _3049_ (.B(_0775_),
    .C(_0779_),
    .A(_0773_),
    .Y(_0780_));
 sg13g2_a21o_1 _3050_ (.A2(_0775_),
    .A1(_0773_),
    .B1(_0779_),
    .X(_0781_));
 sg13g2_and3_1 _3051_ (.X(_0782_),
    .A(net675),
    .B(_0780_),
    .C(_0781_));
 sg13g2_nor2b_1 _3052_ (.A(_0782_),
    .B_N(_0613_),
    .Y(_0783_));
 sg13g2_o21ai_1 _3053_ (.B1(net744),
    .Y(_0784_),
    .A1(net398),
    .A2(net680));
 sg13g2_nor2_1 _3054_ (.A(_0783_),
    .B(_0784_),
    .Y(_0088_));
 sg13g2_mux2_1 _3055_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][15] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][15] ),
    .S(net736),
    .X(_0785_));
 sg13g2_xor2_1 _3056_ (.B(_0785_),
    .A(net590),
    .X(_0786_));
 sg13g2_nand3_1 _3057_ (.B(_0781_),
    .C(_0786_),
    .A(_0777_),
    .Y(_0787_));
 sg13g2_a21o_1 _3058_ (.A2(_0781_),
    .A1(_0777_),
    .B1(_0786_),
    .X(_0788_));
 sg13g2_nand3_1 _3059_ (.B(_0787_),
    .C(_0788_),
    .A(net675),
    .Y(_0789_));
 sg13g2_o21ai_1 _3060_ (.B1(net770),
    .Y(_0790_),
    .A1(net515),
    .A2(net680));
 sg13g2_a21oi_1 _3061_ (.A1(net680),
    .A2(_0789_),
    .Y(_0089_),
    .B1(_0790_));
 sg13g2_and2_2 _3062_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[2] ),
    .B(_0448_),
    .X(_0791_));
 sg13g2_nand2_2 _3063_ (.Y(_0792_),
    .A(net722),
    .B(_0448_));
 sg13g2_nand2_1 _3064_ (.Y(_0793_),
    .A(\cpu_instance.mem_instance.mem_ctrl_instance.stall_txn ),
    .B(net713));
 sg13g2_a21oi_1 _3065_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.stall_txn ),
    .A2(net712),
    .Y(_0794_),
    .B1(\cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[0] ));
 sg13g2_nor2_2 _3066_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[1] ),
    .B(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[0] ),
    .Y(_0795_));
 sg13g2_nor3_2 _3067_ (.A(net500),
    .B(net561),
    .C(net810),
    .Y(_0796_));
 sg13g2_nand2b_2 _3068_ (.Y(_0797_),
    .B(_0795_),
    .A_N(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[2] ));
 sg13g2_and2_1 _3069_ (.A(_0025_),
    .B(net712),
    .X(_0798_));
 sg13g2_o21ai_1 _3070_ (.B1(net712),
    .Y(_0799_),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[1] ),
    .A2(_0025_));
 sg13g2_nor2_1 _3071_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[0] ),
    .B(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ),
    .Y(_0800_));
 sg13g2_nor2_1 _3072_ (.A(_0799_),
    .B(_0800_),
    .Y(_0801_));
 sg13g2_a21oi_2 _3073_ (.B1(_0801_),
    .Y(_0802_),
    .A2(_0799_),
    .A1(_0024_));
 sg13g2_nand2_1 _3074_ (.Y(_0803_),
    .A(_0796_),
    .B(_0802_));
 sg13g2_nand2_1 _3075_ (.Y(_0804_),
    .A(net722),
    .B(_0479_));
 sg13g2_a21oi_2 _3076_ (.B1(_0803_),
    .Y(_0805_),
    .A2(_0804_),
    .A1(_0793_));
 sg13g2_nand2b_1 _3077_ (.Y(_0806_),
    .B(_0805_),
    .A_N(_0794_));
 sg13g2_o21ai_1 _3078_ (.B1(_1306_),
    .Y(_0807_),
    .A1(_0803_),
    .A2(_0804_));
 sg13g2_a21oi_1 _3079_ (.A1(_0806_),
    .A2(_0807_),
    .Y(_0808_),
    .B1(_0791_));
 sg13g2_nor2_1 _3080_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ),
    .B(\cpu_instance.mem_instance.mem_ctrl_instance.stall_txn ),
    .Y(_0809_));
 sg13g2_nor2_1 _3081_ (.A(net720),
    .B(_0792_),
    .Y(_0810_));
 sg13g2_and2_1 _3082_ (.A(_0809_),
    .B(_0810_),
    .X(_0811_));
 sg13g2_nand2_2 _3083_ (.Y(_0812_),
    .A(_0475_),
    .B(_0481_));
 sg13g2_nor2_1 _3084_ (.A(_0792_),
    .B(_0809_),
    .Y(_0813_));
 sg13g2_nor3_1 _3085_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[0] ),
    .B(_0792_),
    .C(_0809_),
    .Y(_0814_));
 sg13g2_a21o_1 _3086_ (.A2(_0811_),
    .A1(net489),
    .B1(_0814_),
    .X(_0815_));
 sg13g2_nor3_1 _3087_ (.A(_0808_),
    .B(_0812_),
    .C(_0815_),
    .Y(_0816_));
 sg13g2_a21oi_1 _3088_ (.A1(_1306_),
    .A2(_0812_),
    .Y(_0090_),
    .B1(_0816_));
 sg13g2_nand2_1 _3089_ (.Y(_0817_),
    .A(net553),
    .B(_0805_));
 sg13g2_nand3b_1 _3090_ (.B(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ),
    .C(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[0] ),
    .Y(_0818_),
    .A_N(_0805_));
 sg13g2_nor2b_1 _3091_ (.A(_0812_),
    .B_N(_0818_),
    .Y(_0819_));
 sg13g2_a22oi_1 _3092_ (.Y(_0091_),
    .B1(_0817_),
    .B2(_0819_),
    .A2(_0812_),
    .A1(_1307_));
 sg13g2_nor3_1 _3093_ (.A(net720),
    .B(net849),
    .C(_0803_),
    .Y(_0820_));
 sg13g2_a21oi_1 _3094_ (.A1(net712),
    .A2(_0820_),
    .Y(_0821_),
    .B1(_0811_));
 sg13g2_nor2_1 _3095_ (.A(_0812_),
    .B(_0821_),
    .Y(_0092_));
 sg13g2_nor2_1 _3096_ (.A(net737),
    .B(\cpu_instance.mem_instance.qspi_ctrl_instance.last_ram_a_sel ),
    .Y(_0822_));
 sg13g2_nor2_1 _3097_ (.A(_0482_),
    .B(_0822_),
    .Y(_0823_));
 sg13g2_nor2_2 _3098_ (.A(_0481_),
    .B(_0823_),
    .Y(_0824_));
 sg13g2_nor2_2 _3099_ (.A(_0480_),
    .B(_0791_),
    .Y(_0825_));
 sg13g2_nand2b_1 _3100_ (.Y(_0826_),
    .B(_0825_),
    .A_N(_0802_));
 sg13g2_nand2b_2 _3101_ (.Y(_0827_),
    .B(_0826_),
    .A_N(_0824_));
 sg13g2_nand2_2 _3102_ (.Y(_0828_),
    .A(_0792_),
    .B(_0796_));
 sg13g2_or3_1 _3103_ (.A(_0023_),
    .B(net713),
    .C(_0828_),
    .X(_0829_));
 sg13g2_nor2_1 _3104_ (.A(net722),
    .B(_0829_),
    .Y(_0830_));
 sg13g2_nor3_2 _3105_ (.A(_0791_),
    .B(_0827_),
    .C(_0830_),
    .Y(_0831_));
 sg13g2_or3_1 _3106_ (.A(_0791_),
    .B(_0827_),
    .C(_0830_),
    .X(_0832_));
 sg13g2_nor2_1 _3107_ (.A(_0480_),
    .B(_0832_),
    .Y(_0833_));
 sg13g2_o21ai_1 _3108_ (.B1(_0475_),
    .Y(_0834_),
    .A1(net810),
    .A2(_0831_));
 sg13g2_a21oi_1 _3109_ (.A1(net810),
    .A2(_0833_),
    .Y(_0093_),
    .B1(_0834_));
 sg13g2_a21oi_1 _3110_ (.A1(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ),
    .A2(_1284_),
    .Y(_0835_),
    .B1(_0456_));
 sg13g2_nor3_1 _3111_ (.A(net713),
    .B(_0454_),
    .C(_0835_),
    .Y(_0836_));
 sg13g2_o21ai_1 _3112_ (.B1(_0795_),
    .Y(_0837_),
    .A1(net500),
    .A2(_0836_));
 sg13g2_nand2_1 _3113_ (.Y(_0838_),
    .A(net561),
    .B(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[0] ));
 sg13g2_nand2_1 _3114_ (.Y(_0839_),
    .A(_0837_),
    .B(_0838_));
 sg13g2_a22oi_1 _3115_ (.Y(_0840_),
    .B1(_0833_),
    .B2(_0839_),
    .A2(_0832_),
    .A1(net561));
 sg13g2_nor2_1 _3116_ (.A(_0476_),
    .B(net562),
    .Y(_0094_));
 sg13g2_o21ai_1 _3117_ (.B1(_0831_),
    .Y(_0841_),
    .A1(_0480_),
    .A2(_0795_));
 sg13g2_nor3_1 _3118_ (.A(net722),
    .B(_0444_),
    .C(_0797_),
    .Y(_0842_));
 sg13g2_a21o_1 _3119_ (.A2(_0480_),
    .A1(net737),
    .B1(_0842_),
    .X(_0843_));
 sg13g2_a22oi_1 _3120_ (.Y(_0844_),
    .B1(_0843_),
    .B2(_0831_),
    .A2(_0841_),
    .A1(net500));
 sg13g2_nor2_1 _3121_ (.A(_0476_),
    .B(_0844_),
    .Y(_0095_));
 sg13g2_nand3_1 _3122_ (.B(_0446_),
    .C(_0796_),
    .A(net720),
    .Y(_0845_));
 sg13g2_nor3_1 _3123_ (.A(_0476_),
    .B(_0802_),
    .C(_0845_),
    .Y(_0096_));
 sg13g2_and3_2 _3124_ (.X(_0846_),
    .A(_1306_),
    .B(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ),
    .C(_0810_));
 sg13g2_mux2_1 _3125_ (.A0(net332),
    .A1(net7),
    .S(_0846_),
    .X(_0097_));
 sg13g2_mux2_1 _3126_ (.A0(net366),
    .A1(net8),
    .S(_0846_),
    .X(_0098_));
 sg13g2_mux2_1 _3127_ (.A0(net368),
    .A1(net9),
    .S(_0846_),
    .X(_0099_));
 sg13g2_mux2_1 _3128_ (.A0(net345),
    .A1(net10),
    .S(_0846_),
    .X(_0100_));
 sg13g2_nand3_1 _3129_ (.B(_0802_),
    .C(_0825_),
    .A(_0797_),
    .Y(_0847_));
 sg13g2_a21oi_1 _3130_ (.A1(net723),
    .A2(net713),
    .Y(_0848_),
    .B1(_0847_));
 sg13g2_nor3_2 _3131_ (.A(_0813_),
    .B(_0827_),
    .C(_0848_),
    .Y(_0849_));
 sg13g2_a21oi_1 _3132_ (.A1(_0030_),
    .A2(_0456_),
    .Y(_0850_),
    .B1(_0835_));
 sg13g2_a21oi_1 _3133_ (.A1(_0029_),
    .A2(net712),
    .Y(_0851_),
    .B1(_0828_));
 sg13g2_inv_1 _3134_ (.Y(_0852_),
    .A(_0851_));
 sg13g2_o21ai_1 _3135_ (.B1(_0851_),
    .Y(_0853_),
    .A1(net713),
    .A2(_0850_));
 sg13g2_nand2_1 _3136_ (.Y(_0854_),
    .A(_0481_),
    .B(_0853_));
 sg13g2_o21ai_1 _3137_ (.B1(_0854_),
    .Y(_0855_),
    .A1(_1283_),
    .A2(_0481_));
 sg13g2_mux2_1 _3138_ (.A0(net724),
    .A1(_0855_),
    .S(_0849_),
    .X(_0856_));
 sg13g2_and2_1 _3139_ (.A(_0475_),
    .B(_0856_),
    .X(_0101_));
 sg13g2_o21ai_1 _3140_ (.B1(_0023_),
    .Y(_0857_),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ),
    .A2(net720));
 sg13g2_a221oi_1 _3141_ (.B2(_0857_),
    .C1(_0443_),
    .B1(_0448_),
    .A1(net722),
    .Y(_0858_),
    .A2(net724));
 sg13g2_nor2_1 _3142_ (.A(_0852_),
    .B(_0858_),
    .Y(_0859_));
 sg13g2_a221oi_1 _3143_ (.B2(net553),
    .C1(_0859_),
    .B1(_0810_),
    .A1(net737),
    .Y(_0860_),
    .A2(_0480_));
 sg13g2_o21ai_1 _3144_ (.B1(_0475_),
    .Y(_0861_),
    .A1(net723),
    .A2(_0849_));
 sg13g2_a21oi_1 _3145_ (.A1(_0849_),
    .A2(_0860_),
    .Y(_0102_),
    .B1(_0861_));
 sg13g2_a21oi_1 _3146_ (.A1(net723),
    .A2(net724),
    .Y(_0862_),
    .B1(_0023_));
 sg13g2_nor3_1 _3147_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ),
    .B(net720),
    .C(net724),
    .Y(_0863_));
 sg13g2_nor2_1 _3148_ (.A(_0454_),
    .B(_0863_),
    .Y(_0864_));
 sg13g2_nor4_1 _3149_ (.A(net713),
    .B(_0828_),
    .C(_0862_),
    .D(_0864_),
    .Y(_0865_));
 sg13g2_o21ai_1 _3150_ (.B1(_0849_),
    .Y(_0866_),
    .A1(_0480_),
    .A2(_0865_));
 sg13g2_o21ai_1 _3151_ (.B1(_0866_),
    .Y(_0867_),
    .A1(net722),
    .A2(_0849_));
 sg13g2_nor2_1 _3152_ (.A(_0476_),
    .B(_0867_),
    .Y(_0103_));
 sg13g2_nand2_2 _3153_ (.Y(_0868_),
    .A(_0480_),
    .B(_0823_));
 sg13g2_nor2_1 _3154_ (.A(net737),
    .B(net830),
    .Y(_0869_));
 sg13g2_o21ai_1 _3155_ (.B1(_0475_),
    .Y(_0870_),
    .A1(_0868_),
    .A2(_0869_));
 sg13g2_a21oi_1 _3156_ (.A1(_1284_),
    .A2(_0868_),
    .Y(_0104_),
    .B1(_0870_));
 sg13g2_a22oi_1 _3157_ (.Y(_0871_),
    .B1(_0868_),
    .B2(net354),
    .A2(_0483_),
    .A1(net737));
 sg13g2_nand2_1 _3158_ (.Y(_0105_),
    .A(_0475_),
    .B(_0871_));
 sg13g2_a21oi_1 _3159_ (.A1(net834),
    .A2(_0868_),
    .Y(_0872_),
    .B1(_0476_));
 sg13g2_o21ai_1 _3160_ (.B1(_0872_),
    .Y(_0106_),
    .A1(_1283_),
    .A2(_0868_));
 sg13g2_nor2_1 _3161_ (.A(net789),
    .B(_0825_),
    .Y(_0873_));
 sg13g2_nor2b_1 _3162_ (.A(_0824_),
    .B_N(net789),
    .Y(_0874_));
 sg13g2_nor3_1 _3163_ (.A(_0476_),
    .B(_0873_),
    .C(_0874_),
    .Y(_0107_));
 sg13g2_o21ai_1 _3164_ (.B1(_0025_),
    .Y(_0875_),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ),
    .A2(net720));
 sg13g2_a21oi_1 _3165_ (.A1(_0455_),
    .A2(_0875_),
    .Y(_0876_),
    .B1(net712));
 sg13g2_nor2_1 _3166_ (.A(_0828_),
    .B(_0876_),
    .Y(_0877_));
 sg13g2_o21ai_1 _3167_ (.B1(_0802_),
    .Y(_0878_),
    .A1(_0842_),
    .A2(_0877_));
 sg13g2_and3_1 _3168_ (.X(_0879_),
    .A(_0829_),
    .B(_0847_),
    .C(_0878_));
 sg13g2_a21oi_1 _3169_ (.A1(_0831_),
    .A2(_0879_),
    .Y(_0880_),
    .B1(net322));
 sg13g2_a21oi_1 _3170_ (.A1(_0833_),
    .A2(_0879_),
    .Y(_0881_),
    .B1(_0476_));
 sg13g2_nor2b_1 _3171_ (.A(_0880_),
    .B_N(_0881_),
    .Y(_0108_));
 sg13g2_and2_2 _3172_ (.A(_0446_),
    .B(_0800_),
    .X(_0882_));
 sg13g2_mux2_1 _3173_ (.A0(net332),
    .A1(net7),
    .S(_0882_),
    .X(_0883_));
 sg13g2_nor2_2 _3174_ (.A(_0791_),
    .B(_0796_),
    .Y(_0884_));
 sg13g2_nand2_2 _3175_ (.Y(_0885_),
    .A(_0792_),
    .B(_0797_));
 sg13g2_o21ai_1 _3176_ (.B1(net721),
    .Y(_0886_),
    .A1(net373),
    .A2(_0884_));
 sg13g2_inv_1 _3177_ (.Y(_0887_),
    .A(_0886_));
 sg13g2_o21ai_1 _3178_ (.B1(_0887_),
    .Y(_0888_),
    .A1(net7),
    .A2(_0885_));
 sg13g2_nand3_1 _3179_ (.B(_0447_),
    .C(_0884_),
    .A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_clk_out ),
    .Y(_0889_));
 sg13g2_a21oi_1 _3180_ (.A1(_0024_),
    .A2(_0792_),
    .Y(_0890_),
    .B1(_0025_));
 sg13g2_a22oi_1 _3181_ (.Y(_0891_),
    .B1(_0889_),
    .B2(_0890_),
    .A2(_0800_),
    .A1(_0798_));
 sg13g2_a21oi_1 _3182_ (.A1(_1284_),
    .A2(_0883_),
    .Y(_0892_),
    .B1(net669));
 sg13g2_a22oi_1 _3183_ (.Y(_0109_),
    .B1(_0892_),
    .B2(_0888_),
    .A2(net669),
    .A1(_1314_));
 sg13g2_nand2b_1 _3184_ (.Y(_0893_),
    .B(net366),
    .A_N(_0882_));
 sg13g2_a21oi_1 _3185_ (.A1(net8),
    .A2(_0882_),
    .Y(_0894_),
    .B1(net721));
 sg13g2_nand2_1 _3186_ (.Y(_0895_),
    .A(net357),
    .B(_0885_));
 sg13g2_a21oi_1 _3187_ (.A1(net8),
    .A2(_0884_),
    .Y(_0896_),
    .B1(_1284_));
 sg13g2_a22oi_1 _3188_ (.Y(_0897_),
    .B1(_0895_),
    .B2(_0896_),
    .A2(_0894_),
    .A1(_0893_));
 sg13g2_mux2_1 _3189_ (.A0(_0897_),
    .A1(net535),
    .S(net669),
    .X(_0110_));
 sg13g2_nand2b_1 _3190_ (.Y(_0898_),
    .B(net368),
    .A_N(_0882_));
 sg13g2_a21oi_1 _3191_ (.A1(net9),
    .A2(_0882_),
    .Y(_0899_),
    .B1(net721));
 sg13g2_nand2_1 _3192_ (.Y(_0900_),
    .A(net358),
    .B(_0885_));
 sg13g2_a21oi_1 _3193_ (.A1(net9),
    .A2(_0884_),
    .Y(_0901_),
    .B1(_1284_));
 sg13g2_a22oi_1 _3194_ (.Y(_0902_),
    .B1(_0900_),
    .B2(_0901_),
    .A2(_0899_),
    .A1(_0898_));
 sg13g2_mux2_1 _3195_ (.A0(_0902_),
    .A1(net545),
    .S(net669),
    .X(_0111_));
 sg13g2_nand2b_1 _3196_ (.Y(_0903_),
    .B(net345),
    .A_N(_0882_));
 sg13g2_a21oi_1 _3197_ (.A1(net10),
    .A2(_0882_),
    .Y(_0904_),
    .B1(net720));
 sg13g2_nand2_1 _3198_ (.Y(_0905_),
    .A(net342),
    .B(_0885_));
 sg13g2_a21oi_1 _3199_ (.A1(net10),
    .A2(_0884_),
    .Y(_0906_),
    .B1(_1284_));
 sg13g2_a22oi_1 _3200_ (.Y(_0907_),
    .B1(_0905_),
    .B2(_0906_),
    .A2(_0904_),
    .A1(_0903_));
 sg13g2_mux2_1 _3201_ (.A0(_0907_),
    .A1(net503),
    .S(net669),
    .X(_0112_));
 sg13g2_nor2_2 _3202_ (.A(_1284_),
    .B(_0884_),
    .Y(_0908_));
 sg13g2_nor2b_1 _3203_ (.A(_0908_),
    .B_N(net387),
    .Y(_0909_));
 sg13g2_a21oi_1 _3204_ (.A1(net351),
    .A2(_0908_),
    .Y(_0910_),
    .B1(_0909_));
 sg13g2_nand2_1 _3205_ (.Y(_0911_),
    .A(net399),
    .B(net668));
 sg13g2_o21ai_1 _3206_ (.B1(_0911_),
    .Y(_0113_),
    .A1(net668),
    .A2(_0910_));
 sg13g2_nor2b_1 _3207_ (.A(_0908_),
    .B_N(\cpu_instance.mem_instance.data_qo_mi[1] ),
    .Y(_0912_));
 sg13g2_a21oi_1 _3208_ (.A1(net339),
    .A2(_0908_),
    .Y(_0913_),
    .B1(_0912_));
 sg13g2_nand2_1 _3209_ (.Y(_0914_),
    .A(net377),
    .B(net668));
 sg13g2_o21ai_1 _3210_ (.B1(_0914_),
    .Y(_0114_),
    .A1(net668),
    .A2(_0913_));
 sg13g2_mux2_1 _3211_ (.A0(\cpu_instance.mem_instance.data_qo_mi[2] ),
    .A1(net349),
    .S(_0908_),
    .X(_0915_));
 sg13g2_nor2_1 _3212_ (.A(net668),
    .B(_0915_),
    .Y(_0916_));
 sg13g2_a21oi_1 _3213_ (.A1(_1315_),
    .A2(net668),
    .Y(_0115_),
    .B1(_0916_));
 sg13g2_nor2b_1 _3214_ (.A(_0908_),
    .B_N(\cpu_instance.mem_instance.data_qo_mi[3] ),
    .Y(_0917_));
 sg13g2_a21oi_1 _3215_ (.A1(net363),
    .A2(_0908_),
    .Y(_0918_),
    .B1(_0917_));
 sg13g2_nand2_1 _3216_ (.Y(_0919_),
    .A(net371),
    .B(net668));
 sg13g2_o21ai_1 _3217_ (.B1(_0919_),
    .Y(_0116_),
    .A1(net668),
    .A2(_0918_));
 sg13g2_nand2b_1 _3218_ (.Y(_0117_),
    .B(net771),
    .A_N(net354));
 sg13g2_mux2_1 _3219_ (.A0(net7),
    .A1(net489),
    .S(net771),
    .X(_0118_));
 sg13g2_mux2_1 _3220_ (.A0(net8),
    .A1(net553),
    .S(net771),
    .X(_0119_));
 sg13g2_a22oi_1 _3221_ (.Y(_0920_),
    .B1(net711),
    .B2(net687),
    .A2(net685),
    .A1(net337));
 sg13g2_inv_1 _3222_ (.Y(_0120_),
    .A(_0920_));
 sg13g2_a22oi_1 _3223_ (.Y(_0921_),
    .B1(net707),
    .B2(net688),
    .A2(net685),
    .A1(net348));
 sg13g2_inv_1 _3224_ (.Y(_0121_),
    .A(_0921_));
 sg13g2_a22oi_1 _3225_ (.Y(_0922_),
    .B1(_0639_),
    .B2(net688),
    .A2(net684),
    .A1(net338));
 sg13g2_inv_1 _3226_ (.Y(_0122_),
    .A(_0922_));
 sg13g2_a22oi_1 _3227_ (.Y(_0923_),
    .B1(net362),
    .B2(net687),
    .A2(net684),
    .A1(net352));
 sg13g2_inv_1 _3228_ (.Y(_0123_),
    .A(_0923_));
 sg13g2_nor2_1 _3229_ (.A(net337),
    .B(_0478_),
    .Y(_0924_));
 sg13g2_a221oi_1 _3230_ (.B2(net687),
    .C1(_0924_),
    .B1(_0667_),
    .A1(_1308_),
    .Y(_0124_),
    .A2(net684));
 sg13g2_nor2_1 _3231_ (.A(net348),
    .B(net689),
    .Y(_0925_));
 sg13g2_a221oi_1 _3232_ (.B2(net688),
    .C1(_0925_),
    .B1(_0680_),
    .A1(_1309_),
    .Y(_0125_),
    .A2(net684));
 sg13g2_nor2_1 _3233_ (.A(net374),
    .B(_0486_),
    .Y(_0926_));
 sg13g2_nor2_1 _3234_ (.A(net338),
    .B(net689),
    .Y(_0927_));
 sg13g2_nor2_1 _3235_ (.A(_0484_),
    .B(_0691_),
    .Y(_0928_));
 sg13g2_nor3_1 _3236_ (.A(_0926_),
    .B(_0927_),
    .C(_0928_),
    .Y(_0126_));
 sg13g2_nor2_1 _3237_ (.A(net352),
    .B(net689),
    .Y(_0929_));
 sg13g2_a221oi_1 _3238_ (.B2(net687),
    .C1(_0929_),
    .B1(_0706_),
    .A1(_1310_),
    .Y(_0127_),
    .A2(net684));
 sg13g2_nor2_1 _3239_ (.A(net364),
    .B(net689),
    .Y(_0930_));
 sg13g2_a221oi_1 _3240_ (.B2(net687),
    .C1(_0930_),
    .B1(_0718_),
    .A1(_1311_),
    .Y(_0128_),
    .A2(net684));
 sg13g2_nor2_1 _3241_ (.A(_0484_),
    .B(_0728_),
    .Y(_0931_));
 sg13g2_a221oi_1 _3242_ (.B2(_1312_),
    .C1(_0931_),
    .B1(net684),
    .A1(_1309_),
    .Y(_0129_),
    .A2(net690));
 sg13g2_nor2_1 _3243_ (.A(net346),
    .B(_0486_),
    .Y(_0932_));
 sg13g2_nor2_1 _3244_ (.A(net374),
    .B(net689),
    .Y(_0933_));
 sg13g2_nor2_1 _3245_ (.A(_0484_),
    .B(_0736_),
    .Y(_0934_));
 sg13g2_nor3_1 _3246_ (.A(_0932_),
    .B(_0933_),
    .C(_0934_),
    .Y(_0130_));
 sg13g2_nor2_1 _3247_ (.A(net382),
    .B(net689),
    .Y(_0935_));
 sg13g2_a221oi_1 _3248_ (.B2(net687),
    .C1(_0935_),
    .B1(_0747_),
    .A1(_1313_),
    .Y(_0131_),
    .A2(net684));
 sg13g2_or2_1 _3249_ (.X(_0936_),
    .B(_0758_),
    .A(_0484_));
 sg13g2_o21ai_1 _3250_ (.B1(_0936_),
    .Y(_0937_),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[12] ),
    .A2(_0486_));
 sg13g2_a21oi_1 _3251_ (.A1(_1311_),
    .A2(net690),
    .Y(_0132_),
    .B1(_0937_));
 sg13g2_nand2b_1 _3252_ (.Y(_0938_),
    .B(net687),
    .A_N(_0765_));
 sg13g2_o21ai_1 _3253_ (.B1(_0938_),
    .Y(_0939_),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[13] ),
    .A2(_0486_));
 sg13g2_a21oi_1 _3254_ (.A1(_1312_),
    .A2(net690),
    .Y(_0133_),
    .B1(_0939_));
 sg13g2_nor2_1 _3255_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[14] ),
    .B(_0486_),
    .Y(_0940_));
 sg13g2_nor2_1 _3256_ (.A(_0484_),
    .B(_0776_),
    .Y(_0941_));
 sg13g2_nor2_1 _3257_ (.A(net346),
    .B(net689),
    .Y(_0942_));
 sg13g2_nor3_1 _3258_ (.A(_0940_),
    .B(_0941_),
    .C(_0942_),
    .Y(_0134_));
 sg13g2_nand2b_1 _3259_ (.Y(_0943_),
    .B(net687),
    .A_N(_0785_));
 sg13g2_o21ai_1 _3260_ (.B1(_0943_),
    .Y(_0944_),
    .A1(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[15] ),
    .A2(_0486_));
 sg13g2_a21oi_1 _3261_ (.A1(_1313_),
    .A2(net690),
    .Y(_0135_),
    .B1(_0944_));
 sg13g2_nor2_1 _3262_ (.A(net736),
    .B(_0605_),
    .Y(_0945_));
 sg13g2_a221oi_1 _3263_ (.B2(\cpu_instance.mem_instance.addr[24] ),
    .C1(_0945_),
    .B1(_0612_),
    .A1(_0605_),
    .Y(_0946_),
    .A2(_0610_));
 sg13g2_o21ai_1 _3264_ (.B1(net745),
    .Y(_0947_),
    .A1(net426),
    .A2(net672));
 sg13g2_a21oi_1 _3265_ (.A1(_0622_),
    .A2(net672),
    .Y(_0136_),
    .B1(_0947_));
 sg13g2_o21ai_1 _3266_ (.B1(net745),
    .Y(_0948_),
    .A1(net493),
    .A2(net672));
 sg13g2_a21oi_1 _3267_ (.A1(_0634_),
    .A2(net672),
    .Y(_0137_),
    .B1(_0948_));
 sg13g2_o21ai_1 _3268_ (.B1(net745),
    .Y(_0949_),
    .A1(net520),
    .A2(net672));
 sg13g2_a21oi_1 _3269_ (.A1(_0646_),
    .A2(net672),
    .Y(_0138_),
    .B1(_0949_));
 sg13g2_o21ai_1 _3270_ (.B1(net746),
    .Y(_0950_),
    .A1(net518),
    .A2(net672));
 sg13g2_a21oi_1 _3271_ (.A1(_0659_),
    .A2(net672),
    .Y(_0139_),
    .B1(_0950_));
 sg13g2_o21ai_1 _3272_ (.B1(net769),
    .Y(_0951_),
    .A1(net565),
    .A2(net674));
 sg13g2_a21oi_1 _3273_ (.A1(_0672_),
    .A2(net674),
    .Y(_0140_),
    .B1(_0951_));
 sg13g2_o21ai_1 _3274_ (.B1(net746),
    .Y(_0952_),
    .A1(net427),
    .A2(net674));
 sg13g2_a21oi_1 _3275_ (.A1(_0685_),
    .A2(net674),
    .Y(_0141_),
    .B1(_0952_));
 sg13g2_o21ai_1 _3276_ (.B1(net745),
    .Y(_0953_),
    .A1(net530),
    .A2(net673));
 sg13g2_a21oi_1 _3277_ (.A1(_0700_),
    .A2(net673),
    .Y(_0142_),
    .B1(_0953_));
 sg13g2_o21ai_1 _3278_ (.B1(net746),
    .Y(_0954_),
    .A1(net542),
    .A2(net673));
 sg13g2_a21oi_1 _3279_ (.A1(_0713_),
    .A2(net673),
    .Y(_0143_),
    .B1(_0954_));
 sg13g2_o21ai_1 _3280_ (.B1(net743),
    .Y(_0955_),
    .A1(net468),
    .A2(net673));
 sg13g2_a21oi_1 _3281_ (.A1(_0724_),
    .A2(net670),
    .Y(_0144_),
    .B1(_0955_));
 sg13g2_o21ai_1 _3282_ (.B1(net743),
    .Y(_0956_),
    .A1(net492),
    .A2(net671));
 sg13g2_a21oi_1 _3283_ (.A1(_0734_),
    .A2(net670),
    .Y(_0145_),
    .B1(_0956_));
 sg13g2_o21ai_1 _3284_ (.B1(net743),
    .Y(_0957_),
    .A1(net577),
    .A2(net670));
 sg13g2_a21oi_1 _3285_ (.A1(_0744_),
    .A2(net670),
    .Y(_0146_),
    .B1(_0957_));
 sg13g2_o21ai_1 _3286_ (.B1(net743),
    .Y(_0958_),
    .A1(net458),
    .A2(net670));
 sg13g2_a21oi_1 _3287_ (.A1(_0752_),
    .A2(net670),
    .Y(_0147_),
    .B1(_0958_));
 sg13g2_o21ai_1 _3288_ (.B1(net744),
    .Y(_0959_),
    .A1(net477),
    .A2(net670));
 sg13g2_a21oi_1 _3289_ (.A1(_0763_),
    .A2(net670),
    .Y(_0148_),
    .B1(_0959_));
 sg13g2_o21ai_1 _3290_ (.B1(net744),
    .Y(_0960_),
    .A1(net510),
    .A2(net671));
 sg13g2_a21oi_1 _3291_ (.A1(_0770_),
    .A2(net671),
    .Y(_0149_),
    .B1(_0960_));
 sg13g2_nor2b_1 _3292_ (.A(_0782_),
    .B_N(net671),
    .Y(_0961_));
 sg13g2_o21ai_1 _3293_ (.B1(net744),
    .Y(_0962_),
    .A1(net541),
    .A2(net671));
 sg13g2_nor2_1 _3294_ (.A(_0961_),
    .B(_0962_),
    .Y(_0150_));
 sg13g2_o21ai_1 _3295_ (.B1(net770),
    .Y(_0963_),
    .A1(net568),
    .A2(net671));
 sg13g2_a21oi_1 _3296_ (.A1(_0789_),
    .A2(net671),
    .Y(_0151_),
    .B1(_0963_));
 sg13g2_nor2_1 _3297_ (.A(net600),
    .B(_0576_),
    .Y(_0152_));
 sg13g2_nor2_1 _3298_ (.A(net595),
    .B(_0576_),
    .Y(_0153_));
 sg13g2_nand2_2 _3299_ (.Y(_0964_),
    .A(net708),
    .B(net707));
 sg13g2_nand3_1 _3300_ (.B(net707),
    .C(_0639_),
    .A(net711),
    .Y(_0965_));
 sg13g2_and4_1 _3301_ (.A(net711),
    .B(net707),
    .C(_0639_),
    .D(_0652_),
    .X(_0966_));
 sg13g2_nand4_1 _3302_ (.B(_0679_),
    .C(_0691_),
    .A(_0666_),
    .Y(_0967_),
    .D(_0966_));
 sg13g2_xnor2_1 _3303_ (.Y(_0968_),
    .A(_0705_),
    .B(_0967_));
 sg13g2_xor2_1 _3304_ (.B(_0965_),
    .A(_0652_),
    .X(_0969_));
 sg13g2_nor4_1 _3305_ (.A(_0652_),
    .B(_0666_),
    .C(_0679_),
    .D(_0691_),
    .Y(_0970_));
 sg13g2_nand2b_1 _3306_ (.Y(_0971_),
    .B(_0705_),
    .A_N(_0970_));
 sg13g2_nor3_1 _3307_ (.A(_0765_),
    .B(_0776_),
    .C(_0785_),
    .Y(_0972_));
 sg13g2_nor2b_1 _3308_ (.A(\cpu_instance.mem_instance.addr[24] ),
    .B_N(\cpu_instance.ctrl_instance.mem_ctrl_op[2] ),
    .Y(_0973_));
 sg13g2_nor4_1 _3309_ (.A(_0728_),
    .B(_0736_),
    .C(_0746_),
    .D(_0758_),
    .Y(_0974_));
 sg13g2_and4_1 _3310_ (.A(_0718_),
    .B(_0972_),
    .C(_0973_),
    .D(_0974_),
    .X(_0975_));
 sg13g2_nand4_1 _3311_ (.B(_0969_),
    .C(_0971_),
    .A(_0968_),
    .Y(_0976_),
    .D(_0975_));
 sg13g2_inv_1 _3312_ (.Y(_0977_),
    .A(_0976_));
 sg13g2_nor3_2 _3313_ (.A(net557),
    .B(net819),
    .C(\cpu_instance.mem_instance.mem_ctrl_instance.state[2] ),
    .Y(_0978_));
 sg13g2_a21oi_1 _3314_ (.A1(_1302_),
    .A2(_0420_),
    .Y(_0979_),
    .B1(_0978_));
 sg13g2_o21ai_1 _3315_ (.B1(_0979_),
    .Y(_0980_),
    .A1(_0417_),
    .A2(_0462_));
 sg13g2_nand2_1 _3316_ (.Y(_0981_),
    .A(_0336_),
    .B(_0980_));
 sg13g2_o21ai_1 _3317_ (.B1(_0416_),
    .Y(_0982_),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.state[1] ),
    .A2(_0418_));
 sg13g2_nand2_1 _3318_ (.Y(_0983_),
    .A(_0426_),
    .B(_0982_));
 sg13g2_nand2b_1 _3319_ (.Y(_0984_),
    .B(_0422_),
    .A_N(_0335_));
 sg13g2_a22oi_1 _3320_ (.Y(_0985_),
    .B1(_0984_),
    .B2(_0978_),
    .A2(_0983_),
    .A1(_0335_));
 sg13g2_and3_1 _3321_ (.X(_0986_),
    .A(_0428_),
    .B(_0981_),
    .C(_0985_));
 sg13g2_nand2_1 _3322_ (.Y(_0987_),
    .A(\cpu_instance.mem_instance.data_ready ),
    .B(_0985_));
 sg13g2_a21oi_1 _3323_ (.A1(_0428_),
    .A2(_0981_),
    .Y(_0988_),
    .B1(_0987_));
 sg13g2_nor3_1 _3324_ (.A(_0977_),
    .B(_0986_),
    .C(net630),
    .Y(_0989_));
 sg13g2_inv_2 _3325_ (.Y(_0990_),
    .A(net628));
 sg13g2_a21oi_1 _3326_ (.A1(net387),
    .A2(net630),
    .Y(_0991_),
    .B1(net628));
 sg13g2_xnor2_1 _3327_ (.Y(_0992_),
    .A(_0639_),
    .B(_0964_));
 sg13g2_xor2_1 _3328_ (.B(_0964_),
    .A(_0639_),
    .X(_0993_));
 sg13g2_mux2_1 _3329_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[7] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[6] ),
    .S(net709),
    .X(_0994_));
 sg13g2_xnor2_1 _3330_ (.Y(_0995_),
    .A(net708),
    .B(net707));
 sg13g2_nor2b_1 _3331_ (.A(_0995_),
    .B_N(_0968_),
    .Y(_0996_));
 sg13g2_inv_1 _3332_ (.Y(_0997_),
    .A(_0996_));
 sg13g2_and2_1 _3333_ (.A(_0968_),
    .B(_0995_),
    .X(_0998_));
 sg13g2_inv_1 _3334_ (.Y(_0999_),
    .A(net666));
 sg13g2_mux2_1 _3335_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[5] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[4] ),
    .S(net709),
    .X(_1000_));
 sg13g2_and2_1 _3336_ (.A(_0998_),
    .B(_1000_),
    .X(_1001_));
 sg13g2_a21o_1 _3337_ (.A2(_0996_),
    .A1(_0994_),
    .B1(_1001_),
    .X(_1002_));
 sg13g2_nor2_2 _3338_ (.A(_0976_),
    .B(net631),
    .Y(_1003_));
 sg13g2_mux2_1 _3339_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[3] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[2] ),
    .S(net708),
    .X(_1004_));
 sg13g2_nor2_1 _3340_ (.A(_0995_),
    .B(_1004_),
    .Y(_1005_));
 sg13g2_nor2_1 _3341_ (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[0] ),
    .B(_0964_),
    .Y(_1006_));
 sg13g2_nor3_1 _3342_ (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[1] ),
    .B(net708),
    .C(net707),
    .Y(_1007_));
 sg13g2_nor3_1 _3343_ (.A(_1005_),
    .B(_1006_),
    .C(_1007_),
    .Y(_1008_));
 sg13g2_a21oi_1 _3344_ (.A1(_0968_),
    .A2(_1008_),
    .Y(_1009_),
    .B1(_0992_));
 sg13g2_nor3_1 _3345_ (.A(_0976_),
    .B(net631),
    .C(_1009_),
    .Y(_1010_));
 sg13g2_o21ai_1 _3346_ (.B1(_1010_),
    .Y(_1011_),
    .A1(_0993_),
    .A2(_1002_));
 sg13g2_o21ai_1 _3347_ (.B1(net777),
    .Y(_1012_),
    .A1(net588),
    .A2(_0990_));
 sg13g2_a21oi_1 _3348_ (.A1(_0991_),
    .A2(_1011_),
    .Y(_0154_),
    .B1(_1012_));
 sg13g2_a21oi_1 _3349_ (.A1(net535),
    .A2(net630),
    .Y(_1013_),
    .B1(net628));
 sg13g2_mux2_1 _3350_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[6] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[5] ),
    .S(net709),
    .X(_1014_));
 sg13g2_nand2_1 _3351_ (.Y(_1015_),
    .A(net666),
    .B(_1014_));
 sg13g2_nor2b_1 _3352_ (.A(net708),
    .B_N(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[8] ),
    .Y(_1016_));
 sg13g2_a21oi_1 _3353_ (.A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[7] ),
    .A2(net708),
    .Y(_1017_),
    .B1(_1016_));
 sg13g2_o21ai_1 _3354_ (.B1(_1015_),
    .Y(_1018_),
    .A1(_0997_),
    .A2(_1017_));
 sg13g2_mux2_1 _3355_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[4] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[3] ),
    .S(net708),
    .X(_1019_));
 sg13g2_nor2_1 _3356_ (.A(_0995_),
    .B(_1019_),
    .Y(_1020_));
 sg13g2_nor2_1 _3357_ (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[1] ),
    .B(_0964_),
    .Y(_1021_));
 sg13g2_nor3_1 _3358_ (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[2] ),
    .B(net708),
    .C(net707),
    .Y(_1022_));
 sg13g2_nor3_1 _3359_ (.A(_1020_),
    .B(_1021_),
    .C(_1022_),
    .Y(_1023_));
 sg13g2_a21oi_1 _3360_ (.A1(_0968_),
    .A2(_1023_),
    .Y(_1024_),
    .B1(_0992_));
 sg13g2_nor3_1 _3361_ (.A(_0976_),
    .B(net631),
    .C(_1024_),
    .Y(_1025_));
 sg13g2_o21ai_1 _3362_ (.B1(_1025_),
    .Y(_1026_),
    .A1(_0993_),
    .A2(_1018_));
 sg13g2_o21ai_1 _3363_ (.B1(net777),
    .Y(_1027_),
    .A1(net782),
    .A2(_0990_));
 sg13g2_a21oi_1 _3364_ (.A1(_1013_),
    .A2(_1026_),
    .Y(_0155_),
    .B1(_1027_));
 sg13g2_a21oi_1 _3365_ (.A1(net545),
    .A2(net630),
    .Y(_1028_),
    .B1(net628));
 sg13g2_a221oi_1 _3366_ (.B2(net666),
    .C1(_0992_),
    .B1(_1004_),
    .A1(net667),
    .Y(_1029_),
    .A2(_1000_));
 sg13g2_mux2_1 _3367_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[9] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[8] ),
    .S(net710),
    .X(_1030_));
 sg13g2_a22oi_1 _3368_ (.Y(_1031_),
    .B1(_1030_),
    .B2(net667),
    .A2(_0998_),
    .A1(_0994_));
 sg13g2_nand2_1 _3369_ (.Y(_1032_),
    .A(_0992_),
    .B(_1031_));
 sg13g2_nand3b_1 _3370_ (.B(_1032_),
    .C(_1003_),
    .Y(_1033_),
    .A_N(_1029_));
 sg13g2_o21ai_1 _3371_ (.B1(net777),
    .Y(_1034_),
    .A1(net574),
    .A2(_0990_));
 sg13g2_a21oi_1 _3372_ (.A1(_1028_),
    .A2(_1033_),
    .Y(_0156_),
    .B1(_1034_));
 sg13g2_a21oi_1 _3373_ (.A1(net503),
    .A2(net630),
    .Y(_1035_),
    .B1(net628));
 sg13g2_a221oi_1 _3374_ (.B2(net666),
    .C1(_0992_),
    .B1(_1019_),
    .A1(net667),
    .Y(_1036_),
    .A2(_1014_));
 sg13g2_mux2_1 _3375_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[10] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[9] ),
    .S(net710),
    .X(_1037_));
 sg13g2_nand2_1 _3376_ (.Y(_1038_),
    .A(net667),
    .B(_1037_));
 sg13g2_o21ai_1 _3377_ (.B1(_1038_),
    .Y(_1039_),
    .A1(_0999_),
    .A2(_1017_));
 sg13g2_o21ai_1 _3378_ (.B1(_1003_),
    .Y(_1040_),
    .A1(_0993_),
    .A2(_1039_));
 sg13g2_o21ai_1 _3379_ (.B1(_1035_),
    .Y(_1041_),
    .A1(_1036_),
    .A2(_1040_));
 sg13g2_o21ai_1 _3380_ (.B1(net776),
    .Y(_1042_),
    .A1(net572),
    .A2(_0990_));
 sg13g2_nor2b_1 _3381_ (.A(_1042_),
    .B_N(_1041_),
    .Y(_0157_));
 sg13g2_a21oi_1 _3382_ (.A1(net399),
    .A2(net630),
    .Y(_1043_),
    .B1(net628));
 sg13g2_mux2_1 _3383_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[11] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[10] ),
    .S(net710),
    .X(_1044_));
 sg13g2_a221oi_1 _3384_ (.B2(net667),
    .C1(_0993_),
    .B1(_1044_),
    .A1(net666),
    .Y(_1045_),
    .A2(_1030_));
 sg13g2_nor3_1 _3385_ (.A(_0976_),
    .B(net631),
    .C(_1045_),
    .Y(_1046_));
 sg13g2_o21ai_1 _3386_ (.B1(_1046_),
    .Y(_1047_),
    .A1(_0992_),
    .A2(_1002_));
 sg13g2_o21ai_1 _3387_ (.B1(net776),
    .Y(_1048_),
    .A1(net564),
    .A2(_0990_));
 sg13g2_a21oi_1 _3388_ (.A1(_1043_),
    .A2(_1047_),
    .Y(_0158_),
    .B1(_1048_));
 sg13g2_a21oi_1 _3389_ (.A1(net377),
    .A2(net630),
    .Y(_1049_),
    .B1(net628));
 sg13g2_mux2_1 _3390_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[12] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[11] ),
    .S(net710),
    .X(_1050_));
 sg13g2_a221oi_1 _3391_ (.B2(net667),
    .C1(_0993_),
    .B1(_1050_),
    .A1(net666),
    .Y(_1051_),
    .A2(_1037_));
 sg13g2_o21ai_1 _3392_ (.B1(_1003_),
    .Y(_1052_),
    .A1(_0992_),
    .A2(_1018_));
 sg13g2_o21ai_1 _3393_ (.B1(_1049_),
    .Y(_1053_),
    .A1(_1051_),
    .A2(_1052_));
 sg13g2_o21ai_1 _3394_ (.B1(net777),
    .Y(_1054_),
    .A1(net496),
    .A2(_0990_));
 sg13g2_nor2b_1 _3395_ (.A(_1054_),
    .B_N(_1053_),
    .Y(_0159_));
 sg13g2_mux2_1 _3396_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[13] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[12] ),
    .S(net710),
    .X(_1055_));
 sg13g2_a221oi_1 _3397_ (.B2(net667),
    .C1(_0993_),
    .B1(_1055_),
    .A1(net666),
    .Y(_1056_),
    .A2(_1044_));
 sg13g2_a21oi_2 _3398_ (.B1(_1056_),
    .Y(_1057_),
    .A2(_1031_),
    .A1(_0993_));
 sg13g2_a221oi_1 _3399_ (.B2(_1057_),
    .C1(_0989_),
    .B1(_1003_),
    .A1(net461),
    .Y(_1058_),
    .A2(net631));
 sg13g2_o21ai_1 _3400_ (.B1(net777),
    .Y(_1059_),
    .A1(net466),
    .A2(_0990_));
 sg13g2_nor2_1 _3401_ (.A(_1058_),
    .B(_1059_),
    .Y(_0160_));
 sg13g2_a21oi_1 _3402_ (.A1(net371),
    .A2(net630),
    .Y(_1060_),
    .B1(net628));
 sg13g2_mux2_1 _3403_ (.A0(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[14] ),
    .A1(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[13] ),
    .S(net710),
    .X(_1061_));
 sg13g2_a221oi_1 _3404_ (.B2(net667),
    .C1(_0993_),
    .B1(_1061_),
    .A1(net666),
    .Y(_1062_),
    .A2(_1050_));
 sg13g2_nor3_1 _3405_ (.A(_0976_),
    .B(net631),
    .C(_1062_),
    .Y(_1063_));
 sg13g2_o21ai_1 _3406_ (.B1(_1063_),
    .Y(_1064_),
    .A1(_0992_),
    .A2(_1039_));
 sg13g2_o21ai_1 _3407_ (.B1(net776),
    .Y(_1065_),
    .A1(net429),
    .A2(_0990_));
 sg13g2_a21oi_1 _3408_ (.A1(_1060_),
    .A2(_1064_),
    .Y(_0161_),
    .B1(_1065_));
 sg13g2_and3_1 _3409_ (.X(_0162_),
    .A(net770),
    .B(net825),
    .C(_0978_));
 sg13g2_nor3_1 _3410_ (.A(\cpu_instance.ctrl_instance.mem_ctrl_op[0] ),
    .B(_1305_),
    .C(\cpu_instance.ctrl_instance.mem_ctrl_op[2] ),
    .Y(_1066_));
 sg13g2_a21oi_1 _3411_ (.A1(net557),
    .A2(_1066_),
    .Y(_1067_),
    .B1(_0978_));
 sg13g2_a221oi_1 _3412_ (.B2(net828),
    .C1(net740),
    .B1(_1067_),
    .A1(_0976_),
    .Y(_0163_),
    .A2(_0978_));
 sg13g2_nand3_1 _3413_ (.B(_0425_),
    .C(_0462_),
    .A(net359),
    .Y(_1068_));
 sg13g2_nor2_1 _3414_ (.A(net739),
    .B(net360),
    .Y(_0164_));
 sg13g2_nor4_1 _3415_ (.A(\cpu_instance.mem_instance.mem_ctrl_instance.state[2] ),
    .B(_1302_),
    .C(net738),
    .D(net369),
    .Y(_0165_));
 sg13g2_nor2_1 _3416_ (.A(\cpu_instance.mem_instance.mem_ctrl_instance.state[3] ),
    .B(_1068_),
    .Y(_1069_));
 sg13g2_nor2_2 _3417_ (.A(_0986_),
    .B(net686),
    .Y(_1070_));
 sg13g2_a22oi_1 _3418_ (.Y(_1071_),
    .B1(_1070_),
    .B2(net373),
    .A2(net686),
    .A1(_0539_));
 sg13g2_nor2_1 _3419_ (.A(net740),
    .B(_1071_),
    .Y(_0166_));
 sg13g2_a22oi_1 _3420_ (.Y(_1072_),
    .B1(_1070_),
    .B2(net357),
    .A2(net686),
    .A1(_0505_));
 sg13g2_nor2_1 _3421_ (.A(net739),
    .B(_1072_),
    .Y(_0167_));
 sg13g2_a22oi_1 _3422_ (.Y(_1073_),
    .B1(_1070_),
    .B2(net358),
    .A2(net686),
    .A1(_0524_));
 sg13g2_nor2_1 _3423_ (.A(net739),
    .B(_1073_),
    .Y(_0168_));
 sg13g2_a22oi_1 _3424_ (.Y(_1074_),
    .B1(_1070_),
    .B2(net342),
    .A2(net686),
    .A1(_0559_));
 sg13g2_nor2_1 _3425_ (.A(net739),
    .B(_1074_),
    .Y(_0169_));
 sg13g2_a22oi_1 _3426_ (.Y(_1075_),
    .B1(_1070_),
    .B2(net351),
    .A2(net686),
    .A1(net616));
 sg13g2_nor2_1 _3427_ (.A(net739),
    .B(_1075_),
    .Y(_0170_));
 sg13g2_a22oi_1 _3428_ (.Y(_1076_),
    .B1(_1070_),
    .B2(net339),
    .A2(net686),
    .A1(net602));
 sg13g2_nor2_1 _3429_ (.A(net739),
    .B(_1076_),
    .Y(_0171_));
 sg13g2_a22oi_1 _3430_ (.Y(_1077_),
    .B1(_1070_),
    .B2(net349),
    .A2(_1069_),
    .A1(_0386_));
 sg13g2_nor2_1 _3431_ (.A(net739),
    .B(net350),
    .Y(_0172_));
 sg13g2_a22oi_1 _3432_ (.Y(_1078_),
    .B1(_1070_),
    .B2(net363),
    .A2(net686),
    .A1(net591));
 sg13g2_nor2_1 _3433_ (.A(net739),
    .B(_1078_),
    .Y(_0173_));
 sg13g2_a22oi_1 _3434_ (.Y(_1079_),
    .B1(net685),
    .B2(net326),
    .A2(net690),
    .A1(net324));
 sg13g2_inv_1 _3435_ (.Y(_0174_),
    .A(_1079_));
 sg13g2_mux4_1 _3436_ (.S0(\cpu_instance.ctrl_instance.reg_sel_in[0] ),
    .A0(\cpu_instance.registers_instance.registers[0][0] ),
    .A1(\cpu_instance.registers_instance.registers[1][0] ),
    .A2(\cpu_instance.registers_instance.registers[2][0] ),
    .A3(uo_out[0]),
    .S1(\cpu_instance.ctrl_instance.reg_sel_in[1] ),
    .X(_1080_));
 sg13g2_mux4_1 _3437_ (.S0(\cpu_instance.ctrl_instance.reg_sel_in[0] ),
    .A0(\cpu_instance.registers_instance.registers[0][1] ),
    .A1(\cpu_instance.registers_instance.registers[1][1] ),
    .A2(\cpu_instance.registers_instance.registers[2][1] ),
    .A3(uo_out[1]),
    .S1(\cpu_instance.ctrl_instance.reg_sel_in[1] ),
    .X(_1081_));
 sg13g2_nand2_2 _3438_ (.Y(_1082_),
    .A(_1080_),
    .B(_1081_));
 sg13g2_nand2_2 _3439_ (.Y(_1083_),
    .A(\cpu_instance.ctrl_instance.use_register_bank_in ),
    .B(\cpu_instance.ctrl_instance.reg_op ));
 sg13g2_mux4_1 _3440_ (.S0(\cpu_instance.ctrl_instance.reg_sel_in[0] ),
    .A0(\cpu_instance.registers_instance.registers[2][3] ),
    .A1(_1295_),
    .A2(_1296_),
    .A3(\cpu_instance.registers_instance.registers[1][3] ),
    .S1(_1287_),
    .X(_1084_));
 sg13g2_nor2b_2 _3441_ (.A(_1083_),
    .B_N(_1084_),
    .Y(_1085_));
 sg13g2_mux4_1 _3442_ (.S0(_1288_),
    .A0(uo_out[2]),
    .A1(\cpu_instance.registers_instance.registers[2][2] ),
    .A2(\cpu_instance.registers_instance.registers[1][2] ),
    .A3(_1299_),
    .S1(_1287_),
    .X(_1086_));
 sg13g2_nand2_2 _3443_ (.Y(_1087_),
    .A(_1085_),
    .B(_1086_));
 sg13g2_nor2_1 _3444_ (.A(_1082_),
    .B(_1087_),
    .Y(_1088_));
 sg13g2_o21ai_1 _3445_ (.B1(net750),
    .Y(_1089_),
    .A1(net498),
    .A2(net664));
 sg13g2_a21oi_1 _3446_ (.A1(net621),
    .A2(net664),
    .Y(_0175_),
    .B1(_1089_));
 sg13g2_o21ai_1 _3447_ (.B1(net752),
    .Y(_1090_),
    .A1(net441),
    .A2(net664));
 sg13g2_a21oi_1 _3448_ (.A1(net625),
    .A2(net664),
    .Y(_0176_),
    .B1(_1090_));
 sg13g2_o21ai_1 _3449_ (.B1(net756),
    .Y(_1091_),
    .A1(net502),
    .A2(net665));
 sg13g2_a21oi_1 _3450_ (.A1(net618),
    .A2(net665),
    .Y(_0177_),
    .B1(_1091_));
 sg13g2_o21ai_1 _3451_ (.B1(net763),
    .Y(_1092_),
    .A1(net408),
    .A2(_1088_));
 sg13g2_a21oi_1 _3452_ (.A1(net615),
    .A2(net665),
    .Y(_0178_),
    .B1(_1092_));
 sg13g2_o21ai_1 _3453_ (.B1(net756),
    .Y(_1093_),
    .A1(net435),
    .A2(net665));
 sg13g2_a21oi_1 _3454_ (.A1(net604),
    .A2(net665),
    .Y(_0179_),
    .B1(_1093_));
 sg13g2_o21ai_1 _3455_ (.B1(net764),
    .Y(_1094_),
    .A1(net488),
    .A2(net665));
 sg13g2_a21oi_1 _3456_ (.A1(net607),
    .A2(net665),
    .Y(_0180_),
    .B1(_1094_));
 sg13g2_o21ai_1 _3457_ (.B1(net752),
    .Y(_1095_),
    .A1(net396),
    .A2(net664));
 sg13g2_a21oi_1 _3458_ (.A1(net597),
    .A2(net664),
    .Y(_0181_),
    .B1(_1095_));
 sg13g2_o21ai_1 _3459_ (.B1(net757),
    .Y(_1096_),
    .A1(net531),
    .A2(net664));
 sg13g2_a21oi_1 _3460_ (.A1(net593),
    .A2(net664),
    .Y(_0182_),
    .B1(_1096_));
 sg13g2_nand2b_2 _3461_ (.Y(_1097_),
    .B(_1081_),
    .A_N(_1080_));
 sg13g2_nor2_1 _3462_ (.A(_1087_),
    .B(_1097_),
    .Y(_1098_));
 sg13g2_o21ai_1 _3463_ (.B1(net767),
    .Y(_1099_),
    .A1(net447),
    .A2(net663));
 sg13g2_a21oi_1 _3464_ (.A1(net622),
    .A2(net663),
    .Y(_0183_),
    .B1(_1099_));
 sg13g2_o21ai_1 _3465_ (.B1(net760),
    .Y(_1100_),
    .A1(net410),
    .A2(net663));
 sg13g2_a21oi_1 _3466_ (.A1(net626),
    .A2(net663),
    .Y(_0184_),
    .B1(_1100_));
 sg13g2_o21ai_1 _3467_ (.B1(net765),
    .Y(_1101_),
    .A1(net529),
    .A2(net663));
 sg13g2_a21oi_1 _3468_ (.A1(net618),
    .A2(net663),
    .Y(_0185_),
    .B1(_1101_));
 sg13g2_o21ai_1 _3469_ (.B1(net766),
    .Y(_1102_),
    .A1(net431),
    .A2(_1098_));
 sg13g2_a21oi_1 _3470_ (.A1(net613),
    .A2(net662),
    .Y(_0186_),
    .B1(_1102_));
 sg13g2_o21ai_1 _3471_ (.B1(net767),
    .Y(_1103_),
    .A1(net433),
    .A2(net662));
 sg13g2_a21oi_1 _3472_ (.A1(net604),
    .A2(net662),
    .Y(_0187_),
    .B1(_1103_));
 sg13g2_o21ai_1 _3473_ (.B1(net764),
    .Y(_1104_),
    .A1(net482),
    .A2(net662));
 sg13g2_a21oi_1 _3474_ (.A1(net607),
    .A2(net663),
    .Y(_0188_),
    .B1(_1104_));
 sg13g2_o21ai_1 _3475_ (.B1(net764),
    .Y(_1105_),
    .A1(net475),
    .A2(net662));
 sg13g2_a21oi_1 _3476_ (.A1(net598),
    .A2(net662),
    .Y(_0189_),
    .B1(_1105_));
 sg13g2_o21ai_1 _3477_ (.B1(net763),
    .Y(_1106_),
    .A1(net409),
    .A2(net662));
 sg13g2_a21oi_1 _3478_ (.A1(net594),
    .A2(net662),
    .Y(_0190_),
    .B1(_1106_));
 sg13g2_nand2b_2 _3479_ (.Y(_1107_),
    .B(_1080_),
    .A_N(_1081_));
 sg13g2_nor2_1 _3480_ (.A(_1087_),
    .B(_1107_),
    .Y(_1108_));
 sg13g2_o21ai_1 _3481_ (.B1(net755),
    .Y(_1109_),
    .A1(net494),
    .A2(net660));
 sg13g2_a21oi_1 _3482_ (.A1(net621),
    .A2(net660),
    .Y(_0191_),
    .B1(_1109_));
 sg13g2_o21ai_1 _3483_ (.B1(net766),
    .Y(_1110_),
    .A1(net465),
    .A2(net661));
 sg13g2_a21oi_1 _3484_ (.A1(net627),
    .A2(_1108_),
    .Y(_0192_),
    .B1(_1110_));
 sg13g2_o21ai_1 _3485_ (.B1(net754),
    .Y(_1111_),
    .A1(net460),
    .A2(net660));
 sg13g2_a21oi_1 _3486_ (.A1(net617),
    .A2(net660),
    .Y(_0193_),
    .B1(_1111_));
 sg13g2_o21ai_1 _3487_ (.B1(net753),
    .Y(_1112_),
    .A1(net491),
    .A2(net660));
 sg13g2_a21oi_1 _3488_ (.A1(net614),
    .A2(net660),
    .Y(_0194_),
    .B1(_1112_));
 sg13g2_o21ai_1 _3489_ (.B1(net755),
    .Y(_1113_),
    .A1(net455),
    .A2(net660));
 sg13g2_a21oi_1 _3490_ (.A1(net604),
    .A2(net660),
    .Y(_0195_),
    .B1(_1113_));
 sg13g2_o21ai_1 _3491_ (.B1(net764),
    .Y(_1114_),
    .A1(net514),
    .A2(net661));
 sg13g2_a21oi_1 _3492_ (.A1(net607),
    .A2(net661),
    .Y(_0196_),
    .B1(_1114_));
 sg13g2_o21ai_1 _3493_ (.B1(net763),
    .Y(_1115_),
    .A1(net512),
    .A2(net661));
 sg13g2_a21oi_1 _3494_ (.A1(net599),
    .A2(net661),
    .Y(_0197_),
    .B1(_1115_));
 sg13g2_o21ai_1 _3495_ (.B1(net754),
    .Y(_1116_),
    .A1(net524),
    .A2(net661));
 sg13g2_a21oi_1 _3496_ (.A1(net593),
    .A2(net661),
    .Y(_0198_),
    .B1(_1116_));
 sg13g2_or2_2 _3497_ (.X(_1117_),
    .B(_1081_),
    .A(_1080_));
 sg13g2_nor2_2 _3498_ (.A(_1087_),
    .B(_1117_),
    .Y(_1118_));
 sg13g2_o21ai_1 _3499_ (.B1(net766),
    .Y(_1119_),
    .A1(net404),
    .A2(net659));
 sg13g2_a21oi_1 _3500_ (.A1(net622),
    .A2(net659),
    .Y(_0199_),
    .B1(_1119_));
 sg13g2_o21ai_1 _3501_ (.B1(net767),
    .Y(_1120_),
    .A1(net425),
    .A2(net659));
 sg13g2_a21oi_1 _3502_ (.A1(net626),
    .A2(net659),
    .Y(_0200_),
    .B1(_1120_));
 sg13g2_o21ai_1 _3503_ (.B1(net757),
    .Y(_1121_),
    .A1(net549),
    .A2(net658));
 sg13g2_a21oi_1 _3504_ (.A1(net617),
    .A2(net658),
    .Y(_0201_),
    .B1(_1121_));
 sg13g2_o21ai_1 _3505_ (.B1(net767),
    .Y(_1122_),
    .A1(net573),
    .A2(net659));
 sg13g2_a21oi_1 _3506_ (.A1(net613),
    .A2(net659),
    .Y(_0202_),
    .B1(_1122_));
 sg13g2_o21ai_1 _3507_ (.B1(net756),
    .Y(_1123_),
    .A1(net459),
    .A2(net658));
 sg13g2_a21oi_1 _3508_ (.A1(net603),
    .A2(net658),
    .Y(_0203_),
    .B1(_1123_));
 sg13g2_o21ai_1 _3509_ (.B1(net766),
    .Y(_1124_),
    .A1(net450),
    .A2(net659));
 sg13g2_a21oi_1 _3510_ (.A1(net610),
    .A2(net659),
    .Y(_0204_),
    .B1(_1124_));
 sg13g2_o21ai_1 _3511_ (.B1(net763),
    .Y(_1125_),
    .A1(net480),
    .A2(net658));
 sg13g2_a21oi_1 _3512_ (.A1(net598),
    .A2(net658),
    .Y(_0205_),
    .B1(_1125_));
 sg13g2_o21ai_1 _3513_ (.B1(net757),
    .Y(_1126_),
    .A1(net501),
    .A2(net658));
 sg13g2_a21oi_1 _3514_ (.A1(net592),
    .A2(net658),
    .Y(_0206_),
    .B1(_1126_));
 sg13g2_nand2b_2 _3515_ (.Y(_1127_),
    .B(_1085_),
    .A_N(_1086_));
 sg13g2_nor2_1 _3516_ (.A(_1082_),
    .B(_1127_),
    .Y(_1128_));
 sg13g2_o21ai_1 _3517_ (.B1(net760),
    .Y(_1129_),
    .A1(net474),
    .A2(net655));
 sg13g2_a21oi_1 _3518_ (.A1(net624),
    .A2(net655),
    .Y(_0207_),
    .B1(_1129_));
 sg13g2_o21ai_1 _3519_ (.B1(net764),
    .Y(_1130_),
    .A1(net481),
    .A2(net656));
 sg13g2_a21oi_1 _3520_ (.A1(net627),
    .A2(net656),
    .Y(_0208_),
    .B1(_1130_));
 sg13g2_o21ai_1 _3521_ (.B1(net763),
    .Y(_1131_),
    .A1(net543),
    .A2(net656));
 sg13g2_a21oi_1 _3522_ (.A1(net618),
    .A2(net656),
    .Y(_0209_),
    .B1(_1131_));
 sg13g2_o21ai_1 _3523_ (.B1(net760),
    .Y(_1132_),
    .A1(net507),
    .A2(net655));
 sg13g2_a21oi_1 _3524_ (.A1(net613),
    .A2(net655),
    .Y(_0210_),
    .B1(_1132_));
 sg13g2_o21ai_1 _3525_ (.B1(net749),
    .Y(_1133_),
    .A1(net430),
    .A2(net657));
 sg13g2_a21oi_1 _3526_ (.A1(net603),
    .A2(net657),
    .Y(_0211_),
    .B1(_1133_));
 sg13g2_o21ai_1 _3527_ (.B1(net749),
    .Y(_1134_),
    .A1(net412),
    .A2(net657));
 sg13g2_a21oi_1 _3528_ (.A1(net606),
    .A2(net657),
    .Y(_0212_),
    .B1(_1134_));
 sg13g2_o21ai_1 _3529_ (.B1(net757),
    .Y(_1135_),
    .A1(net486),
    .A2(net655));
 sg13g2_a21oi_1 _3530_ (.A1(net598),
    .A2(net655),
    .Y(_0213_),
    .B1(_1135_));
 sg13g2_o21ai_1 _3531_ (.B1(net757),
    .Y(_1136_),
    .A1(net534),
    .A2(net655));
 sg13g2_a21oi_1 _3532_ (.A1(net593),
    .A2(net655),
    .Y(_0214_),
    .B1(_1136_));
 sg13g2_nor2_1 _3533_ (.A(_1097_),
    .B(_1127_),
    .Y(_1137_));
 sg13g2_o21ai_1 _3534_ (.B1(net753),
    .Y(_1138_),
    .A1(net424),
    .A2(net653));
 sg13g2_a21oi_1 _3535_ (.A1(net621),
    .A2(net653),
    .Y(_0215_),
    .B1(_1138_));
 sg13g2_o21ai_1 _3536_ (.B1(net763),
    .Y(_1139_),
    .A1(net567),
    .A2(net654));
 sg13g2_a21oi_1 _3537_ (.A1(net626),
    .A2(net654),
    .Y(_0216_),
    .B1(_1139_));
 sg13g2_o21ai_1 _3538_ (.B1(net756),
    .Y(_1140_),
    .A1(net483),
    .A2(net654));
 sg13g2_a21oi_1 _3539_ (.A1(net617),
    .A2(net654),
    .Y(_0217_),
    .B1(_1140_));
 sg13g2_o21ai_1 _3540_ (.B1(net754),
    .Y(_1141_),
    .A1(net442),
    .A2(net653));
 sg13g2_a21oi_1 _3541_ (.A1(net614),
    .A2(net653),
    .Y(_0218_),
    .B1(_1141_));
 sg13g2_o21ai_1 _3542_ (.B1(net756),
    .Y(_1142_),
    .A1(net423),
    .A2(net654));
 sg13g2_a21oi_1 _3543_ (.A1(net603),
    .A2(net654),
    .Y(_0219_),
    .B1(_1142_));
 sg13g2_o21ai_1 _3544_ (.B1(net753),
    .Y(_1143_),
    .A1(net417),
    .A2(net653));
 sg13g2_a21oi_1 _3545_ (.A1(net606),
    .A2(net653),
    .Y(_0220_),
    .B1(_1143_));
 sg13g2_o21ai_1 _3546_ (.B1(net757),
    .Y(_1144_),
    .A1(net476),
    .A2(net654));
 sg13g2_a21oi_1 _3547_ (.A1(net598),
    .A2(net654),
    .Y(_0221_),
    .B1(_1144_));
 sg13g2_o21ai_1 _3548_ (.B1(net754),
    .Y(_1145_),
    .A1(net451),
    .A2(net653));
 sg13g2_a21oi_1 _3549_ (.A1(net593),
    .A2(net653),
    .Y(_0222_),
    .B1(_1145_));
 sg13g2_nor2_1 _3550_ (.A(_1107_),
    .B(_1127_),
    .Y(_1146_));
 sg13g2_o21ai_1 _3551_ (.B1(net753),
    .Y(_1147_),
    .A1(net487),
    .A2(net651));
 sg13g2_a21oi_1 _3552_ (.A1(net621),
    .A2(net651),
    .Y(_0223_),
    .B1(_1147_));
 sg13g2_o21ai_1 _3553_ (.B1(net763),
    .Y(_1148_),
    .A1(net454),
    .A2(net652));
 sg13g2_a21oi_1 _3554_ (.A1(net626),
    .A2(net652),
    .Y(_0224_),
    .B1(_1148_));
 sg13g2_o21ai_1 _3555_ (.B1(net756),
    .Y(_1149_),
    .A1(net497),
    .A2(net652));
 sg13g2_a21oi_1 _3556_ (.A1(net617),
    .A2(net652),
    .Y(_0225_),
    .B1(_1149_));
 sg13g2_o21ai_1 _3557_ (.B1(net763),
    .Y(_1150_),
    .A1(net439),
    .A2(net652));
 sg13g2_a21oi_1 _3558_ (.A1(net615),
    .A2(net652),
    .Y(_0226_),
    .B1(_1150_));
 sg13g2_o21ai_1 _3559_ (.B1(net765),
    .Y(_1151_),
    .A1(net517),
    .A2(_1146_));
 sg13g2_a21oi_1 _3560_ (.A1(net605),
    .A2(net652),
    .Y(_0227_),
    .B1(_1151_));
 sg13g2_o21ai_1 _3561_ (.B1(net754),
    .Y(_1152_),
    .A1(net464),
    .A2(net651));
 sg13g2_a21oi_1 _3562_ (.A1(net606),
    .A2(net651),
    .Y(_0228_),
    .B1(_1152_));
 sg13g2_o21ai_1 _3563_ (.B1(net757),
    .Y(_1153_),
    .A1(net422),
    .A2(net651));
 sg13g2_a21oi_1 _3564_ (.A1(net598),
    .A2(net651),
    .Y(_0229_),
    .B1(_1153_));
 sg13g2_o21ai_1 _3565_ (.B1(net754),
    .Y(_1154_),
    .A1(net453),
    .A2(net651));
 sg13g2_a21oi_1 _3566_ (.A1(net592),
    .A2(net651),
    .Y(_0230_),
    .B1(_1154_));
 sg13g2_nor2_2 _3567_ (.A(_1117_),
    .B(_1127_),
    .Y(_1155_));
 sg13g2_o21ai_1 _3568_ (.B1(net753),
    .Y(_1156_),
    .A1(net575),
    .A2(net649));
 sg13g2_a21oi_1 _3569_ (.A1(net621),
    .A2(net649),
    .Y(_0231_),
    .B1(_1156_));
 sg13g2_o21ai_1 _3570_ (.B1(net764),
    .Y(_1157_),
    .A1(net446),
    .A2(_1155_));
 sg13g2_a21oi_1 _3571_ (.A1(net626),
    .A2(_1155_),
    .Y(_0232_),
    .B1(_1157_));
 sg13g2_o21ai_1 _3572_ (.B1(net755),
    .Y(_1158_),
    .A1(net436),
    .A2(net650));
 sg13g2_a21oi_1 _3573_ (.A1(net617),
    .A2(net650),
    .Y(_0233_),
    .B1(_1158_));
 sg13g2_o21ai_1 _3574_ (.B1(net753),
    .Y(_1159_),
    .A1(net448),
    .A2(net649));
 sg13g2_a21oi_1 _3575_ (.A1(net614),
    .A2(net649),
    .Y(_0234_),
    .B1(_1159_));
 sg13g2_o21ai_1 _3576_ (.B1(net753),
    .Y(_1160_),
    .A1(net432),
    .A2(net649));
 sg13g2_a21oi_1 _3577_ (.A1(net603),
    .A2(net649),
    .Y(_0235_),
    .B1(_1160_));
 sg13g2_o21ai_1 _3578_ (.B1(net754),
    .Y(_1161_),
    .A1(net472),
    .A2(net650));
 sg13g2_a21oi_1 _3579_ (.A1(net606),
    .A2(net650),
    .Y(_0236_),
    .B1(_1161_));
 sg13g2_o21ai_1 _3580_ (.B1(net757),
    .Y(_1162_),
    .A1(net511),
    .A2(net650));
 sg13g2_a21oi_1 _3581_ (.A1(net598),
    .A2(net650),
    .Y(_0237_),
    .B1(_1162_));
 sg13g2_o21ai_1 _3582_ (.B1(net754),
    .Y(_1163_),
    .A1(net499),
    .A2(net649));
 sg13g2_a21oi_1 _3583_ (.A1(net592),
    .A2(net649),
    .Y(_0238_),
    .B1(_1163_));
 sg13g2_nor2_1 _3584_ (.A(_1083_),
    .B(_1084_),
    .Y(_1164_));
 sg13g2_nand2_2 _3585_ (.Y(_1165_),
    .A(_1086_),
    .B(_1164_));
 sg13g2_nor2_1 _3586_ (.A(_1082_),
    .B(_1165_),
    .Y(_1166_));
 sg13g2_o21ai_1 _3587_ (.B1(net767),
    .Y(_1167_),
    .A1(net504),
    .A2(net648));
 sg13g2_a21oi_1 _3588_ (.A1(net623),
    .A2(net648),
    .Y(_0239_),
    .B1(_1167_));
 sg13g2_o21ai_1 _3589_ (.B1(net752),
    .Y(_1168_),
    .A1(net522),
    .A2(net647));
 sg13g2_a21oi_1 _3590_ (.A1(net625),
    .A2(net648),
    .Y(_0240_),
    .B1(_1168_));
 sg13g2_o21ai_1 _3591_ (.B1(net756),
    .Y(_1169_),
    .A1(net452),
    .A2(net648));
 sg13g2_a21oi_1 _3592_ (.A1(net617),
    .A2(net647),
    .Y(_0241_),
    .B1(_1169_));
 sg13g2_o21ai_1 _3593_ (.B1(net753),
    .Y(_1170_),
    .A1(net539),
    .A2(net647));
 sg13g2_a21oi_1 _3594_ (.A1(net614),
    .A2(net647),
    .Y(_0242_),
    .B1(_1170_));
 sg13g2_o21ai_1 _3595_ (.B1(net767),
    .Y(_1171_),
    .A1(net532),
    .A2(_1166_));
 sg13g2_a21oi_1 _3596_ (.A1(net604),
    .A2(net648),
    .Y(_0243_),
    .B1(_1171_));
 sg13g2_o21ai_1 _3597_ (.B1(net749),
    .Y(_1172_),
    .A1(net457),
    .A2(net647));
 sg13g2_a21oi_1 _3598_ (.A1(net606),
    .A2(net647),
    .Y(_0244_),
    .B1(_1172_));
 sg13g2_o21ai_1 _3599_ (.B1(net760),
    .Y(_1173_),
    .A1(net569),
    .A2(net648));
 sg13g2_a21oi_1 _3600_ (.A1(net597),
    .A2(net648),
    .Y(_0245_),
    .B1(_1173_));
 sg13g2_o21ai_1 _3601_ (.B1(net752),
    .Y(_1174_),
    .A1(net467),
    .A2(net647));
 sg13g2_a21oi_1 _3602_ (.A1(net592),
    .A2(net647),
    .Y(_0246_),
    .B1(_1174_));
 sg13g2_nor2_2 _3603_ (.A(_1097_),
    .B(_1165_),
    .Y(_1175_));
 sg13g2_o21ai_1 _3604_ (.B1(net750),
    .Y(_1176_),
    .A1(net471),
    .A2(net645));
 sg13g2_a21oi_1 _3605_ (.A1(net621),
    .A2(net645),
    .Y(_0247_),
    .B1(_1176_));
 sg13g2_o21ai_1 _3606_ (.B1(net751),
    .Y(_1177_),
    .A1(net525),
    .A2(net646));
 sg13g2_a21oi_1 _3607_ (.A1(net625),
    .A2(net646),
    .Y(_0248_),
    .B1(_1177_));
 sg13g2_o21ai_1 _3608_ (.B1(net758),
    .Y(_1178_),
    .A1(net555),
    .A2(net646));
 sg13g2_a21oi_1 _3609_ (.A1(net617),
    .A2(net646),
    .Y(_0249_),
    .B1(_1178_));
 sg13g2_o21ai_1 _3610_ (.B1(net751),
    .Y(_1179_),
    .A1(net560),
    .A2(net646));
 sg13g2_a21oi_1 _3611_ (.A1(net614),
    .A2(net646),
    .Y(_0250_),
    .B1(_1179_));
 sg13g2_o21ai_1 _3612_ (.B1(net750),
    .Y(_1180_),
    .A1(net402),
    .A2(net645));
 sg13g2_a21oi_1 _3613_ (.A1(net603),
    .A2(net645),
    .Y(_0251_),
    .B1(_1180_));
 sg13g2_o21ai_1 _3614_ (.B1(net748),
    .Y(_1181_),
    .A1(net397),
    .A2(net645));
 sg13g2_a21oi_1 _3615_ (.A1(net606),
    .A2(net645),
    .Y(_0252_),
    .B1(_1181_));
 sg13g2_o21ai_1 _3616_ (.B1(net751),
    .Y(_1182_),
    .A1(net415),
    .A2(net646));
 sg13g2_a21oi_1 _3617_ (.A1(net597),
    .A2(net646),
    .Y(_0253_),
    .B1(_1182_));
 sg13g2_o21ai_1 _3618_ (.B1(net748),
    .Y(_1183_),
    .A1(net536),
    .A2(net645));
 sg13g2_a21oi_1 _3619_ (.A1(net592),
    .A2(net645),
    .Y(_0254_),
    .B1(_1183_));
 sg13g2_nor2_1 _3620_ (.A(_1107_),
    .B(_1165_),
    .Y(_1184_));
 sg13g2_o21ai_1 _3621_ (.B1(net748),
    .Y(_1185_),
    .A1(net784),
    .A2(net642));
 sg13g2_a21oi_1 _3622_ (.A1(net621),
    .A2(net642),
    .Y(_0255_),
    .B1(_1185_));
 sg13g2_o21ai_1 _3623_ (.B1(net751),
    .Y(_1186_),
    .A1(net470),
    .A2(net644));
 sg13g2_a21oi_1 _3624_ (.A1(net625),
    .A2(net644),
    .Y(_0256_),
    .B1(_1186_));
 sg13g2_o21ai_1 _3625_ (.B1(net748),
    .Y(_1187_),
    .A1(net523),
    .A2(net643));
 sg13g2_a21oi_1 _3626_ (.A1(net618),
    .A2(net643),
    .Y(_0257_),
    .B1(_1187_));
 sg13g2_o21ai_1 _3627_ (.B1(net748),
    .Y(_1188_),
    .A1(net434),
    .A2(net642));
 sg13g2_a21oi_1 _3628_ (.A1(net614),
    .A2(net642),
    .Y(_0258_),
    .B1(_1188_));
 sg13g2_o21ai_1 _3629_ (.B1(net749),
    .Y(_1189_),
    .A1(net469),
    .A2(net643));
 sg13g2_a21oi_1 _3630_ (.A1(net603),
    .A2(net643),
    .Y(_0259_),
    .B1(_1189_));
 sg13g2_o21ai_1 _3631_ (.B1(net749),
    .Y(_1190_),
    .A1(net449),
    .A2(net642));
 sg13g2_a21oi_1 _3632_ (.A1(net606),
    .A2(net642),
    .Y(_0260_),
    .B1(_1190_));
 sg13g2_o21ai_1 _3633_ (.B1(net759),
    .Y(_1191_),
    .A1(net546),
    .A2(net644));
 sg13g2_a21oi_1 _3634_ (.A1(net597),
    .A2(net644),
    .Y(_0261_),
    .B1(_1191_));
 sg13g2_o21ai_1 _3635_ (.B1(net748),
    .Y(_1192_),
    .A1(net416),
    .A2(net642));
 sg13g2_a21oi_1 _3636_ (.A1(net592),
    .A2(net642),
    .Y(_0262_),
    .B1(_1192_));
 sg13g2_nor2_2 _3637_ (.A(_1117_),
    .B(_1165_),
    .Y(_1193_));
 sg13g2_o21ai_1 _3638_ (.B1(net749),
    .Y(_1194_),
    .A1(net579),
    .A2(net640));
 sg13g2_a21oi_1 _3639_ (.A1(net621),
    .A2(net640),
    .Y(_0263_),
    .B1(_1194_));
 sg13g2_o21ai_1 _3640_ (.B1(net752),
    .Y(_1195_),
    .A1(net428),
    .A2(_1193_));
 sg13g2_a21oi_1 _3641_ (.A1(net625),
    .A2(net641),
    .Y(_0264_),
    .B1(_1195_));
 sg13g2_o21ai_1 _3642_ (.B1(net750),
    .Y(_1196_),
    .A1(net407),
    .A2(net641));
 sg13g2_a21oi_1 _3643_ (.A1(net618),
    .A2(net641),
    .Y(_0265_),
    .B1(_1196_));
 sg13g2_o21ai_1 _3644_ (.B1(net748),
    .Y(_1197_),
    .A1(net484),
    .A2(net640));
 sg13g2_a21oi_1 _3645_ (.A1(net614),
    .A2(net640),
    .Y(_0266_),
    .B1(_1197_));
 sg13g2_o21ai_1 _3646_ (.B1(net749),
    .Y(_1198_),
    .A1(net414),
    .A2(net640));
 sg13g2_a21oi_1 _3647_ (.A1(net603),
    .A2(net640),
    .Y(_0267_),
    .B1(_1198_));
 sg13g2_o21ai_1 _3648_ (.B1(net749),
    .Y(_1199_),
    .A1(net495),
    .A2(net640));
 sg13g2_a21oi_1 _3649_ (.A1(net606),
    .A2(net640),
    .Y(_0268_),
    .B1(_1199_));
 sg13g2_o21ai_1 _3650_ (.B1(net751),
    .Y(_1200_),
    .A1(net418),
    .A2(net641));
 sg13g2_a21oi_1 _3651_ (.A1(net597),
    .A2(net641),
    .Y(_0269_),
    .B1(_1200_));
 sg13g2_o21ai_1 _3652_ (.B1(net752),
    .Y(_1201_),
    .A1(net456),
    .A2(net641));
 sg13g2_a21oi_1 _3653_ (.A1(net592),
    .A2(net641),
    .Y(_0270_),
    .B1(_1201_));
 sg13g2_nand2b_2 _3654_ (.Y(_1202_),
    .B(_1164_),
    .A_N(_1086_));
 sg13g2_nor2_1 _3655_ (.A(_1082_),
    .B(_1202_),
    .Y(_1203_));
 sg13g2_o21ai_1 _3656_ (.B1(net760),
    .Y(_1204_),
    .A1(net490),
    .A2(_1203_));
 sg13g2_a21oi_1 _3657_ (.A1(net624),
    .A2(net638),
    .Y(_0271_),
    .B1(_1204_));
 sg13g2_o21ai_1 _3658_ (.B1(net751),
    .Y(_1205_),
    .A1(net438),
    .A2(net639));
 sg13g2_a21oi_1 _3659_ (.A1(net625),
    .A2(net639),
    .Y(_0272_),
    .B1(_1205_));
 sg13g2_o21ai_1 _3660_ (.B1(net759),
    .Y(_1206_),
    .A1(net559),
    .A2(net638));
 sg13g2_a21oi_1 _3661_ (.A1(net618),
    .A2(net638),
    .Y(_0273_),
    .B1(_1206_));
 sg13g2_o21ai_1 _3662_ (.B1(net751),
    .Y(_1207_),
    .A1(net406),
    .A2(net638));
 sg13g2_a21oi_1 _3663_ (.A1(net614),
    .A2(net639),
    .Y(_0274_),
    .B1(_1207_));
 sg13g2_o21ai_1 _3664_ (.B1(net748),
    .Y(_1208_),
    .A1(net485),
    .A2(net639));
 sg13g2_a21oi_1 _3665_ (.A1(net603),
    .A2(net639),
    .Y(_0275_),
    .B1(_1208_));
 sg13g2_o21ai_1 _3666_ (.B1(net759),
    .Y(_1209_),
    .A1(net556),
    .A2(net638));
 sg13g2_a21oi_1 _3667_ (.A1(net607),
    .A2(net638),
    .Y(_0276_),
    .B1(_1209_));
 sg13g2_o21ai_1 _3668_ (.B1(net751),
    .Y(_1210_),
    .A1(net444),
    .A2(net639));
 sg13g2_a21oi_1 _3669_ (.A1(net597),
    .A2(net639),
    .Y(_0277_),
    .B1(_1210_));
 sg13g2_o21ai_1 _3670_ (.B1(net759),
    .Y(_1211_),
    .A1(net513),
    .A2(net638));
 sg13g2_a21oi_1 _3671_ (.A1(net592),
    .A2(net638),
    .Y(_0278_),
    .B1(_1211_));
 sg13g2_nand2b_2 _3672_ (.Y(_1212_),
    .B(\cpu_instance.ctrl_instance.reg_op ),
    .A_N(\cpu_instance.ctrl_instance.use_register_bank_in ));
 sg13g2_nor3_1 _3673_ (.A(\cpu_instance.ctrl_instance.reg_sel_in[1] ),
    .B(\cpu_instance.ctrl_instance.reg_sel_in[0] ),
    .C(_1212_),
    .Y(_1213_));
 sg13g2_o21ai_1 _3674_ (.B1(net774),
    .Y(_1214_),
    .A1(net802),
    .A2(net699));
 sg13g2_a21oi_1 _3675_ (.A1(net623),
    .A2(net699),
    .Y(_0279_),
    .B1(_1214_));
 sg13g2_o21ai_1 _3676_ (.B1(net774),
    .Y(_1215_),
    .A1(net786),
    .A2(net699));
 sg13g2_a21oi_1 _3677_ (.A1(net627),
    .A2(net699),
    .Y(_0280_),
    .B1(_1215_));
 sg13g2_o21ai_1 _3678_ (.B1(net779),
    .Y(_1216_),
    .A1(net795),
    .A2(net699));
 sg13g2_a21oi_1 _3679_ (.A1(net620),
    .A2(net699),
    .Y(_0281_),
    .B1(_1216_));
 sg13g2_o21ai_1 _3680_ (.B1(net774),
    .Y(_1217_),
    .A1(net383),
    .A2(net699));
 sg13g2_a21oi_1 _3681_ (.A1(_0558_),
    .A2(net699),
    .Y(_0282_),
    .B1(_1217_));
 sg13g2_o21ai_1 _3682_ (.B1(net778),
    .Y(_1218_),
    .A1(net386),
    .A2(net700));
 sg13g2_a21oi_1 _3683_ (.A1(net605),
    .A2(net700),
    .Y(_0283_),
    .B1(_1218_));
 sg13g2_o21ai_1 _3684_ (.B1(net779),
    .Y(_1219_),
    .A1(net578),
    .A2(net700));
 sg13g2_a21oi_1 _3685_ (.A1(net611),
    .A2(net700),
    .Y(_0284_),
    .B1(_1219_));
 sg13g2_o21ai_1 _3686_ (.B1(net778),
    .Y(_1220_),
    .A1(net473),
    .A2(net700));
 sg13g2_a21oi_1 _3687_ (.A1(net600),
    .A2(net700),
    .Y(_0285_),
    .B1(_1220_));
 sg13g2_o21ai_1 _3688_ (.B1(net778),
    .Y(_1221_),
    .A1(net783),
    .A2(net700));
 sg13g2_a21oi_1 _3689_ (.A1(net596),
    .A2(net700),
    .Y(_0286_),
    .B1(_1221_));
 sg13g2_nor3_1 _3690_ (.A(\cpu_instance.ctrl_instance.reg_sel_in[1] ),
    .B(_1288_),
    .C(_1212_),
    .Y(_1222_));
 sg13g2_o21ai_1 _3691_ (.B1(net774),
    .Y(_1223_),
    .A1(net815),
    .A2(net698));
 sg13g2_a21oi_1 _3692_ (.A1(net623),
    .A2(net698),
    .Y(_0287_),
    .B1(_1223_));
 sg13g2_o21ai_1 _3693_ (.B1(net774),
    .Y(_1224_),
    .A1(net824),
    .A2(net698));
 sg13g2_a21oi_1 _3694_ (.A1(net627),
    .A2(net698),
    .Y(_0288_),
    .B1(_1224_));
 sg13g2_o21ai_1 _3695_ (.B1(net779),
    .Y(_1225_),
    .A1(net844),
    .A2(net697));
 sg13g2_a21oi_1 _3696_ (.A1(net620),
    .A2(net697),
    .Y(_0289_),
    .B1(_1225_));
 sg13g2_o21ai_1 _3697_ (.B1(net774),
    .Y(_1226_),
    .A1(net818),
    .A2(net698));
 sg13g2_a21oi_1 _3698_ (.A1(net615),
    .A2(net698),
    .Y(_0290_),
    .B1(_1226_));
 sg13g2_o21ai_1 _3699_ (.B1(net779),
    .Y(_1227_),
    .A1(net478),
    .A2(_1222_));
 sg13g2_a21oi_1 _3700_ (.A1(net605),
    .A2(net698),
    .Y(_0291_),
    .B1(net479));
 sg13g2_o21ai_1 _3701_ (.B1(net779),
    .Y(_1228_),
    .A1(net521),
    .A2(net697));
 sg13g2_a21oi_1 _3702_ (.A1(net611),
    .A2(net697),
    .Y(_0292_),
    .B1(_1228_));
 sg13g2_o21ai_1 _3703_ (.B1(net778),
    .Y(_1229_),
    .A1(net571),
    .A2(net697));
 sg13g2_a21oi_1 _3704_ (.A1(net601),
    .A2(net697),
    .Y(_0293_),
    .B1(_1229_));
 sg13g2_o21ai_1 _3705_ (.B1(net778),
    .Y(_1230_),
    .A1(net587),
    .A2(net697));
 sg13g2_a21oi_1 _3706_ (.A1(net595),
    .A2(net697),
    .Y(_0294_),
    .B1(_1230_));
 sg13g2_nor3_1 _3707_ (.A(_1287_),
    .B(\cpu_instance.ctrl_instance.reg_sel_in[0] ),
    .C(_1212_),
    .Y(_1231_));
 sg13g2_o21ai_1 _3708_ (.B1(net775),
    .Y(_1232_),
    .A1(net823),
    .A2(net696));
 sg13g2_a21oi_1 _3709_ (.A1(net623),
    .A2(net696),
    .Y(_0295_),
    .B1(_1232_));
 sg13g2_o21ai_1 _3710_ (.B1(net774),
    .Y(_1233_),
    .A1(net833),
    .A2(net696));
 sg13g2_a21oi_1 _3711_ (.A1(net627),
    .A2(net696),
    .Y(_0296_),
    .B1(_1233_));
 sg13g2_o21ai_1 _3712_ (.B1(net779),
    .Y(_1234_),
    .A1(net841),
    .A2(net695));
 sg13g2_a21oi_1 _3713_ (.A1(net620),
    .A2(net695),
    .Y(_0297_),
    .B1(_1234_));
 sg13g2_o21ai_1 _3714_ (.B1(net774),
    .Y(_1235_),
    .A1(net821),
    .A2(net696));
 sg13g2_a21oi_1 _3715_ (.A1(net615),
    .A2(net696),
    .Y(_0298_),
    .B1(_1235_));
 sg13g2_o21ai_1 _3716_ (.B1(net778),
    .Y(_1236_),
    .A1(net537),
    .A2(_1231_));
 sg13g2_a21oi_1 _3717_ (.A1(net605),
    .A2(net696),
    .Y(_0299_),
    .B1(net538));
 sg13g2_o21ai_1 _3718_ (.B1(net779),
    .Y(_1237_),
    .A1(net792),
    .A2(net695));
 sg13g2_a21oi_1 _3719_ (.A1(net611),
    .A2(net695),
    .Y(_0300_),
    .B1(_1237_));
 sg13g2_o21ai_1 _3720_ (.B1(net778),
    .Y(_1238_),
    .A1(net552),
    .A2(net695));
 sg13g2_a21oi_1 _3721_ (.A1(net600),
    .A2(net695),
    .Y(_0301_),
    .B1(_1238_));
 sg13g2_o21ai_1 _3722_ (.B1(net778),
    .Y(_1239_),
    .A1(net806),
    .A2(net695));
 sg13g2_a21oi_1 _3723_ (.A1(net595),
    .A2(net695),
    .Y(_0302_),
    .B1(_1239_));
 sg13g2_nor3_1 _3724_ (.A(_1287_),
    .B(_1288_),
    .C(_1212_),
    .Y(_1240_));
 sg13g2_o21ai_1 _3725_ (.B1(net773),
    .Y(_1241_),
    .A1(net850),
    .A2(net694));
 sg13g2_a21oi_1 _3726_ (.A1(net623),
    .A2(net694),
    .Y(_0303_),
    .B1(_1241_));
 sg13g2_o21ai_1 _3727_ (.B1(net773),
    .Y(_1242_),
    .A1(net842),
    .A2(net694));
 sg13g2_a21oi_1 _3728_ (.A1(net627),
    .A2(net694),
    .Y(_0304_),
    .B1(_1242_));
 sg13g2_o21ai_1 _3729_ (.B1(net776),
    .Y(_1243_),
    .A1(net851),
    .A2(net693));
 sg13g2_a21oi_1 _3730_ (.A1(net620),
    .A2(net693),
    .Y(_0305_),
    .B1(_1243_));
 sg13g2_o21ai_1 _3731_ (.B1(net776),
    .Y(_1244_),
    .A1(net582),
    .A2(net692));
 sg13g2_a21oi_1 _3732_ (.A1(net615),
    .A2(net692),
    .Y(_0306_),
    .B1(_1244_));
 sg13g2_o21ai_1 _3733_ (.B1(net777),
    .Y(_1245_),
    .A1(net576),
    .A2(net692));
 sg13g2_a21oi_1 _3734_ (.A1(net605),
    .A2(net692),
    .Y(_0307_),
    .B1(_1245_));
 sg13g2_o21ai_1 _3735_ (.B1(net776),
    .Y(_1246_),
    .A1(net843),
    .A2(net693));
 sg13g2_a21oi_1 _3736_ (.A1(net611),
    .A2(net693),
    .Y(_0308_),
    .B1(_1246_));
 sg13g2_o21ai_1 _3737_ (.B1(net776),
    .Y(_1247_),
    .A1(net837),
    .A2(net692));
 sg13g2_a21oi_1 _3738_ (.A1(net601),
    .A2(net692),
    .Y(_0309_),
    .B1(_1247_));
 sg13g2_o21ai_1 _3739_ (.B1(net776),
    .Y(_1248_),
    .A1(net840),
    .A2(net692));
 sg13g2_a21oi_1 _3740_ (.A1(net596),
    .A2(net692),
    .Y(_0310_),
    .B1(_1248_));
 sg13g2_nor2_1 _3741_ (.A(_1117_),
    .B(_1202_),
    .Y(_1249_));
 sg13g2_o21ai_1 _3742_ (.B1(net761),
    .Y(_1250_),
    .A1(net533),
    .A2(net636));
 sg13g2_a21oi_1 _3743_ (.A1(net623),
    .A2(net636),
    .Y(_0311_),
    .B1(_1250_));
 sg13g2_o21ai_1 _3744_ (.B1(net761),
    .Y(_1251_),
    .A1(net801),
    .A2(net637));
 sg13g2_a21oi_1 _3745_ (.A1(_0504_),
    .A2(net637),
    .Y(_0312_),
    .B1(_1251_));
 sg13g2_o21ai_1 _3746_ (.B1(net762),
    .Y(_1252_),
    .A1(net547),
    .A2(net636));
 sg13g2_a21oi_1 _3747_ (.A1(net619),
    .A2(net636),
    .Y(_0313_),
    .B1(_1252_));
 sg13g2_o21ai_1 _3748_ (.B1(net761),
    .Y(_1253_),
    .A1(net516),
    .A2(net636));
 sg13g2_a21oi_1 _3749_ (.A1(net613),
    .A2(net636),
    .Y(_0314_),
    .B1(_1253_));
 sg13g2_o21ai_1 _3750_ (.B1(net761),
    .Y(_1254_),
    .A1(net580),
    .A2(net636));
 sg13g2_a21oi_1 _3751_ (.A1(net604),
    .A2(net636),
    .Y(_0315_),
    .B1(_1254_));
 sg13g2_o21ai_1 _3752_ (.B1(net773),
    .Y(_1255_),
    .A1(net781),
    .A2(net637));
 sg13g2_a21oi_1 _3753_ (.A1(net608),
    .A2(net637),
    .Y(_0316_),
    .B1(_1255_));
 sg13g2_o21ai_1 _3754_ (.B1(net773),
    .Y(_1256_),
    .A1(net817),
    .A2(net637));
 sg13g2_a21oi_1 _3755_ (.A1(net599),
    .A2(net637),
    .Y(_0317_),
    .B1(_1256_));
 sg13g2_o21ai_1 _3756_ (.B1(net773),
    .Y(_1257_),
    .A1(net803),
    .A2(_1249_));
 sg13g2_a21oi_1 _3757_ (.A1(net595),
    .A2(net637),
    .Y(_0318_),
    .B1(_1257_));
 sg13g2_nor2_1 _3758_ (.A(_1107_),
    .B(_1202_),
    .Y(_1258_));
 sg13g2_o21ai_1 _3759_ (.B1(net761),
    .Y(_1259_),
    .A1(net805),
    .A2(net635));
 sg13g2_a21oi_1 _3760_ (.A1(net622),
    .A2(net635),
    .Y(_0319_),
    .B1(_1259_));
 sg13g2_o21ai_1 _3761_ (.B1(net761),
    .Y(_1260_),
    .A1(net788),
    .A2(net635));
 sg13g2_a21oi_1 _3762_ (.A1(net625),
    .A2(net635),
    .Y(_0320_),
    .B1(_1260_));
 sg13g2_o21ai_1 _3763_ (.B1(net759),
    .Y(_1261_),
    .A1(net811),
    .A2(net634));
 sg13g2_a21oi_1 _3764_ (.A1(net619),
    .A2(net634),
    .Y(_0321_),
    .B1(_1261_));
 sg13g2_o21ai_1 _3765_ (.B1(net759),
    .Y(_1262_),
    .A1(net812),
    .A2(net634));
 sg13g2_a21oi_1 _3766_ (.A1(net613),
    .A2(net634),
    .Y(_0322_),
    .B1(_1262_));
 sg13g2_o21ai_1 _3767_ (.B1(net761),
    .Y(_1263_),
    .A1(net785),
    .A2(net635));
 sg13g2_a21oi_1 _3768_ (.A1(net604),
    .A2(net635),
    .Y(_0323_),
    .B1(_1263_));
 sg13g2_o21ai_1 _3769_ (.B1(net761),
    .Y(_1264_),
    .A1(net551),
    .A2(net635));
 sg13g2_a21oi_1 _3770_ (.A1(net607),
    .A2(net635),
    .Y(_0324_),
    .B1(_1264_));
 sg13g2_o21ai_1 _3771_ (.B1(net759),
    .Y(_1265_),
    .A1(net581),
    .A2(net634));
 sg13g2_a21oi_1 _3772_ (.A1(net597),
    .A2(net634),
    .Y(_0325_),
    .B1(_1265_));
 sg13g2_o21ai_1 _3773_ (.B1(net759),
    .Y(_1266_),
    .A1(net413),
    .A2(net634));
 sg13g2_a21oi_1 _3774_ (.A1(net594),
    .A2(net634),
    .Y(_0326_),
    .B1(_1266_));
 sg13g2_nor2_1 _3775_ (.A(_1097_),
    .B(_1202_),
    .Y(_1267_));
 sg13g2_o21ai_1 _3776_ (.B1(net766),
    .Y(_1268_),
    .A1(net540),
    .A2(net632));
 sg13g2_a21oi_1 _3777_ (.A1(net622),
    .A2(net632),
    .Y(_0327_),
    .B1(_1268_));
 sg13g2_o21ai_1 _3778_ (.B1(net767),
    .Y(_1269_),
    .A1(net519),
    .A2(net632));
 sg13g2_a21oi_1 _3779_ (.A1(net626),
    .A2(net632),
    .Y(_0328_),
    .B1(_1269_));
 sg13g2_o21ai_1 _3780_ (.B1(net756),
    .Y(_1270_),
    .A1(net403),
    .A2(net633));
 sg13g2_a21oi_1 _3781_ (.A1(net617),
    .A2(net633),
    .Y(_0329_),
    .B1(_1270_));
 sg13g2_o21ai_1 _3782_ (.B1(net766),
    .Y(_1271_),
    .A1(net550),
    .A2(_1267_));
 sg13g2_a21oi_1 _3783_ (.A1(net613),
    .A2(net632),
    .Y(_0330_),
    .B1(_1271_));
 sg13g2_o21ai_1 _3784_ (.B1(net766),
    .Y(_1272_),
    .A1(net411),
    .A2(net633));
 sg13g2_a21oi_1 _3785_ (.A1(net604),
    .A2(net632),
    .Y(_0331_),
    .B1(_1272_));
 sg13g2_o21ai_1 _3786_ (.B1(net766),
    .Y(_1273_),
    .A1(net544),
    .A2(net632));
 sg13g2_a21oi_1 _3787_ (.A1(net610),
    .A2(net632),
    .Y(_0332_),
    .B1(_1273_));
 sg13g2_o21ai_1 _3788_ (.B1(net760),
    .Y(_1274_),
    .A1(net443),
    .A2(net633));
 sg13g2_a21oi_1 _3789_ (.A1(net597),
    .A2(net633),
    .Y(_0333_),
    .B1(_1274_));
 sg13g2_o21ai_1 _3790_ (.B1(net752),
    .Y(_1275_),
    .A1(net437),
    .A2(net633));
 sg13g2_a21oi_1 _3791_ (.A1(net593),
    .A2(net633),
    .Y(_0334_),
    .B1(_1275_));
 sg13g2_dfrbp_1 _3792_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net17),
    .D(_0047_),
    .Q_N(_1875_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.stop_txn ));
 sg13g2_dfrbp_1 _3793_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net144),
    .D(_0048_),
    .Q_N(_1874_),
    .Q(\cpu_instance.ctrl_instance.reg_op ));
 sg13g2_dfrbp_1 _3794_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net143),
    .D(_0049_),
    .Q_N(_0026_),
    .Q(\cpu_instance.addr_reg_op[2] ));
 sg13g2_dfrbp_1 _3795_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net142),
    .D(net584),
    .Q_N(_1873_),
    .Q(\cpu_instance.addr_reg_op[1] ));
 sg13g2_dfrbp_1 _3796_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net18),
    .D(_0051_),
    .Q_N(_1876_),
    .Q(\cpu_instance.addr_reg_op[0] ));
 sg13g2_dfrbp_1 _3797_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net19),
    .D(_0000_),
    .Q_N(_1877_),
    .Q(\cpu_instance.ctrl_instance.mem_ctrl_op[0] ));
 sg13g2_dfrbp_1 _3798_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net20),
    .D(_0001_),
    .Q_N(_1878_),
    .Q(\cpu_instance.ctrl_instance.mem_ctrl_op[1] ));
 sg13g2_dfrbp_1 _3799_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net21),
    .D(_0002_),
    .Q_N(_1879_),
    .Q(\cpu_instance.ctrl_instance.mem_ctrl_op[2] ));
 sg13g2_dfrbp_1 _3800_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net22),
    .D(_0003_),
    .Q_N(_1880_),
    .Q(\cpu_instance.ctrl_instance.mux_sel[0] ));
 sg13g2_dfrbp_1 _3801_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net23),
    .D(_0004_),
    .Q_N(_1881_),
    .Q(\cpu_instance.ctrl_instance.mux_sel[1] ));
 sg13g2_dfrbp_1 _3802_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net24),
    .D(_0005_),
    .Q_N(_1882_),
    .Q(\cpu_instance.ctrl_instance.mux_sel[2] ));
 sg13g2_dfrbp_1 _3803_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net25),
    .D(_0014_),
    .Q_N(_1883_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.state[0] ));
 sg13g2_dfrbp_1 _3804_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net26),
    .D(_0015_),
    .Q_N(_1884_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.state[1] ));
 sg13g2_dfrbp_1 _3805_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net111),
    .D(_0016_),
    .Q_N(_1885_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.state[2] ));
 sg13g2_dfrbp_1 _3806_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net141),
    .D(_0017_),
    .Q_N(_0022_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.state[3] ));
 sg13g2_dfrbp_1 _3807_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net140),
    .D(net321),
    .Q_N(_1872_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.stop_txn_reg ));
 sg13g2_dfrbp_1 _3808_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net139),
    .D(_0053_),
    .Q_N(_1871_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[16] ));
 sg13g2_dfrbp_1 _3809_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net137),
    .D(_0054_),
    .Q_N(_1870_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[17] ));
 sg13g2_dfrbp_1 _3810_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net133),
    .D(_0055_),
    .Q_N(_1869_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[18] ));
 sg13g2_dfrbp_1 _3811_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net131),
    .D(_0056_),
    .Q_N(_1868_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[19] ));
 sg13g2_dfrbp_1 _3812_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net129),
    .D(_0057_),
    .Q_N(_1867_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[20] ));
 sg13g2_dfrbp_1 _3813_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net127),
    .D(_0058_),
    .Q_N(_1866_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[21] ));
 sg13g2_dfrbp_1 _3814_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net125),
    .D(_0059_),
    .Q_N(_1865_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[22] ));
 sg13g2_dfrbp_1 _3815_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net123),
    .D(net401),
    .Q_N(_1864_),
    .Q(\cpu_instance.ctrl_instance.jmp_op_addr_sel ));
 sg13g2_dfrbp_1 _3816_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net121),
    .D(_0061_),
    .Q_N(\cpu_instance.mem_instance.addr[24] ),
    .Q(\cpu_instance.addr_sel ));
 sg13g2_dfrbp_1 _3817_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net120),
    .D(_0062_),
    .Q_N(_1863_),
    .Q(\cpu_instance.ctrl_instance.reg_sel_1[0] ));
 sg13g2_dfrbp_1 _3818_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net110),
    .D(_0063_),
    .Q_N(_1862_),
    .Q(\cpu_instance.ctrl_instance.reg_sel_1[1] ));
 sg13g2_dfrbp_1 _3819_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net108),
    .D(_0064_),
    .Q_N(_1861_),
    .Q(\cpu_instance.ctrl_instance.reg_sel_in[0] ));
 sg13g2_dfrbp_1 _3820_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net106),
    .D(_0065_),
    .Q_N(_1860_),
    .Q(\cpu_instance.ctrl_instance.reg_sel_in[1] ));
 sg13g2_dfrbp_1 _3821_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net104),
    .D(net385),
    .Q_N(_1859_),
    .Q(\cpu_instance.ctrl_instance.flag_zero ));
 sg13g2_dfrbp_1 _3822_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net102),
    .D(net420),
    .Q_N(_1858_),
    .Q(\cpu_instance.ctrl_instance.flag_carry ));
 sg13g2_dfrbp_1 _3823_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net100),
    .D(net791),
    .Q_N(_1857_),
    .Q(\cpu_instance.alu_instance.op[0] ));
 sg13g2_dfrbp_1 _3824_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net98),
    .D(net794),
    .Q_N(_1856_),
    .Q(\cpu_instance.alu_instance.op[1] ));
 sg13g2_dfrbp_1 _3825_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net96),
    .D(net814),
    .Q_N(_1855_),
    .Q(\cpu_instance.alu_instance.op[2] ));
 sg13g2_dfrbp_1 _3826_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net94),
    .D(net808),
    .Q_N(_1854_),
    .Q(\cpu_instance.alu_instance.op[3] ));
 sg13g2_dfrbp_1 _3827_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net92),
    .D(net797),
    .Q_N(_1853_),
    .Q(\cpu_instance.ctrl_instance.use_register_bank_out_1 ));
 sg13g2_dfrbp_1 _3828_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net90),
    .D(_0073_),
    .Q_N(_1852_),
    .Q(\cpu_instance.ctrl_instance.use_register_bank_in ));
 sg13g2_dfrbp_1 _3829_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net88),
    .D(_0074_),
    .Q_N(_1851_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][0] ));
 sg13g2_dfrbp_1 _3830_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net86),
    .D(_0075_),
    .Q_N(_1850_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][1] ));
 sg13g2_dfrbp_1 _3831_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net84),
    .D(_0076_),
    .Q_N(_1849_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][2] ));
 sg13g2_dfrbp_1 _3832_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net82),
    .D(_0077_),
    .Q_N(_1848_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][3] ));
 sg13g2_dfrbp_1 _3833_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net80),
    .D(_0078_),
    .Q_N(_1847_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][4] ));
 sg13g2_dfrbp_1 _3834_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net78),
    .D(_0079_),
    .Q_N(_1846_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][5] ));
 sg13g2_dfrbp_1 _3835_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net76),
    .D(_0080_),
    .Q_N(_1845_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][6] ));
 sg13g2_dfrbp_1 _3836_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net74),
    .D(_0081_),
    .Q_N(_1844_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][7] ));
 sg13g2_dfrbp_1 _3837_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net72),
    .D(_0082_),
    .Q_N(_1843_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][8] ));
 sg13g2_dfrbp_1 _3838_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net70),
    .D(_0083_),
    .Q_N(_1842_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][9] ));
 sg13g2_dfrbp_1 _3839_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net68),
    .D(_0084_),
    .Q_N(_1841_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][10] ));
 sg13g2_dfrbp_1 _3840_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net66),
    .D(_0085_),
    .Q_N(_1840_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][11] ));
 sg13g2_dfrbp_1 _3841_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net64),
    .D(_0086_),
    .Q_N(_1839_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][12] ));
 sg13g2_dfrbp_1 _3842_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net62),
    .D(_0087_),
    .Q_N(_1838_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][13] ));
 sg13g2_dfrbp_1 _3843_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net60),
    .D(_0088_),
    .Q_N(_1837_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][14] ));
 sg13g2_dfrbp_1 _3844_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net58),
    .D(_0089_),
    .Q_N(_1836_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][15] ));
 sg13g2_dfrbp_1 _3845_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net56),
    .D(_0090_),
    .Q_N(_1835_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[0] ));
 sg13g2_dfrbp_1 _3846_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net55),
    .D(net554),
    .Q_N(_1834_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[1] ));
 sg13g2_dfrbp_1 _3847_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net54),
    .D(_0092_),
    .Q_N(_1833_),
    .Q(\cpu_instance.mem_instance.data_ready ));
 sg13g2_dfrbp_1 _3848_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net53),
    .D(_0093_),
    .Q_N(_1832_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[0] ));
 sg13g2_dfrbp_1 _3849_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net51),
    .D(_0094_),
    .Q_N(_1831_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[1] ));
 sg13g2_dfrbp_1 _3850_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net49),
    .D(_0095_),
    .Q_N(_1830_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[2] ));
 sg13g2_dfrbp_1 _3851_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net47),
    .D(net846),
    .Q_N(_1829_),
    .Q(\cpu_instance.mem_instance.data_req ));
 sg13g2_dfrbp_1 _3852_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net46),
    .D(_0097_),
    .Q_N(_1828_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[0] ));
 sg13g2_dfrbp_1 _3853_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net45),
    .D(_0098_),
    .Q_N(_1827_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[1] ));
 sg13g2_dfrbp_1 _3854_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net44),
    .D(_0099_),
    .Q_N(_1826_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[2] ));
 sg13g2_dfrbp_1 _3855_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net43),
    .D(_0100_),
    .Q_N(_1825_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[3] ));
 sg13g2_dfrbp_1 _3856_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net42),
    .D(_0101_),
    .Q_N(_0030_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[0] ));
 sg13g2_dfrbp_1 _3857_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net40),
    .D(_0102_),
    .Q_N(_1824_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[1] ));
 sg13g2_dfrbp_1 _3858_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net38),
    .D(_0103_),
    .Q_N(_0023_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[2] ));
 sg13g2_dfrbp_1 _3859_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net36),
    .D(net831),
    .Q_N(_0025_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.is_writing ));
 sg13g2_dfrbp_1 _3860_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net34),
    .D(net391),
    .Q_N(_1823_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_ram_a_select ));
 sg13g2_dfrbp_1 _3861_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net32),
    .D(net835),
    .Q_N(_1822_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ));
 sg13g2_dfrbp_1 _3862_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net30),
    .D(_0107_),
    .Q_N(_0024_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_clk_out ));
 sg13g2_dfrbp_1 _3863_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net28),
    .D(net323),
    .Q_N(_1821_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_data_oe[0] ));
 sg13g2_dfrbp_1 _3864_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net16),
    .D(net388),
    .Q_N(_1820_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[0] ));
 sg13g2_dfrbp_1 _3865_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net15),
    .D(_0110_),
    .Q_N(_1819_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[1] ));
 sg13g2_dfrbp_1 _3866_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net14),
    .D(_0111_),
    .Q_N(_1818_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[2] ));
 sg13g2_dfrbp_1 _3867_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net13),
    .D(_0112_),
    .Q_N(_1817_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[3] ));
 sg13g2_dfrbp_1 _3868_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net12),
    .D(_0113_),
    .Q_N(_1816_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[4] ));
 sg13g2_dfrbp_1 _3869_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net319),
    .D(net378),
    .Q_N(_1815_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[5] ));
 sg13g2_dfrbp_1 _3870_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net318),
    .D(net462),
    .Q_N(_1814_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[6] ));
 sg13g2_dfrbp_1 _3871_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net317),
    .D(net372),
    .Q_N(_1813_),
    .Q(\cpu_instance.mem_instance.data_qo_mi[7] ));
 sg13g2_dfrbp_1 _3872_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net316),
    .D(_0117_),
    .Q_N(_1812_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.last_ram_a_sel ));
 sg13g2_dfrbp_1 _3873_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net315),
    .D(_0118_),
    .Q_N(_1811_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[0] ));
 sg13g2_dfrbp_1 _3874_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net314),
    .D(_0119_),
    .Q_N(_1810_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[1] ));
 sg13g2_dfrbp_1 _3875_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net313),
    .D(_0120_),
    .Q_N(_1809_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[0] ));
 sg13g2_dfrbp_1 _3876_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net312),
    .D(_0121_),
    .Q_N(_1808_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[1] ));
 sg13g2_dfrbp_1 _3877_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net311),
    .D(_0122_),
    .Q_N(_1807_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[2] ));
 sg13g2_dfrbp_1 _3878_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net310),
    .D(_0123_),
    .Q_N(_1806_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[3] ));
 sg13g2_dfrbp_1 _3879_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net309),
    .D(net365),
    .Q_N(_1805_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[4] ));
 sg13g2_dfrbp_1 _3880_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net308),
    .D(_0125_),
    .Q_N(_1804_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[5] ));
 sg13g2_dfrbp_1 _3881_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net307),
    .D(net375),
    .Q_N(_1803_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[6] ));
 sg13g2_dfrbp_1 _3882_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net306),
    .D(net353),
    .Q_N(_1802_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[7] ));
 sg13g2_dfrbp_1 _3883_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net305),
    .D(_0128_),
    .Q_N(_1801_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[8] ));
 sg13g2_dfrbp_1 _3884_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net304),
    .D(_0129_),
    .Q_N(_1800_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[9] ));
 sg13g2_dfrbp_1 _3885_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net303),
    .D(_0130_),
    .Q_N(_1799_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[10] ));
 sg13g2_dfrbp_1 _3886_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net302),
    .D(_0131_),
    .Q_N(_1798_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[11] ));
 sg13g2_dfrbp_1 _3887_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net301),
    .D(net341),
    .Q_N(_1797_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[12] ));
 sg13g2_dfrbp_1 _3888_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net300),
    .D(net344),
    .Q_N(_1796_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[13] ));
 sg13g2_dfrbp_1 _3889_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net299),
    .D(net347),
    .Q_N(_1795_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[14] ));
 sg13g2_dfrbp_1 _3890_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net112),
    .D(net334),
    .Q_N(_1886_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[15] ));
 sg13g2_dfrbp_1 _3891_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net113),
    .D(_0006_),
    .Q_N(_1887_),
    .Q(\cpu_instance.ctrl_instance.state[0] ));
 sg13g2_dfrbp_1 _3892_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net114),
    .D(_0007_),
    .Q_N(_1888_),
    .Q(\cpu_instance.ctrl_instance.state[1] ));
 sg13g2_dfrbp_1 _3893_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net115),
    .D(_0008_),
    .Q_N(_1889_),
    .Q(\cpu_instance.ctrl_instance.state[2] ));
 sg13g2_dfrbp_1 _3894_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net116),
    .D(_0009_),
    .Q_N(_0028_),
    .Q(\cpu_instance.ctrl_instance.state[3] ));
 sg13g2_dfrbp_1 _3895_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net117),
    .D(_0010_),
    .Q_N(_1890_),
    .Q(\cpu_instance.ctrl_instance.state[4] ));
 sg13g2_dfrbp_1 _3896_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net118),
    .D(_0011_),
    .Q_N(_0027_),
    .Q(\cpu_instance.ctrl_instance.state[5] ));
 sg13g2_dfrbp_1 _3897_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net135),
    .D(_0012_),
    .Q_N(_1891_),
    .Q(\cpu_instance.ctrl_instance.state[6] ));
 sg13g2_dfrbp_1 _3898_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net298),
    .D(_0013_),
    .Q_N(_1794_),
    .Q(\cpu_instance.ctrl_instance.state[7] ));
 sg13g2_dfrbp_1 _3899_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net297),
    .D(_0136_),
    .Q_N(_1793_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][0] ));
 sg13g2_dfrbp_1 _3900_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net295),
    .D(_0137_),
    .Q_N(_1792_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][1] ));
 sg13g2_dfrbp_1 _3901_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net293),
    .D(_0138_),
    .Q_N(_1791_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][2] ));
 sg13g2_dfrbp_1 _3902_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net291),
    .D(_0139_),
    .Q_N(_1790_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][3] ));
 sg13g2_dfrbp_1 _3903_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net289),
    .D(_0140_),
    .Q_N(_1789_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][4] ));
 sg13g2_dfrbp_1 _3904_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net287),
    .D(_0141_),
    .Q_N(_1788_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][5] ));
 sg13g2_dfrbp_1 _3905_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net285),
    .D(_0142_),
    .Q_N(_1787_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][6] ));
 sg13g2_dfrbp_1 _3906_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net283),
    .D(_0143_),
    .Q_N(_1786_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][7] ));
 sg13g2_dfrbp_1 _3907_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net281),
    .D(_0144_),
    .Q_N(_1785_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][8] ));
 sg13g2_dfrbp_1 _3908_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net279),
    .D(_0145_),
    .Q_N(_1784_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][9] ));
 sg13g2_dfrbp_1 _3909_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net277),
    .D(_0146_),
    .Q_N(_1783_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][10] ));
 sg13g2_dfrbp_1 _3910_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net275),
    .D(_0147_),
    .Q_N(_1782_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][11] ));
 sg13g2_dfrbp_1 _3911_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net273),
    .D(_0148_),
    .Q_N(_1781_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][12] ));
 sg13g2_dfrbp_1 _3912_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net271),
    .D(_0149_),
    .Q_N(_1780_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][13] ));
 sg13g2_dfrbp_1 _3913_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net269),
    .D(_0150_),
    .Q_N(_1779_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][14] ));
 sg13g2_dfrbp_1 _3914_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net136),
    .D(_0151_),
    .Q_N(_1892_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][15] ));
 sg13g2_dfrbp_1 _3915_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net160),
    .D(_0018_),
    .Q_N(_1893_),
    .Q(_0335_));
 sg13g2_dfrbp_1 _3916_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net267),
    .D(_0019_),
    .Q_N(_1778_),
    .Q(_0336_));
 sg13g2_dfrbp_1 _3917_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net265),
    .D(_0152_),
    .Q_N(_1777_),
    .Q(\cpu_instance.ctrl_instance.reg_sel_2[0] ));
 sg13g2_dfrbp_1 _3918_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net264),
    .D(_0153_),
    .Q_N(_1776_),
    .Q(\cpu_instance.ctrl_instance.reg_sel_2[1] ));
 sg13g2_dfrbp_1 _3919_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net263),
    .D(_0154_),
    .Q_N(_1775_),
    .Q(\cpu_instance.mem_instance.bus_data_out[0] ));
 sg13g2_dfrbp_1 _3920_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net261),
    .D(_0155_),
    .Q_N(_1774_),
    .Q(\cpu_instance.mem_instance.bus_data_out[1] ));
 sg13g2_dfrbp_1 _3921_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net259),
    .D(_0156_),
    .Q_N(_1773_),
    .Q(\cpu_instance.mem_instance.bus_data_out[2] ));
 sg13g2_dfrbp_1 _3922_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net257),
    .D(_0157_),
    .Q_N(_1772_),
    .Q(\cpu_instance.mem_instance.bus_data_out[3] ));
 sg13g2_dfrbp_1 _3923_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net255),
    .D(_0158_),
    .Q_N(_1771_),
    .Q(\cpu_instance.mem_instance.bus_data_out[4] ));
 sg13g2_dfrbp_1 _3924_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net253),
    .D(_0159_),
    .Q_N(_1770_),
    .Q(\cpu_instance.mem_instance.bus_data_out[5] ));
 sg13g2_dfrbp_1 _3925_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net251),
    .D(_0160_),
    .Q_N(_1769_),
    .Q(\cpu_instance.mem_instance.bus_data_out[6] ));
 sg13g2_dfrbp_1 _3926_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net249),
    .D(_0161_),
    .Q_N(_1768_),
    .Q(\cpu_instance.mem_instance.bus_data_out[7] ));
 sg13g2_dfrbp_1 _3927_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net247),
    .D(net826),
    .Q_N(_1767_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.start_read ));
 sg13g2_dfrbp_1 _3928_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net246),
    .D(net829),
    .Q_N(_0021_),
    .Q(\cpu_instance.ctrl_instance.mem_op_done ));
 sg13g2_dfrbp_1 _3929_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net245),
    .D(_0164_),
    .Q_N(_1766_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.start_write ));
 sg13g2_dfrbp_1 _3930_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net244),
    .D(net370),
    .Q_N(_0029_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.stall_txn ));
 sg13g2_dfrbp_1 _3931_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net243),
    .D(_0166_),
    .Q_N(_1765_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[0] ));
 sg13g2_dfrbp_1 _3932_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net241),
    .D(_0167_),
    .Q_N(_1764_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[1] ));
 sg13g2_dfrbp_1 _3933_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net239),
    .D(_0168_),
    .Q_N(_1763_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[2] ));
 sg13g2_dfrbp_1 _3934_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net237),
    .D(_0169_),
    .Q_N(_1762_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[3] ));
 sg13g2_dfrbp_1 _3935_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net235),
    .D(_0170_),
    .Q_N(_1761_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[4] ));
 sg13g2_dfrbp_1 _3936_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net233),
    .D(_0171_),
    .Q_N(_1760_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[5] ));
 sg13g2_dfrbp_1 _3937_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net231),
    .D(_0172_),
    .Q_N(_1759_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[6] ));
 sg13g2_dfrbp_1 _3938_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net229),
    .D(_0173_),
    .Q_N(_1758_),
    .Q(\cpu_instance.mem_instance.data_qi_mo[7] ));
 sg13g2_dfrbp_1 _3939_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net227),
    .D(_0174_),
    .Q_N(_1757_),
    .Q(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[23] ));
 sg13g2_dfrbp_1 _3940_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net225),
    .D(_0175_),
    .Q_N(_1756_),
    .Q(\cpu_instance.registers_instance.register_bank[15][0] ));
 sg13g2_dfrbp_1 _3941_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net223),
    .D(_0176_),
    .Q_N(_1755_),
    .Q(\cpu_instance.registers_instance.register_bank[15][1] ));
 sg13g2_dfrbp_1 _3942_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net221),
    .D(_0177_),
    .Q_N(_1754_),
    .Q(\cpu_instance.registers_instance.register_bank[15][2] ));
 sg13g2_dfrbp_1 _3943_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net219),
    .D(_0178_),
    .Q_N(_1753_),
    .Q(\cpu_instance.registers_instance.register_bank[15][3] ));
 sg13g2_dfrbp_1 _3944_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net217),
    .D(_0179_),
    .Q_N(_1752_),
    .Q(\cpu_instance.registers_instance.register_bank[15][4] ));
 sg13g2_dfrbp_1 _3945_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net215),
    .D(_0180_),
    .Q_N(_1751_),
    .Q(\cpu_instance.registers_instance.register_bank[15][5] ));
 sg13g2_dfrbp_1 _3946_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net213),
    .D(_0181_),
    .Q_N(_1750_),
    .Q(\cpu_instance.registers_instance.register_bank[15][6] ));
 sg13g2_dfrbp_1 _3947_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net211),
    .D(_0182_),
    .Q_N(_1749_),
    .Q(\cpu_instance.registers_instance.register_bank[15][7] ));
 sg13g2_dfrbp_1 _3948_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net209),
    .D(_0183_),
    .Q_N(_1748_),
    .Q(\cpu_instance.registers_instance.register_bank[14][0] ));
 sg13g2_dfrbp_1 _3949_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net207),
    .D(_0184_),
    .Q_N(_1747_),
    .Q(\cpu_instance.registers_instance.register_bank[14][1] ));
 sg13g2_dfrbp_1 _3950_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net205),
    .D(_0185_),
    .Q_N(_1746_),
    .Q(\cpu_instance.registers_instance.register_bank[14][2] ));
 sg13g2_dfrbp_1 _3951_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net203),
    .D(_0186_),
    .Q_N(_1745_),
    .Q(\cpu_instance.registers_instance.register_bank[14][3] ));
 sg13g2_dfrbp_1 _3952_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net201),
    .D(_0187_),
    .Q_N(_1744_),
    .Q(\cpu_instance.registers_instance.register_bank[14][4] ));
 sg13g2_dfrbp_1 _3953_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net199),
    .D(_0188_),
    .Q_N(_1743_),
    .Q(\cpu_instance.registers_instance.register_bank[14][5] ));
 sg13g2_dfrbp_1 _3954_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net197),
    .D(_0189_),
    .Q_N(_1742_),
    .Q(\cpu_instance.registers_instance.register_bank[14][6] ));
 sg13g2_dfrbp_1 _3955_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net195),
    .D(_0190_),
    .Q_N(_1741_),
    .Q(\cpu_instance.registers_instance.register_bank[14][7] ));
 sg13g2_dfrbp_1 _3956_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net193),
    .D(_0191_),
    .Q_N(_1740_),
    .Q(\cpu_instance.registers_instance.register_bank[13][0] ));
 sg13g2_dfrbp_1 _3957_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net191),
    .D(_0192_),
    .Q_N(_1739_),
    .Q(\cpu_instance.registers_instance.register_bank[13][1] ));
 sg13g2_dfrbp_1 _3958_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net189),
    .D(_0193_),
    .Q_N(_1738_),
    .Q(\cpu_instance.registers_instance.register_bank[13][2] ));
 sg13g2_dfrbp_1 _3959_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net187),
    .D(_0194_),
    .Q_N(_1737_),
    .Q(\cpu_instance.registers_instance.register_bank[13][3] ));
 sg13g2_dfrbp_1 _3960_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net185),
    .D(_0195_),
    .Q_N(_1736_),
    .Q(\cpu_instance.registers_instance.register_bank[13][4] ));
 sg13g2_dfrbp_1 _3961_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net183),
    .D(_0196_),
    .Q_N(_1735_),
    .Q(\cpu_instance.registers_instance.register_bank[13][5] ));
 sg13g2_dfrbp_1 _3962_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net181),
    .D(_0197_),
    .Q_N(_1734_),
    .Q(\cpu_instance.registers_instance.register_bank[13][6] ));
 sg13g2_dfrbp_1 _3963_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net179),
    .D(_0198_),
    .Q_N(_1733_),
    .Q(\cpu_instance.registers_instance.register_bank[13][7] ));
 sg13g2_dfrbp_1 _3964_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net177),
    .D(_0199_),
    .Q_N(_1732_),
    .Q(\cpu_instance.registers_instance.register_bank[12][0] ));
 sg13g2_dfrbp_1 _3965_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net175),
    .D(_0200_),
    .Q_N(_1731_),
    .Q(\cpu_instance.registers_instance.register_bank[12][1] ));
 sg13g2_dfrbp_1 _3966_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net173),
    .D(_0201_),
    .Q_N(_1730_),
    .Q(\cpu_instance.registers_instance.register_bank[12][2] ));
 sg13g2_dfrbp_1 _3967_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net171),
    .D(_0202_),
    .Q_N(_1729_),
    .Q(\cpu_instance.registers_instance.register_bank[12][3] ));
 sg13g2_dfrbp_1 _3968_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net169),
    .D(_0203_),
    .Q_N(_1728_),
    .Q(\cpu_instance.registers_instance.register_bank[12][4] ));
 sg13g2_dfrbp_1 _3969_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net167),
    .D(_0204_),
    .Q_N(_1727_),
    .Q(\cpu_instance.registers_instance.register_bank[12][5] ));
 sg13g2_dfrbp_1 _3970_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net165),
    .D(_0205_),
    .Q_N(_1726_),
    .Q(\cpu_instance.registers_instance.register_bank[12][6] ));
 sg13g2_dfrbp_1 _3971_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net163),
    .D(_0206_),
    .Q_N(_1725_),
    .Q(\cpu_instance.registers_instance.register_bank[12][7] ));
 sg13g2_dfrbp_1 _3972_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net161),
    .D(_0207_),
    .Q_N(_1724_),
    .Q(\cpu_instance.registers_instance.register_bank[11][0] ));
 sg13g2_dfrbp_1 _3973_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net159),
    .D(_0208_),
    .Q_N(_1723_),
    .Q(\cpu_instance.registers_instance.register_bank[11][1] ));
 sg13g2_dfrbp_1 _3974_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net157),
    .D(_0209_),
    .Q_N(_1722_),
    .Q(\cpu_instance.registers_instance.register_bank[11][2] ));
 sg13g2_dfrbp_1 _3975_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net155),
    .D(_0210_),
    .Q_N(_1721_),
    .Q(\cpu_instance.registers_instance.register_bank[11][3] ));
 sg13g2_dfrbp_1 _3976_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net153),
    .D(_0211_),
    .Q_N(_1720_),
    .Q(\cpu_instance.registers_instance.register_bank[11][4] ));
 sg13g2_dfrbp_1 _3977_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net151),
    .D(_0212_),
    .Q_N(_1719_),
    .Q(\cpu_instance.registers_instance.register_bank[11][5] ));
 sg13g2_dfrbp_1 _3978_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net149),
    .D(_0213_),
    .Q_N(_1718_),
    .Q(\cpu_instance.registers_instance.register_bank[11][6] ));
 sg13g2_dfrbp_1 _3979_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net147),
    .D(_0214_),
    .Q_N(_1717_),
    .Q(\cpu_instance.registers_instance.register_bank[11][7] ));
 sg13g2_dfrbp_1 _3980_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net145),
    .D(_0215_),
    .Q_N(_1716_),
    .Q(\cpu_instance.registers_instance.register_bank[10][0] ));
 sg13g2_dfrbp_1 _3981_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net134),
    .D(_0216_),
    .Q_N(_1715_),
    .Q(\cpu_instance.registers_instance.register_bank[10][1] ));
 sg13g2_dfrbp_1 _3982_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net130),
    .D(_0217_),
    .Q_N(_1714_),
    .Q(\cpu_instance.registers_instance.register_bank[10][2] ));
 sg13g2_dfrbp_1 _3983_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net126),
    .D(_0218_),
    .Q_N(_1713_),
    .Q(\cpu_instance.registers_instance.register_bank[10][3] ));
 sg13g2_dfrbp_1 _3984_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net122),
    .D(_0219_),
    .Q_N(_1712_),
    .Q(\cpu_instance.registers_instance.register_bank[10][4] ));
 sg13g2_dfrbp_1 _3985_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net109),
    .D(_0220_),
    .Q_N(_1711_),
    .Q(\cpu_instance.registers_instance.register_bank[10][5] ));
 sg13g2_dfrbp_1 _3986_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net105),
    .D(_0221_),
    .Q_N(_1710_),
    .Q(\cpu_instance.registers_instance.register_bank[10][6] ));
 sg13g2_dfrbp_1 _3987_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net101),
    .D(_0222_),
    .Q_N(_1709_),
    .Q(\cpu_instance.registers_instance.register_bank[10][7] ));
 sg13g2_dfrbp_1 _3988_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net97),
    .D(_0223_),
    .Q_N(_1708_),
    .Q(\cpu_instance.registers_instance.register_bank[9][0] ));
 sg13g2_dfrbp_1 _3989_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net93),
    .D(_0224_),
    .Q_N(_1707_),
    .Q(\cpu_instance.registers_instance.register_bank[9][1] ));
 sg13g2_dfrbp_1 _3990_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net89),
    .D(_0225_),
    .Q_N(_1706_),
    .Q(\cpu_instance.registers_instance.register_bank[9][2] ));
 sg13g2_dfrbp_1 _3991_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net85),
    .D(_0226_),
    .Q_N(_1705_),
    .Q(\cpu_instance.registers_instance.register_bank[9][3] ));
 sg13g2_dfrbp_1 _3992_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net81),
    .D(_0227_),
    .Q_N(_1704_),
    .Q(\cpu_instance.registers_instance.register_bank[9][4] ));
 sg13g2_dfrbp_1 _3993_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net77),
    .D(_0228_),
    .Q_N(_1703_),
    .Q(\cpu_instance.registers_instance.register_bank[9][5] ));
 sg13g2_dfrbp_1 _3994_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net73),
    .D(_0229_),
    .Q_N(_1702_),
    .Q(\cpu_instance.registers_instance.register_bank[9][6] ));
 sg13g2_dfrbp_1 _3995_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net69),
    .D(_0230_),
    .Q_N(_1701_),
    .Q(\cpu_instance.registers_instance.register_bank[9][7] ));
 sg13g2_dfrbp_1 _3996_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net65),
    .D(_0231_),
    .Q_N(_1700_),
    .Q(\cpu_instance.registers_instance.register_bank[8][0] ));
 sg13g2_dfrbp_1 _3997_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net61),
    .D(_0232_),
    .Q_N(_1699_),
    .Q(\cpu_instance.registers_instance.register_bank[8][1] ));
 sg13g2_dfrbp_1 _3998_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net57),
    .D(_0233_),
    .Q_N(_1698_),
    .Q(\cpu_instance.registers_instance.register_bank[8][2] ));
 sg13g2_dfrbp_1 _3999_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net50),
    .D(_0234_),
    .Q_N(_1697_),
    .Q(\cpu_instance.registers_instance.register_bank[8][3] ));
 sg13g2_dfrbp_1 _4000_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net41),
    .D(_0235_),
    .Q_N(_1696_),
    .Q(\cpu_instance.registers_instance.register_bank[8][4] ));
 sg13g2_dfrbp_1 _4001_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net37),
    .D(_0236_),
    .Q_N(_1695_),
    .Q(\cpu_instance.registers_instance.register_bank[8][5] ));
 sg13g2_dfrbp_1 _4002_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net33),
    .D(_0237_),
    .Q_N(_1694_),
    .Q(\cpu_instance.registers_instance.register_bank[8][6] ));
 sg13g2_dfrbp_1 _4003_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net29),
    .D(_0238_),
    .Q_N(_1693_),
    .Q(\cpu_instance.registers_instance.register_bank[8][7] ));
 sg13g2_dfrbp_1 _4004_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net296),
    .D(_0239_),
    .Q_N(_1692_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[56] ));
 sg13g2_dfrbp_1 _4005_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net292),
    .D(_0240_),
    .Q_N(_1691_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[57] ));
 sg13g2_dfrbp_1 _4006_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net288),
    .D(_0241_),
    .Q_N(_1690_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[58] ));
 sg13g2_dfrbp_1 _4007_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net284),
    .D(_0242_),
    .Q_N(_1689_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[59] ));
 sg13g2_dfrbp_1 _4008_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net280),
    .D(_0243_),
    .Q_N(_1688_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[60] ));
 sg13g2_dfrbp_1 _4009_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net276),
    .D(_0244_),
    .Q_N(_1687_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[61] ));
 sg13g2_dfrbp_1 _4010_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net272),
    .D(_0245_),
    .Q_N(_1686_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[62] ));
 sg13g2_dfrbp_1 _4011_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net268),
    .D(_0246_),
    .Q_N(_1685_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[63] ));
 sg13g2_dfrbp_1 _4012_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net262),
    .D(_0247_),
    .Q_N(_1684_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[48] ));
 sg13g2_dfrbp_1 _4013_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net258),
    .D(_0248_),
    .Q_N(_1683_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[49] ));
 sg13g2_dfrbp_1 _4014_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net254),
    .D(_0249_),
    .Q_N(_1682_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[50] ));
 sg13g2_dfrbp_1 _4015_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net250),
    .D(_0250_),
    .Q_N(_1681_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[51] ));
 sg13g2_dfrbp_1 _4016_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net242),
    .D(_0251_),
    .Q_N(_1680_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[52] ));
 sg13g2_dfrbp_1 _4017_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net238),
    .D(_0252_),
    .Q_N(_1679_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[53] ));
 sg13g2_dfrbp_1 _4018_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net234),
    .D(_0253_),
    .Q_N(_1678_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[54] ));
 sg13g2_dfrbp_1 _4019_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net230),
    .D(_0254_),
    .Q_N(_1677_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[55] ));
 sg13g2_dfrbp_1 _4020_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net226),
    .D(_0255_),
    .Q_N(_1676_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[40] ));
 sg13g2_dfrbp_1 _4021_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net222),
    .D(_0256_),
    .Q_N(_1675_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[41] ));
 sg13g2_dfrbp_1 _4022_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net218),
    .D(_0257_),
    .Q_N(_1674_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[42] ));
 sg13g2_dfrbp_1 _4023_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net214),
    .D(_0258_),
    .Q_N(_1673_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[43] ));
 sg13g2_dfrbp_1 _4024_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net210),
    .D(_0259_),
    .Q_N(_1672_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[44] ));
 sg13g2_dfrbp_1 _4025_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net206),
    .D(_0260_),
    .Q_N(_1671_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[45] ));
 sg13g2_dfrbp_1 _4026_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net202),
    .D(_0261_),
    .Q_N(_1670_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[46] ));
 sg13g2_dfrbp_1 _4027_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net198),
    .D(_0262_),
    .Q_N(_1669_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[47] ));
 sg13g2_dfrbp_1 _4028_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net194),
    .D(_0263_),
    .Q_N(_1668_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[32] ));
 sg13g2_dfrbp_1 _4029_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net190),
    .D(_0264_),
    .Q_N(_1667_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[33] ));
 sg13g2_dfrbp_1 _4030_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net186),
    .D(_0265_),
    .Q_N(_1666_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[34] ));
 sg13g2_dfrbp_1 _4031_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net182),
    .D(_0266_),
    .Q_N(_1665_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[35] ));
 sg13g2_dfrbp_1 _4032_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net178),
    .D(_0267_),
    .Q_N(_1664_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[36] ));
 sg13g2_dfrbp_1 _4033_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net174),
    .D(_0268_),
    .Q_N(_1663_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[37] ));
 sg13g2_dfrbp_1 _4034_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net170),
    .D(_0269_),
    .Q_N(_1662_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[38] ));
 sg13g2_dfrbp_1 _4035_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net166),
    .D(_0270_),
    .Q_N(_1661_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[39] ));
 sg13g2_dfrbp_1 _4036_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net162),
    .D(_0271_),
    .Q_N(_1660_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[24] ));
 sg13g2_dfrbp_1 _4037_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net158),
    .D(_0272_),
    .Q_N(_1659_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[25] ));
 sg13g2_dfrbp_1 _4038_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net154),
    .D(_0273_),
    .Q_N(_1658_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[26] ));
 sg13g2_dfrbp_1 _4039_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net150),
    .D(_0274_),
    .Q_N(_1657_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[27] ));
 sg13g2_dfrbp_1 _4040_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net146),
    .D(_0275_),
    .Q_N(_1656_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[28] ));
 sg13g2_dfrbp_1 _4041_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net132),
    .D(_0276_),
    .Q_N(_1655_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[29] ));
 sg13g2_dfrbp_1 _4042_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net124),
    .D(_0277_),
    .Q_N(_1654_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[30] ));
 sg13g2_dfrbp_1 _4043_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net107),
    .D(_0278_),
    .Q_N(_1653_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[31] ));
 sg13g2_dfrbp_1 _4044_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net99),
    .D(_0279_),
    .Q_N(_0031_),
    .Q(\cpu_instance.registers_instance.registers[0][0] ));
 sg13g2_dfrbp_1 _4045_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net91),
    .D(_0280_),
    .Q_N(_0033_),
    .Q(\cpu_instance.registers_instance.registers[0][1] ));
 sg13g2_dfrbp_1 _4046_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net83),
    .D(_0281_),
    .Q_N(_0044_),
    .Q(\cpu_instance.registers_instance.registers[0][2] ));
 sg13g2_dfrbp_1 _4047_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net75),
    .D(_0282_),
    .Q_N(_0035_),
    .Q(\cpu_instance.registers_instance.registers[0][3] ));
 sg13g2_dfrbp_1 _4048_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net67),
    .D(_0283_),
    .Q_N(_0039_),
    .Q(\cpu_instance.registers_instance.registers[0][4] ));
 sg13g2_dfrbp_1 _4049_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net59),
    .D(_0284_),
    .Q_N(_0038_),
    .Q(\cpu_instance.registers_instance.registers[0][5] ));
 sg13g2_dfrbp_1 _4050_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net48),
    .D(_0285_),
    .Q_N(_0037_),
    .Q(\cpu_instance.registers_instance.registers[0][6] ));
 sg13g2_dfrbp_1 _4051_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net35),
    .D(_0286_),
    .Q_N(_0020_),
    .Q(\cpu_instance.registers_instance.registers[0][7] ));
 sg13g2_dfrbp_1 _4052_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net27),
    .D(_0287_),
    .Q_N(_1652_),
    .Q(\cpu_instance.registers_instance.registers[1][0] ));
 sg13g2_dfrbp_1 _4053_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net290),
    .D(_0288_),
    .Q_N(_1651_),
    .Q(\cpu_instance.registers_instance.registers[1][1] ));
 sg13g2_dfrbp_1 _4054_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net282),
    .D(_0289_),
    .Q_N(_1650_),
    .Q(\cpu_instance.registers_instance.registers[1][2] ));
 sg13g2_dfrbp_1 _4055_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net274),
    .D(_0290_),
    .Q_N(_1649_),
    .Q(\cpu_instance.registers_instance.registers[1][3] ));
 sg13g2_dfrbp_1 _4056_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net266),
    .D(_0291_),
    .Q_N(_1648_),
    .Q(\cpu_instance.registers_instance.registers[1][4] ));
 sg13g2_dfrbp_1 _4057_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net256),
    .D(_0292_),
    .Q_N(_1647_),
    .Q(\cpu_instance.registers_instance.registers[1][5] ));
 sg13g2_dfrbp_1 _4058_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net248),
    .D(_0293_),
    .Q_N(_1646_),
    .Q(\cpu_instance.registers_instance.registers[1][6] ));
 sg13g2_dfrbp_1 _4059_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net236),
    .D(_0294_),
    .Q_N(_1645_),
    .Q(\cpu_instance.registers_instance.registers[1][7] ));
 sg13g2_dfrbp_1 _4060_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net228),
    .D(_0295_),
    .Q_N(_1644_),
    .Q(\cpu_instance.registers_instance.registers[2][0] ));
 sg13g2_dfrbp_1 _4061_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net220),
    .D(_0296_),
    .Q_N(_1643_),
    .Q(\cpu_instance.registers_instance.registers[2][1] ));
 sg13g2_dfrbp_1 _4062_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net212),
    .D(_0297_),
    .Q_N(_1642_),
    .Q(\cpu_instance.registers_instance.registers[2][2] ));
 sg13g2_dfrbp_1 _4063_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net204),
    .D(_0298_),
    .Q_N(_1641_),
    .Q(\cpu_instance.registers_instance.registers[2][3] ));
 sg13g2_dfrbp_1 _4064_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net196),
    .D(_0299_),
    .Q_N(_1640_),
    .Q(\cpu_instance.registers_instance.registers[2][4] ));
 sg13g2_dfrbp_1 _4065_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net188),
    .D(_0300_),
    .Q_N(_1639_),
    .Q(\cpu_instance.registers_instance.registers[2][5] ));
 sg13g2_dfrbp_1 _4066_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net180),
    .D(_0301_),
    .Q_N(_1638_),
    .Q(\cpu_instance.registers_instance.registers[2][6] ));
 sg13g2_dfrbp_1 _4067_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net172),
    .D(_0302_),
    .Q_N(_1637_),
    .Q(\cpu_instance.registers_instance.registers[2][7] ));
 sg13g2_dfrbp_1 _4068_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net164),
    .D(_0303_),
    .Q_N(_0032_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _4069_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net156),
    .D(_0304_),
    .Q_N(_0034_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _4070_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net148),
    .D(_0305_),
    .Q_N(_1636_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _4071_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net128),
    .D(_0306_),
    .Q_N(_0036_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _4072_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net103),
    .D(_0307_),
    .Q_N(_0040_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _4073_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net87),
    .D(_0308_),
    .Q_N(_1635_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _4074_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net71),
    .D(_0309_),
    .Q_N(_1634_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _4075_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net52),
    .D(_0310_),
    .Q_N(_1633_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _4076_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net31),
    .D(_0311_),
    .Q_N(_0046_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[0] ));
 sg13g2_dfrbp_1 _4077_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net286),
    .D(_0312_),
    .Q_N(_0045_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[1] ));
 sg13g2_dfrbp_1 _4078_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net270),
    .D(_0313_),
    .Q_N(_0043_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[2] ));
 sg13g2_dfrbp_1 _4079_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net252),
    .D(_0314_),
    .Q_N(_0042_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[3] ));
 sg13g2_dfrbp_1 _4080_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net232),
    .D(_0315_),
    .Q_N(_0041_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[4] ));
 sg13g2_dfrbp_1 _4081_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net216),
    .D(_0316_),
    .Q_N(_1632_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[5] ));
 sg13g2_dfrbp_1 _4082_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net200),
    .D(_0317_),
    .Q_N(_1631_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[6] ));
 sg13g2_dfrbp_1 _4083_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net184),
    .D(_0318_),
    .Q_N(_1630_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[7] ));
 sg13g2_dfrbp_1 _4084_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net168),
    .D(_0319_),
    .Q_N(_1629_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[8] ));
 sg13g2_dfrbp_1 _4085_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net152),
    .D(_0320_),
    .Q_N(_1628_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[9] ));
 sg13g2_dfrbp_1 _4086_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net119),
    .D(_0321_),
    .Q_N(_1627_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[10] ));
 sg13g2_dfrbp_1 _4087_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net79),
    .D(_0322_),
    .Q_N(_1626_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[11] ));
 sg13g2_dfrbp_1 _4088_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net39),
    .D(_0323_),
    .Q_N(_1625_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[12] ));
 sg13g2_dfrbp_1 _4089_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net278),
    .D(_0324_),
    .Q_N(_1624_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[13] ));
 sg13g2_dfrbp_1 _4090_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net240),
    .D(_0325_),
    .Q_N(_1623_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[14] ));
 sg13g2_dfrbp_1 _4091_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net208),
    .D(_0326_),
    .Q_N(_1622_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[15] ));
 sg13g2_dfrbp_1 _4092_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net176),
    .D(_0327_),
    .Q_N(_1621_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[16] ));
 sg13g2_dfrbp_1 _4093_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net138),
    .D(_0328_),
    .Q_N(_1620_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[17] ));
 sg13g2_dfrbp_1 _4094_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net63),
    .D(_0329_),
    .Q_N(_1619_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[18] ));
 sg13g2_dfrbp_1 _4095_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net260),
    .D(_0330_),
    .Q_N(_1618_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[19] ));
 sg13g2_dfrbp_1 _4096_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net192),
    .D(_0331_),
    .Q_N(_1617_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[20] ));
 sg13g2_dfrbp_1 _4097_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net95),
    .D(_0332_),
    .Q_N(_1616_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[21] ));
 sg13g2_dfrbp_1 _4098_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net224),
    .D(_0333_),
    .Q_N(_1615_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[22] ));
 sg13g2_dfrbp_1 _4099_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net294),
    .D(_0334_),
    .Q_N(_1614_),
    .Q(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[23] ));
 sg13g2_tiehi _3867__13 (.L_HI(net13));
 sg13g2_tiehi _3866__14 (.L_HI(net14));
 sg13g2_tiehi _3865__15 (.L_HI(net15));
 sg13g2_tiehi _3864__16 (.L_HI(net16));
 sg13g2_tiehi _3792__17 (.L_HI(net17));
 sg13g2_tiehi _3796__18 (.L_HI(net18));
 sg13g2_tiehi _3797__19 (.L_HI(net19));
 sg13g2_tiehi _3798__20 (.L_HI(net20));
 sg13g2_tiehi _3799__21 (.L_HI(net21));
 sg13g2_tiehi _3800__22 (.L_HI(net22));
 sg13g2_tiehi _3801__23 (.L_HI(net23));
 sg13g2_tiehi _3802__24 (.L_HI(net24));
 sg13g2_tiehi _3803__25 (.L_HI(net25));
 sg13g2_tiehi _3804__26 (.L_HI(net26));
 sg13g2_tiehi _4052__27 (.L_HI(net27));
 sg13g2_tiehi _3863__28 (.L_HI(net28));
 sg13g2_tiehi _4003__29 (.L_HI(net29));
 sg13g2_tiehi _3862__30 (.L_HI(net30));
 sg13g2_tiehi _4076__31 (.L_HI(net31));
 sg13g2_tiehi _3861__32 (.L_HI(net32));
 sg13g2_tiehi _4002__33 (.L_HI(net33));
 sg13g2_tiehi _3860__34 (.L_HI(net34));
 sg13g2_tiehi _4051__35 (.L_HI(net35));
 sg13g2_tiehi _3859__36 (.L_HI(net36));
 sg13g2_tiehi _4001__37 (.L_HI(net37));
 sg13g2_tiehi _3858__38 (.L_HI(net38));
 sg13g2_tiehi _4088__39 (.L_HI(net39));
 sg13g2_tiehi _3857__40 (.L_HI(net40));
 sg13g2_tiehi _4000__41 (.L_HI(net41));
 sg13g2_tiehi _3856__42 (.L_HI(net42));
 sg13g2_tiehi _3855__43 (.L_HI(net43));
 sg13g2_tiehi _3854__44 (.L_HI(net44));
 sg13g2_tiehi _3853__45 (.L_HI(net45));
 sg13g2_tiehi _3852__46 (.L_HI(net46));
 sg13g2_tiehi _3851__47 (.L_HI(net47));
 sg13g2_tiehi _4050__48 (.L_HI(net48));
 sg13g2_tiehi _3850__49 (.L_HI(net49));
 sg13g2_tiehi _3999__50 (.L_HI(net50));
 sg13g2_tiehi _3849__51 (.L_HI(net51));
 sg13g2_tiehi _4075__52 (.L_HI(net52));
 sg13g2_tiehi _3848__53 (.L_HI(net53));
 sg13g2_tiehi _3847__54 (.L_HI(net54));
 sg13g2_tiehi _3846__55 (.L_HI(net55));
 sg13g2_tiehi _3845__56 (.L_HI(net56));
 sg13g2_tiehi _3998__57 (.L_HI(net57));
 sg13g2_tiehi _3844__58 (.L_HI(net58));
 sg13g2_tiehi _4049__59 (.L_HI(net59));
 sg13g2_tiehi _3843__60 (.L_HI(net60));
 sg13g2_tiehi _3997__61 (.L_HI(net61));
 sg13g2_tiehi _3842__62 (.L_HI(net62));
 sg13g2_tiehi _4094__63 (.L_HI(net63));
 sg13g2_tiehi _3841__64 (.L_HI(net64));
 sg13g2_tiehi _3996__65 (.L_HI(net65));
 sg13g2_tiehi _3840__66 (.L_HI(net66));
 sg13g2_tiehi _4048__67 (.L_HI(net67));
 sg13g2_tiehi _3839__68 (.L_HI(net68));
 sg13g2_tiehi _3995__69 (.L_HI(net69));
 sg13g2_tiehi _3838__70 (.L_HI(net70));
 sg13g2_tiehi _4074__71 (.L_HI(net71));
 sg13g2_tiehi _3837__72 (.L_HI(net72));
 sg13g2_tiehi _3994__73 (.L_HI(net73));
 sg13g2_tiehi _3836__74 (.L_HI(net74));
 sg13g2_tiehi _4047__75 (.L_HI(net75));
 sg13g2_tiehi _3835__76 (.L_HI(net76));
 sg13g2_tiehi _3993__77 (.L_HI(net77));
 sg13g2_tiehi _3834__78 (.L_HI(net78));
 sg13g2_tiehi _4087__79 (.L_HI(net79));
 sg13g2_tiehi _3833__80 (.L_HI(net80));
 sg13g2_tiehi _3992__81 (.L_HI(net81));
 sg13g2_tiehi _3832__82 (.L_HI(net82));
 sg13g2_tiehi _4046__83 (.L_HI(net83));
 sg13g2_tiehi _3831__84 (.L_HI(net84));
 sg13g2_tiehi _3991__85 (.L_HI(net85));
 sg13g2_tiehi _3830__86 (.L_HI(net86));
 sg13g2_tiehi _4073__87 (.L_HI(net87));
 sg13g2_tiehi _3829__88 (.L_HI(net88));
 sg13g2_tiehi _3990__89 (.L_HI(net89));
 sg13g2_tiehi _3828__90 (.L_HI(net90));
 sg13g2_tiehi _4045__91 (.L_HI(net91));
 sg13g2_tiehi _3827__92 (.L_HI(net92));
 sg13g2_tiehi _3989__93 (.L_HI(net93));
 sg13g2_tiehi _3826__94 (.L_HI(net94));
 sg13g2_tiehi _4097__95 (.L_HI(net95));
 sg13g2_tiehi _3825__96 (.L_HI(net96));
 sg13g2_tiehi _3988__97 (.L_HI(net97));
 sg13g2_tiehi _3824__98 (.L_HI(net98));
 sg13g2_tiehi _4044__99 (.L_HI(net99));
 sg13g2_tiehi _3823__100 (.L_HI(net100));
 sg13g2_tiehi _3987__101 (.L_HI(net101));
 sg13g2_tiehi _3822__102 (.L_HI(net102));
 sg13g2_tiehi _4072__103 (.L_HI(net103));
 sg13g2_tiehi _3821__104 (.L_HI(net104));
 sg13g2_tiehi _3986__105 (.L_HI(net105));
 sg13g2_tiehi _3820__106 (.L_HI(net106));
 sg13g2_tiehi _4043__107 (.L_HI(net107));
 sg13g2_tiehi _3819__108 (.L_HI(net108));
 sg13g2_tiehi _3985__109 (.L_HI(net109));
 sg13g2_tiehi _3818__110 (.L_HI(net110));
 sg13g2_tiehi _3805__111 (.L_HI(net111));
 sg13g2_tiehi _3890__112 (.L_HI(net112));
 sg13g2_tiehi _3891__113 (.L_HI(net113));
 sg13g2_tiehi _3892__114 (.L_HI(net114));
 sg13g2_tiehi _3893__115 (.L_HI(net115));
 sg13g2_tiehi _3894__116 (.L_HI(net116));
 sg13g2_tiehi _3895__117 (.L_HI(net117));
 sg13g2_tiehi _3896__118 (.L_HI(net118));
 sg13g2_tiehi _4086__119 (.L_HI(net119));
 sg13g2_tiehi _3817__120 (.L_HI(net120));
 sg13g2_tiehi _3816__121 (.L_HI(net121));
 sg13g2_tiehi _3984__122 (.L_HI(net122));
 sg13g2_tiehi _3815__123 (.L_HI(net123));
 sg13g2_tiehi _4042__124 (.L_HI(net124));
 sg13g2_tiehi _3814__125 (.L_HI(net125));
 sg13g2_tiehi _3983__126 (.L_HI(net126));
 sg13g2_tiehi _3813__127 (.L_HI(net127));
 sg13g2_tiehi _4071__128 (.L_HI(net128));
 sg13g2_tiehi _3812__129 (.L_HI(net129));
 sg13g2_tiehi _3982__130 (.L_HI(net130));
 sg13g2_tiehi _3811__131 (.L_HI(net131));
 sg13g2_tiehi _4041__132 (.L_HI(net132));
 sg13g2_tiehi _3810__133 (.L_HI(net133));
 sg13g2_tiehi _3981__134 (.L_HI(net134));
 sg13g2_tiehi _3897__135 (.L_HI(net135));
 sg13g2_tiehi _3914__136 (.L_HI(net136));
 sg13g2_tiehi _3809__137 (.L_HI(net137));
 sg13g2_tiehi _4093__138 (.L_HI(net138));
 sg13g2_tiehi _3808__139 (.L_HI(net139));
 sg13g2_tiehi _3807__140 (.L_HI(net140));
 sg13g2_tiehi _3806__141 (.L_HI(net141));
 sg13g2_tiehi _3795__142 (.L_HI(net142));
 sg13g2_tiehi _3794__143 (.L_HI(net143));
 sg13g2_tiehi _3793__144 (.L_HI(net144));
 sg13g2_tiehi _3980__145 (.L_HI(net145));
 sg13g2_tiehi _4040__146 (.L_HI(net146));
 sg13g2_tiehi _3979__147 (.L_HI(net147));
 sg13g2_tiehi _4070__148 (.L_HI(net148));
 sg13g2_tiehi _3978__149 (.L_HI(net149));
 sg13g2_tiehi _4039__150 (.L_HI(net150));
 sg13g2_tiehi _3977__151 (.L_HI(net151));
 sg13g2_tiehi _4085__152 (.L_HI(net152));
 sg13g2_tiehi _3976__153 (.L_HI(net153));
 sg13g2_tiehi _4038__154 (.L_HI(net154));
 sg13g2_tiehi _3975__155 (.L_HI(net155));
 sg13g2_tiehi _4069__156 (.L_HI(net156));
 sg13g2_tiehi _3974__157 (.L_HI(net157));
 sg13g2_tiehi _4037__158 (.L_HI(net158));
 sg13g2_tiehi _3973__159 (.L_HI(net159));
 sg13g2_tiehi _3915__160 (.L_HI(net160));
 sg13g2_tiehi _3972__161 (.L_HI(net161));
 sg13g2_tiehi _4036__162 (.L_HI(net162));
 sg13g2_tiehi _3971__163 (.L_HI(net163));
 sg13g2_tiehi _4068__164 (.L_HI(net164));
 sg13g2_tiehi _3970__165 (.L_HI(net165));
 sg13g2_tiehi _4035__166 (.L_HI(net166));
 sg13g2_tiehi _3969__167 (.L_HI(net167));
 sg13g2_tiehi _4084__168 (.L_HI(net168));
 sg13g2_tiehi _3968__169 (.L_HI(net169));
 sg13g2_tiehi _4034__170 (.L_HI(net170));
 sg13g2_tiehi _3967__171 (.L_HI(net171));
 sg13g2_tiehi _4067__172 (.L_HI(net172));
 sg13g2_tiehi _3966__173 (.L_HI(net173));
 sg13g2_tiehi _4033__174 (.L_HI(net174));
 sg13g2_tiehi _3965__175 (.L_HI(net175));
 sg13g2_tiehi _4092__176 (.L_HI(net176));
 sg13g2_tiehi _3964__177 (.L_HI(net177));
 sg13g2_tiehi _4032__178 (.L_HI(net178));
 sg13g2_tiehi _3963__179 (.L_HI(net179));
 sg13g2_tiehi _4066__180 (.L_HI(net180));
 sg13g2_tiehi _3962__181 (.L_HI(net181));
 sg13g2_tiehi _4031__182 (.L_HI(net182));
 sg13g2_tiehi _3961__183 (.L_HI(net183));
 sg13g2_tiehi _4083__184 (.L_HI(net184));
 sg13g2_tiehi _3960__185 (.L_HI(net185));
 sg13g2_tiehi _4030__186 (.L_HI(net186));
 sg13g2_tiehi _3959__187 (.L_HI(net187));
 sg13g2_tiehi _4065__188 (.L_HI(net188));
 sg13g2_tiehi _3958__189 (.L_HI(net189));
 sg13g2_tiehi _4029__190 (.L_HI(net190));
 sg13g2_tiehi _3957__191 (.L_HI(net191));
 sg13g2_tiehi _4096__192 (.L_HI(net192));
 sg13g2_tiehi _3956__193 (.L_HI(net193));
 sg13g2_tiehi _4028__194 (.L_HI(net194));
 sg13g2_tiehi _3955__195 (.L_HI(net195));
 sg13g2_tiehi _4064__196 (.L_HI(net196));
 sg13g2_tiehi _3954__197 (.L_HI(net197));
 sg13g2_tiehi _4027__198 (.L_HI(net198));
 sg13g2_tiehi _3953__199 (.L_HI(net199));
 sg13g2_tiehi _4082__200 (.L_HI(net200));
 sg13g2_tiehi _3952__201 (.L_HI(net201));
 sg13g2_tiehi _4026__202 (.L_HI(net202));
 sg13g2_tiehi _3951__203 (.L_HI(net203));
 sg13g2_tiehi _4063__204 (.L_HI(net204));
 sg13g2_tiehi _3950__205 (.L_HI(net205));
 sg13g2_tiehi _4025__206 (.L_HI(net206));
 sg13g2_tiehi _3949__207 (.L_HI(net207));
 sg13g2_tiehi _4091__208 (.L_HI(net208));
 sg13g2_tiehi _3948__209 (.L_HI(net209));
 sg13g2_tiehi _4024__210 (.L_HI(net210));
 sg13g2_tiehi _3947__211 (.L_HI(net211));
 sg13g2_tiehi _4062__212 (.L_HI(net212));
 sg13g2_tiehi _3946__213 (.L_HI(net213));
 sg13g2_tiehi _4023__214 (.L_HI(net214));
 sg13g2_tiehi _3945__215 (.L_HI(net215));
 sg13g2_tiehi _4081__216 (.L_HI(net216));
 sg13g2_tiehi _3944__217 (.L_HI(net217));
 sg13g2_tiehi _4022__218 (.L_HI(net218));
 sg13g2_tiehi _3943__219 (.L_HI(net219));
 sg13g2_tiehi _4061__220 (.L_HI(net220));
 sg13g2_tiehi _3942__221 (.L_HI(net221));
 sg13g2_tiehi _4021__222 (.L_HI(net222));
 sg13g2_tiehi _3941__223 (.L_HI(net223));
 sg13g2_tiehi _4098__224 (.L_HI(net224));
 sg13g2_tiehi _3940__225 (.L_HI(net225));
 sg13g2_tiehi _4020__226 (.L_HI(net226));
 sg13g2_tiehi _3939__227 (.L_HI(net227));
 sg13g2_tiehi _4060__228 (.L_HI(net228));
 sg13g2_tiehi _3938__229 (.L_HI(net229));
 sg13g2_tiehi _4019__230 (.L_HI(net230));
 sg13g2_tiehi _3937__231 (.L_HI(net231));
 sg13g2_tiehi _4080__232 (.L_HI(net232));
 sg13g2_tiehi _3936__233 (.L_HI(net233));
 sg13g2_tiehi _4018__234 (.L_HI(net234));
 sg13g2_tiehi _3935__235 (.L_HI(net235));
 sg13g2_tiehi _4059__236 (.L_HI(net236));
 sg13g2_tiehi _3934__237 (.L_HI(net237));
 sg13g2_tiehi _4017__238 (.L_HI(net238));
 sg13g2_tiehi _3933__239 (.L_HI(net239));
 sg13g2_tiehi _4090__240 (.L_HI(net240));
 sg13g2_tiehi _3932__241 (.L_HI(net241));
 sg13g2_tiehi _4016__242 (.L_HI(net242));
 sg13g2_tiehi _3931__243 (.L_HI(net243));
 sg13g2_tiehi _3930__244 (.L_HI(net244));
 sg13g2_tiehi _3929__245 (.L_HI(net245));
 sg13g2_tiehi _3928__246 (.L_HI(net246));
 sg13g2_tiehi _3927__247 (.L_HI(net247));
 sg13g2_tiehi _4058__248 (.L_HI(net248));
 sg13g2_tiehi _3926__249 (.L_HI(net249));
 sg13g2_tiehi _4015__250 (.L_HI(net250));
 sg13g2_tiehi _3925__251 (.L_HI(net251));
 sg13g2_tiehi _4079__252 (.L_HI(net252));
 sg13g2_tiehi _3924__253 (.L_HI(net253));
 sg13g2_tiehi _4014__254 (.L_HI(net254));
 sg13g2_tiehi _3923__255 (.L_HI(net255));
 sg13g2_tiehi _4057__256 (.L_HI(net256));
 sg13g2_tiehi _3922__257 (.L_HI(net257));
 sg13g2_tiehi _4013__258 (.L_HI(net258));
 sg13g2_tiehi _3921__259 (.L_HI(net259));
 sg13g2_tiehi _4095__260 (.L_HI(net260));
 sg13g2_tiehi _3920__261 (.L_HI(net261));
 sg13g2_tiehi _4012__262 (.L_HI(net262));
 sg13g2_tiehi _3919__263 (.L_HI(net263));
 sg13g2_tiehi _3918__264 (.L_HI(net264));
 sg13g2_tiehi _3917__265 (.L_HI(net265));
 sg13g2_tiehi _4056__266 (.L_HI(net266));
 sg13g2_tiehi _3916__267 (.L_HI(net267));
 sg13g2_tiehi _4011__268 (.L_HI(net268));
 sg13g2_tiehi _3913__269 (.L_HI(net269));
 sg13g2_tiehi _4078__270 (.L_HI(net270));
 sg13g2_tiehi _3912__271 (.L_HI(net271));
 sg13g2_tiehi _4010__272 (.L_HI(net272));
 sg13g2_tiehi _3911__273 (.L_HI(net273));
 sg13g2_tiehi _4055__274 (.L_HI(net274));
 sg13g2_tiehi _3910__275 (.L_HI(net275));
 sg13g2_tiehi _4009__276 (.L_HI(net276));
 sg13g2_tiehi _3909__277 (.L_HI(net277));
 sg13g2_tiehi _4089__278 (.L_HI(net278));
 sg13g2_tiehi _3908__279 (.L_HI(net279));
 sg13g2_tiehi _4008__280 (.L_HI(net280));
 sg13g2_tiehi _3907__281 (.L_HI(net281));
 sg13g2_tiehi _4054__282 (.L_HI(net282));
 sg13g2_tiehi _3906__283 (.L_HI(net283));
 sg13g2_tiehi _4007__284 (.L_HI(net284));
 sg13g2_tiehi _3905__285 (.L_HI(net285));
 sg13g2_tiehi _4077__286 (.L_HI(net286));
 sg13g2_tiehi _3904__287 (.L_HI(net287));
 sg13g2_tiehi _4006__288 (.L_HI(net288));
 sg13g2_tiehi _3903__289 (.L_HI(net289));
 sg13g2_tiehi _4053__290 (.L_HI(net290));
 sg13g2_tiehi _3902__291 (.L_HI(net291));
 sg13g2_tiehi _4005__292 (.L_HI(net292));
 sg13g2_tiehi _3901__293 (.L_HI(net293));
 sg13g2_tiehi _4099__294 (.L_HI(net294));
 sg13g2_tiehi _3900__295 (.L_HI(net295));
 sg13g2_tiehi _4004__296 (.L_HI(net296));
 sg13g2_tiehi _3899__297 (.L_HI(net297));
 sg13g2_tiehi _3898__298 (.L_HI(net298));
 sg13g2_tiehi _3889__299 (.L_HI(net299));
 sg13g2_tiehi _3888__300 (.L_HI(net300));
 sg13g2_tiehi _3887__301 (.L_HI(net301));
 sg13g2_tiehi _3886__302 (.L_HI(net302));
 sg13g2_tiehi _3885__303 (.L_HI(net303));
 sg13g2_tiehi _3884__304 (.L_HI(net304));
 sg13g2_tiehi _3883__305 (.L_HI(net305));
 sg13g2_tiehi _3882__306 (.L_HI(net306));
 sg13g2_tiehi _3881__307 (.L_HI(net307));
 sg13g2_tiehi _3880__308 (.L_HI(net308));
 sg13g2_tiehi _3879__309 (.L_HI(net309));
 sg13g2_tiehi _3878__310 (.L_HI(net310));
 sg13g2_tiehi _3877__311 (.L_HI(net311));
 sg13g2_tiehi _3876__312 (.L_HI(net312));
 sg13g2_tiehi _3875__313 (.L_HI(net313));
 sg13g2_tiehi _3874__314 (.L_HI(net314));
 sg13g2_tiehi _3873__315 (.L_HI(net315));
 sg13g2_tiehi _3872__316 (.L_HI(net316));
 sg13g2_tiehi _3871__317 (.L_HI(net317));
 sg13g2_tiehi _3870__318 (.L_HI(net318));
 sg13g2_tiehi _3869__319 (.L_HI(net319));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi _3868__12 (.L_HI(net12));
 sg13g2_buf_2 _4409_ (.A(net772),
    .X(uio_oe[0]));
 sg13g2_buf_1 _4410_ (.A(uio_oe[5]),
    .X(uio_oe[1]));
 sg13g2_buf_1 _4411_ (.A(uio_oe[5]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _4412_ (.A(net771),
    .X(uio_oe[3]));
 sg13g2_buf_1 _4413_ (.A(uio_oe[5]),
    .X(uio_oe[4]));
 sg13g2_buf_2 _4414_ (.A(net771),
    .X(uio_oe[6]));
 sg13g2_buf_2 _4415_ (.A(net771),
    .X(uio_oe[7]));
 sg13g2_buf_2 _4416_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ),
    .X(uio_out[0]));
 sg13g2_buf_2 _4417_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_clk_out ),
    .X(uio_out[3]));
 sg13g2_buf_2 _4418_ (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_ram_a_select ),
    .X(uio_out[6]));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(net590));
 sg13g2_buf_2 fanout590 (.A(_0716_),
    .X(net590));
 sg13g2_buf_4 fanout591 (.X(net591),
    .A(_0373_));
 sg13g2_buf_4 fanout592 (.X(net592),
    .A(net594));
 sg13g2_buf_2 fanout593 (.A(net594),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(net596),
    .X(net594));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(net596));
 sg13g2_buf_4 fanout596 (.X(net596),
    .A(_0372_));
 sg13g2_buf_2 fanout597 (.A(net599),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(net599),
    .X(net598));
 sg13g2_buf_4 fanout599 (.X(net599),
    .A(net601));
 sg13g2_buf_4 fanout600 (.X(net600),
    .A(net601));
 sg13g2_buf_2 fanout601 (.A(_0385_),
    .X(net601));
 sg13g2_buf_4 fanout602 (.X(net602),
    .A(_1583_));
 sg13g2_buf_4 fanout603 (.X(net603),
    .A(net604));
 sg13g2_buf_4 fanout604 (.X(net604),
    .A(net605));
 sg13g2_buf_4 fanout605 (.X(net605),
    .A(_1598_));
 sg13g2_buf_2 fanout606 (.A(net612),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(net612),
    .X(net607));
 sg13g2_buf_4 fanout608 (.X(net608),
    .A(net610));
 sg13g2_buf_2 fanout609 (.A(net610),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(net611),
    .X(net610));
 sg13g2_buf_4 fanout611 (.X(net611),
    .A(net612));
 sg13g2_buf_4 fanout612 (.X(net612),
    .A(_1582_));
 sg13g2_buf_4 fanout613 (.X(net613),
    .A(net615));
 sg13g2_buf_4 fanout614 (.X(net614),
    .A(net615));
 sg13g2_buf_8 fanout615 (.A(_0558_),
    .X(net615));
 sg13g2_buf_4 fanout616 (.X(net616),
    .A(_1599_));
 sg13g2_buf_2 fanout617 (.A(net618),
    .X(net617));
 sg13g2_buf_4 fanout618 (.X(net618),
    .A(net619));
 sg13g2_buf_2 fanout619 (.A(_0523_),
    .X(net619));
 sg13g2_buf_4 fanout620 (.X(net620),
    .A(_0523_));
 sg13g2_buf_2 fanout621 (.A(net624),
    .X(net621));
 sg13g2_buf_4 fanout622 (.X(net622),
    .A(net623));
 sg13g2_buf_4 fanout623 (.X(net623),
    .A(net624));
 sg13g2_buf_4 fanout624 (.X(net624),
    .A(_0538_));
 sg13g2_buf_4 fanout625 (.X(net625),
    .A(net626));
 sg13g2_buf_4 fanout626 (.X(net626),
    .A(net627));
 sg13g2_buf_4 fanout627 (.X(net627),
    .A(_0504_));
 sg13g2_buf_2 fanout628 (.A(_0989_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_0341_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(net631),
    .X(net630));
 sg13g2_buf_4 fanout631 (.X(net631),
    .A(_0988_));
 sg13g2_buf_2 fanout632 (.A(net633),
    .X(net632));
 sg13g2_buf_4 fanout633 (.X(net633),
    .A(_1267_));
 sg13g2_buf_2 fanout634 (.A(_1258_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_1258_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(net637),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_1249_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(net639),
    .X(net638));
 sg13g2_buf_4 fanout639 (.X(net639),
    .A(_1203_));
 sg13g2_buf_2 fanout640 (.A(net641),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_1193_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(net643),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(net644),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_1184_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_1175_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_1175_),
    .X(net646));
 sg13g2_buf_4 fanout647 (.X(net647),
    .A(net648));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(_1166_));
 sg13g2_buf_2 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_4 fanout650 (.X(net650),
    .A(_1155_));
 sg13g2_buf_2 fanout651 (.A(net652),
    .X(net651));
 sg13g2_buf_4 fanout652 (.X(net652),
    .A(_1146_));
 sg13g2_buf_4 fanout653 (.X(net653),
    .A(_1137_));
 sg13g2_buf_4 fanout654 (.X(net654),
    .A(_1137_));
 sg13g2_buf_2 fanout655 (.A(net657),
    .X(net655));
 sg13g2_buf_1 fanout656 (.A(net657),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_1128_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_1118_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_1118_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_4 fanout661 (.X(net661),
    .A(_1108_));
 sg13g2_buf_2 fanout662 (.A(net663),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_1098_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net665),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_1088_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_0998_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_0996_),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(_0891_),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(_0891_),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(net671),
    .X(net670));
 sg13g2_buf_4 fanout671 (.X(net671),
    .A(_0946_));
 sg13g2_buf_2 fanout672 (.A(net673),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(net674),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_0946_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_0616_),
    .X(net675));
 sg13g2_buf_1 fanout676 (.A(_0616_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_0615_),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(net680),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_0613_),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(net682),
    .X(net681));
 sg13g2_buf_1 fanout682 (.A(net683),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_0613_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(net685),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(_0485_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(_1069_),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(net688),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_0483_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_0478_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(_0477_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_0477_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_1 fanout693 (.A(net694),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_1240_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_1231_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(net698),
    .X(net697));
 sg13g2_buf_4 fanout698 (.X(net698),
    .A(_1222_));
 sg13g2_buf_2 fanout699 (.A(_1213_),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(_1213_),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(net703),
    .X(net701));
 sg13g2_buf_1 fanout702 (.A(net703),
    .X(net702));
 sg13g2_buf_1 fanout703 (.A(_0609_),
    .X(net703));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(_1361_));
 sg13g2_buf_4 fanout705 (.X(net705),
    .A(_1358_));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(_1343_));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(_0626_));
 sg13g2_buf_2 fanout708 (.A(net709),
    .X(net708));
 sg13g2_buf_1 fanout709 (.A(net710),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(net711),
    .X(net710));
 sg13g2_buf_4 fanout711 (.X(net711),
    .A(_0618_));
 sg13g2_buf_2 fanout712 (.A(net713),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(_0445_),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(_1404_),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(_1316_),
    .X(net715));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(_1289_));
 sg13g2_buf_2 fanout717 (.A(net718),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(net586),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(\cpu_instance.ctrl_instance.state[3] ),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(net845),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.is_writing ),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(net839),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(net836),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[0] ),
    .X(net724));
 sg13g2_buf_4 fanout725 (.X(net725),
    .A(\cpu_instance.ctrl_instance.use_register_bank_out_1 ));
 sg13g2_buf_2 fanout726 (.A(net728),
    .X(net726));
 sg13g2_buf_1 fanout727 (.A(net728),
    .X(net727));
 sg13g2_buf_1 fanout728 (.A(net729),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(net852),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(net732),
    .X(net730));
 sg13g2_buf_1 fanout731 (.A(net732),
    .X(net731));
 sg13g2_buf_1 fanout732 (.A(net733),
    .X(net732));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(net848));
 sg13g2_buf_4 fanout734 (.X(net734),
    .A(net736));
 sg13g2_buf_2 fanout735 (.A(net736),
    .X(net735));
 sg13g2_buf_4 fanout736 (.X(net736),
    .A(net737));
 sg13g2_buf_2 fanout737 (.A(\cpu_instance.addr_sel ),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(net740),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(net740),
    .X(net739));
 sg13g2_buf_1 fanout740 (.A(net742),
    .X(net740));
 sg13g2_buf_4 fanout741 (.X(net741),
    .A(net742));
 sg13g2_buf_1 fanout742 (.A(_1303_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(net747),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(net747),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(net747),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(net747),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(rst_n),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(net750),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(net750),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(net758),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(net752),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(net758),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(net755),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(net755),
    .X(net754));
 sg13g2_buf_1 fanout755 (.A(net758),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(net758),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(net758),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(net768),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(net762),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(net762),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(net762),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(net768),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(net765),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(net765),
    .X(net764));
 sg13g2_buf_1 fanout765 (.A(net768),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(net767),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(net768),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(rst_n),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(net770),
    .X(net769));
 sg13g2_buf_4 fanout770 (.X(net770),
    .A(net772));
 sg13g2_buf_4 fanout771 (.X(net771),
    .A(net772));
 sg13g2_buf_2 fanout772 (.A(net780),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(net775),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_1 fanout775 (.A(net780),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(net777),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(net780),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(net779),
    .X(net778));
 sg13g2_buf_4 fanout779 (.X(net779),
    .A(net780));
 sg13g2_buf_4 fanout780 (.X(net780),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[4]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[5]),
    .X(net10));
 sg13g2_tielo tt_um_strau0106_simple_viii_11 (.L_LO(net11));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_39_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_41_clk));
 sg13g2_inv_8 clkload8 (.A(clknet_leaf_23_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_27_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_5_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_14_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_7_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_8_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_10_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_20_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.stop_txn ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0052_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold3 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_data_oe[0] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0108_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold5 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[19] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0490_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold7 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[23] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold8 (.A(\cpu_instance.ctrl_instance.state[1] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold9 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[16] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0487_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold11 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[18] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0489_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold13 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[0] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold14 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[11] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0135_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold16 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[17] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0488_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold18 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[0] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold19 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[2] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold20 (.A(\cpu_instance.mem_instance.data_qi_mo[5] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold21 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[8] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0132_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold23 (.A(\cpu_instance.mem_instance.data_qi_mo[3] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold24 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[9] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0133_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold26 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[3] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold27 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[10] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0134_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold29 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[1] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold30 (.A(\cpu_instance.mem_instance.data_qi_mo[6] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold31 (.A(_1077_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold32 (.A(\cpu_instance.mem_instance.data_qi_mo[4] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold33 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[3] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0127_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold35 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_ram_a_select ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold36 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[20] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold37 (.A(\cpu_instance.ctrl_instance.state[6] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold38 (.A(\cpu_instance.mem_instance.data_qi_mo[1] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold39 (.A(\cpu_instance.mem_instance.data_qi_mo[2] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0022_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold41 (.A(_1068_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold42 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][3] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0652_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold44 (.A(\cpu_instance.mem_instance.data_qi_mo[7] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold45 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[4] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0124_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold47 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[1] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold48 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[5] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold49 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_in_buffer[2] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold50 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.state[0] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0165_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold52 (.A(\cpu_instance.mem_instance.data_qo_mi[7] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0116_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold54 (.A(\cpu_instance.mem_instance.data_qi_mo[0] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold55 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[6] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0126_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold57 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[21] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold58 (.A(\cpu_instance.mem_instance.data_qo_mi[5] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0114_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold60 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][8] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold61 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][5] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold62 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][10] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold63 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[7] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold64 (.A(\cpu_instance.registers_instance.registers[0][3] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold65 (.A(\cpu_instance.ctrl_instance.flag_zero ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0066_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold67 (.A(\cpu_instance.registers_instance.registers[0][4] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold68 (.A(\cpu_instance.mem_instance.data_qo_mi[0] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0109_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold70 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.addr[22] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.stop_txn_reg ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0105_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold73 (.A(\cpu_instance.mem_instance.addr[24] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold74 (.A(\cpu_instance.ctrl_instance.use_register_bank_in ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold75 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][6] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold76 (.A(\cpu_instance.ctrl_instance.state[4] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold77 (.A(\cpu_instance.registers_instance.register_bank[15][6] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold78 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[53] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold79 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][14] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold80 (.A(\cpu_instance.mem_instance.data_qo_mi[4] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold81 (.A(\cpu_instance.ctrl_instance.jmp_op_addr_sel ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0060_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold83 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[52] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold84 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[18] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold85 (.A(\cpu_instance.registers_instance.register_bank[12][0] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold86 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][2] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold87 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[27] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold88 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[34] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold89 (.A(\cpu_instance.registers_instance.register_bank[15][3] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cpu_instance.registers_instance.register_bank[14][7] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold91 (.A(\cpu_instance.registers_instance.register_bank[14][1] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold92 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[20] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold93 (.A(\cpu_instance.registers_instance.register_bank[11][5] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold94 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[15] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[36] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold96 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[54] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold97 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[47] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold98 (.A(\cpu_instance.registers_instance.register_bank[10][5] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold99 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[38] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold100 (.A(\cpu_instance.ctrl_instance.flag_carry ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0067_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][4] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold103 (.A(\cpu_instance.registers_instance.register_bank[9][6] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cpu_instance.registers_instance.register_bank[10][4] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold105 (.A(\cpu_instance.registers_instance.register_bank[10][0] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cpu_instance.registers_instance.register_bank[12][1] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold107 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][0] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][5] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold109 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[33] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold110 (.A(\cpu_instance.mem_instance.bus_data_out[7] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold111 (.A(\cpu_instance.registers_instance.register_bank[11][4] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold112 (.A(\cpu_instance.registers_instance.register_bank[14][3] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold113 (.A(\cpu_instance.registers_instance.register_bank[8][4] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold114 (.A(\cpu_instance.registers_instance.register_bank[14][4] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold115 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[43] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold116 (.A(\cpu_instance.registers_instance.register_bank[15][4] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold117 (.A(\cpu_instance.registers_instance.register_bank[8][2] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[23] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold119 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[25] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold120 (.A(\cpu_instance.registers_instance.register_bank[9][3] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold121 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][0] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold122 (.A(\cpu_instance.registers_instance.register_bank[15][1] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold123 (.A(\cpu_instance.registers_instance.register_bank[10][3] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[22] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold125 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[30] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold126 (.A(\cpu_instance.ctrl_instance.state[2] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold127 (.A(\cpu_instance.registers_instance.register_bank[8][1] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold128 (.A(\cpu_instance.registers_instance.register_bank[14][0] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold129 (.A(\cpu_instance.registers_instance.register_bank[8][3] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold130 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[45] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold131 (.A(\cpu_instance.registers_instance.register_bank[12][5] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold132 (.A(\cpu_instance.registers_instance.register_bank[10][7] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold133 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[58] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold134 (.A(\cpu_instance.registers_instance.register_bank[9][7] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold135 (.A(\cpu_instance.registers_instance.register_bank[9][1] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold136 (.A(\cpu_instance.registers_instance.register_bank[13][4] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold137 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[39] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold138 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[61] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold139 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][11] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold140 (.A(\cpu_instance.registers_instance.register_bank[12][4] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold141 (.A(\cpu_instance.registers_instance.register_bank[13][2] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold142 (.A(\cpu_instance.mem_instance.data_qo_mi[6] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0115_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold144 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][13] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold145 (.A(\cpu_instance.registers_instance.register_bank[9][5] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold146 (.A(\cpu_instance.registers_instance.register_bank[13][1] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold147 (.A(\cpu_instance.mem_instance.bus_data_out[6] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold148 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[63] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][8] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold150 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[44] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold151 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[41] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[48] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold153 (.A(\cpu_instance.registers_instance.register_bank[8][5] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold154 (.A(\cpu_instance.registers_instance.registers[0][6] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cpu_instance.registers_instance.register_bank[11][0] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold156 (.A(\cpu_instance.registers_instance.register_bank[14][6] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold157 (.A(\cpu_instance.registers_instance.register_bank[10][6] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold158 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][12] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold159 (.A(\cpu_instance.registers_instance.registers[1][4] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold160 (.A(_1227_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold161 (.A(\cpu_instance.registers_instance.register_bank[12][6] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold162 (.A(\cpu_instance.registers_instance.register_bank[11][1] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold163 (.A(\cpu_instance.registers_instance.register_bank[14][5] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold164 (.A(\cpu_instance.registers_instance.register_bank[10][2] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold165 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[35] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold166 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[28] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold167 (.A(\cpu_instance.registers_instance.register_bank[11][6] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold168 (.A(\cpu_instance.registers_instance.register_bank[9][0] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold169 (.A(\cpu_instance.registers_instance.register_bank[15][5] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold170 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[0] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold171 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[24] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold172 (.A(\cpu_instance.registers_instance.register_bank[13][3] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold173 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][9] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold174 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][1] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold175 (.A(\cpu_instance.registers_instance.register_bank[13][0] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold176 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[37] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold177 (.A(\cpu_instance.mem_instance.bus_data_out[5] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold178 (.A(\cpu_instance.registers_instance.register_bank[9][2] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold179 (.A(\cpu_instance.registers_instance.register_bank[15][0] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold180 (.A(\cpu_instance.registers_instance.register_bank[8][7] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold181 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[2] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold182 (.A(\cpu_instance.registers_instance.register_bank[12][7] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold183 (.A(\cpu_instance.registers_instance.register_bank[15][2] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold184 (.A(\cpu_instance.mem_instance.data_qo_mi[3] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold185 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[56] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold186 (.A(\cpu_instance.ctrl_instance.state[0] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0409_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold188 (.A(\cpu_instance.registers_instance.register_bank[11][3] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold189 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][11] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0027_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold191 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][13] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold192 (.A(\cpu_instance.registers_instance.register_bank[8][6] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold193 (.A(\cpu_instance.registers_instance.register_bank[13][6] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold194 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[31] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold195 (.A(\cpu_instance.registers_instance.register_bank[13][5] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold196 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][15] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold197 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[3] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold198 (.A(\cpu_instance.registers_instance.register_bank[9][4] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold199 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][3] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold200 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[17] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold201 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][2] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold202 (.A(\cpu_instance.registers_instance.registers[1][5] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold203 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[57] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold204 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[42] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold205 (.A(\cpu_instance.registers_instance.register_bank[13][7] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold206 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[49] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0028_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0569_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0570_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold210 (.A(\cpu_instance.registers_instance.register_bank[14][2] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold211 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][6] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold212 (.A(\cpu_instance.registers_instance.register_bank[15][7] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold213 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[60] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold214 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[0] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold215 (.A(\cpu_instance.registers_instance.register_bank[11][7] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold216 (.A(\cpu_instance.mem_instance.data_qo_mi[1] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold217 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[55] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold218 (.A(\cpu_instance.registers_instance.registers[2][4] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold219 (.A(_1236_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold220 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[59] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold221 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[16] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold222 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][14] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold223 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][7] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold224 (.A(\cpu_instance.registers_instance.register_bank[11][2] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold225 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[21] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold226 (.A(\cpu_instance.mem_instance.data_qo_mi[2] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold227 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[46] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold228 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[2] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold229 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][9] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold230 (.A(\cpu_instance.registers_instance.register_bank[12][2] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold231 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[19] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold232 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[13] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold233 (.A(\cpu_instance.registers_instance.registers[2][6] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold234 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.delay_cycles_cfg[1] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0091_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold236 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[50] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold237 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[29] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold238 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.state[3] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0421_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold240 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[26] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold241 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[51] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold242 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[1] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0840_),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold244 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][12] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold245 (.A(\cpu_instance.mem_instance.bus_data_out[4] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold246 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][4] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold247 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][1] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold248 (.A(\cpu_instance.registers_instance.register_bank[10][1] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold249 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][15] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold250 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[62] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold251 (.A(\cpu_instance.ctrl_instance.state[5] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold252 (.A(\cpu_instance.registers_instance.registers[1][6] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold253 (.A(\cpu_instance.mem_instance.bus_data_out[3] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold254 (.A(\cpu_instance.registers_instance.register_bank[12][3] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold255 (.A(\cpu_instance.mem_instance.bus_data_out[2] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold256 (.A(\cpu_instance.registers_instance.register_bank[8][0] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold257 (.A(uo_out[4]),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold258 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][10] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold259 (.A(\cpu_instance.registers_instance.registers[0][5] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold260 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[32] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold261 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[4] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold262 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[14] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold263 (.A(uo_out[3]),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0021_),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0050_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold266 (.A(\cpu_instance.ctrl_instance.state[7] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold267 (.A(\cpu_instance.ctrl_instance.mem_op_done ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold268 (.A(\cpu_instance.registers_instance.registers[1][7] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold269 (.A(\cpu_instance.mem_instance.bus_data_out[0] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold270 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[5] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold271 (.A(\cpu_instance.mem_instance.bus_data_out[1] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold272 (.A(\cpu_instance.registers_instance.registers[0][7] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold273 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[40] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold274 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[12] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold275 (.A(\cpu_instance.registers_instance.registers[0][1] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold276 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[0][7] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold277 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[9] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold278 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_clk_out ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold279 (.A(\cpu_instance.alu_instance.op[0] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0068_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold281 (.A(\cpu_instance.registers_instance.registers[2][5] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold282 (.A(\cpu_instance.alu_instance.op[1] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0069_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold284 (.A(\cpu_instance.registers_instance.registers[0][2] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold285 (.A(\cpu_instance.ctrl_instance.use_register_bank_out_1 ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0072_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold287 (.A(\cpu_instance.ctrl_instance.mem_ctrl_op[1] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0416_),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0424_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold290 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[1] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold291 (.A(\cpu_instance.registers_instance.registers[0][0] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold292 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[7] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold293 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.read_cycles_count[0] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold294 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[8] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold295 (.A(\cpu_instance.registers_instance.registers[2][7] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold296 (.A(\cpu_instance.alu_instance.op[3] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0071_),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold298 (.A(\cpu_instance.ctrl_instance.reg_sel_in[1] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold299 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.nibbles_remaining[0] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold300 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[10] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold301 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[11] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold302 (.A(\cpu_instance.alu_instance.op[2] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0070_),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold304 (.A(\cpu_instance.registers_instance.registers[1][0] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold305 (.A(\cpu_instance.mem_instance.data_req ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold306 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.register_bank_in[6] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold307 (.A(\cpu_instance.registers_instance.registers[1][3] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold308 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.state[1] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0429_),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold310 (.A(\cpu_instance.registers_instance.registers[2][3] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold311 (.A(\cpu_instance.ctrl_instance.state[5] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold312 (.A(\cpu_instance.registers_instance.registers[2][0] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold313 (.A(\cpu_instance.registers_instance.registers[1][1] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold314 (.A(\cpu_instance.ctrl_instance.mem_ctrl_op[2] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0162_),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold316 (.A(\cpu_instance.mem_instance.data_ready ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0428_),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0163_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold319 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.start_read ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0104_),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold321 (.A(\cpu_instance.ctrl_instance.state[7] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold322 (.A(\cpu_instance.registers_instance.registers[2][1] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold323 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.spi_flash_select ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0106_),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold325 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[1] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold326 (.A(uo_out[6]),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold327 (.A(\cpu_instance.ctrl_instance.state[3] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold328 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.fsm_state[2] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold329 (.A(uo_out[7]),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold330 (.A(\cpu_instance.registers_instance.registers[2][2] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold331 (.A(uo_out[1]),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold332 (.A(uo_out[5]),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold333 (.A(\cpu_instance.registers_instance.registers[1][2] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold334 (.A(\cpu_instance.mem_instance.qspi_ctrl_instance.is_writing ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0096_),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold336 (.A(\cpu_instance.ctrl_instance.state[0] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold337 (.A(\cpu_instance.ctrl_instance.reg_sel_1[0] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold338 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.stall_txn ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold339 (.A(uo_out[0]),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold340 (.A(uo_out[2]),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold341 (.A(\cpu_instance.ctrl_instance.reg_sel_1[1] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0021_),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold343 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.state[1] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold344 (.A(\cpu_instance.mem_instance.mem_ctrl_instance.addrs[1][10] ),
    .X(net855));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_fill_1 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_297 ();
 sg13g2_fill_1 FILLER_0_304 ();
 sg13g2_fill_1 FILLER_0_340 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_fill_2 FILLER_1_259 ();
 sg13g2_fill_1 FILLER_1_261 ();
 sg13g2_fill_1 FILLER_1_288 ();
 sg13g2_fill_1 FILLER_1_294 ();
 sg13g2_fill_2 FILLER_1_326 ();
 sg13g2_fill_1 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_4 FILLER_2_252 ();
 sg13g2_fill_2 FILLER_2_256 ();
 sg13g2_fill_2 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_4 FILLER_3_259 ();
 sg13g2_fill_1 FILLER_3_272 ();
 sg13g2_fill_2 FILLER_3_278 ();
 sg13g2_fill_2 FILLER_3_303 ();
 sg13g2_fill_1 FILLER_3_305 ();
 sg13g2_fill_2 FILLER_3_320 ();
 sg13g2_fill_1 FILLER_3_322 ();
 sg13g2_fill_1 FILLER_3_349 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_4 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_4 FILLER_4_266 ();
 sg13g2_fill_2 FILLER_4_270 ();
 sg13g2_fill_2 FILLER_4_276 ();
 sg13g2_fill_2 FILLER_4_283 ();
 sg13g2_fill_1 FILLER_4_285 ();
 sg13g2_fill_2 FILLER_4_341 ();
 sg13g2_fill_1 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_386 ();
 sg13g2_decap_8 FILLER_4_393 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_fill_2 FILLER_5_273 ();
 sg13g2_fill_1 FILLER_5_305 ();
 sg13g2_fill_2 FILLER_5_349 ();
 sg13g2_fill_1 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_4 FILLER_6_245 ();
 sg13g2_fill_1 FILLER_6_249 ();
 sg13g2_fill_2 FILLER_6_311 ();
 sg13g2_fill_2 FILLER_6_328 ();
 sg13g2_fill_1 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_decap_8 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_4 FILLER_7_245 ();
 sg13g2_fill_2 FILLER_7_275 ();
 sg13g2_fill_1 FILLER_7_277 ();
 sg13g2_fill_2 FILLER_7_297 ();
 sg13g2_fill_1 FILLER_7_299 ();
 sg13g2_fill_1 FILLER_7_315 ();
 sg13g2_fill_2 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_fill_2 FILLER_8_260 ();
 sg13g2_fill_1 FILLER_8_262 ();
 sg13g2_fill_2 FILLER_8_283 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_149 ();
 sg13g2_decap_8 FILLER_9_156 ();
 sg13g2_decap_8 FILLER_9_163 ();
 sg13g2_decap_8 FILLER_9_170 ();
 sg13g2_decap_8 FILLER_9_177 ();
 sg13g2_decap_8 FILLER_9_184 ();
 sg13g2_decap_8 FILLER_9_191 ();
 sg13g2_decap_8 FILLER_9_198 ();
 sg13g2_decap_8 FILLER_9_205 ();
 sg13g2_decap_8 FILLER_9_212 ();
 sg13g2_decap_8 FILLER_9_219 ();
 sg13g2_decap_8 FILLER_9_226 ();
 sg13g2_decap_8 FILLER_9_233 ();
 sg13g2_decap_8 FILLER_9_240 ();
 sg13g2_decap_4 FILLER_9_252 ();
 sg13g2_fill_2 FILLER_9_256 ();
 sg13g2_decap_8 FILLER_9_267 ();
 sg13g2_decap_8 FILLER_9_274 ();
 sg13g2_fill_1 FILLER_9_281 ();
 sg13g2_fill_1 FILLER_9_313 ();
 sg13g2_fill_2 FILLER_9_328 ();
 sg13g2_fill_2 FILLER_9_360 ();
 sg13g2_fill_1 FILLER_9_362 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_fill_1 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_4 FILLER_10_238 ();
 sg13g2_fill_1 FILLER_10_298 ();
 sg13g2_fill_2 FILLER_10_368 ();
 sg13g2_fill_1 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_fill_1 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_decap_8 FILLER_11_179 ();
 sg13g2_decap_8 FILLER_11_186 ();
 sg13g2_decap_8 FILLER_11_193 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_221 ();
 sg13g2_decap_8 FILLER_11_228 ();
 sg13g2_decap_4 FILLER_11_235 ();
 sg13g2_fill_2 FILLER_11_239 ();
 sg13g2_fill_2 FILLER_11_267 ();
 sg13g2_fill_1 FILLER_11_269 ();
 sg13g2_decap_4 FILLER_11_294 ();
 sg13g2_fill_2 FILLER_11_302 ();
 sg13g2_fill_1 FILLER_11_304 ();
 sg13g2_fill_2 FILLER_11_339 ();
 sg13g2_fill_1 FILLER_11_349 ();
 sg13g2_fill_2 FILLER_11_364 ();
 sg13g2_fill_1 FILLER_11_366 ();
 sg13g2_decap_4 FILLER_11_383 ();
 sg13g2_fill_1 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_fill_1 FILLER_12_98 ();
 sg13g2_fill_2 FILLER_12_125 ();
 sg13g2_decap_8 FILLER_12_164 ();
 sg13g2_decap_8 FILLER_12_171 ();
 sg13g2_decap_8 FILLER_12_178 ();
 sg13g2_decap_8 FILLER_12_185 ();
 sg13g2_decap_8 FILLER_12_192 ();
 sg13g2_decap_8 FILLER_12_199 ();
 sg13g2_decap_8 FILLER_12_206 ();
 sg13g2_decap_8 FILLER_12_213 ();
 sg13g2_decap_8 FILLER_12_220 ();
 sg13g2_decap_8 FILLER_12_227 ();
 sg13g2_decap_8 FILLER_12_234 ();
 sg13g2_decap_8 FILLER_12_241 ();
 sg13g2_decap_4 FILLER_12_248 ();
 sg13g2_fill_2 FILLER_12_265 ();
 sg13g2_fill_1 FILLER_12_267 ();
 sg13g2_decap_4 FILLER_12_303 ();
 sg13g2_fill_1 FILLER_12_307 ();
 sg13g2_decap_4 FILLER_12_313 ();
 sg13g2_fill_2 FILLER_12_317 ();
 sg13g2_decap_4 FILLER_12_328 ();
 sg13g2_fill_1 FILLER_12_344 ();
 sg13g2_fill_2 FILLER_12_350 ();
 sg13g2_fill_1 FILLER_12_352 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_fill_2 FILLER_13_91 ();
 sg13g2_fill_2 FILLER_13_136 ();
 sg13g2_fill_1 FILLER_13_138 ();
 sg13g2_decap_8 FILLER_13_179 ();
 sg13g2_decap_8 FILLER_13_186 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_decap_8 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_214 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_235 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_decap_4 FILLER_13_249 ();
 sg13g2_decap_4 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_fill_1 FILLER_14_112 ();
 sg13g2_fill_2 FILLER_14_132 ();
 sg13g2_decap_8 FILLER_14_183 ();
 sg13g2_decap_8 FILLER_14_190 ();
 sg13g2_decap_8 FILLER_14_197 ();
 sg13g2_decap_8 FILLER_14_204 ();
 sg13g2_decap_8 FILLER_14_211 ();
 sg13g2_decap_8 FILLER_14_218 ();
 sg13g2_decap_8 FILLER_14_225 ();
 sg13g2_decap_8 FILLER_14_232 ();
 sg13g2_decap_4 FILLER_14_239 ();
 sg13g2_fill_1 FILLER_14_243 ();
 sg13g2_fill_1 FILLER_14_275 ();
 sg13g2_fill_2 FILLER_14_286 ();
 sg13g2_fill_1 FILLER_14_288 ();
 sg13g2_fill_2 FILLER_14_339 ();
 sg13g2_fill_1 FILLER_14_341 ();
 sg13g2_fill_2 FILLER_14_351 ();
 sg13g2_fill_1 FILLER_14_353 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_4 FILLER_15_70 ();
 sg13g2_fill_1 FILLER_15_74 ();
 sg13g2_decap_8 FILLER_15_101 ();
 sg13g2_decap_4 FILLER_15_108 ();
 sg13g2_fill_2 FILLER_15_116 ();
 sg13g2_decap_4 FILLER_15_123 ();
 sg13g2_fill_2 FILLER_15_127 ();
 sg13g2_decap_8 FILLER_15_134 ();
 sg13g2_decap_4 FILLER_15_141 ();
 sg13g2_fill_1 FILLER_15_145 ();
 sg13g2_decap_4 FILLER_15_150 ();
 sg13g2_decap_8 FILLER_15_200 ();
 sg13g2_decap_8 FILLER_15_207 ();
 sg13g2_decap_8 FILLER_15_214 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_4 FILLER_15_235 ();
 sg13g2_fill_2 FILLER_15_283 ();
 sg13g2_fill_1 FILLER_15_285 ();
 sg13g2_fill_1 FILLER_15_310 ();
 sg13g2_fill_1 FILLER_15_317 ();
 sg13g2_fill_1 FILLER_15_348 ();
 sg13g2_fill_1 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_4 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_100 ();
 sg13g2_fill_2 FILLER_16_146 ();
 sg13g2_decap_8 FILLER_16_209 ();
 sg13g2_decap_8 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_230 ();
 sg13g2_decap_8 FILLER_16_237 ();
 sg13g2_fill_2 FILLER_16_244 ();
 sg13g2_fill_1 FILLER_16_246 ();
 sg13g2_fill_2 FILLER_16_256 ();
 sg13g2_decap_8 FILLER_16_288 ();
 sg13g2_fill_2 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_4 FILLER_17_63 ();
 sg13g2_fill_1 FILLER_17_90 ();
 sg13g2_fill_2 FILLER_17_128 ();
 sg13g2_fill_1 FILLER_17_254 ();
 sg13g2_fill_2 FILLER_17_265 ();
 sg13g2_fill_2 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_fill_2 FILLER_18_77 ();
 sg13g2_fill_1 FILLER_18_79 ();
 sg13g2_fill_2 FILLER_18_108 ();
 sg13g2_fill_1 FILLER_18_126 ();
 sg13g2_fill_2 FILLER_18_167 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_fill_1 FILLER_18_190 ();
 sg13g2_fill_2 FILLER_18_202 ();
 sg13g2_fill_1 FILLER_18_204 ();
 sg13g2_decap_4 FILLER_18_231 ();
 sg13g2_fill_2 FILLER_18_283 ();
 sg13g2_fill_1 FILLER_18_285 ();
 sg13g2_decap_4 FILLER_18_301 ();
 sg13g2_fill_1 FILLER_18_305 ();
 sg13g2_fill_1 FILLER_18_342 ();
 sg13g2_fill_2 FILLER_18_349 ();
 sg13g2_fill_2 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_fill_1 FILLER_19_70 ();
 sg13g2_fill_2 FILLER_19_120 ();
 sg13g2_fill_1 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_156 ();
 sg13g2_fill_2 FILLER_19_175 ();
 sg13g2_fill_2 FILLER_19_236 ();
 sg13g2_decap_8 FILLER_19_275 ();
 sg13g2_fill_1 FILLER_19_282 ();
 sg13g2_decap_8 FILLER_19_297 ();
 sg13g2_fill_2 FILLER_19_304 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_fill_2 FILLER_19_317 ();
 sg13g2_fill_2 FILLER_19_328 ();
 sg13g2_fill_2 FILLER_19_339 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_70 ();
 sg13g2_fill_2 FILLER_20_108 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_decap_4 FILLER_20_119 ();
 sg13g2_fill_1 FILLER_20_123 ();
 sg13g2_fill_1 FILLER_20_138 ();
 sg13g2_fill_1 FILLER_20_151 ();
 sg13g2_decap_4 FILLER_20_156 ();
 sg13g2_fill_2 FILLER_20_160 ();
 sg13g2_fill_2 FILLER_20_181 ();
 sg13g2_fill_1 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_decap_4 FILLER_20_195 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_260 ();
 sg13g2_fill_1 FILLER_20_271 ();
 sg13g2_fill_2 FILLER_20_276 ();
 sg13g2_fill_1 FILLER_20_278 ();
 sg13g2_decap_8 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_fill_2 FILLER_20_362 ();
 sg13g2_fill_2 FILLER_20_388 ();
 sg13g2_fill_1 FILLER_20_390 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_fill_2 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_112 ();
 sg13g2_fill_1 FILLER_21_114 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_fill_1 FILLER_21_146 ();
 sg13g2_fill_2 FILLER_21_157 ();
 sg13g2_fill_1 FILLER_21_164 ();
 sg13g2_decap_4 FILLER_21_213 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_decap_4 FILLER_21_227 ();
 sg13g2_fill_1 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_258 ();
 sg13g2_fill_1 FILLER_21_260 ();
 sg13g2_fill_1 FILLER_21_297 ();
 sg13g2_fill_1 FILLER_21_304 ();
 sg13g2_fill_1 FILLER_21_331 ();
 sg13g2_fill_2 FILLER_21_338 ();
 sg13g2_fill_1 FILLER_21_340 ();
 sg13g2_fill_2 FILLER_21_346 ();
 sg13g2_fill_1 FILLER_21_348 ();
 sg13g2_fill_2 FILLER_21_379 ();
 sg13g2_fill_1 FILLER_21_381 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_fill_2 FILLER_22_91 ();
 sg13g2_fill_1 FILLER_22_93 ();
 sg13g2_fill_2 FILLER_22_99 ();
 sg13g2_fill_1 FILLER_22_108 ();
 sg13g2_fill_2 FILLER_22_147 ();
 sg13g2_fill_2 FILLER_22_164 ();
 sg13g2_fill_1 FILLER_22_166 ();
 sg13g2_fill_2 FILLER_22_217 ();
 sg13g2_decap_4 FILLER_22_232 ();
 sg13g2_fill_2 FILLER_22_236 ();
 sg13g2_fill_1 FILLER_22_246 ();
 sg13g2_fill_1 FILLER_22_293 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_4 FILLER_23_70 ();
 sg13g2_fill_1 FILLER_23_74 ();
 sg13g2_decap_4 FILLER_23_84 ();
 sg13g2_fill_1 FILLER_23_106 ();
 sg13g2_fill_2 FILLER_23_122 ();
 sg13g2_fill_2 FILLER_23_132 ();
 sg13g2_fill_2 FILLER_23_142 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_fill_2 FILLER_23_152 ();
 sg13g2_fill_1 FILLER_23_154 ();
 sg13g2_fill_2 FILLER_23_174 ();
 sg13g2_fill_1 FILLER_23_176 ();
 sg13g2_fill_1 FILLER_23_193 ();
 sg13g2_decap_4 FILLER_23_247 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_fill_1 FILLER_23_324 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_fill_2 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_86 ();
 sg13g2_fill_2 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_138 ();
 sg13g2_fill_2 FILLER_24_188 ();
 sg13g2_fill_2 FILLER_24_239 ();
 sg13g2_fill_1 FILLER_24_302 ();
 sg13g2_fill_2 FILLER_24_326 ();
 sg13g2_fill_1 FILLER_24_328 ();
 sg13g2_fill_1 FILLER_24_335 ();
 sg13g2_fill_1 FILLER_24_355 ();
 sg13g2_fill_2 FILLER_24_366 ();
 sg13g2_fill_1 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_63 ();
 sg13g2_fill_2 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_111 ();
 sg13g2_decap_4 FILLER_25_118 ();
 sg13g2_fill_2 FILLER_25_122 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_207 ();
 sg13g2_decap_4 FILLER_25_237 ();
 sg13g2_fill_1 FILLER_25_241 ();
 sg13g2_fill_2 FILLER_25_258 ();
 sg13g2_fill_2 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_118 ();
 sg13g2_decap_4 FILLER_26_125 ();
 sg13g2_fill_2 FILLER_26_129 ();
 sg13g2_fill_2 FILLER_26_135 ();
 sg13g2_fill_1 FILLER_26_137 ();
 sg13g2_fill_2 FILLER_26_142 ();
 sg13g2_fill_1 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_150 ();
 sg13g2_fill_2 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_177 ();
 sg13g2_fill_2 FILLER_26_223 ();
 sg13g2_fill_1 FILLER_26_225 ();
 sg13g2_fill_2 FILLER_26_326 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_fill_2 FILLER_26_352 ();
 sg13g2_fill_1 FILLER_26_354 ();
 sg13g2_fill_1 FILLER_26_381 ();
 sg13g2_fill_1 FILLER_26_396 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_4 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_67 ();
 sg13g2_fill_1 FILLER_27_86 ();
 sg13g2_decap_8 FILLER_27_113 ();
 sg13g2_fill_2 FILLER_27_120 ();
 sg13g2_fill_1 FILLER_27_122 ();
 sg13g2_decap_8 FILLER_27_134 ();
 sg13g2_fill_2 FILLER_27_141 ();
 sg13g2_decap_4 FILLER_27_181 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_decap_8 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_260 ();
 sg13g2_fill_2 FILLER_27_286 ();
 sg13g2_fill_1 FILLER_27_288 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_297 ();
 sg13g2_fill_1 FILLER_27_332 ();
 sg13g2_fill_1 FILLER_27_368 ();
 sg13g2_fill_2 FILLER_27_380 ();
 sg13g2_fill_1 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_4 FILLER_28_77 ();
 sg13g2_fill_2 FILLER_28_81 ();
 sg13g2_fill_2 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_decap_8 FILLER_28_181 ();
 sg13g2_decap_4 FILLER_28_188 ();
 sg13g2_fill_2 FILLER_28_192 ();
 sg13g2_decap_8 FILLER_28_198 ();
 sg13g2_decap_8 FILLER_28_205 ();
 sg13g2_fill_2 FILLER_28_212 ();
 sg13g2_decap_8 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_226 ();
 sg13g2_fill_2 FILLER_28_268 ();
 sg13g2_fill_2 FILLER_28_306 ();
 sg13g2_fill_2 FILLER_28_371 ();
 sg13g2_fill_1 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_4 FILLER_29_56 ();
 sg13g2_fill_1 FILLER_29_60 ();
 sg13g2_fill_1 FILLER_29_87 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_fill_1 FILLER_29_154 ();
 sg13g2_fill_2 FILLER_29_174 ();
 sg13g2_fill_1 FILLER_29_191 ();
 sg13g2_fill_2 FILLER_29_202 ();
 sg13g2_decap_4 FILLER_29_219 ();
 sg13g2_fill_2 FILLER_29_231 ();
 sg13g2_fill_1 FILLER_29_342 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_1 FILLER_30_92 ();
 sg13g2_fill_2 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_157 ();
 sg13g2_fill_2 FILLER_30_169 ();
 sg13g2_fill_1 FILLER_30_171 ();
 sg13g2_fill_2 FILLER_30_196 ();
 sg13g2_fill_1 FILLER_30_198 ();
 sg13g2_fill_1 FILLER_30_302 ();
 sg13g2_decap_4 FILLER_30_320 ();
 sg13g2_fill_1 FILLER_30_324 ();
 sg13g2_fill_2 FILLER_30_330 ();
 sg13g2_fill_1 FILLER_30_332 ();
 sg13g2_fill_1 FILLER_30_342 ();
 sg13g2_fill_2 FILLER_30_348 ();
 sg13g2_fill_2 FILLER_30_356 ();
 sg13g2_fill_2 FILLER_30_372 ();
 sg13g2_fill_1 FILLER_30_374 ();
 sg13g2_fill_1 FILLER_30_386 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_4 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_60 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_fill_1 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_113 ();
 sg13g2_fill_1 FILLER_31_135 ();
 sg13g2_fill_1 FILLER_31_148 ();
 sg13g2_fill_2 FILLER_31_168 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_decap_4 FILLER_31_225 ();
 sg13g2_fill_1 FILLER_31_234 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_fill_1 FILLER_31_246 ();
 sg13g2_fill_2 FILLER_31_252 ();
 sg13g2_fill_2 FILLER_31_263 ();
 sg13g2_fill_2 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_278 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_decap_8 FILLER_31_320 ();
 sg13g2_fill_2 FILLER_31_380 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_fill_2 FILLER_32_70 ();
 sg13g2_fill_1 FILLER_32_76 ();
 sg13g2_fill_2 FILLER_32_126 ();
 sg13g2_fill_2 FILLER_32_153 ();
 sg13g2_fill_2 FILLER_32_163 ();
 sg13g2_fill_2 FILLER_32_170 ();
 sg13g2_fill_1 FILLER_32_172 ();
 sg13g2_fill_2 FILLER_32_178 ();
 sg13g2_fill_1 FILLER_32_180 ();
 sg13g2_fill_2 FILLER_32_189 ();
 sg13g2_fill_1 FILLER_32_191 ();
 sg13g2_decap_4 FILLER_32_197 ();
 sg13g2_decap_8 FILLER_32_220 ();
 sg13g2_fill_1 FILLER_32_227 ();
 sg13g2_fill_1 FILLER_32_233 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_4 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_268 ();
 sg13g2_decap_4 FILLER_32_275 ();
 sg13g2_decap_4 FILLER_32_283 ();
 sg13g2_fill_1 FILLER_32_287 ();
 sg13g2_fill_1 FILLER_32_297 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_350 ();
 sg13g2_fill_2 FILLER_32_387 ();
 sg13g2_fill_1 FILLER_32_389 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_4 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_60 ();
 sg13g2_fill_2 FILLER_33_87 ();
 sg13g2_fill_1 FILLER_33_124 ();
 sg13g2_decap_4 FILLER_33_147 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_fill_2 FILLER_33_160 ();
 sg13g2_fill_1 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_decap_4 FILLER_33_186 ();
 sg13g2_decap_4 FILLER_33_195 ();
 sg13g2_fill_2 FILLER_33_199 ();
 sg13g2_fill_2 FILLER_33_210 ();
 sg13g2_fill_1 FILLER_33_212 ();
 sg13g2_decap_4 FILLER_33_219 ();
 sg13g2_fill_1 FILLER_33_223 ();
 sg13g2_decap_8 FILLER_33_250 ();
 sg13g2_fill_2 FILLER_33_257 ();
 sg13g2_fill_2 FILLER_33_269 ();
 sg13g2_fill_1 FILLER_33_271 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_287 ();
 sg13g2_fill_1 FILLER_33_289 ();
 sg13g2_fill_1 FILLER_33_303 ();
 sg13g2_fill_2 FILLER_33_350 ();
 sg13g2_fill_2 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_fill_2 FILLER_34_63 ();
 sg13g2_fill_1 FILLER_34_65 ();
 sg13g2_fill_1 FILLER_34_104 ();
 sg13g2_fill_1 FILLER_34_159 ();
 sg13g2_fill_2 FILLER_34_178 ();
 sg13g2_fill_1 FILLER_34_180 ();
 sg13g2_decap_4 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_decap_4 FILLER_34_236 ();
 sg13g2_fill_2 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_fill_2 FILLER_35_70 ();
 sg13g2_fill_1 FILLER_35_76 ();
 sg13g2_fill_1 FILLER_35_81 ();
 sg13g2_fill_2 FILLER_35_105 ();
 sg13g2_fill_1 FILLER_35_156 ();
 sg13g2_fill_2 FILLER_35_174 ();
 sg13g2_fill_1 FILLER_35_176 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_fill_2 FILLER_35_318 ();
 sg13g2_fill_1 FILLER_35_320 ();
 sg13g2_fill_1 FILLER_35_397 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_4 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_67 ();
 sg13g2_fill_1 FILLER_36_93 ();
 sg13g2_fill_1 FILLER_36_132 ();
 sg13g2_fill_1 FILLER_36_150 ();
 sg13g2_fill_2 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_239 ();
 sg13g2_fill_2 FILLER_36_266 ();
 sg13g2_fill_1 FILLER_36_333 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_fill_2 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_183 ();
 sg13g2_decap_8 FILLER_37_206 ();
 sg13g2_decap_8 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_220 ();
 sg13g2_fill_1 FILLER_37_222 ();
 sg13g2_fill_2 FILLER_37_233 ();
 sg13g2_fill_2 FILLER_37_296 ();
 sg13g2_fill_2 FILLER_37_308 ();
 sg13g2_fill_2 FILLER_37_314 ();
 sg13g2_fill_2 FILLER_37_346 ();
 sg13g2_fill_1 FILLER_37_348 ();
 sg13g2_fill_2 FILLER_37_364 ();
 sg13g2_fill_1 FILLER_37_366 ();
 sg13g2_fill_2 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_4 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_53 ();
 sg13g2_fill_1 FILLER_38_120 ();
 sg13g2_fill_2 FILLER_38_170 ();
 sg13g2_fill_1 FILLER_38_184 ();
 sg13g2_decap_8 FILLER_38_195 ();
 sg13g2_decap_4 FILLER_38_202 ();
 sg13g2_fill_2 FILLER_38_206 ();
 sg13g2_decap_4 FILLER_38_214 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_fill_2 FILLER_38_245 ();
 sg13g2_fill_2 FILLER_38_262 ();
 sg13g2_fill_2 FILLER_38_282 ();
 sg13g2_decap_8 FILLER_38_305 ();
 sg13g2_fill_2 FILLER_38_346 ();
 sg13g2_fill_2 FILLER_38_358 ();
 sg13g2_fill_1 FILLER_38_360 ();
 sg13g2_fill_2 FILLER_38_370 ();
 sg13g2_fill_1 FILLER_38_372 ();
 sg13g2_fill_2 FILLER_38_392 ();
 sg13g2_fill_1 FILLER_38_394 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_4 FILLER_39_49 ();
 sg13g2_fill_2 FILLER_39_53 ();
 sg13g2_fill_2 FILLER_39_131 ();
 sg13g2_fill_1 FILLER_39_133 ();
 sg13g2_fill_1 FILLER_39_174 ();
 sg13g2_fill_1 FILLER_39_179 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_fill_2 FILLER_39_203 ();
 sg13g2_fill_1 FILLER_39_205 ();
 sg13g2_fill_1 FILLER_39_239 ();
 sg13g2_fill_2 FILLER_39_253 ();
 sg13g2_fill_1 FILLER_39_255 ();
 sg13g2_decap_8 FILLER_39_282 ();
 sg13g2_decap_4 FILLER_39_289 ();
 sg13g2_fill_1 FILLER_39_293 ();
 sg13g2_fill_2 FILLER_39_369 ();
 sg13g2_fill_1 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_fill_1 FILLER_40_82 ();
 sg13g2_fill_1 FILLER_40_128 ();
 sg13g2_fill_1 FILLER_40_133 ();
 sg13g2_decap_4 FILLER_40_160 ();
 sg13g2_decap_8 FILLER_40_190 ();
 sg13g2_fill_2 FILLER_40_217 ();
 sg13g2_fill_1 FILLER_40_219 ();
 sg13g2_fill_2 FILLER_40_344 ();
 sg13g2_fill_1 FILLER_40_346 ();
 sg13g2_fill_1 FILLER_40_394 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_fill_2 FILLER_41_56 ();
 sg13g2_fill_2 FILLER_41_84 ();
 sg13g2_fill_2 FILLER_41_138 ();
 sg13g2_fill_2 FILLER_41_160 ();
 sg13g2_decap_8 FILLER_41_188 ();
 sg13g2_decap_4 FILLER_41_195 ();
 sg13g2_decap_4 FILLER_41_215 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_4 FILLER_41_245 ();
 sg13g2_fill_1 FILLER_41_249 ();
 sg13g2_decap_4 FILLER_41_259 ();
 sg13g2_decap_4 FILLER_41_284 ();
 sg13g2_fill_2 FILLER_41_288 ();
 sg13g2_fill_2 FILLER_41_295 ();
 sg13g2_fill_1 FILLER_41_297 ();
 sg13g2_fill_1 FILLER_41_318 ();
 sg13g2_fill_2 FILLER_41_331 ();
 sg13g2_fill_2 FILLER_41_345 ();
 sg13g2_fill_1 FILLER_41_347 ();
 sg13g2_fill_2 FILLER_41_353 ();
 sg13g2_fill_2 FILLER_41_381 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_fill_2 FILLER_42_63 ();
 sg13g2_fill_1 FILLER_42_65 ();
 sg13g2_fill_2 FILLER_42_73 ();
 sg13g2_fill_1 FILLER_42_114 ();
 sg13g2_decap_4 FILLER_42_141 ();
 sg13g2_decap_4 FILLER_42_149 ();
 sg13g2_decap_4 FILLER_42_158 ();
 sg13g2_decap_4 FILLER_42_194 ();
 sg13g2_fill_1 FILLER_42_198 ();
 sg13g2_fill_1 FILLER_42_207 ();
 sg13g2_fill_2 FILLER_42_221 ();
 sg13g2_fill_1 FILLER_42_223 ();
 sg13g2_fill_1 FILLER_42_230 ();
 sg13g2_decap_8 FILLER_42_241 ();
 sg13g2_fill_1 FILLER_42_248 ();
 sg13g2_decap_8 FILLER_42_285 ();
 sg13g2_fill_2 FILLER_42_292 ();
 sg13g2_fill_1 FILLER_42_294 ();
 sg13g2_decap_8 FILLER_42_299 ();
 sg13g2_decap_4 FILLER_42_306 ();
 sg13g2_decap_8 FILLER_42_314 ();
 sg13g2_decap_8 FILLER_42_321 ();
 sg13g2_decap_4 FILLER_42_328 ();
 sg13g2_fill_1 FILLER_42_366 ();
 sg13g2_fill_1 FILLER_42_382 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_fill_2 FILLER_43_77 ();
 sg13g2_decap_4 FILLER_43_108 ();
 sg13g2_fill_1 FILLER_43_112 ();
 sg13g2_fill_2 FILLER_43_131 ();
 sg13g2_decap_8 FILLER_43_142 ();
 sg13g2_decap_8 FILLER_43_149 ();
 sg13g2_fill_2 FILLER_43_156 ();
 sg13g2_decap_8 FILLER_43_163 ();
 sg13g2_fill_2 FILLER_43_170 ();
 sg13g2_decap_8 FILLER_43_180 ();
 sg13g2_decap_8 FILLER_43_187 ();
 sg13g2_fill_1 FILLER_43_199 ();
 sg13g2_decap_4 FILLER_43_246 ();
 sg13g2_fill_1 FILLER_43_250 ();
 sg13g2_fill_1 FILLER_43_256 ();
 sg13g2_fill_1 FILLER_43_283 ();
 sg13g2_fill_1 FILLER_43_301 ();
 sg13g2_decap_8 FILLER_43_306 ();
 sg13g2_decap_8 FILLER_43_321 ();
 sg13g2_fill_2 FILLER_43_369 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_fill_2 FILLER_44_63 ();
 sg13g2_fill_1 FILLER_44_75 ();
 sg13g2_decap_8 FILLER_44_117 ();
 sg13g2_fill_2 FILLER_44_124 ();
 sg13g2_decap_8 FILLER_44_135 ();
 sg13g2_fill_1 FILLER_44_142 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_fill_2 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_176 ();
 sg13g2_decap_4 FILLER_44_183 ();
 sg13g2_fill_2 FILLER_44_249 ();
 sg13g2_fill_1 FILLER_44_256 ();
 sg13g2_fill_2 FILLER_44_313 ();
 sg13g2_fill_1 FILLER_44_315 ();
 sg13g2_fill_1 FILLER_44_335 ();
 sg13g2_fill_2 FILLER_44_345 ();
 sg13g2_fill_1 FILLER_44_347 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_4 FILLER_45_56 ();
 sg13g2_fill_2 FILLER_45_129 ();
 sg13g2_fill_1 FILLER_45_131 ();
 sg13g2_fill_1 FILLER_45_158 ();
 sg13g2_fill_1 FILLER_45_185 ();
 sg13g2_decap_8 FILLER_45_244 ();
 sg13g2_fill_2 FILLER_45_251 ();
 sg13g2_fill_1 FILLER_45_253 ();
 sg13g2_fill_2 FILLER_45_264 ();
 sg13g2_fill_1 FILLER_45_266 ();
 sg13g2_fill_1 FILLER_45_280 ();
 sg13g2_fill_2 FILLER_45_300 ();
 sg13g2_decap_4 FILLER_45_323 ();
 sg13g2_fill_2 FILLER_45_327 ();
 sg13g2_fill_2 FILLER_45_368 ();
 sg13g2_fill_2 FILLER_45_381 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_101 ();
 sg13g2_fill_1 FILLER_46_164 ();
 sg13g2_fill_2 FILLER_46_196 ();
 sg13g2_fill_1 FILLER_46_220 ();
 sg13g2_decap_4 FILLER_46_230 ();
 sg13g2_decap_8 FILLER_46_244 ();
 sg13g2_decap_4 FILLER_46_256 ();
 sg13g2_fill_1 FILLER_46_265 ();
 sg13g2_fill_1 FILLER_46_284 ();
 sg13g2_fill_2 FILLER_46_289 ();
 sg13g2_fill_1 FILLER_46_308 ();
 sg13g2_fill_2 FILLER_46_353 ();
 sg13g2_fill_2 FILLER_46_363 ();
 sg13g2_fill_1 FILLER_46_365 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_fill_2 FILLER_47_56 ();
 sg13g2_fill_1 FILLER_47_58 ();
 sg13g2_decap_4 FILLER_47_70 ();
 sg13g2_fill_2 FILLER_47_79 ();
 sg13g2_decap_8 FILLER_47_89 ();
 sg13g2_fill_2 FILLER_47_96 ();
 sg13g2_fill_1 FILLER_47_124 ();
 sg13g2_fill_2 FILLER_47_190 ();
 sg13g2_fill_1 FILLER_47_192 ();
 sg13g2_fill_1 FILLER_47_208 ();
 sg13g2_fill_1 FILLER_47_212 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_4 FILLER_47_224 ();
 sg13g2_fill_1 FILLER_47_228 ();
 sg13g2_fill_1 FILLER_47_238 ();
 sg13g2_fill_2 FILLER_47_249 ();
 sg13g2_decap_8 FILLER_47_290 ();
 sg13g2_decap_8 FILLER_47_297 ();
 sg13g2_decap_8 FILLER_47_304 ();
 sg13g2_fill_1 FILLER_47_311 ();
 sg13g2_fill_1 FILLER_47_330 ();
 sg13g2_fill_2 FILLER_47_365 ();
 sg13g2_fill_1 FILLER_47_367 ();
 sg13g2_fill_1 FILLER_47_373 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_4 FILLER_48_49 ();
 sg13g2_fill_2 FILLER_48_53 ();
 sg13g2_fill_1 FILLER_48_116 ();
 sg13g2_fill_1 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_fill_1 FILLER_48_217 ();
 sg13g2_fill_1 FILLER_48_300 ();
 sg13g2_decap_8 FILLER_48_306 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_fill_2 FILLER_48_336 ();
 sg13g2_fill_2 FILLER_48_351 ();
 sg13g2_fill_1 FILLER_48_353 ();
 sg13g2_fill_1 FILLER_48_380 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_fill_2 FILLER_49_63 ();
 sg13g2_fill_1 FILLER_49_65 ();
 sg13g2_fill_2 FILLER_49_78 ();
 sg13g2_fill_1 FILLER_49_80 ();
 sg13g2_fill_1 FILLER_49_107 ();
 sg13g2_fill_2 FILLER_49_190 ();
 sg13g2_decap_8 FILLER_49_209 ();
 sg13g2_decap_8 FILLER_49_221 ();
 sg13g2_fill_1 FILLER_49_228 ();
 sg13g2_decap_4 FILLER_49_244 ();
 sg13g2_fill_1 FILLER_49_283 ();
 sg13g2_decap_8 FILLER_49_325 ();
 sg13g2_fill_1 FILLER_49_332 ();
 sg13g2_decap_8 FILLER_49_339 ();
 sg13g2_fill_1 FILLER_49_346 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_fill_2 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_62 ();
 sg13g2_fill_1 FILLER_50_69 ();
 sg13g2_fill_2 FILLER_50_74 ();
 sg13g2_fill_2 FILLER_50_140 ();
 sg13g2_fill_1 FILLER_50_188 ();
 sg13g2_fill_2 FILLER_50_199 ();
 sg13g2_fill_1 FILLER_50_201 ();
 sg13g2_fill_2 FILLER_50_228 ();
 sg13g2_fill_2 FILLER_50_256 ();
 sg13g2_fill_1 FILLER_50_258 ();
 sg13g2_fill_1 FILLER_50_278 ();
 sg13g2_fill_2 FILLER_50_302 ();
 sg13g2_decap_8 FILLER_50_318 ();
 sg13g2_decap_4 FILLER_50_325 ();
 sg13g2_fill_2 FILLER_50_329 ();
 sg13g2_decap_8 FILLER_50_343 ();
 sg13g2_decap_4 FILLER_50_350 ();
 sg13g2_fill_2 FILLER_50_354 ();
 sg13g2_fill_2 FILLER_50_368 ();
 sg13g2_fill_2 FILLER_50_381 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_4 FILLER_51_35 ();
 sg13g2_decap_4 FILLER_51_44 ();
 sg13g2_fill_1 FILLER_51_79 ();
 sg13g2_fill_1 FILLER_51_165 ();
 sg13g2_fill_1 FILLER_51_175 ();
 sg13g2_fill_1 FILLER_51_190 ();
 sg13g2_fill_2 FILLER_51_215 ();
 sg13g2_decap_8 FILLER_51_234 ();
 sg13g2_decap_4 FILLER_51_245 ();
 sg13g2_decap_8 FILLER_51_267 ();
 sg13g2_decap_8 FILLER_51_282 ();
 sg13g2_decap_8 FILLER_51_289 ();
 sg13g2_fill_1 FILLER_51_331 ();
 sg13g2_fill_2 FILLER_51_367 ();
 sg13g2_fill_1 FILLER_51_369 ();
 sg13g2_fill_1 FILLER_51_390 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_4 FILLER_52_28 ();
 sg13g2_fill_2 FILLER_52_32 ();
 sg13g2_fill_1 FILLER_52_48 ();
 sg13g2_fill_2 FILLER_52_110 ();
 sg13g2_fill_1 FILLER_52_112 ();
 sg13g2_fill_2 FILLER_52_138 ();
 sg13g2_fill_2 FILLER_52_167 ();
 sg13g2_fill_1 FILLER_52_178 ();
 sg13g2_fill_1 FILLER_52_184 ();
 sg13g2_fill_1 FILLER_52_243 ();
 sg13g2_decap_8 FILLER_52_250 ();
 sg13g2_fill_2 FILLER_52_257 ();
 sg13g2_decap_8 FILLER_52_277 ();
 sg13g2_decap_8 FILLER_52_284 ();
 sg13g2_decap_8 FILLER_52_291 ();
 sg13g2_fill_2 FILLER_52_298 ();
 sg13g2_decap_4 FILLER_52_304 ();
 sg13g2_fill_2 FILLER_52_308 ();
 sg13g2_fill_1 FILLER_52_322 ();
 sg13g2_fill_2 FILLER_52_331 ();
 sg13g2_fill_1 FILLER_52_349 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_4 FILLER_53_28 ();
 sg13g2_fill_1 FILLER_53_32 ();
 sg13g2_fill_1 FILLER_53_91 ();
 sg13g2_fill_1 FILLER_53_127 ();
 sg13g2_fill_1 FILLER_53_241 ();
 sg13g2_fill_2 FILLER_53_280 ();
 sg13g2_decap_4 FILLER_53_337 ();
 sg13g2_fill_2 FILLER_53_349 ();
 sg13g2_fill_1 FILLER_53_351 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_4 FILLER_54_28 ();
 sg13g2_fill_1 FILLER_54_32 ();
 sg13g2_fill_2 FILLER_54_181 ();
 sg13g2_fill_2 FILLER_54_201 ();
 sg13g2_fill_1 FILLER_54_203 ();
 sg13g2_fill_1 FILLER_54_230 ();
 sg13g2_fill_2 FILLER_54_244 ();
 sg13g2_decap_4 FILLER_54_251 ();
 sg13g2_decap_4 FILLER_54_260 ();
 sg13g2_fill_2 FILLER_54_300 ();
 sg13g2_fill_1 FILLER_54_302 ();
 sg13g2_fill_1 FILLER_54_319 ();
 sg13g2_fill_2 FILLER_54_335 ();
 sg13g2_fill_1 FILLER_54_337 ();
 sg13g2_decap_8 FILLER_54_346 ();
 sg13g2_fill_2 FILLER_54_353 ();
 sg13g2_fill_1 FILLER_54_355 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_4 FILLER_55_21 ();
 sg13g2_fill_1 FILLER_55_25 ();
 sg13g2_fill_2 FILLER_55_52 ();
 sg13g2_fill_1 FILLER_55_63 ();
 sg13g2_fill_2 FILLER_55_119 ();
 sg13g2_fill_2 FILLER_55_145 ();
 sg13g2_fill_1 FILLER_55_147 ();
 sg13g2_fill_1 FILLER_55_201 ();
 sg13g2_decap_4 FILLER_55_211 ();
 sg13g2_fill_2 FILLER_55_222 ();
 sg13g2_fill_2 FILLER_55_328 ();
 sg13g2_fill_1 FILLER_55_330 ();
 sg13g2_decap_4 FILLER_55_357 ();
 sg13g2_fill_2 FILLER_55_361 ();
 sg13g2_decap_4 FILLER_55_367 ();
 sg13g2_fill_1 FILLER_55_371 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_4 FILLER_56_21 ();
 sg13g2_fill_2 FILLER_56_25 ();
 sg13g2_fill_2 FILLER_56_45 ();
 sg13g2_fill_1 FILLER_56_124 ();
 sg13g2_fill_1 FILLER_56_142 ();
 sg13g2_fill_2 FILLER_56_161 ();
 sg13g2_fill_1 FILLER_56_163 ();
 sg13g2_fill_1 FILLER_56_195 ();
 sg13g2_fill_2 FILLER_56_199 ();
 sg13g2_decap_8 FILLER_56_209 ();
 sg13g2_fill_2 FILLER_56_216 ();
 sg13g2_fill_1 FILLER_56_218 ();
 sg13g2_decap_4 FILLER_56_228 ();
 sg13g2_fill_1 FILLER_56_232 ();
 sg13g2_fill_2 FILLER_56_252 ();
 sg13g2_fill_2 FILLER_56_263 ();
 sg13g2_fill_1 FILLER_56_265 ();
 sg13g2_fill_1 FILLER_56_287 ();
 sg13g2_decap_4 FILLER_56_293 ();
 sg13g2_fill_1 FILLER_56_297 ();
 sg13g2_fill_1 FILLER_56_316 ();
 sg13g2_decap_4 FILLER_56_333 ();
 sg13g2_fill_2 FILLER_56_337 ();
 sg13g2_decap_8 FILLER_56_351 ();
 sg13g2_decap_8 FILLER_56_358 ();
 sg13g2_decap_8 FILLER_56_365 ();
 sg13g2_decap_8 FILLER_56_372 ();
 sg13g2_fill_2 FILLER_56_379 ();
 sg13g2_decap_8 FILLER_56_389 ();
 sg13g2_decap_8 FILLER_56_396 ();
 sg13g2_decap_4 FILLER_56_403 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_4 FILLER_57_21 ();
 sg13g2_fill_1 FILLER_57_63 ();
 sg13g2_fill_2 FILLER_57_78 ();
 sg13g2_fill_1 FILLER_57_80 ();
 sg13g2_fill_1 FILLER_57_86 ();
 sg13g2_fill_2 FILLER_57_128 ();
 sg13g2_fill_1 FILLER_57_160 ();
 sg13g2_fill_1 FILLER_57_176 ();
 sg13g2_fill_2 FILLER_57_191 ();
 sg13g2_fill_2 FILLER_57_214 ();
 sg13g2_fill_2 FILLER_57_236 ();
 sg13g2_fill_2 FILLER_57_317 ();
 sg13g2_fill_2 FILLER_57_340 ();
 sg13g2_decap_8 FILLER_57_360 ();
 sg13g2_decap_8 FILLER_57_367 ();
 sg13g2_decap_8 FILLER_57_374 ();
 sg13g2_decap_8 FILLER_57_381 ();
 sg13g2_decap_8 FILLER_57_388 ();
 sg13g2_decap_8 FILLER_57_395 ();
 sg13g2_decap_8 FILLER_57_402 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_fill_1 FILLER_58_28 ();
 sg13g2_fill_2 FILLER_58_42 ();
 sg13g2_fill_2 FILLER_58_62 ();
 sg13g2_fill_1 FILLER_58_64 ();
 sg13g2_fill_1 FILLER_58_75 ();
 sg13g2_decap_4 FILLER_58_81 ();
 sg13g2_fill_1 FILLER_58_98 ();
 sg13g2_fill_2 FILLER_58_136 ();
 sg13g2_decap_8 FILLER_58_371 ();
 sg13g2_decap_8 FILLER_58_378 ();
 sg13g2_decap_8 FILLER_58_385 ();
 sg13g2_decap_4 FILLER_58_392 ();
 sg13g2_decap_8 FILLER_58_399 ();
 sg13g2_fill_2 FILLER_58_406 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_4 FILLER_59_35 ();
 sg13g2_fill_1 FILLER_59_39 ();
 sg13g2_decap_8 FILLER_59_45 ();
 sg13g2_decap_4 FILLER_59_52 ();
 sg13g2_fill_2 FILLER_59_56 ();
 sg13g2_decap_4 FILLER_59_76 ();
 sg13g2_fill_1 FILLER_59_80 ();
 sg13g2_fill_1 FILLER_59_85 ();
 sg13g2_fill_2 FILLER_59_152 ();
 sg13g2_fill_2 FILLER_59_218 ();
 sg13g2_fill_1 FILLER_59_220 ();
 sg13g2_fill_1 FILLER_59_236 ();
 sg13g2_fill_2 FILLER_59_246 ();
 sg13g2_fill_1 FILLER_59_248 ();
 sg13g2_fill_2 FILLER_59_254 ();
 sg13g2_fill_1 FILLER_59_256 ();
 sg13g2_decap_4 FILLER_59_275 ();
 sg13g2_fill_2 FILLER_59_310 ();
 sg13g2_fill_2 FILLER_59_322 ();
 sg13g2_decap_4 FILLER_59_335 ();
 sg13g2_fill_1 FILLER_59_339 ();
 sg13g2_decap_4 FILLER_59_381 ();
 sg13g2_fill_1 FILLER_59_390 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_4 FILLER_60_28 ();
 sg13g2_fill_2 FILLER_60_58 ();
 sg13g2_fill_1 FILLER_60_69 ();
 sg13g2_fill_2 FILLER_60_116 ();
 sg13g2_decap_8 FILLER_60_235 ();
 sg13g2_fill_2 FILLER_60_242 ();
 sg13g2_fill_2 FILLER_60_270 ();
 sg13g2_fill_2 FILLER_60_316 ();
 sg13g2_fill_2 FILLER_60_330 ();
 sg13g2_fill_1 FILLER_60_332 ();
 sg13g2_fill_2 FILLER_60_343 ();
 sg13g2_fill_2 FILLER_60_350 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_4 FILLER_61_35 ();
 sg13g2_fill_2 FILLER_61_39 ();
 sg13g2_decap_4 FILLER_61_55 ();
 sg13g2_decap_4 FILLER_61_74 ();
 sg13g2_fill_2 FILLER_61_83 ();
 sg13g2_fill_1 FILLER_61_85 ();
 sg13g2_fill_2 FILLER_61_117 ();
 sg13g2_fill_1 FILLER_61_119 ();
 sg13g2_fill_1 FILLER_61_148 ();
 sg13g2_fill_2 FILLER_61_153 ();
 sg13g2_fill_2 FILLER_61_173 ();
 sg13g2_fill_1 FILLER_61_175 ();
 sg13g2_fill_1 FILLER_61_193 ();
 sg13g2_decap_4 FILLER_61_207 ();
 sg13g2_fill_2 FILLER_61_211 ();
 sg13g2_fill_1 FILLER_61_222 ();
 sg13g2_decap_8 FILLER_61_227 ();
 sg13g2_fill_1 FILLER_61_234 ();
 sg13g2_decap_8 FILLER_61_243 ();
 sg13g2_fill_1 FILLER_61_255 ();
 sg13g2_fill_2 FILLER_61_348 ();
 sg13g2_fill_1 FILLER_61_386 ();
 sg13g2_fill_1 FILLER_61_394 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_4 FILLER_62_42 ();
 sg13g2_fill_1 FILLER_62_46 ();
 sg13g2_fill_2 FILLER_62_57 ();
 sg13g2_fill_1 FILLER_62_78 ();
 sg13g2_fill_1 FILLER_62_92 ();
 sg13g2_fill_1 FILLER_62_144 ();
 sg13g2_decap_4 FILLER_62_210 ();
 sg13g2_decap_4 FILLER_62_217 ();
 sg13g2_fill_2 FILLER_62_225 ();
 sg13g2_fill_1 FILLER_62_227 ();
 sg13g2_fill_1 FILLER_62_262 ();
 sg13g2_decap_4 FILLER_62_293 ();
 sg13g2_fill_2 FILLER_62_304 ();
 sg13g2_decap_8 FILLER_62_310 ();
 sg13g2_fill_1 FILLER_62_317 ();
 sg13g2_decap_4 FILLER_62_331 ();
 sg13g2_fill_2 FILLER_62_335 ();
 sg13g2_fill_2 FILLER_62_342 ();
 sg13g2_fill_1 FILLER_62_344 ();
 sg13g2_fill_2 FILLER_62_375 ();
 sg13g2_fill_1 FILLER_62_377 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_fill_1 FILLER_63_63 ();
 sg13g2_fill_2 FILLER_63_98 ();
 sg13g2_fill_1 FILLER_63_100 ();
 sg13g2_fill_2 FILLER_63_198 ();
 sg13g2_fill_1 FILLER_63_200 ();
 sg13g2_decap_4 FILLER_63_217 ();
 sg13g2_fill_1 FILLER_63_221 ();
 sg13g2_fill_1 FILLER_63_254 ();
 sg13g2_decap_4 FILLER_63_301 ();
 sg13g2_fill_2 FILLER_63_305 ();
 sg13g2_fill_2 FILLER_63_313 ();
 sg13g2_decap_8 FILLER_63_323 ();
 sg13g2_decap_8 FILLER_63_330 ();
 sg13g2_decap_4 FILLER_63_337 ();
 sg13g2_decap_4 FILLER_63_349 ();
 sg13g2_fill_2 FILLER_63_353 ();
 sg13g2_fill_2 FILLER_63_361 ();
 sg13g2_decap_4 FILLER_63_380 ();
 sg13g2_fill_1 FILLER_63_392 ();
 sg13g2_fill_2 FILLER_63_406 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_4 FILLER_64_21 ();
 sg13g2_fill_1 FILLER_64_25 ();
 sg13g2_fill_2 FILLER_64_52 ();
 sg13g2_fill_2 FILLER_64_64 ();
 sg13g2_fill_2 FILLER_64_80 ();
 sg13g2_fill_1 FILLER_64_82 ();
 sg13g2_fill_1 FILLER_64_111 ();
 sg13g2_fill_2 FILLER_64_124 ();
 sg13g2_fill_1 FILLER_64_141 ();
 sg13g2_fill_1 FILLER_64_148 ();
 sg13g2_fill_2 FILLER_64_158 ();
 sg13g2_decap_4 FILLER_64_183 ();
 sg13g2_fill_1 FILLER_64_187 ();
 sg13g2_fill_2 FILLER_64_209 ();
 sg13g2_fill_1 FILLER_64_211 ();
 sg13g2_decap_8 FILLER_64_220 ();
 sg13g2_fill_2 FILLER_64_249 ();
 sg13g2_fill_1 FILLER_64_251 ();
 sg13g2_fill_2 FILLER_64_271 ();
 sg13g2_fill_1 FILLER_64_273 ();
 sg13g2_fill_2 FILLER_64_299 ();
 sg13g2_fill_1 FILLER_64_346 ();
 sg13g2_fill_1 FILLER_64_351 ();
 sg13g2_decap_8 FILLER_64_373 ();
 sg13g2_fill_2 FILLER_64_380 ();
 sg13g2_decap_4 FILLER_64_392 ();
 sg13g2_decap_4 FILLER_64_405 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_fill_1 FILLER_65_32 ();
 sg13g2_fill_1 FILLER_65_63 ();
 sg13g2_fill_1 FILLER_65_87 ();
 sg13g2_fill_2 FILLER_65_115 ();
 sg13g2_fill_1 FILLER_65_117 ();
 sg13g2_decap_8 FILLER_65_122 ();
 sg13g2_fill_2 FILLER_65_142 ();
 sg13g2_fill_2 FILLER_65_163 ();
 sg13g2_fill_2 FILLER_65_173 ();
 sg13g2_fill_1 FILLER_65_175 ();
 sg13g2_decap_8 FILLER_65_194 ();
 sg13g2_fill_1 FILLER_65_201 ();
 sg13g2_decap_8 FILLER_65_223 ();
 sg13g2_decap_8 FILLER_65_247 ();
 sg13g2_decap_8 FILLER_65_254 ();
 sg13g2_fill_1 FILLER_65_261 ();
 sg13g2_fill_1 FILLER_65_277 ();
 sg13g2_fill_2 FILLER_65_320 ();
 sg13g2_fill_2 FILLER_65_343 ();
 sg13g2_fill_1 FILLER_65_363 ();
 sg13g2_fill_1 FILLER_65_388 ();
 sg13g2_decap_8 FILLER_65_401 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_fill_2 FILLER_66_14 ();
 sg13g2_fill_1 FILLER_66_16 ();
 sg13g2_decap_4 FILLER_66_47 ();
 sg13g2_fill_1 FILLER_66_51 ();
 sg13g2_fill_1 FILLER_66_63 ();
 sg13g2_fill_2 FILLER_66_68 ();
 sg13g2_fill_2 FILLER_66_105 ();
 sg13g2_fill_2 FILLER_66_139 ();
 sg13g2_decap_8 FILLER_66_194 ();
 sg13g2_decap_8 FILLER_66_206 ();
 sg13g2_decap_8 FILLER_66_225 ();
 sg13g2_decap_8 FILLER_66_232 ();
 sg13g2_decap_8 FILLER_66_239 ();
 sg13g2_decap_4 FILLER_66_246 ();
 sg13g2_fill_2 FILLER_66_250 ();
 sg13g2_fill_1 FILLER_66_256 ();
 sg13g2_fill_2 FILLER_66_289 ();
 sg13g2_fill_1 FILLER_66_291 ();
 sg13g2_decap_8 FILLER_66_315 ();
 sg13g2_fill_2 FILLER_66_322 ();
 sg13g2_fill_1 FILLER_66_324 ();
 sg13g2_fill_2 FILLER_66_338 ();
 sg13g2_fill_1 FILLER_66_340 ();
 sg13g2_fill_2 FILLER_66_345 ();
 sg13g2_fill_1 FILLER_66_347 ();
 sg13g2_fill_2 FILLER_66_376 ();
 sg13g2_fill_1 FILLER_66_378 ();
 sg13g2_decap_8 FILLER_66_394 ();
 sg13g2_decap_8 FILLER_66_401 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_fill_2 FILLER_67_14 ();
 sg13g2_fill_1 FILLER_67_34 ();
 sg13g2_fill_2 FILLER_67_55 ();
 sg13g2_fill_1 FILLER_67_57 ();
 sg13g2_decap_4 FILLER_67_77 ();
 sg13g2_fill_1 FILLER_67_81 ();
 sg13g2_fill_2 FILLER_67_175 ();
 sg13g2_fill_1 FILLER_67_203 ();
 sg13g2_fill_2 FILLER_67_209 ();
 sg13g2_fill_1 FILLER_67_211 ();
 sg13g2_fill_1 FILLER_67_230 ();
 sg13g2_fill_1 FILLER_67_265 ();
 sg13g2_fill_1 FILLER_67_275 ();
 sg13g2_fill_2 FILLER_67_297 ();
 sg13g2_fill_1 FILLER_67_299 ();
 sg13g2_decap_4 FILLER_67_360 ();
 sg13g2_fill_2 FILLER_67_364 ();
 sg13g2_decap_8 FILLER_67_377 ();
 sg13g2_decap_4 FILLER_67_387 ();
 sg13g2_fill_1 FILLER_67_391 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_fill_2 FILLER_68_40 ();
 sg13g2_fill_2 FILLER_68_51 ();
 sg13g2_fill_1 FILLER_68_53 ();
 sg13g2_decap_4 FILLER_68_72 ();
 sg13g2_fill_1 FILLER_68_76 ();
 sg13g2_fill_2 FILLER_68_91 ();
 sg13g2_fill_1 FILLER_68_106 ();
 sg13g2_fill_1 FILLER_68_157 ();
 sg13g2_fill_2 FILLER_68_176 ();
 sg13g2_fill_1 FILLER_68_222 ();
 sg13g2_fill_2 FILLER_68_239 ();
 sg13g2_fill_1 FILLER_68_241 ();
 sg13g2_decap_4 FILLER_68_297 ();
 sg13g2_decap_4 FILLER_68_320 ();
 sg13g2_decap_8 FILLER_68_328 ();
 sg13g2_decap_8 FILLER_68_335 ();
 sg13g2_decap_8 FILLER_68_342 ();
 sg13g2_decap_8 FILLER_68_349 ();
 sg13g2_decap_8 FILLER_68_356 ();
 sg13g2_decap_8 FILLER_68_363 ();
 sg13g2_decap_4 FILLER_68_370 ();
 sg13g2_decap_4 FILLER_68_377 ();
 sg13g2_fill_2 FILLER_68_381 ();
 sg13g2_fill_2 FILLER_68_393 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_4 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_54 ();
 sg13g2_fill_2 FILLER_69_74 ();
 sg13g2_fill_1 FILLER_69_81 ();
 sg13g2_fill_2 FILLER_69_101 ();
 sg13g2_fill_1 FILLER_69_103 ();
 sg13g2_fill_2 FILLER_69_118 ();
 sg13g2_fill_1 FILLER_69_154 ();
 sg13g2_fill_1 FILLER_69_198 ();
 sg13g2_fill_2 FILLER_69_209 ();
 sg13g2_fill_1 FILLER_69_211 ();
 sg13g2_fill_2 FILLER_69_218 ();
 sg13g2_decap_4 FILLER_69_238 ();
 sg13g2_fill_1 FILLER_69_242 ();
 sg13g2_fill_2 FILLER_69_252 ();
 sg13g2_fill_1 FILLER_69_254 ();
 sg13g2_fill_1 FILLER_69_260 ();
 sg13g2_decap_4 FILLER_69_296 ();
 sg13g2_fill_1 FILLER_69_300 ();
 sg13g2_fill_2 FILLER_69_306 ();
 sg13g2_fill_1 FILLER_69_308 ();
 sg13g2_fill_2 FILLER_69_319 ();
 sg13g2_decap_8 FILLER_69_326 ();
 sg13g2_fill_1 FILLER_69_333 ();
 sg13g2_fill_1 FILLER_69_351 ();
 sg13g2_decap_4 FILLER_69_356 ();
 sg13g2_fill_1 FILLER_69_360 ();
 sg13g2_fill_2 FILLER_69_373 ();
 sg13g2_fill_1 FILLER_69_381 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_fill_2 FILLER_70_45 ();
 sg13g2_fill_2 FILLER_70_68 ();
 sg13g2_fill_2 FILLER_70_84 ();
 sg13g2_fill_1 FILLER_70_86 ();
 sg13g2_fill_2 FILLER_70_107 ();
 sg13g2_fill_2 FILLER_70_125 ();
 sg13g2_fill_2 FILLER_70_150 ();
 sg13g2_fill_2 FILLER_70_232 ();
 sg13g2_decap_4 FILLER_70_246 ();
 sg13g2_fill_1 FILLER_70_250 ();
 sg13g2_fill_1 FILLER_70_270 ();
 sg13g2_fill_2 FILLER_70_292 ();
 sg13g2_fill_1 FILLER_70_294 ();
 sg13g2_fill_2 FILLER_70_303 ();
 sg13g2_fill_2 FILLER_70_343 ();
 sg13g2_fill_1 FILLER_70_345 ();
 sg13g2_fill_1 FILLER_70_387 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_fill_2 FILLER_71_14 ();
 sg13g2_fill_2 FILLER_71_74 ();
 sg13g2_decap_4 FILLER_71_100 ();
 sg13g2_fill_1 FILLER_71_119 ();
 sg13g2_fill_2 FILLER_71_188 ();
 sg13g2_fill_2 FILLER_71_195 ();
 sg13g2_fill_1 FILLER_71_197 ();
 sg13g2_decap_4 FILLER_71_202 ();
 sg13g2_fill_1 FILLER_71_206 ();
 sg13g2_fill_2 FILLER_71_258 ();
 sg13g2_fill_1 FILLER_71_341 ();
 sg13g2_fill_1 FILLER_71_356 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_fill_1 FILLER_72_21 ();
 sg13g2_fill_1 FILLER_72_40 ();
 sg13g2_fill_2 FILLER_72_59 ();
 sg13g2_decap_8 FILLER_72_89 ();
 sg13g2_decap_4 FILLER_72_96 ();
 sg13g2_fill_1 FILLER_72_100 ();
 sg13g2_fill_2 FILLER_72_161 ();
 sg13g2_fill_1 FILLER_72_163 ();
 sg13g2_fill_2 FILLER_72_177 ();
 sg13g2_decap_4 FILLER_72_189 ();
 sg13g2_fill_2 FILLER_72_202 ();
 sg13g2_fill_1 FILLER_72_204 ();
 sg13g2_fill_2 FILLER_72_210 ();
 sg13g2_fill_1 FILLER_72_212 ();
 sg13g2_fill_2 FILLER_72_270 ();
 sg13g2_fill_1 FILLER_72_272 ();
 sg13g2_fill_1 FILLER_72_356 ();
 sg13g2_decap_8 FILLER_72_376 ();
 sg13g2_fill_1 FILLER_72_383 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_fill_2 FILLER_73_21 ();
 sg13g2_fill_1 FILLER_73_23 ();
 sg13g2_fill_1 FILLER_73_67 ();
 sg13g2_decap_4 FILLER_73_95 ();
 sg13g2_decap_4 FILLER_73_116 ();
 sg13g2_fill_1 FILLER_73_120 ();
 sg13g2_fill_1 FILLER_73_129 ();
 sg13g2_fill_2 FILLER_73_188 ();
 sg13g2_fill_2 FILLER_73_225 ();
 sg13g2_fill_1 FILLER_73_227 ();
 sg13g2_fill_1 FILLER_73_236 ();
 sg13g2_decap_4 FILLER_73_350 ();
 sg13g2_fill_2 FILLER_73_387 ();
 sg13g2_fill_1 FILLER_73_389 ();
 sg13g2_fill_1 FILLER_73_394 ();
 sg13g2_decap_8 FILLER_73_398 ();
 sg13g2_decap_4 FILLER_73_405 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_fill_2 FILLER_74_28 ();
 sg13g2_fill_1 FILLER_74_79 ();
 sg13g2_fill_2 FILLER_74_90 ();
 sg13g2_decap_8 FILLER_74_102 ();
 sg13g2_fill_1 FILLER_74_109 ();
 sg13g2_fill_2 FILLER_74_164 ();
 sg13g2_fill_2 FILLER_74_192 ();
 sg13g2_fill_1 FILLER_74_233 ();
 sg13g2_decap_8 FILLER_74_330 ();
 sg13g2_decap_4 FILLER_74_337 ();
 sg13g2_fill_1 FILLER_74_341 ();
 sg13g2_fill_1 FILLER_74_358 ();
 sg13g2_fill_1 FILLER_74_365 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_4 FILLER_75_35 ();
 sg13g2_fill_1 FILLER_75_39 ();
 sg13g2_decap_4 FILLER_75_44 ();
 sg13g2_decap_4 FILLER_75_52 ();
 sg13g2_fill_1 FILLER_75_56 ();
 sg13g2_fill_2 FILLER_75_83 ();
 sg13g2_fill_1 FILLER_75_85 ();
 sg13g2_fill_1 FILLER_75_121 ();
 sg13g2_decap_4 FILLER_75_128 ();
 sg13g2_fill_2 FILLER_75_138 ();
 sg13g2_fill_1 FILLER_75_140 ();
 sg13g2_fill_1 FILLER_75_151 ();
 sg13g2_fill_2 FILLER_75_178 ();
 sg13g2_fill_1 FILLER_75_180 ();
 sg13g2_fill_1 FILLER_75_200 ();
 sg13g2_fill_2 FILLER_75_214 ();
 sg13g2_fill_2 FILLER_75_226 ();
 sg13g2_fill_2 FILLER_75_237 ();
 sg13g2_fill_1 FILLER_75_239 ();
 sg13g2_fill_2 FILLER_75_245 ();
 sg13g2_fill_1 FILLER_75_252 ();
 sg13g2_fill_2 FILLER_75_270 ();
 sg13g2_fill_1 FILLER_75_272 ();
 sg13g2_fill_2 FILLER_75_300 ();
 sg13g2_fill_2 FILLER_75_315 ();
 sg13g2_decap_4 FILLER_75_327 ();
 sg13g2_fill_2 FILLER_75_331 ();
 sg13g2_decap_4 FILLER_75_342 ();
 sg13g2_fill_1 FILLER_75_346 ();
 sg13g2_fill_1 FILLER_75_351 ();
 sg13g2_decap_4 FILLER_75_404 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_4 FILLER_76_63 ();
 sg13g2_fill_1 FILLER_76_67 ();
 sg13g2_decap_8 FILLER_76_74 ();
 sg13g2_fill_1 FILLER_76_81 ();
 sg13g2_fill_1 FILLER_76_91 ();
 sg13g2_fill_1 FILLER_76_171 ();
 sg13g2_fill_1 FILLER_76_206 ();
 sg13g2_fill_1 FILLER_76_212 ();
 sg13g2_fill_2 FILLER_76_283 ();
 sg13g2_fill_1 FILLER_76_285 ();
 sg13g2_fill_2 FILLER_76_300 ();
 sg13g2_fill_1 FILLER_76_311 ();
 sg13g2_fill_2 FILLER_76_361 ();
 sg13g2_fill_1 FILLER_76_377 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_fill_2 FILLER_76_406 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_4 FILLER_77_42 ();
 sg13g2_fill_1 FILLER_77_83 ();
 sg13g2_decap_4 FILLER_77_109 ();
 sg13g2_decap_4 FILLER_77_122 ();
 sg13g2_fill_1 FILLER_77_177 ();
 sg13g2_fill_2 FILLER_77_182 ();
 sg13g2_fill_1 FILLER_77_184 ();
 sg13g2_fill_1 FILLER_77_189 ();
 sg13g2_fill_2 FILLER_77_242 ();
 sg13g2_fill_2 FILLER_77_285 ();
 sg13g2_fill_2 FILLER_77_313 ();
 sg13g2_fill_1 FILLER_77_320 ();
 sg13g2_fill_1 FILLER_77_390 ();
 sg13g2_decap_4 FILLER_77_404 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_fill_1 FILLER_78_49 ();
 sg13g2_fill_2 FILLER_78_126 ();
 sg13g2_fill_1 FILLER_78_209 ();
 sg13g2_fill_2 FILLER_78_272 ();
 sg13g2_fill_1 FILLER_78_326 ();
 sg13g2_fill_2 FILLER_78_380 ();
 sg13g2_fill_1 FILLER_78_382 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_fill_1 FILLER_79_56 ();
 sg13g2_fill_1 FILLER_79_86 ();
 sg13g2_fill_1 FILLER_79_91 ();
 sg13g2_fill_2 FILLER_79_239 ();
 sg13g2_fill_2 FILLER_79_250 ();
 sg13g2_fill_2 FILLER_79_345 ();
 sg13g2_fill_1 FILLER_79_347 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_1 FILLER_80_70 ();
 sg13g2_decap_8 FILLER_80_80 ();
 sg13g2_decap_8 FILLER_80_87 ();
 sg13g2_decap_4 FILLER_80_94 ();
 sg13g2_fill_2 FILLER_80_98 ();
 sg13g2_fill_1 FILLER_80_109 ();
 sg13g2_fill_1 FILLER_80_119 ();
 sg13g2_decap_8 FILLER_80_124 ();
 sg13g2_fill_1 FILLER_80_131 ();
 sg13g2_decap_4 FILLER_80_145 ();
 sg13g2_decap_8 FILLER_80_175 ();
 sg13g2_decap_4 FILLER_80_182 ();
 sg13g2_fill_1 FILLER_80_186 ();
 sg13g2_decap_8 FILLER_80_191 ();
 sg13g2_decap_8 FILLER_80_198 ();
 sg13g2_fill_1 FILLER_80_205 ();
 sg13g2_decap_8 FILLER_80_214 ();
 sg13g2_decap_8 FILLER_80_221 ();
 sg13g2_decap_8 FILLER_80_228 ();
 sg13g2_decap_8 FILLER_80_235 ();
 sg13g2_decap_8 FILLER_80_242 ();
 sg13g2_fill_1 FILLER_80_249 ();
 sg13g2_fill_1 FILLER_80_287 ();
 sg13g2_fill_2 FILLER_80_293 ();
 sg13g2_fill_1 FILLER_80_295 ();
 sg13g2_fill_2 FILLER_80_309 ();
 sg13g2_fill_2 FILLER_80_324 ();
 sg13g2_fill_2 FILLER_80_351 ();
 sg13g2_fill_1 FILLER_80_353 ();
 sg13g2_fill_1 FILLER_80_370 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_out[7] = net11;
endmodule

module tt_um_urish_sic1 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \A[0] ;
 wire \A[1] ;
 wire \A[2] ;
 wire \A[3] ;
 wire \A[4] ;
 wire \A[5] ;
 wire \A[6] ;
 wire \A[7] ;
 wire \B[0] ;
 wire \B[1] ;
 wire \B[2] ;
 wire \B[3] ;
 wire \B[4] ;
 wire \B[5] ;
 wire \B[6] ;
 wire \B[7] ;
 wire \C[0] ;
 wire \C[1] ;
 wire \C[2] ;
 wire \C[3] ;
 wire \C[4] ;
 wire \C[5] ;
 wire \C[6] ;
 wire \C[7] ;
 wire \PC[0] ;
 wire \PC[1] ;
 wire \PC[2] ;
 wire \PC[3] ;
 wire \PC[4] ;
 wire \PC[5] ;
 wire \PC[6] ;
 wire \PC[7] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire halted;
 wire \mem.addr[0] ;
 wire \mem.addr[1] ;
 wire \mem.addr[2] ;
 wire \mem.addr[3] ;
 wire \mem.addr[4] ;
 wire \mem.addr[5] ;
 wire \mem.addr[6] ;
 wire \mem.addr[7] ;
 wire \mem.data_in[0] ;
 wire \mem.data_in[1] ;
 wire \mem.data_in[2] ;
 wire \mem.data_in[3] ;
 wire \mem.data_in[4] ;
 wire \mem.data_in[5] ;
 wire \mem.data_in[6] ;
 wire \mem.data_in[7] ;
 wire \mem.mem[0][0] ;
 wire \mem.mem[0][1] ;
 wire \mem.mem[0][2] ;
 wire \mem.mem[0][3] ;
 wire \mem.mem[0][4] ;
 wire \mem.mem[0][5] ;
 wire \mem.mem[0][6] ;
 wire \mem.mem[0][7] ;
 wire \mem.mem[100][0] ;
 wire \mem.mem[100][1] ;
 wire \mem.mem[100][2] ;
 wire \mem.mem[100][3] ;
 wire \mem.mem[100][4] ;
 wire \mem.mem[100][5] ;
 wire \mem.mem[100][6] ;
 wire \mem.mem[100][7] ;
 wire \mem.mem[101][0] ;
 wire \mem.mem[101][1] ;
 wire \mem.mem[101][2] ;
 wire \mem.mem[101][3] ;
 wire \mem.mem[101][4] ;
 wire \mem.mem[101][5] ;
 wire \mem.mem[101][6] ;
 wire \mem.mem[101][7] ;
 wire \mem.mem[102][0] ;
 wire \mem.mem[102][1] ;
 wire \mem.mem[102][2] ;
 wire \mem.mem[102][3] ;
 wire \mem.mem[102][4] ;
 wire \mem.mem[102][5] ;
 wire \mem.mem[102][6] ;
 wire \mem.mem[102][7] ;
 wire \mem.mem[103][0] ;
 wire \mem.mem[103][1] ;
 wire \mem.mem[103][2] ;
 wire \mem.mem[103][3] ;
 wire \mem.mem[103][4] ;
 wire \mem.mem[103][5] ;
 wire \mem.mem[103][6] ;
 wire \mem.mem[103][7] ;
 wire \mem.mem[104][0] ;
 wire \mem.mem[104][1] ;
 wire \mem.mem[104][2] ;
 wire \mem.mem[104][3] ;
 wire \mem.mem[104][4] ;
 wire \mem.mem[104][5] ;
 wire \mem.mem[104][6] ;
 wire \mem.mem[104][7] ;
 wire \mem.mem[105][0] ;
 wire \mem.mem[105][1] ;
 wire \mem.mem[105][2] ;
 wire \mem.mem[105][3] ;
 wire \mem.mem[105][4] ;
 wire \mem.mem[105][5] ;
 wire \mem.mem[105][6] ;
 wire \mem.mem[105][7] ;
 wire \mem.mem[106][0] ;
 wire \mem.mem[106][1] ;
 wire \mem.mem[106][2] ;
 wire \mem.mem[106][3] ;
 wire \mem.mem[106][4] ;
 wire \mem.mem[106][5] ;
 wire \mem.mem[106][6] ;
 wire \mem.mem[106][7] ;
 wire \mem.mem[107][0] ;
 wire \mem.mem[107][1] ;
 wire \mem.mem[107][2] ;
 wire \mem.mem[107][3] ;
 wire \mem.mem[107][4] ;
 wire \mem.mem[107][5] ;
 wire \mem.mem[107][6] ;
 wire \mem.mem[107][7] ;
 wire \mem.mem[108][0] ;
 wire \mem.mem[108][1] ;
 wire \mem.mem[108][2] ;
 wire \mem.mem[108][3] ;
 wire \mem.mem[108][4] ;
 wire \mem.mem[108][5] ;
 wire \mem.mem[108][6] ;
 wire \mem.mem[108][7] ;
 wire \mem.mem[109][0] ;
 wire \mem.mem[109][1] ;
 wire \mem.mem[109][2] ;
 wire \mem.mem[109][3] ;
 wire \mem.mem[109][4] ;
 wire \mem.mem[109][5] ;
 wire \mem.mem[109][6] ;
 wire \mem.mem[109][7] ;
 wire \mem.mem[10][0] ;
 wire \mem.mem[10][1] ;
 wire \mem.mem[10][2] ;
 wire \mem.mem[10][3] ;
 wire \mem.mem[10][4] ;
 wire \mem.mem[10][5] ;
 wire \mem.mem[10][6] ;
 wire \mem.mem[10][7] ;
 wire \mem.mem[110][0] ;
 wire \mem.mem[110][1] ;
 wire \mem.mem[110][2] ;
 wire \mem.mem[110][3] ;
 wire \mem.mem[110][4] ;
 wire \mem.mem[110][5] ;
 wire \mem.mem[110][6] ;
 wire \mem.mem[110][7] ;
 wire \mem.mem[111][0] ;
 wire \mem.mem[111][1] ;
 wire \mem.mem[111][2] ;
 wire \mem.mem[111][3] ;
 wire \mem.mem[111][4] ;
 wire \mem.mem[111][5] ;
 wire \mem.mem[111][6] ;
 wire \mem.mem[111][7] ;
 wire \mem.mem[112][0] ;
 wire \mem.mem[112][1] ;
 wire \mem.mem[112][2] ;
 wire \mem.mem[112][3] ;
 wire \mem.mem[112][4] ;
 wire \mem.mem[112][5] ;
 wire \mem.mem[112][6] ;
 wire \mem.mem[112][7] ;
 wire \mem.mem[113][0] ;
 wire \mem.mem[113][1] ;
 wire \mem.mem[113][2] ;
 wire \mem.mem[113][3] ;
 wire \mem.mem[113][4] ;
 wire \mem.mem[113][5] ;
 wire \mem.mem[113][6] ;
 wire \mem.mem[113][7] ;
 wire \mem.mem[114][0] ;
 wire \mem.mem[114][1] ;
 wire \mem.mem[114][2] ;
 wire \mem.mem[114][3] ;
 wire \mem.mem[114][4] ;
 wire \mem.mem[114][5] ;
 wire \mem.mem[114][6] ;
 wire \mem.mem[114][7] ;
 wire \mem.mem[115][0] ;
 wire \mem.mem[115][1] ;
 wire \mem.mem[115][2] ;
 wire \mem.mem[115][3] ;
 wire \mem.mem[115][4] ;
 wire \mem.mem[115][5] ;
 wire \mem.mem[115][6] ;
 wire \mem.mem[115][7] ;
 wire \mem.mem[116][0] ;
 wire \mem.mem[116][1] ;
 wire \mem.mem[116][2] ;
 wire \mem.mem[116][3] ;
 wire \mem.mem[116][4] ;
 wire \mem.mem[116][5] ;
 wire \mem.mem[116][6] ;
 wire \mem.mem[116][7] ;
 wire \mem.mem[117][0] ;
 wire \mem.mem[117][1] ;
 wire \mem.mem[117][2] ;
 wire \mem.mem[117][3] ;
 wire \mem.mem[117][4] ;
 wire \mem.mem[117][5] ;
 wire \mem.mem[117][6] ;
 wire \mem.mem[117][7] ;
 wire \mem.mem[118][0] ;
 wire \mem.mem[118][1] ;
 wire \mem.mem[118][2] ;
 wire \mem.mem[118][3] ;
 wire \mem.mem[118][4] ;
 wire \mem.mem[118][5] ;
 wire \mem.mem[118][6] ;
 wire \mem.mem[118][7] ;
 wire \mem.mem[119][0] ;
 wire \mem.mem[119][1] ;
 wire \mem.mem[119][2] ;
 wire \mem.mem[119][3] ;
 wire \mem.mem[119][4] ;
 wire \mem.mem[119][5] ;
 wire \mem.mem[119][6] ;
 wire \mem.mem[119][7] ;
 wire \mem.mem[11][0] ;
 wire \mem.mem[11][1] ;
 wire \mem.mem[11][2] ;
 wire \mem.mem[11][3] ;
 wire \mem.mem[11][4] ;
 wire \mem.mem[11][5] ;
 wire \mem.mem[11][6] ;
 wire \mem.mem[11][7] ;
 wire \mem.mem[120][0] ;
 wire \mem.mem[120][1] ;
 wire \mem.mem[120][2] ;
 wire \mem.mem[120][3] ;
 wire \mem.mem[120][4] ;
 wire \mem.mem[120][5] ;
 wire \mem.mem[120][6] ;
 wire \mem.mem[120][7] ;
 wire \mem.mem[121][0] ;
 wire \mem.mem[121][1] ;
 wire \mem.mem[121][2] ;
 wire \mem.mem[121][3] ;
 wire \mem.mem[121][4] ;
 wire \mem.mem[121][5] ;
 wire \mem.mem[121][6] ;
 wire \mem.mem[121][7] ;
 wire \mem.mem[122][0] ;
 wire \mem.mem[122][1] ;
 wire \mem.mem[122][2] ;
 wire \mem.mem[122][3] ;
 wire \mem.mem[122][4] ;
 wire \mem.mem[122][5] ;
 wire \mem.mem[122][6] ;
 wire \mem.mem[122][7] ;
 wire \mem.mem[123][0] ;
 wire \mem.mem[123][1] ;
 wire \mem.mem[123][2] ;
 wire \mem.mem[123][3] ;
 wire \mem.mem[123][4] ;
 wire \mem.mem[123][5] ;
 wire \mem.mem[123][6] ;
 wire \mem.mem[123][7] ;
 wire \mem.mem[124][0] ;
 wire \mem.mem[124][1] ;
 wire \mem.mem[124][2] ;
 wire \mem.mem[124][3] ;
 wire \mem.mem[124][4] ;
 wire \mem.mem[124][5] ;
 wire \mem.mem[124][6] ;
 wire \mem.mem[124][7] ;
 wire \mem.mem[125][0] ;
 wire \mem.mem[125][1] ;
 wire \mem.mem[125][2] ;
 wire \mem.mem[125][3] ;
 wire \mem.mem[125][4] ;
 wire \mem.mem[125][5] ;
 wire \mem.mem[125][6] ;
 wire \mem.mem[125][7] ;
 wire \mem.mem[126][0] ;
 wire \mem.mem[126][1] ;
 wire \mem.mem[126][2] ;
 wire \mem.mem[126][3] ;
 wire \mem.mem[126][4] ;
 wire \mem.mem[126][5] ;
 wire \mem.mem[126][6] ;
 wire \mem.mem[126][7] ;
 wire \mem.mem[127][0] ;
 wire \mem.mem[127][1] ;
 wire \mem.mem[127][2] ;
 wire \mem.mem[127][3] ;
 wire \mem.mem[127][4] ;
 wire \mem.mem[127][5] ;
 wire \mem.mem[127][6] ;
 wire \mem.mem[127][7] ;
 wire \mem.mem[128][0] ;
 wire \mem.mem[128][1] ;
 wire \mem.mem[128][2] ;
 wire \mem.mem[128][3] ;
 wire \mem.mem[128][4] ;
 wire \mem.mem[128][5] ;
 wire \mem.mem[128][6] ;
 wire \mem.mem[128][7] ;
 wire \mem.mem[129][0] ;
 wire \mem.mem[129][1] ;
 wire \mem.mem[129][2] ;
 wire \mem.mem[129][3] ;
 wire \mem.mem[129][4] ;
 wire \mem.mem[129][5] ;
 wire \mem.mem[129][6] ;
 wire \mem.mem[129][7] ;
 wire \mem.mem[12][0] ;
 wire \mem.mem[12][1] ;
 wire \mem.mem[12][2] ;
 wire \mem.mem[12][3] ;
 wire \mem.mem[12][4] ;
 wire \mem.mem[12][5] ;
 wire \mem.mem[12][6] ;
 wire \mem.mem[12][7] ;
 wire \mem.mem[130][0] ;
 wire \mem.mem[130][1] ;
 wire \mem.mem[130][2] ;
 wire \mem.mem[130][3] ;
 wire \mem.mem[130][4] ;
 wire \mem.mem[130][5] ;
 wire \mem.mem[130][6] ;
 wire \mem.mem[130][7] ;
 wire \mem.mem[131][0] ;
 wire \mem.mem[131][1] ;
 wire \mem.mem[131][2] ;
 wire \mem.mem[131][3] ;
 wire \mem.mem[131][4] ;
 wire \mem.mem[131][5] ;
 wire \mem.mem[131][6] ;
 wire \mem.mem[131][7] ;
 wire \mem.mem[132][0] ;
 wire \mem.mem[132][1] ;
 wire \mem.mem[132][2] ;
 wire \mem.mem[132][3] ;
 wire \mem.mem[132][4] ;
 wire \mem.mem[132][5] ;
 wire \mem.mem[132][6] ;
 wire \mem.mem[132][7] ;
 wire \mem.mem[133][0] ;
 wire \mem.mem[133][1] ;
 wire \mem.mem[133][2] ;
 wire \mem.mem[133][3] ;
 wire \mem.mem[133][4] ;
 wire \mem.mem[133][5] ;
 wire \mem.mem[133][6] ;
 wire \mem.mem[133][7] ;
 wire \mem.mem[134][0] ;
 wire \mem.mem[134][1] ;
 wire \mem.mem[134][2] ;
 wire \mem.mem[134][3] ;
 wire \mem.mem[134][4] ;
 wire \mem.mem[134][5] ;
 wire \mem.mem[134][6] ;
 wire \mem.mem[134][7] ;
 wire \mem.mem[135][0] ;
 wire \mem.mem[135][1] ;
 wire \mem.mem[135][2] ;
 wire \mem.mem[135][3] ;
 wire \mem.mem[135][4] ;
 wire \mem.mem[135][5] ;
 wire \mem.mem[135][6] ;
 wire \mem.mem[135][7] ;
 wire \mem.mem[136][0] ;
 wire \mem.mem[136][1] ;
 wire \mem.mem[136][2] ;
 wire \mem.mem[136][3] ;
 wire \mem.mem[136][4] ;
 wire \mem.mem[136][5] ;
 wire \mem.mem[136][6] ;
 wire \mem.mem[136][7] ;
 wire \mem.mem[137][0] ;
 wire \mem.mem[137][1] ;
 wire \mem.mem[137][2] ;
 wire \mem.mem[137][3] ;
 wire \mem.mem[137][4] ;
 wire \mem.mem[137][5] ;
 wire \mem.mem[137][6] ;
 wire \mem.mem[137][7] ;
 wire \mem.mem[138][0] ;
 wire \mem.mem[138][1] ;
 wire \mem.mem[138][2] ;
 wire \mem.mem[138][3] ;
 wire \mem.mem[138][4] ;
 wire \mem.mem[138][5] ;
 wire \mem.mem[138][6] ;
 wire \mem.mem[138][7] ;
 wire \mem.mem[139][0] ;
 wire \mem.mem[139][1] ;
 wire \mem.mem[139][2] ;
 wire \mem.mem[139][3] ;
 wire \mem.mem[139][4] ;
 wire \mem.mem[139][5] ;
 wire \mem.mem[139][6] ;
 wire \mem.mem[139][7] ;
 wire \mem.mem[13][0] ;
 wire \mem.mem[13][1] ;
 wire \mem.mem[13][2] ;
 wire \mem.mem[13][3] ;
 wire \mem.mem[13][4] ;
 wire \mem.mem[13][5] ;
 wire \mem.mem[13][6] ;
 wire \mem.mem[13][7] ;
 wire \mem.mem[140][0] ;
 wire \mem.mem[140][1] ;
 wire \mem.mem[140][2] ;
 wire \mem.mem[140][3] ;
 wire \mem.mem[140][4] ;
 wire \mem.mem[140][5] ;
 wire \mem.mem[140][6] ;
 wire \mem.mem[140][7] ;
 wire \mem.mem[141][0] ;
 wire \mem.mem[141][1] ;
 wire \mem.mem[141][2] ;
 wire \mem.mem[141][3] ;
 wire \mem.mem[141][4] ;
 wire \mem.mem[141][5] ;
 wire \mem.mem[141][6] ;
 wire \mem.mem[141][7] ;
 wire \mem.mem[142][0] ;
 wire \mem.mem[142][1] ;
 wire \mem.mem[142][2] ;
 wire \mem.mem[142][3] ;
 wire \mem.mem[142][4] ;
 wire \mem.mem[142][5] ;
 wire \mem.mem[142][6] ;
 wire \mem.mem[142][7] ;
 wire \mem.mem[143][0] ;
 wire \mem.mem[143][1] ;
 wire \mem.mem[143][2] ;
 wire \mem.mem[143][3] ;
 wire \mem.mem[143][4] ;
 wire \mem.mem[143][5] ;
 wire \mem.mem[143][6] ;
 wire \mem.mem[143][7] ;
 wire \mem.mem[144][0] ;
 wire \mem.mem[144][1] ;
 wire \mem.mem[144][2] ;
 wire \mem.mem[144][3] ;
 wire \mem.mem[144][4] ;
 wire \mem.mem[144][5] ;
 wire \mem.mem[144][6] ;
 wire \mem.mem[144][7] ;
 wire \mem.mem[145][0] ;
 wire \mem.mem[145][1] ;
 wire \mem.mem[145][2] ;
 wire \mem.mem[145][3] ;
 wire \mem.mem[145][4] ;
 wire \mem.mem[145][5] ;
 wire \mem.mem[145][6] ;
 wire \mem.mem[145][7] ;
 wire \mem.mem[146][0] ;
 wire \mem.mem[146][1] ;
 wire \mem.mem[146][2] ;
 wire \mem.mem[146][3] ;
 wire \mem.mem[146][4] ;
 wire \mem.mem[146][5] ;
 wire \mem.mem[146][6] ;
 wire \mem.mem[146][7] ;
 wire \mem.mem[147][0] ;
 wire \mem.mem[147][1] ;
 wire \mem.mem[147][2] ;
 wire \mem.mem[147][3] ;
 wire \mem.mem[147][4] ;
 wire \mem.mem[147][5] ;
 wire \mem.mem[147][6] ;
 wire \mem.mem[147][7] ;
 wire \mem.mem[148][0] ;
 wire \mem.mem[148][1] ;
 wire \mem.mem[148][2] ;
 wire \mem.mem[148][3] ;
 wire \mem.mem[148][4] ;
 wire \mem.mem[148][5] ;
 wire \mem.mem[148][6] ;
 wire \mem.mem[148][7] ;
 wire \mem.mem[149][0] ;
 wire \mem.mem[149][1] ;
 wire \mem.mem[149][2] ;
 wire \mem.mem[149][3] ;
 wire \mem.mem[149][4] ;
 wire \mem.mem[149][5] ;
 wire \mem.mem[149][6] ;
 wire \mem.mem[149][7] ;
 wire \mem.mem[14][0] ;
 wire \mem.mem[14][1] ;
 wire \mem.mem[14][2] ;
 wire \mem.mem[14][3] ;
 wire \mem.mem[14][4] ;
 wire \mem.mem[14][5] ;
 wire \mem.mem[14][6] ;
 wire \mem.mem[14][7] ;
 wire \mem.mem[150][0] ;
 wire \mem.mem[150][1] ;
 wire \mem.mem[150][2] ;
 wire \mem.mem[150][3] ;
 wire \mem.mem[150][4] ;
 wire \mem.mem[150][5] ;
 wire \mem.mem[150][6] ;
 wire \mem.mem[150][7] ;
 wire \mem.mem[151][0] ;
 wire \mem.mem[151][1] ;
 wire \mem.mem[151][2] ;
 wire \mem.mem[151][3] ;
 wire \mem.mem[151][4] ;
 wire \mem.mem[151][5] ;
 wire \mem.mem[151][6] ;
 wire \mem.mem[151][7] ;
 wire \mem.mem[152][0] ;
 wire \mem.mem[152][1] ;
 wire \mem.mem[152][2] ;
 wire \mem.mem[152][3] ;
 wire \mem.mem[152][4] ;
 wire \mem.mem[152][5] ;
 wire \mem.mem[152][6] ;
 wire \mem.mem[152][7] ;
 wire \mem.mem[153][0] ;
 wire \mem.mem[153][1] ;
 wire \mem.mem[153][2] ;
 wire \mem.mem[153][3] ;
 wire \mem.mem[153][4] ;
 wire \mem.mem[153][5] ;
 wire \mem.mem[153][6] ;
 wire \mem.mem[153][7] ;
 wire \mem.mem[154][0] ;
 wire \mem.mem[154][1] ;
 wire \mem.mem[154][2] ;
 wire \mem.mem[154][3] ;
 wire \mem.mem[154][4] ;
 wire \mem.mem[154][5] ;
 wire \mem.mem[154][6] ;
 wire \mem.mem[154][7] ;
 wire \mem.mem[155][0] ;
 wire \mem.mem[155][1] ;
 wire \mem.mem[155][2] ;
 wire \mem.mem[155][3] ;
 wire \mem.mem[155][4] ;
 wire \mem.mem[155][5] ;
 wire \mem.mem[155][6] ;
 wire \mem.mem[155][7] ;
 wire \mem.mem[156][0] ;
 wire \mem.mem[156][1] ;
 wire \mem.mem[156][2] ;
 wire \mem.mem[156][3] ;
 wire \mem.mem[156][4] ;
 wire \mem.mem[156][5] ;
 wire \mem.mem[156][6] ;
 wire \mem.mem[156][7] ;
 wire \mem.mem[157][0] ;
 wire \mem.mem[157][1] ;
 wire \mem.mem[157][2] ;
 wire \mem.mem[157][3] ;
 wire \mem.mem[157][4] ;
 wire \mem.mem[157][5] ;
 wire \mem.mem[157][6] ;
 wire \mem.mem[157][7] ;
 wire \mem.mem[158][0] ;
 wire \mem.mem[158][1] ;
 wire \mem.mem[158][2] ;
 wire \mem.mem[158][3] ;
 wire \mem.mem[158][4] ;
 wire \mem.mem[158][5] ;
 wire \mem.mem[158][6] ;
 wire \mem.mem[158][7] ;
 wire \mem.mem[159][0] ;
 wire \mem.mem[159][1] ;
 wire \mem.mem[159][2] ;
 wire \mem.mem[159][3] ;
 wire \mem.mem[159][4] ;
 wire \mem.mem[159][5] ;
 wire \mem.mem[159][6] ;
 wire \mem.mem[159][7] ;
 wire \mem.mem[15][0] ;
 wire \mem.mem[15][1] ;
 wire \mem.mem[15][2] ;
 wire \mem.mem[15][3] ;
 wire \mem.mem[15][4] ;
 wire \mem.mem[15][5] ;
 wire \mem.mem[15][6] ;
 wire \mem.mem[15][7] ;
 wire \mem.mem[160][0] ;
 wire \mem.mem[160][1] ;
 wire \mem.mem[160][2] ;
 wire \mem.mem[160][3] ;
 wire \mem.mem[160][4] ;
 wire \mem.mem[160][5] ;
 wire \mem.mem[160][6] ;
 wire \mem.mem[160][7] ;
 wire \mem.mem[161][0] ;
 wire \mem.mem[161][1] ;
 wire \mem.mem[161][2] ;
 wire \mem.mem[161][3] ;
 wire \mem.mem[161][4] ;
 wire \mem.mem[161][5] ;
 wire \mem.mem[161][6] ;
 wire \mem.mem[161][7] ;
 wire \mem.mem[162][0] ;
 wire \mem.mem[162][1] ;
 wire \mem.mem[162][2] ;
 wire \mem.mem[162][3] ;
 wire \mem.mem[162][4] ;
 wire \mem.mem[162][5] ;
 wire \mem.mem[162][6] ;
 wire \mem.mem[162][7] ;
 wire \mem.mem[163][0] ;
 wire \mem.mem[163][1] ;
 wire \mem.mem[163][2] ;
 wire \mem.mem[163][3] ;
 wire \mem.mem[163][4] ;
 wire \mem.mem[163][5] ;
 wire \mem.mem[163][6] ;
 wire \mem.mem[163][7] ;
 wire \mem.mem[164][0] ;
 wire \mem.mem[164][1] ;
 wire \mem.mem[164][2] ;
 wire \mem.mem[164][3] ;
 wire \mem.mem[164][4] ;
 wire \mem.mem[164][5] ;
 wire \mem.mem[164][6] ;
 wire \mem.mem[164][7] ;
 wire \mem.mem[165][0] ;
 wire \mem.mem[165][1] ;
 wire \mem.mem[165][2] ;
 wire \mem.mem[165][3] ;
 wire \mem.mem[165][4] ;
 wire \mem.mem[165][5] ;
 wire \mem.mem[165][6] ;
 wire \mem.mem[165][7] ;
 wire \mem.mem[166][0] ;
 wire \mem.mem[166][1] ;
 wire \mem.mem[166][2] ;
 wire \mem.mem[166][3] ;
 wire \mem.mem[166][4] ;
 wire \mem.mem[166][5] ;
 wire \mem.mem[166][6] ;
 wire \mem.mem[166][7] ;
 wire \mem.mem[167][0] ;
 wire \mem.mem[167][1] ;
 wire \mem.mem[167][2] ;
 wire \mem.mem[167][3] ;
 wire \mem.mem[167][4] ;
 wire \mem.mem[167][5] ;
 wire \mem.mem[167][6] ;
 wire \mem.mem[167][7] ;
 wire \mem.mem[168][0] ;
 wire \mem.mem[168][1] ;
 wire \mem.mem[168][2] ;
 wire \mem.mem[168][3] ;
 wire \mem.mem[168][4] ;
 wire \mem.mem[168][5] ;
 wire \mem.mem[168][6] ;
 wire \mem.mem[168][7] ;
 wire \mem.mem[169][0] ;
 wire \mem.mem[169][1] ;
 wire \mem.mem[169][2] ;
 wire \mem.mem[169][3] ;
 wire \mem.mem[169][4] ;
 wire \mem.mem[169][5] ;
 wire \mem.mem[169][6] ;
 wire \mem.mem[169][7] ;
 wire \mem.mem[16][0] ;
 wire \mem.mem[16][1] ;
 wire \mem.mem[16][2] ;
 wire \mem.mem[16][3] ;
 wire \mem.mem[16][4] ;
 wire \mem.mem[16][5] ;
 wire \mem.mem[16][6] ;
 wire \mem.mem[16][7] ;
 wire \mem.mem[170][0] ;
 wire \mem.mem[170][1] ;
 wire \mem.mem[170][2] ;
 wire \mem.mem[170][3] ;
 wire \mem.mem[170][4] ;
 wire \mem.mem[170][5] ;
 wire \mem.mem[170][6] ;
 wire \mem.mem[170][7] ;
 wire \mem.mem[171][0] ;
 wire \mem.mem[171][1] ;
 wire \mem.mem[171][2] ;
 wire \mem.mem[171][3] ;
 wire \mem.mem[171][4] ;
 wire \mem.mem[171][5] ;
 wire \mem.mem[171][6] ;
 wire \mem.mem[171][7] ;
 wire \mem.mem[172][0] ;
 wire \mem.mem[172][1] ;
 wire \mem.mem[172][2] ;
 wire \mem.mem[172][3] ;
 wire \mem.mem[172][4] ;
 wire \mem.mem[172][5] ;
 wire \mem.mem[172][6] ;
 wire \mem.mem[172][7] ;
 wire \mem.mem[173][0] ;
 wire \mem.mem[173][1] ;
 wire \mem.mem[173][2] ;
 wire \mem.mem[173][3] ;
 wire \mem.mem[173][4] ;
 wire \mem.mem[173][5] ;
 wire \mem.mem[173][6] ;
 wire \mem.mem[173][7] ;
 wire \mem.mem[174][0] ;
 wire \mem.mem[174][1] ;
 wire \mem.mem[174][2] ;
 wire \mem.mem[174][3] ;
 wire \mem.mem[174][4] ;
 wire \mem.mem[174][5] ;
 wire \mem.mem[174][6] ;
 wire \mem.mem[174][7] ;
 wire \mem.mem[175][0] ;
 wire \mem.mem[175][1] ;
 wire \mem.mem[175][2] ;
 wire \mem.mem[175][3] ;
 wire \mem.mem[175][4] ;
 wire \mem.mem[175][5] ;
 wire \mem.mem[175][6] ;
 wire \mem.mem[175][7] ;
 wire \mem.mem[176][0] ;
 wire \mem.mem[176][1] ;
 wire \mem.mem[176][2] ;
 wire \mem.mem[176][3] ;
 wire \mem.mem[176][4] ;
 wire \mem.mem[176][5] ;
 wire \mem.mem[176][6] ;
 wire \mem.mem[176][7] ;
 wire \mem.mem[177][0] ;
 wire \mem.mem[177][1] ;
 wire \mem.mem[177][2] ;
 wire \mem.mem[177][3] ;
 wire \mem.mem[177][4] ;
 wire \mem.mem[177][5] ;
 wire \mem.mem[177][6] ;
 wire \mem.mem[177][7] ;
 wire \mem.mem[178][0] ;
 wire \mem.mem[178][1] ;
 wire \mem.mem[178][2] ;
 wire \mem.mem[178][3] ;
 wire \mem.mem[178][4] ;
 wire \mem.mem[178][5] ;
 wire \mem.mem[178][6] ;
 wire \mem.mem[178][7] ;
 wire \mem.mem[179][0] ;
 wire \mem.mem[179][1] ;
 wire \mem.mem[179][2] ;
 wire \mem.mem[179][3] ;
 wire \mem.mem[179][4] ;
 wire \mem.mem[179][5] ;
 wire \mem.mem[179][6] ;
 wire \mem.mem[179][7] ;
 wire \mem.mem[17][0] ;
 wire \mem.mem[17][1] ;
 wire \mem.mem[17][2] ;
 wire \mem.mem[17][3] ;
 wire \mem.mem[17][4] ;
 wire \mem.mem[17][5] ;
 wire \mem.mem[17][6] ;
 wire \mem.mem[17][7] ;
 wire \mem.mem[180][0] ;
 wire \mem.mem[180][1] ;
 wire \mem.mem[180][2] ;
 wire \mem.mem[180][3] ;
 wire \mem.mem[180][4] ;
 wire \mem.mem[180][5] ;
 wire \mem.mem[180][6] ;
 wire \mem.mem[180][7] ;
 wire \mem.mem[181][0] ;
 wire \mem.mem[181][1] ;
 wire \mem.mem[181][2] ;
 wire \mem.mem[181][3] ;
 wire \mem.mem[181][4] ;
 wire \mem.mem[181][5] ;
 wire \mem.mem[181][6] ;
 wire \mem.mem[181][7] ;
 wire \mem.mem[182][0] ;
 wire \mem.mem[182][1] ;
 wire \mem.mem[182][2] ;
 wire \mem.mem[182][3] ;
 wire \mem.mem[182][4] ;
 wire \mem.mem[182][5] ;
 wire \mem.mem[182][6] ;
 wire \mem.mem[182][7] ;
 wire \mem.mem[183][0] ;
 wire \mem.mem[183][1] ;
 wire \mem.mem[183][2] ;
 wire \mem.mem[183][3] ;
 wire \mem.mem[183][4] ;
 wire \mem.mem[183][5] ;
 wire \mem.mem[183][6] ;
 wire \mem.mem[183][7] ;
 wire \mem.mem[184][0] ;
 wire \mem.mem[184][1] ;
 wire \mem.mem[184][2] ;
 wire \mem.mem[184][3] ;
 wire \mem.mem[184][4] ;
 wire \mem.mem[184][5] ;
 wire \mem.mem[184][6] ;
 wire \mem.mem[184][7] ;
 wire \mem.mem[185][0] ;
 wire \mem.mem[185][1] ;
 wire \mem.mem[185][2] ;
 wire \mem.mem[185][3] ;
 wire \mem.mem[185][4] ;
 wire \mem.mem[185][5] ;
 wire \mem.mem[185][6] ;
 wire \mem.mem[185][7] ;
 wire \mem.mem[186][0] ;
 wire \mem.mem[186][1] ;
 wire \mem.mem[186][2] ;
 wire \mem.mem[186][3] ;
 wire \mem.mem[186][4] ;
 wire \mem.mem[186][5] ;
 wire \mem.mem[186][6] ;
 wire \mem.mem[186][7] ;
 wire \mem.mem[187][0] ;
 wire \mem.mem[187][1] ;
 wire \mem.mem[187][2] ;
 wire \mem.mem[187][3] ;
 wire \mem.mem[187][4] ;
 wire \mem.mem[187][5] ;
 wire \mem.mem[187][6] ;
 wire \mem.mem[187][7] ;
 wire \mem.mem[188][0] ;
 wire \mem.mem[188][1] ;
 wire \mem.mem[188][2] ;
 wire \mem.mem[188][3] ;
 wire \mem.mem[188][4] ;
 wire \mem.mem[188][5] ;
 wire \mem.mem[188][6] ;
 wire \mem.mem[188][7] ;
 wire \mem.mem[189][0] ;
 wire \mem.mem[189][1] ;
 wire \mem.mem[189][2] ;
 wire \mem.mem[189][3] ;
 wire \mem.mem[189][4] ;
 wire \mem.mem[189][5] ;
 wire \mem.mem[189][6] ;
 wire \mem.mem[189][7] ;
 wire \mem.mem[18][0] ;
 wire \mem.mem[18][1] ;
 wire \mem.mem[18][2] ;
 wire \mem.mem[18][3] ;
 wire \mem.mem[18][4] ;
 wire \mem.mem[18][5] ;
 wire \mem.mem[18][6] ;
 wire \mem.mem[18][7] ;
 wire \mem.mem[190][0] ;
 wire \mem.mem[190][1] ;
 wire \mem.mem[190][2] ;
 wire \mem.mem[190][3] ;
 wire \mem.mem[190][4] ;
 wire \mem.mem[190][5] ;
 wire \mem.mem[190][6] ;
 wire \mem.mem[190][7] ;
 wire \mem.mem[191][0] ;
 wire \mem.mem[191][1] ;
 wire \mem.mem[191][2] ;
 wire \mem.mem[191][3] ;
 wire \mem.mem[191][4] ;
 wire \mem.mem[191][5] ;
 wire \mem.mem[191][6] ;
 wire \mem.mem[191][7] ;
 wire \mem.mem[192][0] ;
 wire \mem.mem[192][1] ;
 wire \mem.mem[192][2] ;
 wire \mem.mem[192][3] ;
 wire \mem.mem[192][4] ;
 wire \mem.mem[192][5] ;
 wire \mem.mem[192][6] ;
 wire \mem.mem[192][7] ;
 wire \mem.mem[193][0] ;
 wire \mem.mem[193][1] ;
 wire \mem.mem[193][2] ;
 wire \mem.mem[193][3] ;
 wire \mem.mem[193][4] ;
 wire \mem.mem[193][5] ;
 wire \mem.mem[193][6] ;
 wire \mem.mem[193][7] ;
 wire \mem.mem[194][0] ;
 wire \mem.mem[194][1] ;
 wire \mem.mem[194][2] ;
 wire \mem.mem[194][3] ;
 wire \mem.mem[194][4] ;
 wire \mem.mem[194][5] ;
 wire \mem.mem[194][6] ;
 wire \mem.mem[194][7] ;
 wire \mem.mem[195][0] ;
 wire \mem.mem[195][1] ;
 wire \mem.mem[195][2] ;
 wire \mem.mem[195][3] ;
 wire \mem.mem[195][4] ;
 wire \mem.mem[195][5] ;
 wire \mem.mem[195][6] ;
 wire \mem.mem[195][7] ;
 wire \mem.mem[196][0] ;
 wire \mem.mem[196][1] ;
 wire \mem.mem[196][2] ;
 wire \mem.mem[196][3] ;
 wire \mem.mem[196][4] ;
 wire \mem.mem[196][5] ;
 wire \mem.mem[196][6] ;
 wire \mem.mem[196][7] ;
 wire \mem.mem[197][0] ;
 wire \mem.mem[197][1] ;
 wire \mem.mem[197][2] ;
 wire \mem.mem[197][3] ;
 wire \mem.mem[197][4] ;
 wire \mem.mem[197][5] ;
 wire \mem.mem[197][6] ;
 wire \mem.mem[197][7] ;
 wire \mem.mem[198][0] ;
 wire \mem.mem[198][1] ;
 wire \mem.mem[198][2] ;
 wire \mem.mem[198][3] ;
 wire \mem.mem[198][4] ;
 wire \mem.mem[198][5] ;
 wire \mem.mem[198][6] ;
 wire \mem.mem[198][7] ;
 wire \mem.mem[199][0] ;
 wire \mem.mem[199][1] ;
 wire \mem.mem[199][2] ;
 wire \mem.mem[199][3] ;
 wire \mem.mem[199][4] ;
 wire \mem.mem[199][5] ;
 wire \mem.mem[199][6] ;
 wire \mem.mem[199][7] ;
 wire \mem.mem[19][0] ;
 wire \mem.mem[19][1] ;
 wire \mem.mem[19][2] ;
 wire \mem.mem[19][3] ;
 wire \mem.mem[19][4] ;
 wire \mem.mem[19][5] ;
 wire \mem.mem[19][6] ;
 wire \mem.mem[19][7] ;
 wire \mem.mem[1][0] ;
 wire \mem.mem[1][1] ;
 wire \mem.mem[1][2] ;
 wire \mem.mem[1][3] ;
 wire \mem.mem[1][4] ;
 wire \mem.mem[1][5] ;
 wire \mem.mem[1][6] ;
 wire \mem.mem[1][7] ;
 wire \mem.mem[200][0] ;
 wire \mem.mem[200][1] ;
 wire \mem.mem[200][2] ;
 wire \mem.mem[200][3] ;
 wire \mem.mem[200][4] ;
 wire \mem.mem[200][5] ;
 wire \mem.mem[200][6] ;
 wire \mem.mem[200][7] ;
 wire \mem.mem[201][0] ;
 wire \mem.mem[201][1] ;
 wire \mem.mem[201][2] ;
 wire \mem.mem[201][3] ;
 wire \mem.mem[201][4] ;
 wire \mem.mem[201][5] ;
 wire \mem.mem[201][6] ;
 wire \mem.mem[201][7] ;
 wire \mem.mem[202][0] ;
 wire \mem.mem[202][1] ;
 wire \mem.mem[202][2] ;
 wire \mem.mem[202][3] ;
 wire \mem.mem[202][4] ;
 wire \mem.mem[202][5] ;
 wire \mem.mem[202][6] ;
 wire \mem.mem[202][7] ;
 wire \mem.mem[203][0] ;
 wire \mem.mem[203][1] ;
 wire \mem.mem[203][2] ;
 wire \mem.mem[203][3] ;
 wire \mem.mem[203][4] ;
 wire \mem.mem[203][5] ;
 wire \mem.mem[203][6] ;
 wire \mem.mem[203][7] ;
 wire \mem.mem[204][0] ;
 wire \mem.mem[204][1] ;
 wire \mem.mem[204][2] ;
 wire \mem.mem[204][3] ;
 wire \mem.mem[204][4] ;
 wire \mem.mem[204][5] ;
 wire \mem.mem[204][6] ;
 wire \mem.mem[204][7] ;
 wire \mem.mem[205][0] ;
 wire \mem.mem[205][1] ;
 wire \mem.mem[205][2] ;
 wire \mem.mem[205][3] ;
 wire \mem.mem[205][4] ;
 wire \mem.mem[205][5] ;
 wire \mem.mem[205][6] ;
 wire \mem.mem[205][7] ;
 wire \mem.mem[206][0] ;
 wire \mem.mem[206][1] ;
 wire \mem.mem[206][2] ;
 wire \mem.mem[206][3] ;
 wire \mem.mem[206][4] ;
 wire \mem.mem[206][5] ;
 wire \mem.mem[206][6] ;
 wire \mem.mem[206][7] ;
 wire \mem.mem[207][0] ;
 wire \mem.mem[207][1] ;
 wire \mem.mem[207][2] ;
 wire \mem.mem[207][3] ;
 wire \mem.mem[207][4] ;
 wire \mem.mem[207][5] ;
 wire \mem.mem[207][6] ;
 wire \mem.mem[207][7] ;
 wire \mem.mem[208][0] ;
 wire \mem.mem[208][1] ;
 wire \mem.mem[208][2] ;
 wire \mem.mem[208][3] ;
 wire \mem.mem[208][4] ;
 wire \mem.mem[208][5] ;
 wire \mem.mem[208][6] ;
 wire \mem.mem[208][7] ;
 wire \mem.mem[209][0] ;
 wire \mem.mem[209][1] ;
 wire \mem.mem[209][2] ;
 wire \mem.mem[209][3] ;
 wire \mem.mem[209][4] ;
 wire \mem.mem[209][5] ;
 wire \mem.mem[209][6] ;
 wire \mem.mem[209][7] ;
 wire \mem.mem[20][0] ;
 wire \mem.mem[20][1] ;
 wire \mem.mem[20][2] ;
 wire \mem.mem[20][3] ;
 wire \mem.mem[20][4] ;
 wire \mem.mem[20][5] ;
 wire \mem.mem[20][6] ;
 wire \mem.mem[20][7] ;
 wire \mem.mem[210][0] ;
 wire \mem.mem[210][1] ;
 wire \mem.mem[210][2] ;
 wire \mem.mem[210][3] ;
 wire \mem.mem[210][4] ;
 wire \mem.mem[210][5] ;
 wire \mem.mem[210][6] ;
 wire \mem.mem[210][7] ;
 wire \mem.mem[211][0] ;
 wire \mem.mem[211][1] ;
 wire \mem.mem[211][2] ;
 wire \mem.mem[211][3] ;
 wire \mem.mem[211][4] ;
 wire \mem.mem[211][5] ;
 wire \mem.mem[211][6] ;
 wire \mem.mem[211][7] ;
 wire \mem.mem[212][0] ;
 wire \mem.mem[212][1] ;
 wire \mem.mem[212][2] ;
 wire \mem.mem[212][3] ;
 wire \mem.mem[212][4] ;
 wire \mem.mem[212][5] ;
 wire \mem.mem[212][6] ;
 wire \mem.mem[212][7] ;
 wire \mem.mem[213][0] ;
 wire \mem.mem[213][1] ;
 wire \mem.mem[213][2] ;
 wire \mem.mem[213][3] ;
 wire \mem.mem[213][4] ;
 wire \mem.mem[213][5] ;
 wire \mem.mem[213][6] ;
 wire \mem.mem[213][7] ;
 wire \mem.mem[214][0] ;
 wire \mem.mem[214][1] ;
 wire \mem.mem[214][2] ;
 wire \mem.mem[214][3] ;
 wire \mem.mem[214][4] ;
 wire \mem.mem[214][5] ;
 wire \mem.mem[214][6] ;
 wire \mem.mem[214][7] ;
 wire \mem.mem[215][0] ;
 wire \mem.mem[215][1] ;
 wire \mem.mem[215][2] ;
 wire \mem.mem[215][3] ;
 wire \mem.mem[215][4] ;
 wire \mem.mem[215][5] ;
 wire \mem.mem[215][6] ;
 wire \mem.mem[215][7] ;
 wire \mem.mem[216][0] ;
 wire \mem.mem[216][1] ;
 wire \mem.mem[216][2] ;
 wire \mem.mem[216][3] ;
 wire \mem.mem[216][4] ;
 wire \mem.mem[216][5] ;
 wire \mem.mem[216][6] ;
 wire \mem.mem[216][7] ;
 wire \mem.mem[217][0] ;
 wire \mem.mem[217][1] ;
 wire \mem.mem[217][2] ;
 wire \mem.mem[217][3] ;
 wire \mem.mem[217][4] ;
 wire \mem.mem[217][5] ;
 wire \mem.mem[217][6] ;
 wire \mem.mem[217][7] ;
 wire \mem.mem[218][0] ;
 wire \mem.mem[218][1] ;
 wire \mem.mem[218][2] ;
 wire \mem.mem[218][3] ;
 wire \mem.mem[218][4] ;
 wire \mem.mem[218][5] ;
 wire \mem.mem[218][6] ;
 wire \mem.mem[218][7] ;
 wire \mem.mem[219][0] ;
 wire \mem.mem[219][1] ;
 wire \mem.mem[219][2] ;
 wire \mem.mem[219][3] ;
 wire \mem.mem[219][4] ;
 wire \mem.mem[219][5] ;
 wire \mem.mem[219][6] ;
 wire \mem.mem[219][7] ;
 wire \mem.mem[21][0] ;
 wire \mem.mem[21][1] ;
 wire \mem.mem[21][2] ;
 wire \mem.mem[21][3] ;
 wire \mem.mem[21][4] ;
 wire \mem.mem[21][5] ;
 wire \mem.mem[21][6] ;
 wire \mem.mem[21][7] ;
 wire \mem.mem[220][0] ;
 wire \mem.mem[220][1] ;
 wire \mem.mem[220][2] ;
 wire \mem.mem[220][3] ;
 wire \mem.mem[220][4] ;
 wire \mem.mem[220][5] ;
 wire \mem.mem[220][6] ;
 wire \mem.mem[220][7] ;
 wire \mem.mem[221][0] ;
 wire \mem.mem[221][1] ;
 wire \mem.mem[221][2] ;
 wire \mem.mem[221][3] ;
 wire \mem.mem[221][4] ;
 wire \mem.mem[221][5] ;
 wire \mem.mem[221][6] ;
 wire \mem.mem[221][7] ;
 wire \mem.mem[222][0] ;
 wire \mem.mem[222][1] ;
 wire \mem.mem[222][2] ;
 wire \mem.mem[222][3] ;
 wire \mem.mem[222][4] ;
 wire \mem.mem[222][5] ;
 wire \mem.mem[222][6] ;
 wire \mem.mem[222][7] ;
 wire \mem.mem[223][0] ;
 wire \mem.mem[223][1] ;
 wire \mem.mem[223][2] ;
 wire \mem.mem[223][3] ;
 wire \mem.mem[223][4] ;
 wire \mem.mem[223][5] ;
 wire \mem.mem[223][6] ;
 wire \mem.mem[223][7] ;
 wire \mem.mem[224][0] ;
 wire \mem.mem[224][1] ;
 wire \mem.mem[224][2] ;
 wire \mem.mem[224][3] ;
 wire \mem.mem[224][4] ;
 wire \mem.mem[224][5] ;
 wire \mem.mem[224][6] ;
 wire \mem.mem[224][7] ;
 wire \mem.mem[225][0] ;
 wire \mem.mem[225][1] ;
 wire \mem.mem[225][2] ;
 wire \mem.mem[225][3] ;
 wire \mem.mem[225][4] ;
 wire \mem.mem[225][5] ;
 wire \mem.mem[225][6] ;
 wire \mem.mem[225][7] ;
 wire \mem.mem[226][0] ;
 wire \mem.mem[226][1] ;
 wire \mem.mem[226][2] ;
 wire \mem.mem[226][3] ;
 wire \mem.mem[226][4] ;
 wire \mem.mem[226][5] ;
 wire \mem.mem[226][6] ;
 wire \mem.mem[226][7] ;
 wire \mem.mem[227][0] ;
 wire \mem.mem[227][1] ;
 wire \mem.mem[227][2] ;
 wire \mem.mem[227][3] ;
 wire \mem.mem[227][4] ;
 wire \mem.mem[227][5] ;
 wire \mem.mem[227][6] ;
 wire \mem.mem[227][7] ;
 wire \mem.mem[228][0] ;
 wire \mem.mem[228][1] ;
 wire \mem.mem[228][2] ;
 wire \mem.mem[228][3] ;
 wire \mem.mem[228][4] ;
 wire \mem.mem[228][5] ;
 wire \mem.mem[228][6] ;
 wire \mem.mem[228][7] ;
 wire \mem.mem[229][0] ;
 wire \mem.mem[229][1] ;
 wire \mem.mem[229][2] ;
 wire \mem.mem[229][3] ;
 wire \mem.mem[229][4] ;
 wire \mem.mem[229][5] ;
 wire \mem.mem[229][6] ;
 wire \mem.mem[229][7] ;
 wire \mem.mem[22][0] ;
 wire \mem.mem[22][1] ;
 wire \mem.mem[22][2] ;
 wire \mem.mem[22][3] ;
 wire \mem.mem[22][4] ;
 wire \mem.mem[22][5] ;
 wire \mem.mem[22][6] ;
 wire \mem.mem[22][7] ;
 wire \mem.mem[230][0] ;
 wire \mem.mem[230][1] ;
 wire \mem.mem[230][2] ;
 wire \mem.mem[230][3] ;
 wire \mem.mem[230][4] ;
 wire \mem.mem[230][5] ;
 wire \mem.mem[230][6] ;
 wire \mem.mem[230][7] ;
 wire \mem.mem[231][0] ;
 wire \mem.mem[231][1] ;
 wire \mem.mem[231][2] ;
 wire \mem.mem[231][3] ;
 wire \mem.mem[231][4] ;
 wire \mem.mem[231][5] ;
 wire \mem.mem[231][6] ;
 wire \mem.mem[231][7] ;
 wire \mem.mem[232][0] ;
 wire \mem.mem[232][1] ;
 wire \mem.mem[232][2] ;
 wire \mem.mem[232][3] ;
 wire \mem.mem[232][4] ;
 wire \mem.mem[232][5] ;
 wire \mem.mem[232][6] ;
 wire \mem.mem[232][7] ;
 wire \mem.mem[233][0] ;
 wire \mem.mem[233][1] ;
 wire \mem.mem[233][2] ;
 wire \mem.mem[233][3] ;
 wire \mem.mem[233][4] ;
 wire \mem.mem[233][5] ;
 wire \mem.mem[233][6] ;
 wire \mem.mem[233][7] ;
 wire \mem.mem[234][0] ;
 wire \mem.mem[234][1] ;
 wire \mem.mem[234][2] ;
 wire \mem.mem[234][3] ;
 wire \mem.mem[234][4] ;
 wire \mem.mem[234][5] ;
 wire \mem.mem[234][6] ;
 wire \mem.mem[234][7] ;
 wire \mem.mem[235][0] ;
 wire \mem.mem[235][1] ;
 wire \mem.mem[235][2] ;
 wire \mem.mem[235][3] ;
 wire \mem.mem[235][4] ;
 wire \mem.mem[235][5] ;
 wire \mem.mem[235][6] ;
 wire \mem.mem[235][7] ;
 wire \mem.mem[236][0] ;
 wire \mem.mem[236][1] ;
 wire \mem.mem[236][2] ;
 wire \mem.mem[236][3] ;
 wire \mem.mem[236][4] ;
 wire \mem.mem[236][5] ;
 wire \mem.mem[236][6] ;
 wire \mem.mem[236][7] ;
 wire \mem.mem[237][0] ;
 wire \mem.mem[237][1] ;
 wire \mem.mem[237][2] ;
 wire \mem.mem[237][3] ;
 wire \mem.mem[237][4] ;
 wire \mem.mem[237][5] ;
 wire \mem.mem[237][6] ;
 wire \mem.mem[237][7] ;
 wire \mem.mem[238][0] ;
 wire \mem.mem[238][1] ;
 wire \mem.mem[238][2] ;
 wire \mem.mem[238][3] ;
 wire \mem.mem[238][4] ;
 wire \mem.mem[238][5] ;
 wire \mem.mem[238][6] ;
 wire \mem.mem[238][7] ;
 wire \mem.mem[239][0] ;
 wire \mem.mem[239][1] ;
 wire \mem.mem[239][2] ;
 wire \mem.mem[239][3] ;
 wire \mem.mem[239][4] ;
 wire \mem.mem[239][5] ;
 wire \mem.mem[239][6] ;
 wire \mem.mem[239][7] ;
 wire \mem.mem[23][0] ;
 wire \mem.mem[23][1] ;
 wire \mem.mem[23][2] ;
 wire \mem.mem[23][3] ;
 wire \mem.mem[23][4] ;
 wire \mem.mem[23][5] ;
 wire \mem.mem[23][6] ;
 wire \mem.mem[23][7] ;
 wire \mem.mem[240][0] ;
 wire \mem.mem[240][1] ;
 wire \mem.mem[240][2] ;
 wire \mem.mem[240][3] ;
 wire \mem.mem[240][4] ;
 wire \mem.mem[240][5] ;
 wire \mem.mem[240][6] ;
 wire \mem.mem[240][7] ;
 wire \mem.mem[241][0] ;
 wire \mem.mem[241][1] ;
 wire \mem.mem[241][2] ;
 wire \mem.mem[241][3] ;
 wire \mem.mem[241][4] ;
 wire \mem.mem[241][5] ;
 wire \mem.mem[241][6] ;
 wire \mem.mem[241][7] ;
 wire \mem.mem[242][0] ;
 wire \mem.mem[242][1] ;
 wire \mem.mem[242][2] ;
 wire \mem.mem[242][3] ;
 wire \mem.mem[242][4] ;
 wire \mem.mem[242][5] ;
 wire \mem.mem[242][6] ;
 wire \mem.mem[242][7] ;
 wire \mem.mem[243][0] ;
 wire \mem.mem[243][1] ;
 wire \mem.mem[243][2] ;
 wire \mem.mem[243][3] ;
 wire \mem.mem[243][4] ;
 wire \mem.mem[243][5] ;
 wire \mem.mem[243][6] ;
 wire \mem.mem[243][7] ;
 wire \mem.mem[244][0] ;
 wire \mem.mem[244][1] ;
 wire \mem.mem[244][2] ;
 wire \mem.mem[244][3] ;
 wire \mem.mem[244][4] ;
 wire \mem.mem[244][5] ;
 wire \mem.mem[244][6] ;
 wire \mem.mem[244][7] ;
 wire \mem.mem[245][0] ;
 wire \mem.mem[245][1] ;
 wire \mem.mem[245][2] ;
 wire \mem.mem[245][3] ;
 wire \mem.mem[245][4] ;
 wire \mem.mem[245][5] ;
 wire \mem.mem[245][6] ;
 wire \mem.mem[245][7] ;
 wire \mem.mem[246][0] ;
 wire \mem.mem[246][1] ;
 wire \mem.mem[246][2] ;
 wire \mem.mem[246][3] ;
 wire \mem.mem[246][4] ;
 wire \mem.mem[246][5] ;
 wire \mem.mem[246][6] ;
 wire \mem.mem[246][7] ;
 wire \mem.mem[247][0] ;
 wire \mem.mem[247][1] ;
 wire \mem.mem[247][2] ;
 wire \mem.mem[247][3] ;
 wire \mem.mem[247][4] ;
 wire \mem.mem[247][5] ;
 wire \mem.mem[247][6] ;
 wire \mem.mem[247][7] ;
 wire \mem.mem[248][0] ;
 wire \mem.mem[248][1] ;
 wire \mem.mem[248][2] ;
 wire \mem.mem[248][3] ;
 wire \mem.mem[248][4] ;
 wire \mem.mem[248][5] ;
 wire \mem.mem[248][6] ;
 wire \mem.mem[248][7] ;
 wire \mem.mem[249][0] ;
 wire \mem.mem[249][1] ;
 wire \mem.mem[249][2] ;
 wire \mem.mem[249][3] ;
 wire \mem.mem[249][4] ;
 wire \mem.mem[249][5] ;
 wire \mem.mem[249][6] ;
 wire \mem.mem[249][7] ;
 wire \mem.mem[24][0] ;
 wire \mem.mem[24][1] ;
 wire \mem.mem[24][2] ;
 wire \mem.mem[24][3] ;
 wire \mem.mem[24][4] ;
 wire \mem.mem[24][5] ;
 wire \mem.mem[24][6] ;
 wire \mem.mem[24][7] ;
 wire \mem.mem[250][0] ;
 wire \mem.mem[250][1] ;
 wire \mem.mem[250][2] ;
 wire \mem.mem[250][3] ;
 wire \mem.mem[250][4] ;
 wire \mem.mem[250][5] ;
 wire \mem.mem[250][6] ;
 wire \mem.mem[250][7] ;
 wire \mem.mem[251][0] ;
 wire \mem.mem[251][1] ;
 wire \mem.mem[251][2] ;
 wire \mem.mem[251][3] ;
 wire \mem.mem[251][4] ;
 wire \mem.mem[251][5] ;
 wire \mem.mem[251][6] ;
 wire \mem.mem[251][7] ;
 wire \mem.mem[252][0] ;
 wire \mem.mem[252][1] ;
 wire \mem.mem[252][2] ;
 wire \mem.mem[252][3] ;
 wire \mem.mem[252][4] ;
 wire \mem.mem[252][5] ;
 wire \mem.mem[252][6] ;
 wire \mem.mem[252][7] ;
 wire \mem.mem[25][0] ;
 wire \mem.mem[25][1] ;
 wire \mem.mem[25][2] ;
 wire \mem.mem[25][3] ;
 wire \mem.mem[25][4] ;
 wire \mem.mem[25][5] ;
 wire \mem.mem[25][6] ;
 wire \mem.mem[25][7] ;
 wire \mem.mem[26][0] ;
 wire \mem.mem[26][1] ;
 wire \mem.mem[26][2] ;
 wire \mem.mem[26][3] ;
 wire \mem.mem[26][4] ;
 wire \mem.mem[26][5] ;
 wire \mem.mem[26][6] ;
 wire \mem.mem[26][7] ;
 wire \mem.mem[27][0] ;
 wire \mem.mem[27][1] ;
 wire \mem.mem[27][2] ;
 wire \mem.mem[27][3] ;
 wire \mem.mem[27][4] ;
 wire \mem.mem[27][5] ;
 wire \mem.mem[27][6] ;
 wire \mem.mem[27][7] ;
 wire \mem.mem[28][0] ;
 wire \mem.mem[28][1] ;
 wire \mem.mem[28][2] ;
 wire \mem.mem[28][3] ;
 wire \mem.mem[28][4] ;
 wire \mem.mem[28][5] ;
 wire \mem.mem[28][6] ;
 wire \mem.mem[28][7] ;
 wire \mem.mem[29][0] ;
 wire \mem.mem[29][1] ;
 wire \mem.mem[29][2] ;
 wire \mem.mem[29][3] ;
 wire \mem.mem[29][4] ;
 wire \mem.mem[29][5] ;
 wire \mem.mem[29][6] ;
 wire \mem.mem[29][7] ;
 wire \mem.mem[2][0] ;
 wire \mem.mem[2][1] ;
 wire \mem.mem[2][2] ;
 wire \mem.mem[2][3] ;
 wire \mem.mem[2][4] ;
 wire \mem.mem[2][5] ;
 wire \mem.mem[2][6] ;
 wire \mem.mem[2][7] ;
 wire \mem.mem[30][0] ;
 wire \mem.mem[30][1] ;
 wire \mem.mem[30][2] ;
 wire \mem.mem[30][3] ;
 wire \mem.mem[30][4] ;
 wire \mem.mem[30][5] ;
 wire \mem.mem[30][6] ;
 wire \mem.mem[30][7] ;
 wire \mem.mem[31][0] ;
 wire \mem.mem[31][1] ;
 wire \mem.mem[31][2] ;
 wire \mem.mem[31][3] ;
 wire \mem.mem[31][4] ;
 wire \mem.mem[31][5] ;
 wire \mem.mem[31][6] ;
 wire \mem.mem[31][7] ;
 wire \mem.mem[32][0] ;
 wire \mem.mem[32][1] ;
 wire \mem.mem[32][2] ;
 wire \mem.mem[32][3] ;
 wire \mem.mem[32][4] ;
 wire \mem.mem[32][5] ;
 wire \mem.mem[32][6] ;
 wire \mem.mem[32][7] ;
 wire \mem.mem[33][0] ;
 wire \mem.mem[33][1] ;
 wire \mem.mem[33][2] ;
 wire \mem.mem[33][3] ;
 wire \mem.mem[33][4] ;
 wire \mem.mem[33][5] ;
 wire \mem.mem[33][6] ;
 wire \mem.mem[33][7] ;
 wire \mem.mem[34][0] ;
 wire \mem.mem[34][1] ;
 wire \mem.mem[34][2] ;
 wire \mem.mem[34][3] ;
 wire \mem.mem[34][4] ;
 wire \mem.mem[34][5] ;
 wire \mem.mem[34][6] ;
 wire \mem.mem[34][7] ;
 wire \mem.mem[35][0] ;
 wire \mem.mem[35][1] ;
 wire \mem.mem[35][2] ;
 wire \mem.mem[35][3] ;
 wire \mem.mem[35][4] ;
 wire \mem.mem[35][5] ;
 wire \mem.mem[35][6] ;
 wire \mem.mem[35][7] ;
 wire \mem.mem[36][0] ;
 wire \mem.mem[36][1] ;
 wire \mem.mem[36][2] ;
 wire \mem.mem[36][3] ;
 wire \mem.mem[36][4] ;
 wire \mem.mem[36][5] ;
 wire \mem.mem[36][6] ;
 wire \mem.mem[36][7] ;
 wire \mem.mem[37][0] ;
 wire \mem.mem[37][1] ;
 wire \mem.mem[37][2] ;
 wire \mem.mem[37][3] ;
 wire \mem.mem[37][4] ;
 wire \mem.mem[37][5] ;
 wire \mem.mem[37][6] ;
 wire \mem.mem[37][7] ;
 wire \mem.mem[38][0] ;
 wire \mem.mem[38][1] ;
 wire \mem.mem[38][2] ;
 wire \mem.mem[38][3] ;
 wire \mem.mem[38][4] ;
 wire \mem.mem[38][5] ;
 wire \mem.mem[38][6] ;
 wire \mem.mem[38][7] ;
 wire \mem.mem[39][0] ;
 wire \mem.mem[39][1] ;
 wire \mem.mem[39][2] ;
 wire \mem.mem[39][3] ;
 wire \mem.mem[39][4] ;
 wire \mem.mem[39][5] ;
 wire \mem.mem[39][6] ;
 wire \mem.mem[39][7] ;
 wire \mem.mem[3][0] ;
 wire \mem.mem[3][1] ;
 wire \mem.mem[3][2] ;
 wire \mem.mem[3][3] ;
 wire \mem.mem[3][4] ;
 wire \mem.mem[3][5] ;
 wire \mem.mem[3][6] ;
 wire \mem.mem[3][7] ;
 wire \mem.mem[40][0] ;
 wire \mem.mem[40][1] ;
 wire \mem.mem[40][2] ;
 wire \mem.mem[40][3] ;
 wire \mem.mem[40][4] ;
 wire \mem.mem[40][5] ;
 wire \mem.mem[40][6] ;
 wire \mem.mem[40][7] ;
 wire \mem.mem[41][0] ;
 wire \mem.mem[41][1] ;
 wire \mem.mem[41][2] ;
 wire \mem.mem[41][3] ;
 wire \mem.mem[41][4] ;
 wire \mem.mem[41][5] ;
 wire \mem.mem[41][6] ;
 wire \mem.mem[41][7] ;
 wire \mem.mem[42][0] ;
 wire \mem.mem[42][1] ;
 wire \mem.mem[42][2] ;
 wire \mem.mem[42][3] ;
 wire \mem.mem[42][4] ;
 wire \mem.mem[42][5] ;
 wire \mem.mem[42][6] ;
 wire \mem.mem[42][7] ;
 wire \mem.mem[43][0] ;
 wire \mem.mem[43][1] ;
 wire \mem.mem[43][2] ;
 wire \mem.mem[43][3] ;
 wire \mem.mem[43][4] ;
 wire \mem.mem[43][5] ;
 wire \mem.mem[43][6] ;
 wire \mem.mem[43][7] ;
 wire \mem.mem[44][0] ;
 wire \mem.mem[44][1] ;
 wire \mem.mem[44][2] ;
 wire \mem.mem[44][3] ;
 wire \mem.mem[44][4] ;
 wire \mem.mem[44][5] ;
 wire \mem.mem[44][6] ;
 wire \mem.mem[44][7] ;
 wire \mem.mem[45][0] ;
 wire \mem.mem[45][1] ;
 wire \mem.mem[45][2] ;
 wire \mem.mem[45][3] ;
 wire \mem.mem[45][4] ;
 wire \mem.mem[45][5] ;
 wire \mem.mem[45][6] ;
 wire \mem.mem[45][7] ;
 wire \mem.mem[46][0] ;
 wire \mem.mem[46][1] ;
 wire \mem.mem[46][2] ;
 wire \mem.mem[46][3] ;
 wire \mem.mem[46][4] ;
 wire \mem.mem[46][5] ;
 wire \mem.mem[46][6] ;
 wire \mem.mem[46][7] ;
 wire \mem.mem[47][0] ;
 wire \mem.mem[47][1] ;
 wire \mem.mem[47][2] ;
 wire \mem.mem[47][3] ;
 wire \mem.mem[47][4] ;
 wire \mem.mem[47][5] ;
 wire \mem.mem[47][6] ;
 wire \mem.mem[47][7] ;
 wire \mem.mem[48][0] ;
 wire \mem.mem[48][1] ;
 wire \mem.mem[48][2] ;
 wire \mem.mem[48][3] ;
 wire \mem.mem[48][4] ;
 wire \mem.mem[48][5] ;
 wire \mem.mem[48][6] ;
 wire \mem.mem[48][7] ;
 wire \mem.mem[49][0] ;
 wire \mem.mem[49][1] ;
 wire \mem.mem[49][2] ;
 wire \mem.mem[49][3] ;
 wire \mem.mem[49][4] ;
 wire \mem.mem[49][5] ;
 wire \mem.mem[49][6] ;
 wire \mem.mem[49][7] ;
 wire \mem.mem[4][0] ;
 wire \mem.mem[4][1] ;
 wire \mem.mem[4][2] ;
 wire \mem.mem[4][3] ;
 wire \mem.mem[4][4] ;
 wire \mem.mem[4][5] ;
 wire \mem.mem[4][6] ;
 wire \mem.mem[4][7] ;
 wire \mem.mem[50][0] ;
 wire \mem.mem[50][1] ;
 wire \mem.mem[50][2] ;
 wire \mem.mem[50][3] ;
 wire \mem.mem[50][4] ;
 wire \mem.mem[50][5] ;
 wire \mem.mem[50][6] ;
 wire \mem.mem[50][7] ;
 wire \mem.mem[51][0] ;
 wire \mem.mem[51][1] ;
 wire \mem.mem[51][2] ;
 wire \mem.mem[51][3] ;
 wire \mem.mem[51][4] ;
 wire \mem.mem[51][5] ;
 wire \mem.mem[51][6] ;
 wire \mem.mem[51][7] ;
 wire \mem.mem[52][0] ;
 wire \mem.mem[52][1] ;
 wire \mem.mem[52][2] ;
 wire \mem.mem[52][3] ;
 wire \mem.mem[52][4] ;
 wire \mem.mem[52][5] ;
 wire \mem.mem[52][6] ;
 wire \mem.mem[52][7] ;
 wire \mem.mem[53][0] ;
 wire \mem.mem[53][1] ;
 wire \mem.mem[53][2] ;
 wire \mem.mem[53][3] ;
 wire \mem.mem[53][4] ;
 wire \mem.mem[53][5] ;
 wire \mem.mem[53][6] ;
 wire \mem.mem[53][7] ;
 wire \mem.mem[54][0] ;
 wire \mem.mem[54][1] ;
 wire \mem.mem[54][2] ;
 wire \mem.mem[54][3] ;
 wire \mem.mem[54][4] ;
 wire \mem.mem[54][5] ;
 wire \mem.mem[54][6] ;
 wire \mem.mem[54][7] ;
 wire \mem.mem[55][0] ;
 wire \mem.mem[55][1] ;
 wire \mem.mem[55][2] ;
 wire \mem.mem[55][3] ;
 wire \mem.mem[55][4] ;
 wire \mem.mem[55][5] ;
 wire \mem.mem[55][6] ;
 wire \mem.mem[55][7] ;
 wire \mem.mem[56][0] ;
 wire \mem.mem[56][1] ;
 wire \mem.mem[56][2] ;
 wire \mem.mem[56][3] ;
 wire \mem.mem[56][4] ;
 wire \mem.mem[56][5] ;
 wire \mem.mem[56][6] ;
 wire \mem.mem[56][7] ;
 wire \mem.mem[57][0] ;
 wire \mem.mem[57][1] ;
 wire \mem.mem[57][2] ;
 wire \mem.mem[57][3] ;
 wire \mem.mem[57][4] ;
 wire \mem.mem[57][5] ;
 wire \mem.mem[57][6] ;
 wire \mem.mem[57][7] ;
 wire \mem.mem[58][0] ;
 wire \mem.mem[58][1] ;
 wire \mem.mem[58][2] ;
 wire \mem.mem[58][3] ;
 wire \mem.mem[58][4] ;
 wire \mem.mem[58][5] ;
 wire \mem.mem[58][6] ;
 wire \mem.mem[58][7] ;
 wire \mem.mem[59][0] ;
 wire \mem.mem[59][1] ;
 wire \mem.mem[59][2] ;
 wire \mem.mem[59][3] ;
 wire \mem.mem[59][4] ;
 wire \mem.mem[59][5] ;
 wire \mem.mem[59][6] ;
 wire \mem.mem[59][7] ;
 wire \mem.mem[5][0] ;
 wire \mem.mem[5][1] ;
 wire \mem.mem[5][2] ;
 wire \mem.mem[5][3] ;
 wire \mem.mem[5][4] ;
 wire \mem.mem[5][5] ;
 wire \mem.mem[5][6] ;
 wire \mem.mem[5][7] ;
 wire \mem.mem[60][0] ;
 wire \mem.mem[60][1] ;
 wire \mem.mem[60][2] ;
 wire \mem.mem[60][3] ;
 wire \mem.mem[60][4] ;
 wire \mem.mem[60][5] ;
 wire \mem.mem[60][6] ;
 wire \mem.mem[60][7] ;
 wire \mem.mem[61][0] ;
 wire \mem.mem[61][1] ;
 wire \mem.mem[61][2] ;
 wire \mem.mem[61][3] ;
 wire \mem.mem[61][4] ;
 wire \mem.mem[61][5] ;
 wire \mem.mem[61][6] ;
 wire \mem.mem[61][7] ;
 wire \mem.mem[62][0] ;
 wire \mem.mem[62][1] ;
 wire \mem.mem[62][2] ;
 wire \mem.mem[62][3] ;
 wire \mem.mem[62][4] ;
 wire \mem.mem[62][5] ;
 wire \mem.mem[62][6] ;
 wire \mem.mem[62][7] ;
 wire \mem.mem[63][0] ;
 wire \mem.mem[63][1] ;
 wire \mem.mem[63][2] ;
 wire \mem.mem[63][3] ;
 wire \mem.mem[63][4] ;
 wire \mem.mem[63][5] ;
 wire \mem.mem[63][6] ;
 wire \mem.mem[63][7] ;
 wire \mem.mem[64][0] ;
 wire \mem.mem[64][1] ;
 wire \mem.mem[64][2] ;
 wire \mem.mem[64][3] ;
 wire \mem.mem[64][4] ;
 wire \mem.mem[64][5] ;
 wire \mem.mem[64][6] ;
 wire \mem.mem[64][7] ;
 wire \mem.mem[65][0] ;
 wire \mem.mem[65][1] ;
 wire \mem.mem[65][2] ;
 wire \mem.mem[65][3] ;
 wire \mem.mem[65][4] ;
 wire \mem.mem[65][5] ;
 wire \mem.mem[65][6] ;
 wire \mem.mem[65][7] ;
 wire \mem.mem[66][0] ;
 wire \mem.mem[66][1] ;
 wire \mem.mem[66][2] ;
 wire \mem.mem[66][3] ;
 wire \mem.mem[66][4] ;
 wire \mem.mem[66][5] ;
 wire \mem.mem[66][6] ;
 wire \mem.mem[66][7] ;
 wire \mem.mem[67][0] ;
 wire \mem.mem[67][1] ;
 wire \mem.mem[67][2] ;
 wire \mem.mem[67][3] ;
 wire \mem.mem[67][4] ;
 wire \mem.mem[67][5] ;
 wire \mem.mem[67][6] ;
 wire \mem.mem[67][7] ;
 wire \mem.mem[68][0] ;
 wire \mem.mem[68][1] ;
 wire \mem.mem[68][2] ;
 wire \mem.mem[68][3] ;
 wire \mem.mem[68][4] ;
 wire \mem.mem[68][5] ;
 wire \mem.mem[68][6] ;
 wire \mem.mem[68][7] ;
 wire \mem.mem[69][0] ;
 wire \mem.mem[69][1] ;
 wire \mem.mem[69][2] ;
 wire \mem.mem[69][3] ;
 wire \mem.mem[69][4] ;
 wire \mem.mem[69][5] ;
 wire \mem.mem[69][6] ;
 wire \mem.mem[69][7] ;
 wire \mem.mem[6][0] ;
 wire \mem.mem[6][1] ;
 wire \mem.mem[6][2] ;
 wire \mem.mem[6][3] ;
 wire \mem.mem[6][4] ;
 wire \mem.mem[6][5] ;
 wire \mem.mem[6][6] ;
 wire \mem.mem[6][7] ;
 wire \mem.mem[70][0] ;
 wire \mem.mem[70][1] ;
 wire \mem.mem[70][2] ;
 wire \mem.mem[70][3] ;
 wire \mem.mem[70][4] ;
 wire \mem.mem[70][5] ;
 wire \mem.mem[70][6] ;
 wire \mem.mem[70][7] ;
 wire \mem.mem[71][0] ;
 wire \mem.mem[71][1] ;
 wire \mem.mem[71][2] ;
 wire \mem.mem[71][3] ;
 wire \mem.mem[71][4] ;
 wire \mem.mem[71][5] ;
 wire \mem.mem[71][6] ;
 wire \mem.mem[71][7] ;
 wire \mem.mem[72][0] ;
 wire \mem.mem[72][1] ;
 wire \mem.mem[72][2] ;
 wire \mem.mem[72][3] ;
 wire \mem.mem[72][4] ;
 wire \mem.mem[72][5] ;
 wire \mem.mem[72][6] ;
 wire \mem.mem[72][7] ;
 wire \mem.mem[73][0] ;
 wire \mem.mem[73][1] ;
 wire \mem.mem[73][2] ;
 wire \mem.mem[73][3] ;
 wire \mem.mem[73][4] ;
 wire \mem.mem[73][5] ;
 wire \mem.mem[73][6] ;
 wire \mem.mem[73][7] ;
 wire \mem.mem[74][0] ;
 wire \mem.mem[74][1] ;
 wire \mem.mem[74][2] ;
 wire \mem.mem[74][3] ;
 wire \mem.mem[74][4] ;
 wire \mem.mem[74][5] ;
 wire \mem.mem[74][6] ;
 wire \mem.mem[74][7] ;
 wire \mem.mem[75][0] ;
 wire \mem.mem[75][1] ;
 wire \mem.mem[75][2] ;
 wire \mem.mem[75][3] ;
 wire \mem.mem[75][4] ;
 wire \mem.mem[75][5] ;
 wire \mem.mem[75][6] ;
 wire \mem.mem[75][7] ;
 wire \mem.mem[76][0] ;
 wire \mem.mem[76][1] ;
 wire \mem.mem[76][2] ;
 wire \mem.mem[76][3] ;
 wire \mem.mem[76][4] ;
 wire \mem.mem[76][5] ;
 wire \mem.mem[76][6] ;
 wire \mem.mem[76][7] ;
 wire \mem.mem[77][0] ;
 wire \mem.mem[77][1] ;
 wire \mem.mem[77][2] ;
 wire \mem.mem[77][3] ;
 wire \mem.mem[77][4] ;
 wire \mem.mem[77][5] ;
 wire \mem.mem[77][6] ;
 wire \mem.mem[77][7] ;
 wire \mem.mem[78][0] ;
 wire \mem.mem[78][1] ;
 wire \mem.mem[78][2] ;
 wire \mem.mem[78][3] ;
 wire \mem.mem[78][4] ;
 wire \mem.mem[78][5] ;
 wire \mem.mem[78][6] ;
 wire \mem.mem[78][7] ;
 wire \mem.mem[79][0] ;
 wire \mem.mem[79][1] ;
 wire \mem.mem[79][2] ;
 wire \mem.mem[79][3] ;
 wire \mem.mem[79][4] ;
 wire \mem.mem[79][5] ;
 wire \mem.mem[79][6] ;
 wire \mem.mem[79][7] ;
 wire \mem.mem[7][0] ;
 wire \mem.mem[7][1] ;
 wire \mem.mem[7][2] ;
 wire \mem.mem[7][3] ;
 wire \mem.mem[7][4] ;
 wire \mem.mem[7][5] ;
 wire \mem.mem[7][6] ;
 wire \mem.mem[7][7] ;
 wire \mem.mem[80][0] ;
 wire \mem.mem[80][1] ;
 wire \mem.mem[80][2] ;
 wire \mem.mem[80][3] ;
 wire \mem.mem[80][4] ;
 wire \mem.mem[80][5] ;
 wire \mem.mem[80][6] ;
 wire \mem.mem[80][7] ;
 wire \mem.mem[81][0] ;
 wire \mem.mem[81][1] ;
 wire \mem.mem[81][2] ;
 wire \mem.mem[81][3] ;
 wire \mem.mem[81][4] ;
 wire \mem.mem[81][5] ;
 wire \mem.mem[81][6] ;
 wire \mem.mem[81][7] ;
 wire \mem.mem[82][0] ;
 wire \mem.mem[82][1] ;
 wire \mem.mem[82][2] ;
 wire \mem.mem[82][3] ;
 wire \mem.mem[82][4] ;
 wire \mem.mem[82][5] ;
 wire \mem.mem[82][6] ;
 wire \mem.mem[82][7] ;
 wire \mem.mem[83][0] ;
 wire \mem.mem[83][1] ;
 wire \mem.mem[83][2] ;
 wire \mem.mem[83][3] ;
 wire \mem.mem[83][4] ;
 wire \mem.mem[83][5] ;
 wire \mem.mem[83][6] ;
 wire \mem.mem[83][7] ;
 wire \mem.mem[84][0] ;
 wire \mem.mem[84][1] ;
 wire \mem.mem[84][2] ;
 wire \mem.mem[84][3] ;
 wire \mem.mem[84][4] ;
 wire \mem.mem[84][5] ;
 wire \mem.mem[84][6] ;
 wire \mem.mem[84][7] ;
 wire \mem.mem[85][0] ;
 wire \mem.mem[85][1] ;
 wire \mem.mem[85][2] ;
 wire \mem.mem[85][3] ;
 wire \mem.mem[85][4] ;
 wire \mem.mem[85][5] ;
 wire \mem.mem[85][6] ;
 wire \mem.mem[85][7] ;
 wire \mem.mem[86][0] ;
 wire \mem.mem[86][1] ;
 wire \mem.mem[86][2] ;
 wire \mem.mem[86][3] ;
 wire \mem.mem[86][4] ;
 wire \mem.mem[86][5] ;
 wire \mem.mem[86][6] ;
 wire \mem.mem[86][7] ;
 wire \mem.mem[87][0] ;
 wire \mem.mem[87][1] ;
 wire \mem.mem[87][2] ;
 wire \mem.mem[87][3] ;
 wire \mem.mem[87][4] ;
 wire \mem.mem[87][5] ;
 wire \mem.mem[87][6] ;
 wire \mem.mem[87][7] ;
 wire \mem.mem[88][0] ;
 wire \mem.mem[88][1] ;
 wire \mem.mem[88][2] ;
 wire \mem.mem[88][3] ;
 wire \mem.mem[88][4] ;
 wire \mem.mem[88][5] ;
 wire \mem.mem[88][6] ;
 wire \mem.mem[88][7] ;
 wire \mem.mem[89][0] ;
 wire \mem.mem[89][1] ;
 wire \mem.mem[89][2] ;
 wire \mem.mem[89][3] ;
 wire \mem.mem[89][4] ;
 wire \mem.mem[89][5] ;
 wire \mem.mem[89][6] ;
 wire \mem.mem[89][7] ;
 wire \mem.mem[8][0] ;
 wire \mem.mem[8][1] ;
 wire \mem.mem[8][2] ;
 wire \mem.mem[8][3] ;
 wire \mem.mem[8][4] ;
 wire \mem.mem[8][5] ;
 wire \mem.mem[8][6] ;
 wire \mem.mem[8][7] ;
 wire \mem.mem[90][0] ;
 wire \mem.mem[90][1] ;
 wire \mem.mem[90][2] ;
 wire \mem.mem[90][3] ;
 wire \mem.mem[90][4] ;
 wire \mem.mem[90][5] ;
 wire \mem.mem[90][6] ;
 wire \mem.mem[90][7] ;
 wire \mem.mem[91][0] ;
 wire \mem.mem[91][1] ;
 wire \mem.mem[91][2] ;
 wire \mem.mem[91][3] ;
 wire \mem.mem[91][4] ;
 wire \mem.mem[91][5] ;
 wire \mem.mem[91][6] ;
 wire \mem.mem[91][7] ;
 wire \mem.mem[92][0] ;
 wire \mem.mem[92][1] ;
 wire \mem.mem[92][2] ;
 wire \mem.mem[92][3] ;
 wire \mem.mem[92][4] ;
 wire \mem.mem[92][5] ;
 wire \mem.mem[92][6] ;
 wire \mem.mem[92][7] ;
 wire \mem.mem[93][0] ;
 wire \mem.mem[93][1] ;
 wire \mem.mem[93][2] ;
 wire \mem.mem[93][3] ;
 wire \mem.mem[93][4] ;
 wire \mem.mem[93][5] ;
 wire \mem.mem[93][6] ;
 wire \mem.mem[93][7] ;
 wire \mem.mem[94][0] ;
 wire \mem.mem[94][1] ;
 wire \mem.mem[94][2] ;
 wire \mem.mem[94][3] ;
 wire \mem.mem[94][4] ;
 wire \mem.mem[94][5] ;
 wire \mem.mem[94][6] ;
 wire \mem.mem[94][7] ;
 wire \mem.mem[95][0] ;
 wire \mem.mem[95][1] ;
 wire \mem.mem[95][2] ;
 wire \mem.mem[95][3] ;
 wire \mem.mem[95][4] ;
 wire \mem.mem[95][5] ;
 wire \mem.mem[95][6] ;
 wire \mem.mem[95][7] ;
 wire \mem.mem[96][0] ;
 wire \mem.mem[96][1] ;
 wire \mem.mem[96][2] ;
 wire \mem.mem[96][3] ;
 wire \mem.mem[96][4] ;
 wire \mem.mem[96][5] ;
 wire \mem.mem[96][6] ;
 wire \mem.mem[96][7] ;
 wire \mem.mem[97][0] ;
 wire \mem.mem[97][1] ;
 wire \mem.mem[97][2] ;
 wire \mem.mem[97][3] ;
 wire \mem.mem[97][4] ;
 wire \mem.mem[97][5] ;
 wire \mem.mem[97][6] ;
 wire \mem.mem[97][7] ;
 wire \mem.mem[98][0] ;
 wire \mem.mem[98][1] ;
 wire \mem.mem[98][2] ;
 wire \mem.mem[98][3] ;
 wire \mem.mem[98][4] ;
 wire \mem.mem[98][5] ;
 wire \mem.mem[98][6] ;
 wire \mem.mem[98][7] ;
 wire \mem.mem[99][0] ;
 wire \mem.mem[99][1] ;
 wire \mem.mem[99][2] ;
 wire \mem.mem[99][3] ;
 wire \mem.mem[99][4] ;
 wire \mem.mem[99][5] ;
 wire \mem.mem[99][6] ;
 wire \mem.mem[99][7] ;
 wire \mem.mem[9][0] ;
 wire \mem.mem[9][1] ;
 wire \mem.mem[9][2] ;
 wire \mem.mem[9][3] ;
 wire \mem.mem[9][4] ;
 wire \mem.mem[9][5] ;
 wire \mem.mem[9][6] ;
 wire \mem.mem[9][7] ;
 wire \mem.out_strobe ;
 wire \mem.wr_en ;
 wire \mem_A[0] ;
 wire \mem_A[1] ;
 wire \mem_A[2] ;
 wire \mem_A[3] ;
 wire \mem_A[4] ;
 wire \mem_A[5] ;
 wire \mem_A[6] ;
 wire \mem_A[7] ;
 wire prev_run;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \state[5] ;
 wire \state[6] ;
 wire net13;
 wire net2131;
 wire net14;
 wire net15;
 wire clknet_leaf_0_clk;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net5488;
 wire net5489;
 wire net5490;
 wire net5491;
 wire net5492;
 wire net5493;
 wire net5494;
 wire net5495;
 wire net5496;
 wire net5497;
 wire net5498;
 wire net5499;
 wire net5500;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5507;
 wire net5508;
 wire net5509;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5514;
 wire net5515;
 wire net5516;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5523;
 wire net5524;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net5530;
 wire net5531;
 wire net5532;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net5540;
 wire net5541;
 wire net5542;
 wire net5543;
 wire net5544;
 wire net5545;
 wire net5546;
 wire net5547;
 wire net5548;
 wire net5549;
 wire net5550;
 wire net5551;
 wire net5552;
 wire net5553;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5574;
 wire net5575;
 wire net5576;
 wire net5577;
 wire net5578;
 wire net5579;
 wire net5580;
 wire net5581;
 wire net5582;
 wire net5583;
 wire net5584;
 wire net5585;
 wire net5586;
 wire net5587;
 wire net5588;
 wire net5589;
 wire net5590;
 wire net5591;
 wire net5592;
 wire net5593;
 wire net5594;
 wire net5595;
 wire net5596;
 wire net5597;
 wire net5598;
 wire net5599;
 wire net5600;
 wire net5601;
 wire net5602;
 wire net5603;
 wire net5604;
 wire net5605;
 wire net5606;
 wire net5607;
 wire net5608;
 wire net5609;
 wire net5610;
 wire net5611;
 wire net5612;
 wire net5613;
 wire net5614;
 wire net5615;
 wire net5616;
 wire net5617;
 wire net5618;
 wire net5619;
 wire net5620;
 wire net5621;
 wire net5622;
 wire net5623;
 wire net5624;
 wire net5625;
 wire net5626;
 wire net5627;
 wire net5628;
 wire net5629;
 wire net5630;
 wire net5631;
 wire net5632;
 wire net5633;
 wire net5634;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5638;
 wire net5639;
 wire net5640;
 wire net5641;
 wire net5642;
 wire net5643;
 wire net5644;
 wire net5645;
 wire net5646;
 wire net5647;
 wire net5648;
 wire net5649;
 wire net5650;
 wire net5651;
 wire net5652;
 wire net5653;
 wire net5654;
 wire net5655;
 wire net5656;
 wire net5657;
 wire net5658;
 wire net5659;
 wire net5660;
 wire net5661;
 wire net5662;
 wire net5663;
 wire net5664;
 wire net5665;
 wire net5666;
 wire net5667;
 wire net5668;
 wire net5669;
 wire net5670;
 wire net5671;
 wire net5672;
 wire net5673;
 wire net5674;
 wire net5675;
 wire net5676;
 wire net5677;
 wire net5678;
 wire net5679;
 wire net5680;
 wire net5681;
 wire net5682;
 wire net5683;
 wire net5684;
 wire net5685;
 wire net5686;
 wire net5687;
 wire net5688;
 wire net5689;
 wire net5690;
 wire net5691;
 wire net5692;
 wire net5693;
 wire net5694;
 wire net5695;
 wire net5696;
 wire net5697;
 wire net5698;
 wire net5699;
 wire net5700;
 wire net5701;
 wire net5702;
 wire net5703;
 wire net5704;
 wire net5705;
 wire net5706;
 wire net5707;
 wire net5708;
 wire net5709;
 wire net5710;
 wire net5711;
 wire net5712;
 wire net5713;
 wire net5714;
 wire net5715;
 wire net5716;
 wire net5717;
 wire net5718;
 wire net5719;
 wire net5720;
 wire net5721;
 wire net5722;
 wire net5723;
 wire net5724;
 wire net5725;
 wire net5726;
 wire net5727;
 wire net5728;
 wire net5729;
 wire net5730;
 wire net5731;
 wire net5732;
 wire net5733;
 wire net5734;
 wire net5735;
 wire net5736;
 wire net5737;
 wire net5738;
 wire net5739;
 wire net5740;
 wire net5741;
 wire net5742;
 wire net5743;
 wire net5744;
 wire net5745;
 wire net5746;
 wire net5747;
 wire net5748;
 wire net5749;
 wire net5750;
 wire net5751;
 wire net5752;
 wire net5753;
 wire net5754;
 wire net5755;
 wire net5756;
 wire net5757;
 wire net5758;
 wire net5759;
 wire net5760;
 wire net5761;
 wire net5762;
 wire net5763;
 wire net5764;
 wire net5765;
 wire net5766;
 wire net5767;
 wire net5768;
 wire net5769;
 wire net5770;
 wire net5771;
 wire net5772;
 wire net5773;
 wire net5774;
 wire net5775;
 wire net5776;
 wire net5777;
 wire net5778;
 wire net5779;
 wire net5780;
 wire net5781;
 wire net5782;
 wire net5783;
 wire net5784;
 wire net5785;
 wire net5786;
 wire net5787;
 wire net5788;
 wire net5789;
 wire net5790;
 wire net5791;
 wire net5792;
 wire net5793;
 wire net5794;
 wire net5795;
 wire net5796;
 wire net5797;
 wire net5798;
 wire net5799;
 wire net5800;
 wire net5801;
 wire net5802;
 wire net5803;
 wire net5804;
 wire net5805;
 wire net5806;
 wire net5807;
 wire net5808;
 wire net5809;
 wire net5810;
 wire net5811;
 wire net5812;
 wire net5813;
 wire net5814;
 wire net5815;
 wire net5816;
 wire net5817;
 wire net5818;
 wire net5819;
 wire net5820;
 wire net5821;
 wire net5822;
 wire net5823;
 wire net5824;
 wire net5825;
 wire net5826;
 wire net5827;
 wire net5828;
 wire net5829;
 wire net5830;
 wire net5831;
 wire net5832;
 wire net5833;
 wire net5834;
 wire net5835;
 wire net5836;
 wire net5837;
 wire net5838;
 wire net5839;
 wire net5840;
 wire net5841;
 wire net5842;
 wire net5843;
 wire net5844;
 wire net5845;
 wire net5846;
 wire net5847;
 wire net5848;
 wire net5849;
 wire net5850;
 wire net5851;
 wire net5852;
 wire net5853;
 wire net5854;
 wire net5855;
 wire net5856;
 wire net5857;
 wire net5858;
 wire net5859;
 wire net5860;
 wire net5861;
 wire net5862;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5866;
 wire net5867;
 wire net5868;
 wire net5869;
 wire net5870;
 wire net5871;
 wire net5872;
 wire net5873;
 wire net5874;
 wire net5875;
 wire net5876;
 wire net5877;
 wire net5878;
 wire net5879;
 wire net5880;
 wire net5881;
 wire net5882;
 wire net5883;
 wire net5884;
 wire net5885;
 wire net5886;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net5890;
 wire net5891;
 wire net5892;
 wire net5893;
 wire net5894;
 wire net5895;
 wire net5896;
 wire net5897;
 wire net5898;
 wire net5899;
 wire net5900;
 wire net5901;
 wire net5902;
 wire net5903;
 wire net5904;
 wire net5905;
 wire net5906;
 wire net5907;
 wire net5908;
 wire net5909;
 wire net5910;
 wire net5911;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5915;
 wire net5916;
 wire net5917;
 wire net5918;
 wire net5919;
 wire net5920;
 wire net5921;
 wire net5922;
 wire net5923;
 wire net5924;
 wire net5925;
 wire net5926;
 wire net5927;
 wire net5928;
 wire net5929;
 wire net5930;
 wire net5931;
 wire net5932;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net5940;
 wire net5941;
 wire net5942;
 wire net5943;
 wire net5944;
 wire net5945;
 wire net5946;
 wire net5947;
 wire net5948;
 wire net5949;
 wire net5950;
 wire net5951;
 wire net5952;
 wire net5953;
 wire net5954;
 wire net5955;
 wire net5956;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net5960;
 wire net5961;
 wire net5962;
 wire net5963;
 wire net5964;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5969;
 wire net5970;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5989;
 wire net5990;
 wire net5991;
 wire net5992;
 wire net5993;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6000;
 wire net6001;
 wire net6002;
 wire net6003;
 wire net6004;
 wire net6005;
 wire net6006;
 wire net6007;
 wire net6008;
 wire net6009;
 wire net6010;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6016;
 wire net6017;
 wire net6018;
 wire net6019;
 wire net6020;
 wire net6021;
 wire net6022;
 wire net6023;
 wire net6024;
 wire net6025;
 wire net6026;
 wire net6027;
 wire net6028;
 wire net6029;
 wire net6030;
 wire net6031;
 wire net6032;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6038;
 wire net6039;
 wire net6040;
 wire net6041;
 wire net6042;
 wire net6043;
 wire net6044;
 wire net6045;
 wire net6046;
 wire net6047;
 wire net6048;
 wire net6049;
 wire net6050;
 wire net6051;
 wire net6052;
 wire net6053;
 wire net6054;
 wire net6055;
 wire net6056;
 wire net6057;
 wire net6058;
 wire net6059;
 wire net6060;
 wire net6061;
 wire net6062;
 wire net6063;
 wire net6064;
 wire net6065;
 wire net6066;
 wire net6067;
 wire net6068;
 wire net6069;
 wire net6070;
 wire net6071;
 wire net6072;
 wire net6073;
 wire net6074;
 wire net6075;
 wire net6076;
 wire net6077;
 wire net6078;
 wire net6079;
 wire net6080;
 wire net6081;
 wire net6082;
 wire net6083;
 wire net6084;
 wire net6085;
 wire net6086;
 wire net6087;
 wire net6088;
 wire net6089;
 wire net6090;
 wire net6091;
 wire net6092;
 wire net6093;
 wire net6094;
 wire net6095;
 wire net6096;
 wire net6097;
 wire net6098;
 wire net6099;
 wire net6100;
 wire net6101;
 wire net6102;
 wire net6103;
 wire net6104;
 wire net6105;
 wire net6106;
 wire net6107;
 wire net6108;
 wire net6109;
 wire net6110;
 wire net6111;
 wire net6112;
 wire net6113;
 wire net6114;
 wire net6115;
 wire net6116;
 wire net6117;
 wire net6118;
 wire net6119;
 wire net6120;
 wire net6121;
 wire net6122;
 wire net6123;
 wire net6124;
 wire net6125;
 wire net6126;
 wire net6127;
 wire net6128;
 wire net6129;
 wire net6130;
 wire net6131;
 wire net6132;
 wire net6133;
 wire net6134;
 wire net6135;
 wire net6136;
 wire net6137;
 wire net6138;
 wire net6139;
 wire net6140;
 wire net6141;
 wire net6142;
 wire net6143;
 wire net6144;
 wire net6145;
 wire net6146;
 wire net6147;
 wire net6148;
 wire net6149;
 wire net6150;
 wire net6151;
 wire net6152;
 wire net6153;
 wire net6154;
 wire net6155;
 wire net6156;
 wire net6157;
 wire net6158;
 wire net6159;
 wire net6160;
 wire net6161;
 wire net6162;
 wire net6163;
 wire net6164;
 wire net6165;
 wire net6166;
 wire net6167;
 wire net6168;
 wire net6169;
 wire net6170;
 wire net6171;
 wire net6172;
 wire net6173;
 wire net6174;
 wire net6175;
 wire net6176;
 wire net6177;
 wire net6178;
 wire net6179;
 wire net6180;
 wire net6181;
 wire net6182;
 wire net6183;
 wire net6184;
 wire net6185;
 wire net6186;
 wire net6187;
 wire net6188;
 wire net6189;
 wire net6190;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0_0_clk;
 wire clknet_6_1_0_clk;
 wire clknet_6_2_0_clk;
 wire clknet_6_3_0_clk;
 wire clknet_6_4_0_clk;
 wire clknet_6_5_0_clk;
 wire clknet_6_6_0_clk;
 wire clknet_6_7_0_clk;
 wire clknet_6_8_0_clk;
 wire clknet_6_9_0_clk;
 wire clknet_6_10_0_clk;
 wire clknet_6_11_0_clk;
 wire clknet_6_12_0_clk;
 wire clknet_6_13_0_clk;
 wire clknet_6_14_0_clk;
 wire clknet_6_15_0_clk;
 wire clknet_6_16_0_clk;
 wire clknet_6_17_0_clk;
 wire clknet_6_18_0_clk;
 wire clknet_6_19_0_clk;
 wire clknet_6_20_0_clk;
 wire clknet_6_21_0_clk;
 wire clknet_6_22_0_clk;
 wire clknet_6_23_0_clk;
 wire clknet_6_24_0_clk;
 wire clknet_6_25_0_clk;
 wire clknet_6_26_0_clk;
 wire clknet_6_27_0_clk;
 wire clknet_6_28_0_clk;
 wire clknet_6_29_0_clk;
 wire clknet_6_30_0_clk;
 wire clknet_6_31_0_clk;
 wire clknet_6_32_0_clk;
 wire clknet_6_33_0_clk;
 wire clknet_6_34_0_clk;
 wire clknet_6_35_0_clk;
 wire clknet_6_36_0_clk;
 wire clknet_6_37_0_clk;
 wire clknet_6_38_0_clk;
 wire clknet_6_39_0_clk;
 wire clknet_6_40_0_clk;
 wire clknet_6_41_0_clk;
 wire clknet_6_42_0_clk;
 wire clknet_6_43_0_clk;
 wire clknet_6_44_0_clk;
 wire clknet_6_45_0_clk;
 wire clknet_6_46_0_clk;
 wire clknet_6_47_0_clk;
 wire clknet_6_48_0_clk;
 wire clknet_6_49_0_clk;
 wire clknet_6_50_0_clk;
 wire clknet_6_51_0_clk;
 wire clknet_6_52_0_clk;
 wire clknet_6_53_0_clk;
 wire clknet_6_54_0_clk;
 wire clknet_6_55_0_clk;
 wire clknet_6_56_0_clk;
 wire clknet_6_57_0_clk;
 wire clknet_6_58_0_clk;
 wire clknet_6_59_0_clk;
 wire clknet_6_60_0_clk;
 wire clknet_6_61_0_clk;
 wire clknet_6_62_0_clk;
 wire clknet_6_63_0_clk;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;

 sg13g2_inv_1 _11302_ (.Y(_02820_),
    .A(\mem.data_in[7] ));
 sg13g2_inv_1 _11303_ (.Y(_02821_),
    .A(\mem.data_in[6] ));
 sg13g2_inv_1 _11304_ (.Y(_02822_),
    .A(\mem.data_in[5] ));
 sg13g2_inv_4 _11305_ (.A(\mem.data_in[4] ),
    .Y(_02823_));
 sg13g2_inv_1 _11306_ (.Y(_02824_),
    .A(\mem.data_in[3] ));
 sg13g2_inv_1 _11307_ (.Y(_02825_),
    .A(\mem.data_in[2] ));
 sg13g2_inv_1 _11308_ (.Y(_02826_),
    .A(\mem.data_in[1] ));
 sg13g2_inv_1 _11309_ (.Y(_02827_),
    .A(\mem.data_in[0] ));
 sg13g2_inv_1 _11310_ (.Y(_02828_),
    .A(\mem_A[0] ));
 sg13g2_inv_2 _11311_ (.Y(_02829_),
    .A(net4253));
 sg13g2_inv_2 _11312_ (.Y(_02830_),
    .A(\mem.addr[2] ));
 sg13g2_inv_1 _11313_ (.Y(_02831_),
    .A(net4234));
 sg13g2_inv_1 _11314_ (.Y(_02832_),
    .A(net4219));
 sg13g2_inv_4 _11315_ (.A(net6018),
    .Y(_02833_));
 sg13g2_inv_1 _11316_ (.Y(_02834_),
    .A(net5918));
 sg13g2_inv_1 _11317_ (.Y(_02835_),
    .A(net5857));
 sg13g2_inv_2 _11318_ (.Y(_02836_),
    .A(net5833));
 sg13g2_inv_4 _11319_ (.A(net5816),
    .Y(_02837_));
 sg13g2_inv_1 _11320_ (.Y(_02838_),
    .A(net5810));
 sg13g2_inv_4 _11321_ (.A(net5808),
    .Y(_02839_));
 sg13g2_inv_4 _11322_ (.A(_00007_),
    .Y(_02840_));
 sg13g2_inv_2 _11323_ (.Y(_02841_),
    .A(net3));
 sg13g2_inv_1 _11324_ (.Y(_02842_),
    .A(net4239));
 sg13g2_inv_1 _11325_ (.Y(_02843_),
    .A(net4));
 sg13g2_inv_1 _11326_ (.Y(_02844_),
    .A(\mem.mem[4][2] ));
 sg13g2_inv_1 _11327_ (.Y(_02845_),
    .A(\mem.mem[22][2] ));
 sg13g2_inv_1 _11328_ (.Y(_02846_),
    .A(\mem.mem[36][2] ));
 sg13g2_inv_1 _11329_ (.Y(_02847_),
    .A(net3712));
 sg13g2_inv_1 _11330_ (.Y(_02848_),
    .A(\mem.mem[100][2] ));
 sg13g2_inv_1 _11331_ (.Y(_02849_),
    .A(\mem.mem[126][2] ));
 sg13g2_inv_1 _11332_ (.Y(_02850_),
    .A(\mem.mem[221][2] ));
 sg13g2_inv_1 _11333_ (.Y(_02851_),
    .A(\mem.mem[237][2] ));
 sg13g2_inv_1 _11334_ (.Y(_02852_),
    .A(net5));
 sg13g2_inv_1 _11335_ (.Y(_02853_),
    .A(\mem.mem[36][3] ));
 sg13g2_inv_1 _11336_ (.Y(_02854_),
    .A(\mem.mem[78][3] ));
 sg13g2_inv_1 _11337_ (.Y(_02855_),
    .A(\mem.mem[94][3] ));
 sg13g2_inv_1 _11338_ (.Y(_02856_),
    .A(net3904));
 sg13g2_inv_1 _11339_ (.Y(_02857_),
    .A(net6));
 sg13g2_inv_1 _11340_ (.Y(_02858_),
    .A(\mem.mem[20][4] ));
 sg13g2_inv_1 _11341_ (.Y(_02859_),
    .A(\mem.mem[36][4] ));
 sg13g2_inv_1 _11342_ (.Y(_02860_),
    .A(net3969));
 sg13g2_inv_1 _11343_ (.Y(_02861_),
    .A(\mem.mem[110][4] ));
 sg13g2_inv_1 _11344_ (.Y(_02862_),
    .A(\mem.mem[116][4] ));
 sg13g2_inv_1 _11345_ (.Y(_02863_),
    .A(\mem.mem[204][4] ));
 sg13g2_inv_1 _11346_ (.Y(_02864_),
    .A(\mem.mem[222][4] ));
 sg13g2_inv_1 _11347_ (.Y(_02865_),
    .A(net7));
 sg13g2_inv_1 _11348_ (.Y(_02866_),
    .A(\mem.mem[14][5] ));
 sg13g2_inv_1 _11349_ (.Y(_02867_),
    .A(\mem.mem[110][5] ));
 sg13g2_inv_1 _11350_ (.Y(_02868_),
    .A(net8));
 sg13g2_inv_1 _11351_ (.Y(_02869_),
    .A(\mem.mem[4][6] ));
 sg13g2_inv_1 _11352_ (.Y(_02870_),
    .A(\mem.mem[14][6] ));
 sg13g2_inv_1 _11353_ (.Y(_02871_),
    .A(net4146));
 sg13g2_inv_1 _11354_ (.Y(_02872_),
    .A(\mem.mem[102][6] ));
 sg13g2_inv_1 _11355_ (.Y(_02873_),
    .A(\mem.mem[116][6] ));
 sg13g2_inv_1 _11356_ (.Y(_02874_),
    .A(\mem.mem[222][6] ));
 sg13g2_inv_1 _11357_ (.Y(_02875_),
    .A(net9));
 sg13g2_inv_1 _11358_ (.Y(_02876_),
    .A(\mem.mem[22][7] ));
 sg13g2_inv_1 _11359_ (.Y(_02877_),
    .A(net3893));
 sg13g2_inv_1 _11360_ (.Y(_02878_),
    .A(\mem.mem[126][7] ));
 sg13g2_inv_1 _11361_ (.Y(_02879_),
    .A(net3385));
 sg13g2_inv_2 _11362_ (.Y(_02880_),
    .A(net2));
 sg13g2_inv_2 _11363_ (.Y(_02881_),
    .A(net6180));
 sg13g2_inv_1 _11364_ (.Y(_02882_),
    .A(net5793));
 sg13g2_inv_1 _11365_ (.Y(_02883_),
    .A(net6182));
 sg13g2_inv_1 _11366_ (.Y(_02884_),
    .A(halted));
 sg13g2_inv_1 _11367_ (.Y(_02885_),
    .A(net3335));
 sg13g2_inv_1 _11368_ (.Y(_02886_),
    .A(net3401));
 sg13g2_inv_1 _11369_ (.Y(_02887_),
    .A(net3091));
 sg13g2_inv_1 _11370_ (.Y(_02888_),
    .A(\mem.mem[174][0] ));
 sg13g2_inv_1 _11371_ (.Y(_02889_),
    .A(net3505));
 sg13g2_inv_1 _11372_ (.Y(_02890_),
    .A(\mem.mem[142][1] ));
 sg13g2_and2_1 _11373_ (.A(net5787),
    .B(net6185),
    .X(_00009_));
 sg13g2_and2_1 _11374_ (.A(net5797),
    .B(net6182),
    .X(_00011_));
 sg13g2_and2_1 _11375_ (.A(net5786),
    .B(net6182),
    .X(_00008_));
 sg13g2_nor2_1 _11376_ (.A(net5261),
    .B(net6176),
    .Y(_00010_));
 sg13g2_and2_1 _11377_ (.A(net5794),
    .B(net6183),
    .X(_00012_));
 sg13g2_or2_1 _11378_ (.X(_02891_),
    .B(\PC[0] ),
    .A(\PC[1] ));
 sg13g2_nand3_1 _11379_ (.B(\PC[2] ),
    .C(_02891_),
    .A(\PC[3] ),
    .Y(_02892_));
 sg13g2_nand2_1 _11380_ (.Y(_02893_),
    .A(\PC[5] ),
    .B(\PC[4] ));
 sg13g2_nor2_1 _11381_ (.A(_02892_),
    .B(_02893_),
    .Y(_02894_));
 sg13g2_nor3_1 _11382_ (.A(_00017_),
    .B(_02892_),
    .C(_02893_),
    .Y(_02895_));
 sg13g2_nor3_1 _11383_ (.A(\mem.data_in[2] ),
    .B(\mem.data_in[1] ),
    .C(\mem.data_in[0] ),
    .Y(_02896_));
 sg13g2_nor4_1 _11384_ (.A(\mem.data_in[6] ),
    .B(\mem.data_in[5] ),
    .C(\mem.data_in[4] ),
    .D(\mem.data_in[3] ),
    .Y(_02897_));
 sg13g2_a21oi_1 _11385_ (.A1(_02896_),
    .A2(_02897_),
    .Y(_02898_),
    .B1(\mem.data_in[7] ));
 sg13g2_xnor2_1 _11386_ (.Y(_02899_),
    .A(_02831_),
    .B(_02895_));
 sg13g2_nor2_1 _11387_ (.A(_00020_),
    .B(net5256),
    .Y(_02900_));
 sg13g2_a21oi_1 _11388_ (.A1(net5256),
    .A2(_02899_),
    .Y(_02901_),
    .B1(_02900_));
 sg13g2_nand2_1 _11389_ (.Y(_02902_),
    .A(_00018_),
    .B(_02892_));
 sg13g2_or2_1 _11390_ (.X(_02903_),
    .B(_02892_),
    .A(_00018_));
 sg13g2_nand3_1 _11391_ (.B(_02902_),
    .C(_02903_),
    .A(net5256),
    .Y(_02904_));
 sg13g2_o21ai_1 _11392_ (.B1(_02904_),
    .Y(_02905_),
    .A1(_00023_),
    .A2(net5256));
 sg13g2_mux2_1 _11393_ (.A0(net4185),
    .A1(_00019_),
    .S(net5255),
    .X(_02906_));
 sg13g2_nor2_1 _11394_ (.A(_00026_),
    .B(net5255),
    .Y(_02907_));
 sg13g2_nand2_1 _11395_ (.Y(_02908_),
    .A(\PC[1] ),
    .B(\PC[0] ));
 sg13g2_nand2_1 _11396_ (.Y(_02909_),
    .A(_02891_),
    .B(_02908_));
 sg13g2_a21oi_1 _11397_ (.A1(net5255),
    .A2(_02909_),
    .Y(_02910_),
    .B1(_02907_));
 sg13g2_inv_1 _11398_ (.Y(_02911_),
    .A(_02910_));
 sg13g2_nand2b_1 _11399_ (.Y(_02912_),
    .B(_02910_),
    .A_N(_02906_));
 sg13g2_a21o_1 _11400_ (.A2(_02891_),
    .A1(\PC[2] ),
    .B1(\PC[3] ),
    .X(_02913_));
 sg13g2_nand3_1 _11401_ (.B(net5255),
    .C(_02913_),
    .A(_02892_),
    .Y(_02914_));
 sg13g2_o21ai_1 _11402_ (.B1(_02914_),
    .Y(_02915_),
    .A1(_00024_),
    .A2(net5255));
 sg13g2_xor2_1 _11403_ (.B(_02891_),
    .A(\PC[2] ),
    .X(_02916_));
 sg13g2_nand2_1 _11404_ (.Y(_02917_),
    .A(net5255),
    .B(_02916_));
 sg13g2_o21ai_1 _11405_ (.B1(_02917_),
    .Y(_02918_),
    .A1(net4236),
    .A2(net5255));
 sg13g2_and4_1 _11406_ (.A(_02905_),
    .B(_02912_),
    .C(_02915_),
    .D(_02918_),
    .X(_02919_));
 sg13g2_xnor2_1 _11407_ (.Y(_02920_),
    .A(\PC[5] ),
    .B(_02903_));
 sg13g2_nand2_1 _11408_ (.Y(_02921_),
    .A(net5256),
    .B(_02920_));
 sg13g2_o21ai_1 _11409_ (.B1(_02921_),
    .Y(_02922_),
    .A1(_00022_),
    .A2(net5256));
 sg13g2_o21ai_1 _11410_ (.B1(_00017_),
    .Y(_02923_),
    .A1(_02892_),
    .A2(_02893_));
 sg13g2_nand3b_1 _11411_ (.B(net5256),
    .C(_02923_),
    .Y(_02924_),
    .A_N(_02895_));
 sg13g2_o21ai_1 _11412_ (.B1(_02924_),
    .Y(_02925_),
    .A1(_00021_),
    .A2(net5255));
 sg13g2_nand3_1 _11413_ (.B(_02922_),
    .C(_02925_),
    .A(_02919_),
    .Y(_02926_));
 sg13g2_o21ai_1 _11414_ (.B1(net10),
    .Y(_02927_),
    .A1(_02901_),
    .A2(_02926_));
 sg13g2_inv_1 _11415_ (.Y(_02928_),
    .A(_02927_));
 sg13g2_nand3_1 _11416_ (.B(\PC[6] ),
    .C(_02894_),
    .A(\PC[7] ),
    .Y(_02929_));
 sg13g2_nand3b_1 _11417_ (.B(_02929_),
    .C(net10),
    .Y(_02930_),
    .A_N(net4227));
 sg13g2_inv_1 _11418_ (.Y(_02931_),
    .A(_02930_));
 sg13g2_a22oi_1 _11419_ (.Y(_02932_),
    .B1(_02931_),
    .B2(net4216),
    .A2(_02928_),
    .A1(net5793));
 sg13g2_nor2_1 _11420_ (.A(net6176),
    .B(net4217),
    .Y(_00014_));
 sg13g2_a22oi_1 _11421_ (.Y(_02933_),
    .B1(_02930_),
    .B2(net4216),
    .A2(_02927_),
    .A1(net5792));
 sg13g2_nand2_1 _11422_ (.Y(_00013_),
    .A(net6190),
    .B(_02933_));
 sg13g2_nor2_2 _11423_ (.A(\mem.addr[1] ),
    .B(\mem.addr[0] ),
    .Y(_02934_));
 sg13g2_or2_2 _11424_ (.X(_02935_),
    .B(\mem.addr[0] ),
    .A(net5805));
 sg13g2_nor2_2 _11425_ (.A(_02829_),
    .B(\mem.addr[2] ),
    .Y(_02936_));
 sg13g2_nand2_2 _11426_ (.Y(_02937_),
    .A(\mem.addr[3] ),
    .B(_02830_));
 sg13g2_nor2_2 _11427_ (.A(_02935_),
    .B(_02937_),
    .Y(_02938_));
 sg13g2_nand2_2 _11428_ (.Y(_02939_),
    .A(_02934_),
    .B(_02936_));
 sg13g2_nand2_2 _11429_ (.Y(_02940_),
    .A(\mem.addr[7] ),
    .B(net5803));
 sg13g2_nand4_1 _11430_ (.B(net5802),
    .C(\mem.addr[5] ),
    .A(net5801),
    .Y(_02941_),
    .D(\mem.addr[4] ));
 sg13g2_nor2_2 _11431_ (.A(_02829_),
    .B(_02830_),
    .Y(_02942_));
 sg13g2_nand2_2 _11432_ (.Y(_02943_),
    .A(\mem.addr[3] ),
    .B(\mem.addr[2] ));
 sg13g2_nor3_2 _11433_ (.A(_02934_),
    .B(_02941_),
    .C(_02943_),
    .Y(_02944_));
 sg13g2_nand3b_1 _11434_ (.B(_02942_),
    .C(_02935_),
    .Y(_02945_),
    .A_N(_02941_));
 sg13g2_nor3_2 _11435_ (.A(net6177),
    .B(_00015_),
    .C(_02944_),
    .Y(_02946_));
 sg13g2_nand3b_1 _11436_ (.B(_02945_),
    .C(net6187),
    .Y(_02947_),
    .A_N(_00015_));
 sg13g2_nand3b_1 _11437_ (.B(net5804),
    .C(_02946_),
    .Y(_02948_),
    .A_N(\mem.addr[5] ));
 sg13g2_nor2b_2 _11438_ (.A(net5801),
    .B_N(net5802),
    .Y(_02949_));
 sg13g2_nand2b_1 _11439_ (.Y(_02950_),
    .B(net5802),
    .A_N(net5801));
 sg13g2_nor2_1 _11440_ (.A(net5229),
    .B(net5259),
    .Y(_02951_));
 sg13g2_nand2_1 _11441_ (.Y(_02952_),
    .A(net5244),
    .B(net5224));
 sg13g2_nand2_1 _11442_ (.Y(_02953_),
    .A(net3190),
    .B(net5160));
 sg13g2_o21ai_1 _11443_ (.B1(_02953_),
    .Y(_00027_),
    .A1(net5429),
    .A2(net5160));
 sg13g2_nand2_1 _11444_ (.Y(_02954_),
    .A(net2186),
    .B(net5161));
 sg13g2_o21ai_1 _11445_ (.B1(_02954_),
    .Y(_00028_),
    .A1(net5474),
    .A2(net5161));
 sg13g2_nand2_1 _11446_ (.Y(_02955_),
    .A(net2675),
    .B(net5161));
 sg13g2_o21ai_1 _11447_ (.B1(_02955_),
    .Y(_00029_),
    .A1(net5520),
    .A2(net5161));
 sg13g2_nand2_1 _11448_ (.Y(_02956_),
    .A(net3093),
    .B(net5161));
 sg13g2_o21ai_1 _11449_ (.B1(_02956_),
    .Y(_00030_),
    .A1(net5563),
    .A2(_02952_));
 sg13g2_nand2_1 _11450_ (.Y(_02957_),
    .A(net3068),
    .B(net5160));
 sg13g2_o21ai_1 _11451_ (.B1(_02957_),
    .Y(_00031_),
    .A1(net5610),
    .A2(net5160));
 sg13g2_nand2_1 _11452_ (.Y(_02958_),
    .A(net3248),
    .B(net5161));
 sg13g2_o21ai_1 _11453_ (.B1(_02958_),
    .Y(_00032_),
    .A1(net5656),
    .A2(net5161));
 sg13g2_nand2_1 _11454_ (.Y(_02959_),
    .A(net3647),
    .B(net5160));
 sg13g2_o21ai_1 _11455_ (.B1(_02959_),
    .Y(_00033_),
    .A1(net5701),
    .A2(net5160));
 sg13g2_nand2_1 _11456_ (.Y(_02960_),
    .A(net2225),
    .B(net5160));
 sg13g2_o21ai_1 _11457_ (.B1(_02960_),
    .Y(_00034_),
    .A1(net5746),
    .A2(net5160));
 sg13g2_and2_2 _11458_ (.A(net5805),
    .B(net5806),
    .X(_02961_));
 sg13g2_nand2_2 _11459_ (.Y(_02962_),
    .A(net5805),
    .B(net5806));
 sg13g2_nor2_2 _11460_ (.A(_02937_),
    .B(_02962_),
    .Y(_02963_));
 sg13g2_nand2_2 _11461_ (.Y(_02964_),
    .A(_02936_),
    .B(_02961_));
 sg13g2_nand3b_1 _11462_ (.B(_02946_),
    .C(\mem.addr[5] ),
    .Y(_02965_),
    .A_N(net5804));
 sg13g2_nor2_2 _11463_ (.A(\mem.addr[7] ),
    .B(net5803),
    .Y(_02966_));
 sg13g2_nor2b_2 _11464_ (.A(net5228),
    .B_N(_02966_),
    .Y(_02967_));
 sg13g2_nand2b_2 _11465_ (.Y(_02968_),
    .B(_02966_),
    .A_N(net5228));
 sg13g2_nand2_2 _11466_ (.Y(_02969_),
    .A(_02963_),
    .B(_02967_));
 sg13g2_nand2_1 _11467_ (.Y(_02970_),
    .A(net3234),
    .B(net5158));
 sg13g2_o21ai_1 _11468_ (.B1(_02970_),
    .Y(_00035_),
    .A1(net5463),
    .A2(net5158));
 sg13g2_nand2_1 _11469_ (.Y(_02971_),
    .A(net2260),
    .B(net5159));
 sg13g2_o21ai_1 _11470_ (.B1(_02971_),
    .Y(_00036_),
    .A1(net5509),
    .A2(net5159));
 sg13g2_nand2_1 _11471_ (.Y(_02972_),
    .A(net3156),
    .B(net5159));
 sg13g2_o21ai_1 _11472_ (.B1(_02972_),
    .Y(_00037_),
    .A1(net5555),
    .A2(net5159));
 sg13g2_nand2_1 _11473_ (.Y(_02973_),
    .A(net3143),
    .B(net5159));
 sg13g2_o21ai_1 _11474_ (.B1(_02973_),
    .Y(_00038_),
    .A1(net5601),
    .A2(net5159));
 sg13g2_nand2_1 _11475_ (.Y(_02974_),
    .A(net3034),
    .B(net5158));
 sg13g2_o21ai_1 _11476_ (.B1(_02974_),
    .Y(_00039_),
    .A1(net5647),
    .A2(net5158));
 sg13g2_nand2_1 _11477_ (.Y(_02975_),
    .A(net2423),
    .B(net5158));
 sg13g2_o21ai_1 _11478_ (.B1(_02975_),
    .Y(_00040_),
    .A1(net5691),
    .A2(net5158));
 sg13g2_nand2_1 _11479_ (.Y(_02976_),
    .A(net3062),
    .B(net5158));
 sg13g2_o21ai_1 _11480_ (.B1(_02976_),
    .Y(_00041_),
    .A1(net5735),
    .A2(net5158));
 sg13g2_nand2_1 _11481_ (.Y(_02977_),
    .A(net3087),
    .B(net5159));
 sg13g2_o21ai_1 _11482_ (.B1(_02977_),
    .Y(_00042_),
    .A1(net5781),
    .A2(net5159));
 sg13g2_nor2b_2 _11483_ (.A(net5806),
    .B_N(net5805),
    .Y(_02978_));
 sg13g2_nand2b_2 _11484_ (.Y(_02979_),
    .B(net5805),
    .A_N(net5806));
 sg13g2_nor2_2 _11485_ (.A(_02937_),
    .B(_02979_),
    .Y(_02980_));
 sg13g2_nand2_2 _11486_ (.Y(_02981_),
    .A(_02936_),
    .B(_02978_));
 sg13g2_nor2_2 _11487_ (.A(net5222),
    .B(_02981_),
    .Y(_02982_));
 sg13g2_nor2_1 _11488_ (.A(net4088),
    .B(net5156),
    .Y(_02983_));
 sg13g2_a21oi_1 _11489_ (.A1(net5463),
    .A2(net5156),
    .Y(_00043_),
    .B1(_02983_));
 sg13g2_nor2_1 _11490_ (.A(net4117),
    .B(net5157),
    .Y(_02984_));
 sg13g2_a21oi_1 _11491_ (.A1(net5509),
    .A2(net5157),
    .Y(_00044_),
    .B1(_02984_));
 sg13g2_nor2_1 _11492_ (.A(net3560),
    .B(net5156),
    .Y(_02985_));
 sg13g2_a21oi_1 _11493_ (.A1(net5555),
    .A2(net5156),
    .Y(_00045_),
    .B1(_02985_));
 sg13g2_nor2_1 _11494_ (.A(net3262),
    .B(net5157),
    .Y(_02986_));
 sg13g2_a21oi_1 _11495_ (.A1(net5601),
    .A2(net5157),
    .Y(_00046_),
    .B1(_02986_));
 sg13g2_nor2_1 _11496_ (.A(net3622),
    .B(net5156),
    .Y(_02987_));
 sg13g2_a21oi_1 _11497_ (.A1(net5646),
    .A2(net5156),
    .Y(_00047_),
    .B1(_02987_));
 sg13g2_nor2_1 _11498_ (.A(net4119),
    .B(net5157),
    .Y(_02988_));
 sg13g2_a21oi_1 _11499_ (.A1(net5691),
    .A2(net5157),
    .Y(_00048_),
    .B1(_02988_));
 sg13g2_nor2_1 _11500_ (.A(net3167),
    .B(net5157),
    .Y(_02989_));
 sg13g2_a21oi_1 _11501_ (.A1(net5735),
    .A2(net5157),
    .Y(_00049_),
    .B1(_02989_));
 sg13g2_nor2_1 _11502_ (.A(net3549),
    .B(net5156),
    .Y(_02990_));
 sg13g2_a21oi_1 _11503_ (.A1(net5781),
    .A2(net5156),
    .Y(_00050_),
    .B1(_02990_));
 sg13g2_nor3_1 _11504_ (.A(\mem.addr[5] ),
    .B(net5804),
    .C(_02947_),
    .Y(_02991_));
 sg13g2_nand2_1 _11505_ (.Y(_02992_),
    .A(_02949_),
    .B(net5221));
 sg13g2_nor2_1 _11506_ (.A(_02981_),
    .B(net5155),
    .Y(_02993_));
 sg13g2_nor2_1 _11507_ (.A(net2910),
    .B(net4788),
    .Y(_02994_));
 sg13g2_a21oi_1 _11508_ (.A1(net5428),
    .A2(net4788),
    .Y(_00051_),
    .B1(_02994_));
 sg13g2_nor2_1 _11509_ (.A(net3611),
    .B(net4789),
    .Y(_02995_));
 sg13g2_a21oi_1 _11510_ (.A1(net5475),
    .A2(net4789),
    .Y(_00052_),
    .B1(_02995_));
 sg13g2_nor2_1 _11511_ (.A(net3571),
    .B(net4789),
    .Y(_02996_));
 sg13g2_a21oi_1 _11512_ (.A1(net5518),
    .A2(net4789),
    .Y(_00053_),
    .B1(_02996_));
 sg13g2_nor2_1 _11513_ (.A(net3556),
    .B(net4789),
    .Y(_02997_));
 sg13g2_a21oi_1 _11514_ (.A1(net5565),
    .A2(net4789),
    .Y(_00054_),
    .B1(_02997_));
 sg13g2_nor2_1 _11515_ (.A(net3342),
    .B(net4789),
    .Y(_02998_));
 sg13g2_a21oi_1 _11516_ (.A1(net5610),
    .A2(net4789),
    .Y(_00055_),
    .B1(_02998_));
 sg13g2_nor2_1 _11517_ (.A(net3244),
    .B(net4788),
    .Y(_02999_));
 sg13g2_a21oi_1 _11518_ (.A1(net5655),
    .A2(net4788),
    .Y(_00056_),
    .B1(_02999_));
 sg13g2_nor2_1 _11519_ (.A(net3695),
    .B(net4788),
    .Y(_03000_));
 sg13g2_a21oi_1 _11520_ (.A1(net5700),
    .A2(net4788),
    .Y(_00057_),
    .B1(_03000_));
 sg13g2_nor2_1 _11521_ (.A(net3995),
    .B(net4788),
    .Y(_03001_));
 sg13g2_a21oi_1 _11522_ (.A1(net5745),
    .A2(net4788),
    .Y(_00058_),
    .B1(_03001_));
 sg13g2_nand2_1 _11523_ (.Y(_03002_),
    .A(\mem.addr[2] ),
    .B(_02961_));
 sg13g2_nand2_2 _11524_ (.Y(_03003_),
    .A(_02942_),
    .B(_02961_));
 sg13g2_inv_1 _11525_ (.Y(_03004_),
    .A(net5241));
 sg13g2_nor2_2 _11526_ (.A(net5222),
    .B(net5241),
    .Y(_03005_));
 sg13g2_nor2_1 _11527_ (.A(net3878),
    .B(net5152),
    .Y(_03006_));
 sg13g2_a21oi_1 _11528_ (.A1(net5461),
    .A2(net5152),
    .Y(_00059_),
    .B1(_03006_));
 sg13g2_nor2_1 _11529_ (.A(net3802),
    .B(net5152),
    .Y(_03007_));
 sg13g2_a21oi_1 _11530_ (.A1(net5507),
    .A2(net5152),
    .Y(_00060_),
    .B1(_03007_));
 sg13g2_nor2_1 _11531_ (.A(net3982),
    .B(net5153),
    .Y(_03008_));
 sg13g2_a21oi_1 _11532_ (.A1(net5554),
    .A2(_03005_),
    .Y(_00061_),
    .B1(_03008_));
 sg13g2_nor2_1 _11533_ (.A(net4007),
    .B(net5153),
    .Y(_03009_));
 sg13g2_a21oi_1 _11534_ (.A1(net5601),
    .A2(net5153),
    .Y(_00062_),
    .B1(_03009_));
 sg13g2_nor2_1 _11535_ (.A(net3430),
    .B(net5153),
    .Y(_03010_));
 sg13g2_a21oi_1 _11536_ (.A1(net5644),
    .A2(net5152),
    .Y(_00063_),
    .B1(_03010_));
 sg13g2_nor2_1 _11537_ (.A(net3509),
    .B(net5152),
    .Y(_03011_));
 sg13g2_a21oi_1 _11538_ (.A1(net5688),
    .A2(net5152),
    .Y(_00064_),
    .B1(_03011_));
 sg13g2_nor2_1 _11539_ (.A(net4018),
    .B(net5153),
    .Y(_03012_));
 sg13g2_a21oi_1 _11540_ (.A1(net5734),
    .A2(net5152),
    .Y(_00065_),
    .B1(_03012_));
 sg13g2_nor2_1 _11541_ (.A(net3576),
    .B(net5153),
    .Y(_03013_));
 sg13g2_a21oi_1 _11542_ (.A1(net5782),
    .A2(net5153),
    .Y(_00066_),
    .B1(_03013_));
 sg13g2_nor2b_2 _11543_ (.A(net5805),
    .B_N(net5806),
    .Y(_03014_));
 sg13g2_nand2b_2 _11544_ (.Y(_03015_),
    .B(net5806),
    .A_N(net5805));
 sg13g2_nor2_2 _11545_ (.A(_02937_),
    .B(_03015_),
    .Y(_03016_));
 sg13g2_nand2_2 _11546_ (.Y(_03017_),
    .A(_02936_),
    .B(_03014_));
 sg13g2_nor2_2 _11547_ (.A(net5222),
    .B(_03017_),
    .Y(_03018_));
 sg13g2_nor2_1 _11548_ (.A(net4076),
    .B(net5150),
    .Y(_03019_));
 sg13g2_a21oi_1 _11549_ (.A1(net5463),
    .A2(net5150),
    .Y(_00067_),
    .B1(_03019_));
 sg13g2_nor2_1 _11550_ (.A(net3958),
    .B(net5150),
    .Y(_03020_));
 sg13g2_a21oi_1 _11551_ (.A1(net5509),
    .A2(net5150),
    .Y(_00068_),
    .B1(_03020_));
 sg13g2_nor2_1 _11552_ (.A(net4067),
    .B(net5151),
    .Y(_03021_));
 sg13g2_a21oi_1 _11553_ (.A1(net5555),
    .A2(_03018_),
    .Y(_00069_),
    .B1(_03021_));
 sg13g2_nor2_1 _11554_ (.A(net3880),
    .B(net5151),
    .Y(_03022_));
 sg13g2_a21oi_1 _11555_ (.A1(net5602),
    .A2(net5151),
    .Y(_00070_),
    .B1(_03022_));
 sg13g2_nor2_1 _11556_ (.A(net3717),
    .B(net5151),
    .Y(_03023_));
 sg13g2_a21oi_1 _11557_ (.A1(net5646),
    .A2(net5151),
    .Y(_00071_),
    .B1(_03023_));
 sg13g2_nor2_1 _11558_ (.A(net3889),
    .B(net5150),
    .Y(_03024_));
 sg13g2_a21oi_1 _11559_ (.A1(net5691),
    .A2(net5150),
    .Y(_00072_),
    .B1(_03024_));
 sg13g2_nor2_1 _11560_ (.A(net3289),
    .B(net5150),
    .Y(_03025_));
 sg13g2_a21oi_1 _11561_ (.A1(net5735),
    .A2(net5150),
    .Y(_00073_),
    .B1(_03025_));
 sg13g2_nor2_1 _11562_ (.A(net3786),
    .B(net5151),
    .Y(_03026_));
 sg13g2_a21oi_1 _11563_ (.A1(net5781),
    .A2(net5151),
    .Y(_00074_),
    .B1(_03026_));
 sg13g2_nor2_1 _11564_ (.A(net5154),
    .B(_03017_),
    .Y(_03027_));
 sg13g2_nor2_1 _11565_ (.A(net3748),
    .B(net4786),
    .Y(_03028_));
 sg13g2_a21oi_1 _11566_ (.A1(net5428),
    .A2(net4786),
    .Y(_00075_),
    .B1(_03028_));
 sg13g2_nor2_1 _11567_ (.A(net3781),
    .B(net4787),
    .Y(_03029_));
 sg13g2_a21oi_1 _11568_ (.A1(net5475),
    .A2(net4787),
    .Y(_00076_),
    .B1(_03029_));
 sg13g2_nor2_1 _11569_ (.A(net3765),
    .B(net4787),
    .Y(_03030_));
 sg13g2_a21oi_1 _11570_ (.A1(net5518),
    .A2(net4787),
    .Y(_00077_),
    .B1(_03030_));
 sg13g2_nor2_1 _11571_ (.A(net3399),
    .B(net4787),
    .Y(_03031_));
 sg13g2_a21oi_1 _11572_ (.A1(net5565),
    .A2(net4787),
    .Y(_00078_),
    .B1(_03031_));
 sg13g2_nor2_1 _11573_ (.A(net3752),
    .B(net4787),
    .Y(_03032_));
 sg13g2_a21oi_1 _11574_ (.A1(net5610),
    .A2(net4787),
    .Y(_00079_),
    .B1(_03032_));
 sg13g2_nor2_1 _11575_ (.A(net3665),
    .B(net4786),
    .Y(_03033_));
 sg13g2_a21oi_1 _11576_ (.A1(net5655),
    .A2(net4786),
    .Y(_00080_),
    .B1(_03033_));
 sg13g2_nor2_1 _11577_ (.A(net3607),
    .B(net4786),
    .Y(_03034_));
 sg13g2_a21oi_1 _11578_ (.A1(net5700),
    .A2(net4786),
    .Y(_00081_),
    .B1(_03034_));
 sg13g2_nor2_1 _11579_ (.A(net3796),
    .B(net4786),
    .Y(_03035_));
 sg13g2_a21oi_1 _11580_ (.A1(net5745),
    .A2(net4786),
    .Y(_00082_),
    .B1(_03035_));
 sg13g2_nor2_1 _11581_ (.A(_02939_),
    .B(net5154),
    .Y(_03036_));
 sg13g2_nor2_1 _11582_ (.A(net3606),
    .B(net4784),
    .Y(_03037_));
 sg13g2_a21oi_1 _11583_ (.A1(net5428),
    .A2(net4784),
    .Y(_00083_),
    .B1(_03037_));
 sg13g2_nor2_1 _11584_ (.A(net3867),
    .B(net4785),
    .Y(_03038_));
 sg13g2_a21oi_1 _11585_ (.A1(net5475),
    .A2(net4785),
    .Y(_00084_),
    .B1(_03038_));
 sg13g2_nor2_1 _11586_ (.A(net3780),
    .B(net4785),
    .Y(_03039_));
 sg13g2_a21oi_1 _11587_ (.A1(net5518),
    .A2(net4785),
    .Y(_00085_),
    .B1(_03039_));
 sg13g2_nor2_1 _11588_ (.A(net3446),
    .B(net4785),
    .Y(_03040_));
 sg13g2_a21oi_1 _11589_ (.A1(net5565),
    .A2(net4785),
    .Y(_00086_),
    .B1(_03040_));
 sg13g2_nor2_1 _11590_ (.A(net3804),
    .B(net4785),
    .Y(_03041_));
 sg13g2_a21oi_1 _11591_ (.A1(net5610),
    .A2(net4785),
    .Y(_00087_),
    .B1(_03041_));
 sg13g2_nor2_1 _11592_ (.A(net3734),
    .B(net4784),
    .Y(_03042_));
 sg13g2_a21oi_1 _11593_ (.A1(net5655),
    .A2(net4784),
    .Y(_00088_),
    .B1(_03042_));
 sg13g2_nor2_1 _11594_ (.A(net3226),
    .B(net4784),
    .Y(_03043_));
 sg13g2_a21oi_1 _11595_ (.A1(net5700),
    .A2(net4784),
    .Y(_00089_),
    .B1(_03043_));
 sg13g2_nor2_1 _11596_ (.A(net3455),
    .B(net4784),
    .Y(_03044_));
 sg13g2_a21oi_1 _11597_ (.A1(net5745),
    .A2(net4784),
    .Y(_00090_),
    .B1(_03044_));
 sg13g2_nor2_2 _11598_ (.A(\mem.addr[3] ),
    .B(_02830_),
    .Y(_03045_));
 sg13g2_nand2_2 _11599_ (.Y(_03046_),
    .A(_02829_),
    .B(\mem.addr[2] ));
 sg13g2_nor2_2 _11600_ (.A(_02962_),
    .B(_03046_),
    .Y(_03047_));
 sg13g2_nand2_1 _11601_ (.Y(_03048_),
    .A(net5223),
    .B(net5237));
 sg13g2_nand2_1 _11602_ (.Y(_03049_),
    .A(net3140),
    .B(net5148));
 sg13g2_o21ai_1 _11603_ (.B1(_03049_),
    .Y(_00091_),
    .A1(net5423),
    .A2(net5148));
 sg13g2_nand2_1 _11604_ (.Y(_03050_),
    .A(net2892),
    .B(net5149));
 sg13g2_o21ai_1 _11605_ (.B1(_03050_),
    .Y(_00092_),
    .A1(net5468),
    .A2(net5149));
 sg13g2_nand2_1 _11606_ (.Y(_03051_),
    .A(net2872),
    .B(net5148));
 sg13g2_o21ai_1 _11607_ (.B1(_03051_),
    .Y(_00093_),
    .A1(net5513),
    .A2(net5148));
 sg13g2_nand2_1 _11608_ (.Y(_03052_),
    .A(net3201),
    .B(net5148));
 sg13g2_o21ai_1 _11609_ (.B1(_03052_),
    .Y(_00094_),
    .A1(net5558),
    .A2(net5148));
 sg13g2_nand2_1 _11610_ (.Y(_03053_),
    .A(net3057),
    .B(net5149));
 sg13g2_o21ai_1 _11611_ (.B1(_03053_),
    .Y(_00095_),
    .A1(net5605),
    .A2(_03048_));
 sg13g2_nand2_1 _11612_ (.Y(_03054_),
    .A(net2839),
    .B(net5148));
 sg13g2_o21ai_1 _11613_ (.B1(_03054_),
    .Y(_00096_),
    .A1(net5649),
    .A2(net5148));
 sg13g2_nand2_1 _11614_ (.Y(_03055_),
    .A(net3270),
    .B(net5149));
 sg13g2_o21ai_1 _11615_ (.B1(_03055_),
    .Y(_00097_),
    .A1(net5694),
    .A2(net5149));
 sg13g2_nand2_1 _11616_ (.Y(_03056_),
    .A(net3296),
    .B(net5149));
 sg13g2_o21ai_1 _11617_ (.B1(_03056_),
    .Y(_00098_),
    .A1(net5742),
    .A2(net5149));
 sg13g2_nand3_1 _11618_ (.B(net5221),
    .C(net5237),
    .A(_02949_),
    .Y(_03057_));
 sg13g2_nand2_1 _11619_ (.Y(_03058_),
    .A(net2211),
    .B(net5147));
 sg13g2_o21ai_1 _11620_ (.B1(_03058_),
    .Y(_00099_),
    .A1(net5429),
    .A2(net5147));
 sg13g2_nand2_1 _11621_ (.Y(_03059_),
    .A(net2882),
    .B(net5147));
 sg13g2_o21ai_1 _11622_ (.B1(_03059_),
    .Y(_00100_),
    .A1(net5473),
    .A2(_03057_));
 sg13g2_nand2_1 _11623_ (.Y(_03060_),
    .A(net2219),
    .B(net5147));
 sg13g2_o21ai_1 _11624_ (.B1(_03060_),
    .Y(_00101_),
    .A1(net5520),
    .A2(net5147));
 sg13g2_nand2_1 _11625_ (.Y(_03061_),
    .A(net2515),
    .B(net5147));
 sg13g2_o21ai_1 _11626_ (.B1(_03061_),
    .Y(_00102_),
    .A1(net5562),
    .A2(net5147));
 sg13g2_nand2_1 _11627_ (.Y(_03062_),
    .A(net2597),
    .B(net5146));
 sg13g2_o21ai_1 _11628_ (.B1(_03062_),
    .Y(_00103_),
    .A1(net5609),
    .A2(net5146));
 sg13g2_nand2_1 _11629_ (.Y(_03063_),
    .A(net2399),
    .B(net5146));
 sg13g2_o21ai_1 _11630_ (.B1(_03063_),
    .Y(_00104_),
    .A1(net5654),
    .A2(net5146));
 sg13g2_nand2_1 _11631_ (.Y(_03064_),
    .A(net2583),
    .B(net5146));
 sg13g2_o21ai_1 _11632_ (.B1(_03064_),
    .Y(_00105_),
    .A1(net5700),
    .A2(net5146));
 sg13g2_nand2_1 _11633_ (.Y(_03065_),
    .A(net3283),
    .B(net5146));
 sg13g2_o21ai_1 _11634_ (.B1(_03065_),
    .Y(_00106_),
    .A1(net5742),
    .A2(net5146));
 sg13g2_nor2_2 _11635_ (.A(_02979_),
    .B(_03046_),
    .Y(_03066_));
 sg13g2_nand2_2 _11636_ (.Y(_03067_),
    .A(_02978_),
    .B(_03045_));
 sg13g2_nand2_1 _11637_ (.Y(_03068_),
    .A(net5223),
    .B(net5236));
 sg13g2_nand2_1 _11638_ (.Y(_03069_),
    .A(net2160),
    .B(net5145));
 sg13g2_o21ai_1 _11639_ (.B1(_03069_),
    .Y(_00107_),
    .A1(net5423),
    .A2(net5144));
 sg13g2_nand2_1 _11640_ (.Y(_03070_),
    .A(net2309),
    .B(net5145));
 sg13g2_o21ai_1 _11641_ (.B1(_03070_),
    .Y(_00108_),
    .A1(net5468),
    .A2(net5144));
 sg13g2_nand2_1 _11642_ (.Y(_03071_),
    .A(net2947),
    .B(net5144));
 sg13g2_o21ai_1 _11643_ (.B1(_03071_),
    .Y(_00109_),
    .A1(net5513),
    .A2(net5144));
 sg13g2_nand2_1 _11644_ (.Y(_03072_),
    .A(net2467),
    .B(net5144));
 sg13g2_o21ai_1 _11645_ (.B1(_03072_),
    .Y(_00110_),
    .A1(net5558),
    .A2(net5144));
 sg13g2_nand2_1 _11646_ (.Y(_03073_),
    .A(net2314),
    .B(net5145));
 sg13g2_o21ai_1 _11647_ (.B1(_03073_),
    .Y(_00111_),
    .A1(net5605),
    .A2(net5145));
 sg13g2_nand2_1 _11648_ (.Y(_03074_),
    .A(net2362),
    .B(net5144));
 sg13g2_o21ai_1 _11649_ (.B1(_03074_),
    .Y(_00112_),
    .A1(net5649),
    .A2(net5144));
 sg13g2_nand2_1 _11650_ (.Y(_03075_),
    .A(net3481),
    .B(net5145));
 sg13g2_o21ai_1 _11651_ (.B1(_03075_),
    .Y(_00113_),
    .A1(net5694),
    .A2(net5145));
 sg13g2_nand2_1 _11652_ (.Y(_03076_),
    .A(net2167),
    .B(net5145));
 sg13g2_o21ai_1 _11653_ (.B1(_03076_),
    .Y(_00114_),
    .A1(net5742),
    .A2(net5145));
 sg13g2_nand2_1 _11654_ (.Y(_03077_),
    .A(_02966_),
    .B(net5220));
 sg13g2_nor2_2 _11655_ (.A(\mem.addr[3] ),
    .B(\mem.addr[2] ),
    .Y(_03078_));
 sg13g2_and2_2 _11656_ (.A(_02978_),
    .B(_03078_),
    .X(_03079_));
 sg13g2_nand2_2 _11657_ (.Y(_03080_),
    .A(_02978_),
    .B(_03078_));
 sg13g2_nor2_1 _11658_ (.A(net5142),
    .B(net5254),
    .Y(_03081_));
 sg13g2_nor2_1 _11659_ (.A(net3631),
    .B(net4782),
    .Y(_03082_));
 sg13g2_a21oi_1 _11660_ (.A1(net5438),
    .A2(net4782),
    .Y(_00115_),
    .B1(_03082_));
 sg13g2_nor2_1 _11661_ (.A(net3831),
    .B(net4782),
    .Y(_03083_));
 sg13g2_a21oi_1 _11662_ (.A1(net5483),
    .A2(net4782),
    .Y(_00116_),
    .B1(_03083_));
 sg13g2_nor2_1 _11663_ (.A(net3900),
    .B(net4782),
    .Y(_03084_));
 sg13g2_a21oi_1 _11664_ (.A1(net5529),
    .A2(net4782),
    .Y(_00117_),
    .B1(_03084_));
 sg13g2_nor2_1 _11665_ (.A(net3977),
    .B(net4783),
    .Y(_03085_));
 sg13g2_a21oi_1 _11666_ (.A1(net5573),
    .A2(net4783),
    .Y(_00118_),
    .B1(_03085_));
 sg13g2_nor2_1 _11667_ (.A(net3760),
    .B(net4783),
    .Y(_03086_));
 sg13g2_a21oi_1 _11668_ (.A1(net5618),
    .A2(net4783),
    .Y(_00119_),
    .B1(_03086_));
 sg13g2_nor2_1 _11669_ (.A(net3846),
    .B(net4783),
    .Y(_03087_));
 sg13g2_a21oi_1 _11670_ (.A1(net5671),
    .A2(net4783),
    .Y(_00120_),
    .B1(_03087_));
 sg13g2_nor2_1 _11671_ (.A(net3948),
    .B(net4782),
    .Y(_03088_));
 sg13g2_a21oi_1 _11672_ (.A1(net5707),
    .A2(net4782),
    .Y(_00121_),
    .B1(_03088_));
 sg13g2_nor2_1 _11673_ (.A(net4130),
    .B(net4783),
    .Y(_03089_));
 sg13g2_a21oi_1 _11674_ (.A1(net5753),
    .A2(net4783),
    .Y(_00122_),
    .B1(_03089_));
 sg13g2_nor2_1 _11675_ (.A(net5154),
    .B(_03067_),
    .Y(_03090_));
 sg13g2_nor2_1 _11676_ (.A(net3990),
    .B(net4781),
    .Y(_03091_));
 sg13g2_a21oi_1 _11677_ (.A1(net5428),
    .A2(_03090_),
    .Y(_00123_),
    .B1(_03091_));
 sg13g2_nor2_1 _11678_ (.A(net3539),
    .B(net4781),
    .Y(_03092_));
 sg13g2_a21oi_1 _11679_ (.A1(net5473),
    .A2(net4781),
    .Y(_00124_),
    .B1(_03092_));
 sg13g2_nor2_1 _11680_ (.A(net3801),
    .B(net4781),
    .Y(_03093_));
 sg13g2_a21oi_1 _11681_ (.A1(net5520),
    .A2(net4781),
    .Y(_00125_),
    .B1(_03093_));
 sg13g2_nor2_1 _11682_ (.A(net3452),
    .B(net4781),
    .Y(_03094_));
 sg13g2_a21oi_1 _11683_ (.A1(net5562),
    .A2(net4781),
    .Y(_00126_),
    .B1(_03094_));
 sg13g2_nor2_1 _11684_ (.A(net3725),
    .B(net4780),
    .Y(_03095_));
 sg13g2_a21oi_1 _11685_ (.A1(net5609),
    .A2(net4780),
    .Y(_00127_),
    .B1(_03095_));
 sg13g2_nor2_1 _11686_ (.A(net3769),
    .B(net4780),
    .Y(_03096_));
 sg13g2_a21oi_1 _11687_ (.A1(net5654),
    .A2(net4780),
    .Y(_00128_),
    .B1(_03096_));
 sg13g2_nor2_1 _11688_ (.A(net3947),
    .B(net4780),
    .Y(_03097_));
 sg13g2_a21oi_1 _11689_ (.A1(net5700),
    .A2(net4780),
    .Y(_00129_),
    .B1(_03097_));
 sg13g2_nor2_1 _11690_ (.A(net3541),
    .B(net4780),
    .Y(_03098_));
 sg13g2_a21oi_1 _11691_ (.A1(net5746),
    .A2(net4780),
    .Y(_00130_),
    .B1(_03098_));
 sg13g2_nor2_1 _11692_ (.A(_03067_),
    .B(net5142),
    .Y(_03099_));
 sg13g2_nor2_1 _11693_ (.A(net3440),
    .B(net4778),
    .Y(_03100_));
 sg13g2_a21oi_1 _11694_ (.A1(net5438),
    .A2(net4778),
    .Y(_00131_),
    .B1(_03100_));
 sg13g2_nor2_1 _11695_ (.A(net4124),
    .B(_03099_),
    .Y(_03101_));
 sg13g2_a21oi_1 _11696_ (.A1(net5483),
    .A2(net4779),
    .Y(_00132_),
    .B1(_03101_));
 sg13g2_nor2_1 _11697_ (.A(net4162),
    .B(net4779),
    .Y(_03102_));
 sg13g2_a21oi_1 _11698_ (.A1(net5527),
    .A2(net4778),
    .Y(_00133_),
    .B1(_03102_));
 sg13g2_nor2_1 _11699_ (.A(net3823),
    .B(net4778),
    .Y(_03103_));
 sg13g2_a21oi_1 _11700_ (.A1(net5571),
    .A2(net4778),
    .Y(_00134_),
    .B1(_03103_));
 sg13g2_nor2_1 _11701_ (.A(net3756),
    .B(net4779),
    .Y(_03104_));
 sg13g2_a21oi_1 _11702_ (.A1(net5629),
    .A2(net4778),
    .Y(_00135_),
    .B1(_03104_));
 sg13g2_nor2_1 _11703_ (.A(net3484),
    .B(net4779),
    .Y(_03105_));
 sg13g2_a21oi_1 _11704_ (.A1(net5670),
    .A2(net4779),
    .Y(_00136_),
    .B1(_03105_));
 sg13g2_nor2_1 _11705_ (.A(net4161),
    .B(net4778),
    .Y(_03106_));
 sg13g2_a21oi_1 _11706_ (.A1(net5717),
    .A2(net4778),
    .Y(_00137_),
    .B1(_03106_));
 sg13g2_nor2_1 _11707_ (.A(net3835),
    .B(net4779),
    .Y(_03107_));
 sg13g2_a21oi_1 _11708_ (.A1(net5762),
    .A2(net4779),
    .Y(_00138_),
    .B1(_03107_));
 sg13g2_nor2_2 _11709_ (.A(_02935_),
    .B(_03046_),
    .Y(_03108_));
 sg13g2_nand2_2 _11710_ (.Y(_03109_),
    .A(_02934_),
    .B(_03045_));
 sg13g2_nor2_1 _11711_ (.A(net5155),
    .B(_03109_),
    .Y(_03110_));
 sg13g2_nor2_1 _11712_ (.A(net3405),
    .B(net4777),
    .Y(_03111_));
 sg13g2_a21oi_1 _11713_ (.A1(net5428),
    .A2(net4777),
    .Y(_00139_),
    .B1(_03111_));
 sg13g2_nor2_1 _11714_ (.A(net3985),
    .B(_03110_),
    .Y(_03112_));
 sg13g2_a21oi_1 _11715_ (.A1(net5473),
    .A2(net4777),
    .Y(_00140_),
    .B1(_03112_));
 sg13g2_nor2_1 _11716_ (.A(net3898),
    .B(net4776),
    .Y(_03113_));
 sg13g2_a21oi_1 _11717_ (.A1(net5520),
    .A2(net4776),
    .Y(_00141_),
    .B1(_03113_));
 sg13g2_nor2_1 _11718_ (.A(net4052),
    .B(net4777),
    .Y(_03114_));
 sg13g2_a21oi_1 _11719_ (.A1(net5562),
    .A2(net4777),
    .Y(_00142_),
    .B1(_03114_));
 sg13g2_nor2_1 _11720_ (.A(net3511),
    .B(net4776),
    .Y(_03115_));
 sg13g2_a21oi_1 _11721_ (.A1(net5609),
    .A2(net4776),
    .Y(_00143_),
    .B1(_03115_));
 sg13g2_nor2_1 _11722_ (.A(net3689),
    .B(net4776),
    .Y(_03116_));
 sg13g2_a21oi_1 _11723_ (.A1(net5654),
    .A2(net4777),
    .Y(_00144_),
    .B1(_03116_));
 sg13g2_nor2_1 _11724_ (.A(net4046),
    .B(net4776),
    .Y(_03117_));
 sg13g2_a21oi_1 _11725_ (.A1(net5700),
    .A2(net4777),
    .Y(_00145_),
    .B1(_03117_));
 sg13g2_nor2_1 _11726_ (.A(net4027),
    .B(net4776),
    .Y(_03118_));
 sg13g2_a21oi_1 _11727_ (.A1(net5746),
    .A2(net4776),
    .Y(_00146_),
    .B1(_03118_));
 sg13g2_and2_2 _11728_ (.A(_02961_),
    .B(_03078_),
    .X(_03119_));
 sg13g2_nand2_2 _11729_ (.Y(_03120_),
    .A(_02961_),
    .B(_03078_));
 sg13g2_nor2_2 _11730_ (.A(net5154),
    .B(_03120_),
    .Y(_03121_));
 sg13g2_nor2_1 _11731_ (.A(net3974),
    .B(_03121_),
    .Y(_03122_));
 sg13g2_a21oi_1 _11732_ (.A1(net5429),
    .A2(net4775),
    .Y(_00147_),
    .B1(_03122_));
 sg13g2_nor2_1 _11733_ (.A(net3836),
    .B(net4775),
    .Y(_03123_));
 sg13g2_a21oi_1 _11734_ (.A1(net5473),
    .A2(net4775),
    .Y(_00148_),
    .B1(_03123_));
 sg13g2_nor2_1 _11735_ (.A(net3733),
    .B(net4775),
    .Y(_03124_));
 sg13g2_a21oi_1 _11736_ (.A1(net5514),
    .A2(net4775),
    .Y(_00149_),
    .B1(_03124_));
 sg13g2_nor2_1 _11737_ (.A(net3957),
    .B(net4775),
    .Y(_03125_));
 sg13g2_a21oi_1 _11738_ (.A1(net5562),
    .A2(net4775),
    .Y(_00150_),
    .B1(_03125_));
 sg13g2_nor2_1 _11739_ (.A(net3940),
    .B(net4774),
    .Y(_03126_));
 sg13g2_a21oi_1 _11740_ (.A1(net5609),
    .A2(net4774),
    .Y(_00151_),
    .B1(_03126_));
 sg13g2_nor2_1 _11741_ (.A(net3491),
    .B(net4774),
    .Y(_03127_));
 sg13g2_a21oi_1 _11742_ (.A1(net5651),
    .A2(net4774),
    .Y(_00152_),
    .B1(_03127_));
 sg13g2_nor2_1 _11743_ (.A(net3820),
    .B(net4774),
    .Y(_03128_));
 sg13g2_a21oi_1 _11744_ (.A1(net5694),
    .A2(net4774),
    .Y(_00153_),
    .B1(_03128_));
 sg13g2_nor2_1 _11745_ (.A(net3528),
    .B(net4774),
    .Y(_03129_));
 sg13g2_a21oi_1 _11746_ (.A1(net5740),
    .A2(net4774),
    .Y(_00154_),
    .B1(_03129_));
 sg13g2_nor2_2 _11747_ (.A(net5154),
    .B(net5254),
    .Y(_03130_));
 sg13g2_nor2_1 _11748_ (.A(net3287),
    .B(net4773),
    .Y(_03131_));
 sg13g2_a21oi_1 _11749_ (.A1(net5429),
    .A2(net4773),
    .Y(_00155_),
    .B1(_03131_));
 sg13g2_nor2_1 _11750_ (.A(net4044),
    .B(net4773),
    .Y(_03132_));
 sg13g2_a21oi_1 _11751_ (.A1(net5473),
    .A2(net4773),
    .Y(_00156_),
    .B1(_03132_));
 sg13g2_nor2_1 _11752_ (.A(net3943),
    .B(net4772),
    .Y(_03133_));
 sg13g2_a21oi_1 _11753_ (.A1(net5514),
    .A2(net4772),
    .Y(_00157_),
    .B1(_03133_));
 sg13g2_nor2_1 _11754_ (.A(net3534),
    .B(_03130_),
    .Y(_03134_));
 sg13g2_a21oi_1 _11755_ (.A1(net5562),
    .A2(net4773),
    .Y(_00158_),
    .B1(_03134_));
 sg13g2_nor2_1 _11756_ (.A(net4163),
    .B(net4773),
    .Y(_03135_));
 sg13g2_a21oi_1 _11757_ (.A1(net5604),
    .A2(net4773),
    .Y(_00159_),
    .B1(_03135_));
 sg13g2_nor2_1 _11758_ (.A(net3507),
    .B(net4772),
    .Y(_03136_));
 sg13g2_a21oi_1 _11759_ (.A1(net5651),
    .A2(net4772),
    .Y(_00160_),
    .B1(_03136_));
 sg13g2_nor2_1 _11760_ (.A(net3346),
    .B(net4772),
    .Y(_03137_));
 sg13g2_a21oi_1 _11761_ (.A1(net5694),
    .A2(net4772),
    .Y(_00161_),
    .B1(_03137_));
 sg13g2_nor2_1 _11762_ (.A(net3810),
    .B(net4772),
    .Y(_03138_));
 sg13g2_a21oi_1 _11763_ (.A1(net5740),
    .A2(net4772),
    .Y(_00162_),
    .B1(_03138_));
 sg13g2_and2_2 _11764_ (.A(_03014_),
    .B(_03078_),
    .X(_03139_));
 sg13g2_nand2_2 _11765_ (.Y(_03140_),
    .A(_03014_),
    .B(_03078_));
 sg13g2_nor2_2 _11766_ (.A(net5154),
    .B(net5252),
    .Y(_03141_));
 sg13g2_nor2_1 _11767_ (.A(net3923),
    .B(net4771),
    .Y(_03142_));
 sg13g2_a21oi_1 _11768_ (.A1(net5429),
    .A2(net4771),
    .Y(_00163_),
    .B1(_03142_));
 sg13g2_nor2_1 _11769_ (.A(net3627),
    .B(net4771),
    .Y(_03143_));
 sg13g2_a21oi_1 _11770_ (.A1(net5473),
    .A2(net4771),
    .Y(_00164_),
    .B1(_03143_));
 sg13g2_nor2_1 _11771_ (.A(net4159),
    .B(net4770),
    .Y(_03144_));
 sg13g2_a21oi_1 _11772_ (.A1(net5514),
    .A2(net4770),
    .Y(_00165_),
    .B1(_03144_));
 sg13g2_nor2_1 _11773_ (.A(net4006),
    .B(net4771),
    .Y(_03145_));
 sg13g2_a21oi_1 _11774_ (.A1(net5562),
    .A2(_03141_),
    .Y(_00166_),
    .B1(_03145_));
 sg13g2_nor2_1 _11775_ (.A(net3812),
    .B(net4770),
    .Y(_03146_));
 sg13g2_a21oi_1 _11776_ (.A1(net5604),
    .A2(net4770),
    .Y(_00167_),
    .B1(_03146_));
 sg13g2_nor2_1 _11777_ (.A(net3978),
    .B(net4771),
    .Y(_03147_));
 sg13g2_a21oi_1 _11778_ (.A1(net5651),
    .A2(net4771),
    .Y(_00168_),
    .B1(_03147_));
 sg13g2_nor2_1 _11779_ (.A(net3660),
    .B(net4770),
    .Y(_03148_));
 sg13g2_a21oi_1 _11780_ (.A1(net5694),
    .A2(net4770),
    .Y(_00169_),
    .B1(_03148_));
 sg13g2_nor2_1 _11781_ (.A(net3441),
    .B(net4770),
    .Y(_03149_));
 sg13g2_a21oi_1 _11782_ (.A1(net5740),
    .A2(net4770),
    .Y(_00170_),
    .B1(_03149_));
 sg13g2_nor2_2 _11783_ (.A(_02939_),
    .B(net5222),
    .Y(_03150_));
 sg13g2_nor2_1 _11784_ (.A(net4015),
    .B(net5141),
    .Y(_03151_));
 sg13g2_a21oi_1 _11785_ (.A1(net5463),
    .A2(net5141),
    .Y(_00171_),
    .B1(_03151_));
 sg13g2_nor2_1 _11786_ (.A(net3992),
    .B(net5140),
    .Y(_03152_));
 sg13g2_a21oi_1 _11787_ (.A1(net5508),
    .A2(net5140),
    .Y(_00172_),
    .B1(_03152_));
 sg13g2_nor2_1 _11788_ (.A(net3973),
    .B(net5140),
    .Y(_03153_));
 sg13g2_a21oi_1 _11789_ (.A1(net5555),
    .A2(net5140),
    .Y(_00173_),
    .B1(_03153_));
 sg13g2_nor2_1 _11790_ (.A(net4078),
    .B(net5140),
    .Y(_03154_));
 sg13g2_a21oi_1 _11791_ (.A1(net5601),
    .A2(net5140),
    .Y(_00174_),
    .B1(_03154_));
 sg13g2_nor2_1 _11792_ (.A(net3425),
    .B(net5140),
    .Y(_03155_));
 sg13g2_a21oi_1 _11793_ (.A1(net5646),
    .A2(net5140),
    .Y(_00175_),
    .B1(_03155_));
 sg13g2_nor2_1 _11794_ (.A(net3777),
    .B(net5141),
    .Y(_03156_));
 sg13g2_a21oi_1 _11795_ (.A1(net5691),
    .A2(net5141),
    .Y(_00176_),
    .B1(_03156_));
 sg13g2_nor2_1 _11796_ (.A(net3463),
    .B(net5141),
    .Y(_03157_));
 sg13g2_a21oi_1 _11797_ (.A1(net5735),
    .A2(net5141),
    .Y(_00177_),
    .B1(_03157_));
 sg13g2_nor2_1 _11798_ (.A(net4167),
    .B(net5141),
    .Y(_03158_));
 sg13g2_a21oi_1 _11799_ (.A1(net5781),
    .A2(_03150_),
    .Y(_00178_),
    .B1(_03158_));
 sg13g2_nor2b_1 _11800_ (.A(net5803),
    .B_N(\mem.addr[7] ),
    .Y(_03159_));
 sg13g2_nand2b_1 _11801_ (.Y(_03160_),
    .B(net5801),
    .A_N(net5803));
 sg13g2_nand2_1 _11802_ (.Y(_03161_),
    .A(net5221),
    .B(_03159_));
 sg13g2_nor2_2 _11803_ (.A(_03140_),
    .B(net5138),
    .Y(_03162_));
 sg13g2_nor2_1 _11804_ (.A(net3768),
    .B(_03162_),
    .Y(_03163_));
 sg13g2_a21oi_1 _11805_ (.A1(net5450),
    .A2(net4768),
    .Y(_00179_),
    .B1(_03163_));
 sg13g2_nor2_1 _11806_ (.A(net3788),
    .B(net4769),
    .Y(_03164_));
 sg13g2_a21oi_1 _11807_ (.A1(net5495),
    .A2(net4769),
    .Y(_00180_),
    .B1(_03164_));
 sg13g2_nor2_1 _11808_ (.A(net3830),
    .B(net4769),
    .Y(_03165_));
 sg13g2_a21oi_1 _11809_ (.A1(net5540),
    .A2(net4768),
    .Y(_00181_),
    .B1(_03165_));
 sg13g2_nor2_1 _11810_ (.A(net4025),
    .B(net4768),
    .Y(_03166_));
 sg13g2_a21oi_1 _11811_ (.A1(net5584),
    .A2(net4768),
    .Y(_00182_),
    .B1(_03166_));
 sg13g2_nor2_1 _11812_ (.A(net3994),
    .B(net4769),
    .Y(_03167_));
 sg13g2_a21oi_1 _11813_ (.A1(net5626),
    .A2(net4769),
    .Y(_00183_),
    .B1(_03167_));
 sg13g2_nor2_1 _11814_ (.A(net3527),
    .B(net4769),
    .Y(_03168_));
 sg13g2_a21oi_1 _11815_ (.A1(net5675),
    .A2(net4769),
    .Y(_00184_),
    .B1(_03168_));
 sg13g2_nor2_1 _11816_ (.A(net3881),
    .B(net4768),
    .Y(_03169_));
 sg13g2_a21oi_1 _11817_ (.A1(net5720),
    .A2(net4768),
    .Y(_00185_),
    .B1(_03169_));
 sg13g2_nor2_1 _11818_ (.A(net4145),
    .B(net4768),
    .Y(_03170_));
 sg13g2_a21oi_1 _11819_ (.A1(net5768),
    .A2(net4768),
    .Y(_00186_),
    .B1(_03170_));
 sg13g2_nor2_1 _11820_ (.A(net5142),
    .B(_03120_),
    .Y(_03171_));
 sg13g2_nor2_1 _11821_ (.A(net4158),
    .B(net4766),
    .Y(_03172_));
 sg13g2_a21oi_1 _11822_ (.A1(net5437),
    .A2(net4766),
    .Y(_00187_),
    .B1(_03172_));
 sg13g2_nor2_1 _11823_ (.A(net3803),
    .B(net4766),
    .Y(_03173_));
 sg13g2_a21oi_1 _11824_ (.A1(net5482),
    .A2(net4766),
    .Y(_00188_),
    .B1(_03173_));
 sg13g2_nor2_1 _11825_ (.A(net3339),
    .B(net4766),
    .Y(_03174_));
 sg13g2_a21oi_1 _11826_ (.A1(net5529),
    .A2(net4766),
    .Y(_00189_),
    .B1(_03174_));
 sg13g2_nor2_1 _11827_ (.A(net4173),
    .B(net4767),
    .Y(_03175_));
 sg13g2_a21oi_1 _11828_ (.A1(net5573),
    .A2(net4767),
    .Y(_00190_),
    .B1(_03175_));
 sg13g2_nor2_1 _11829_ (.A(net4127),
    .B(net4767),
    .Y(_03176_));
 sg13g2_a21oi_1 _11830_ (.A1(net5628),
    .A2(net4767),
    .Y(_00191_),
    .B1(_03176_));
 sg13g2_nor2_1 _11831_ (.A(net3858),
    .B(net4767),
    .Y(_03177_));
 sg13g2_a21oi_1 _11832_ (.A1(net5671),
    .A2(net4767),
    .Y(_00192_),
    .B1(_03177_));
 sg13g2_nor2_1 _11833_ (.A(net3613),
    .B(net4766),
    .Y(_03178_));
 sg13g2_a21oi_1 _11834_ (.A1(net5722),
    .A2(net4766),
    .Y(_00193_),
    .B1(_03178_));
 sg13g2_nor2_1 _11835_ (.A(net4143),
    .B(net4767),
    .Y(_03179_));
 sg13g2_a21oi_1 _11836_ (.A1(net5753),
    .A2(net4767),
    .Y(_00194_),
    .B1(_03179_));
 sg13g2_nand3_1 _11837_ (.B(net5804),
    .C(_02946_),
    .A(\mem.addr[5] ),
    .Y(_03180_));
 sg13g2_nor3_1 _11838_ (.A(net5801),
    .B(net5802),
    .C(_03180_),
    .Y(_03181_));
 sg13g2_nand2_1 _11839_ (.Y(_03182_),
    .A(net5243),
    .B(net5218));
 sg13g2_nand2_1 _11840_ (.Y(_03183_),
    .A(net3141),
    .B(net5136));
 sg13g2_o21ai_1 _11841_ (.B1(_03183_),
    .Y(_00195_),
    .A1(net5426),
    .A2(net5136));
 sg13g2_nand2_1 _11842_ (.Y(_03184_),
    .A(net2732),
    .B(net5136));
 sg13g2_o21ai_1 _11843_ (.B1(_03184_),
    .Y(_00196_),
    .A1(net5472),
    .A2(net5136));
 sg13g2_nand2_1 _11844_ (.Y(_03185_),
    .A(net2944),
    .B(net5136));
 sg13g2_o21ai_1 _11845_ (.B1(_03185_),
    .Y(_00197_),
    .A1(net5516),
    .A2(net5136));
 sg13g2_nand2_1 _11846_ (.Y(_03186_),
    .A(net2382),
    .B(net5137));
 sg13g2_o21ai_1 _11847_ (.B1(_03186_),
    .Y(_00198_),
    .A1(net5560),
    .A2(_03182_));
 sg13g2_nand2_1 _11848_ (.Y(_03187_),
    .A(net2255),
    .B(net5137));
 sg13g2_o21ai_1 _11849_ (.B1(_03187_),
    .Y(_00199_),
    .A1(net5607),
    .A2(net5137));
 sg13g2_nand2_1 _11850_ (.Y(_03188_),
    .A(net2737),
    .B(net5136));
 sg13g2_o21ai_1 _11851_ (.B1(_03188_),
    .Y(_00200_),
    .A1(net5653),
    .A2(net5137));
 sg13g2_nand2_1 _11852_ (.Y(_03189_),
    .A(net2677),
    .B(net5136));
 sg13g2_o21ai_1 _11853_ (.B1(_03189_),
    .Y(_00201_),
    .A1(net5698),
    .A2(net5137));
 sg13g2_nand2_1 _11854_ (.Y(_03190_),
    .A(net3454),
    .B(net5137));
 sg13g2_o21ai_1 _11855_ (.B1(_03190_),
    .Y(_00202_),
    .A1(net5744),
    .A2(net5137));
 sg13g2_nor2_1 _11856_ (.A(net5222),
    .B(_03067_),
    .Y(_03191_));
 sg13g2_nor2_1 _11857_ (.A(net3451),
    .B(net5135),
    .Y(_03192_));
 sg13g2_a21oi_1 _11858_ (.A1(net5460),
    .A2(net5135),
    .Y(_00203_),
    .B1(_03192_));
 sg13g2_nor2_1 _11859_ (.A(net3770),
    .B(net5135),
    .Y(_03193_));
 sg13g2_a21oi_1 _11860_ (.A1(net5508),
    .A2(net5135),
    .Y(_00204_),
    .B1(_03193_));
 sg13g2_nor2_1 _11861_ (.A(net3950),
    .B(net5135),
    .Y(_03194_));
 sg13g2_a21oi_1 _11862_ (.A1(net5553),
    .A2(net5135),
    .Y(_00205_),
    .B1(_03194_));
 sg13g2_nor2_1 _11863_ (.A(net3747),
    .B(net5134),
    .Y(_03195_));
 sg13g2_a21oi_1 _11864_ (.A1(net5597),
    .A2(net5134),
    .Y(_00206_),
    .B1(_03195_));
 sg13g2_nor2_1 _11865_ (.A(net3901),
    .B(net5134),
    .Y(_03196_));
 sg13g2_a21oi_1 _11866_ (.A1(net5646),
    .A2(net5134),
    .Y(_00207_),
    .B1(_03196_));
 sg13g2_nor2_1 _11867_ (.A(net3639),
    .B(net5134),
    .Y(_03197_));
 sg13g2_a21oi_1 _11868_ (.A1(net5690),
    .A2(net5134),
    .Y(_00208_),
    .B1(_03197_));
 sg13g2_nor2_1 _11869_ (.A(net3813),
    .B(net5134),
    .Y(_03198_));
 sg13g2_a21oi_1 _11870_ (.A1(net5736),
    .A2(net5134),
    .Y(_00209_),
    .B1(_03198_));
 sg13g2_nor2_1 _11871_ (.A(net3960),
    .B(net5135),
    .Y(_03199_));
 sg13g2_a21oi_1 _11872_ (.A1(net5780),
    .A2(_03191_),
    .Y(_00210_),
    .B1(_03199_));
 sg13g2_nor2_2 _11873_ (.A(_03015_),
    .B(_03046_),
    .Y(_03200_));
 sg13g2_nand2_2 _11874_ (.Y(_03201_),
    .A(_03014_),
    .B(_03045_));
 sg13g2_nor2_1 _11875_ (.A(net5222),
    .B(_03201_),
    .Y(_03202_));
 sg13g2_nor2_1 _11876_ (.A(net4104),
    .B(net5133),
    .Y(_03203_));
 sg13g2_a21oi_1 _11877_ (.A1(net5463),
    .A2(net5132),
    .Y(_00211_),
    .B1(_03203_));
 sg13g2_nor2_1 _11878_ (.A(net3433),
    .B(net5133),
    .Y(_03204_));
 sg13g2_a21oi_1 _11879_ (.A1(net5508),
    .A2(net5133),
    .Y(_00212_),
    .B1(_03204_));
 sg13g2_nor2_1 _11880_ (.A(net4156),
    .B(net5132),
    .Y(_03205_));
 sg13g2_a21oi_1 _11881_ (.A1(net5551),
    .A2(net5132),
    .Y(_00213_),
    .B1(_03205_));
 sg13g2_nor2_1 _11882_ (.A(net3934),
    .B(net5132),
    .Y(_03206_));
 sg13g2_a21oi_1 _11883_ (.A1(net5597),
    .A2(net5132),
    .Y(_00214_),
    .B1(_03206_));
 sg13g2_nor2_1 _11884_ (.A(net3470),
    .B(net5132),
    .Y(_03207_));
 sg13g2_a21oi_1 _11885_ (.A1(net5646),
    .A2(net5132),
    .Y(_00215_),
    .B1(_03207_));
 sg13g2_nor2_1 _11886_ (.A(net3565),
    .B(net5133),
    .Y(_03208_));
 sg13g2_a21oi_1 _11887_ (.A1(net5690),
    .A2(net5133),
    .Y(_00216_),
    .B1(_03208_));
 sg13g2_nor2_1 _11888_ (.A(net3912),
    .B(net5133),
    .Y(_03209_));
 sg13g2_a21oi_1 _11889_ (.A1(net5735),
    .A2(net5133),
    .Y(_00217_),
    .B1(_03209_));
 sg13g2_nor2_1 _11890_ (.A(net3389),
    .B(_03202_),
    .Y(_03210_));
 sg13g2_a21oi_1 _11891_ (.A1(net5780),
    .A2(net5132),
    .Y(_00218_),
    .B1(_03210_));
 sg13g2_nor2_2 _11892_ (.A(_02943_),
    .B(_03015_),
    .Y(_03211_));
 sg13g2_nand2_2 _11893_ (.Y(_03212_),
    .A(_02942_),
    .B(_03014_));
 sg13g2_nor2_1 _11894_ (.A(_02950_),
    .B(net5227),
    .Y(_03213_));
 sg13g2_nand2_1 _11895_ (.Y(_03214_),
    .A(net5251),
    .B(net5215));
 sg13g2_nand2_1 _11896_ (.Y(_03215_),
    .A(net3317),
    .B(net5131));
 sg13g2_o21ai_1 _11897_ (.B1(_03215_),
    .Y(_00219_),
    .A1(net5436),
    .A2(net5131));
 sg13g2_nand2_1 _11898_ (.Y(_03216_),
    .A(net2995),
    .B(net5130));
 sg13g2_o21ai_1 _11899_ (.B1(_03216_),
    .Y(_00220_),
    .A1(net5477),
    .A2(net5130));
 sg13g2_nand2_1 _11900_ (.Y(_03217_),
    .A(net2373),
    .B(net5131));
 sg13g2_o21ai_1 _11901_ (.B1(_03217_),
    .Y(_00221_),
    .A1(net5526),
    .A2(net5131));
 sg13g2_nand2_1 _11902_ (.Y(_03218_),
    .A(net2277),
    .B(net5130));
 sg13g2_o21ai_1 _11903_ (.B1(_03218_),
    .Y(_00222_),
    .A1(net5572),
    .A2(net5130));
 sg13g2_nand2_1 _11904_ (.Y(_03219_),
    .A(net3274),
    .B(net5130));
 sg13g2_o21ai_1 _11905_ (.B1(_03219_),
    .Y(_00223_),
    .A1(net5616),
    .A2(net5130));
 sg13g2_nand2_1 _11906_ (.Y(_03220_),
    .A(net3216),
    .B(net5130));
 sg13g2_o21ai_1 _11907_ (.B1(_03220_),
    .Y(_00224_),
    .A1(net5659),
    .A2(net5130));
 sg13g2_nand2_1 _11908_ (.Y(_03221_),
    .A(net3282),
    .B(net5131));
 sg13g2_o21ai_1 _11909_ (.B1(_03221_),
    .Y(_00225_),
    .A1(net5708),
    .A2(net5131));
 sg13g2_nand2_1 _11910_ (.Y(_03222_),
    .A(net2823),
    .B(net5131));
 sg13g2_o21ai_1 _11911_ (.B1(_03222_),
    .Y(_00226_),
    .A1(net5754),
    .A2(net5131));
 sg13g2_nor2_1 _11912_ (.A(net5259),
    .B(_03180_),
    .Y(_03223_));
 sg13g2_nand2_1 _11913_ (.Y(_03224_),
    .A(net5237),
    .B(net5213));
 sg13g2_nand2_1 _11914_ (.Y(_03225_),
    .A(net2421),
    .B(net5128));
 sg13g2_o21ai_1 _11915_ (.B1(_03225_),
    .Y(_00227_),
    .A1(net5434),
    .A2(net5128));
 sg13g2_nand2_1 _11916_ (.Y(_03226_),
    .A(net2591),
    .B(net5128));
 sg13g2_o21ai_1 _11917_ (.B1(_03226_),
    .Y(_00228_),
    .A1(net5480),
    .A2(net5128));
 sg13g2_nand2_1 _11918_ (.Y(_03227_),
    .A(net2714),
    .B(net5129));
 sg13g2_o21ai_1 _11919_ (.B1(_03227_),
    .Y(_00229_),
    .A1(net5518),
    .A2(net5129));
 sg13g2_nand2_1 _11920_ (.Y(_03228_),
    .A(net2435),
    .B(net5129));
 sg13g2_o21ai_1 _11921_ (.B1(_03228_),
    .Y(_00230_),
    .A1(net5565),
    .A2(net5129));
 sg13g2_nand2_1 _11922_ (.Y(_03229_),
    .A(net2577),
    .B(net5128));
 sg13g2_o21ai_1 _11923_ (.B1(_03229_),
    .Y(_00231_),
    .A1(net5614),
    .A2(net5128));
 sg13g2_nand2_1 _11924_ (.Y(_03230_),
    .A(net2221),
    .B(net5129));
 sg13g2_o21ai_1 _11925_ (.B1(_03230_),
    .Y(_00232_),
    .A1(net5654),
    .A2(net5129));
 sg13g2_nand2_1 _11926_ (.Y(_03231_),
    .A(net2523),
    .B(_03224_));
 sg13g2_o21ai_1 _11927_ (.B1(_03231_),
    .Y(_00233_),
    .A1(net5704),
    .A2(net5129));
 sg13g2_nand2_1 _11928_ (.Y(_03232_),
    .A(net2895),
    .B(net5128));
 sg13g2_o21ai_1 _11929_ (.B1(_03232_),
    .Y(_00234_),
    .A1(net5751),
    .A2(net5128));
 sg13g2_nor2_1 _11930_ (.A(net5222),
    .B(_03109_),
    .Y(_03233_));
 sg13g2_nor2_1 _11931_ (.A(net3356),
    .B(net5127),
    .Y(_03234_));
 sg13g2_a21oi_1 _11932_ (.A1(net5459),
    .A2(net5127),
    .Y(_00235_),
    .B1(_03234_));
 sg13g2_nor2_1 _11933_ (.A(net3779),
    .B(net5127),
    .Y(_03235_));
 sg13g2_a21oi_1 _11934_ (.A1(net5507),
    .A2(net5127),
    .Y(_00236_),
    .B1(_03235_));
 sg13g2_nor2_1 _11935_ (.A(net3569),
    .B(net5126),
    .Y(_03236_));
 sg13g2_a21oi_1 _11936_ (.A1(net5553),
    .A2(net5126),
    .Y(_00237_),
    .B1(_03236_));
 sg13g2_nor2_1 _11937_ (.A(net3474),
    .B(net5126),
    .Y(_03237_));
 sg13g2_a21oi_1 _11938_ (.A1(net5597),
    .A2(net5126),
    .Y(_00238_),
    .B1(_03237_));
 sg13g2_nor2_1 _11939_ (.A(net4122),
    .B(net5126),
    .Y(_03238_));
 sg13g2_a21oi_1 _11940_ (.A1(net5641),
    .A2(net5126),
    .Y(_00239_),
    .B1(_03238_));
 sg13g2_nor2_1 _11941_ (.A(net4121),
    .B(net5126),
    .Y(_03239_));
 sg13g2_a21oi_1 _11942_ (.A1(net5690),
    .A2(net5126),
    .Y(_00240_),
    .B1(_03239_));
 sg13g2_nor2_1 _11943_ (.A(net3566),
    .B(net5127),
    .Y(_03240_));
 sg13g2_a21oi_1 _11944_ (.A1(net5736),
    .A2(net5127),
    .Y(_00241_),
    .B1(_03240_));
 sg13g2_nor2_1 _11945_ (.A(net3862),
    .B(net5127),
    .Y(_03241_));
 sg13g2_a21oi_1 _11946_ (.A1(net5780),
    .A2(net5127),
    .Y(_00242_),
    .B1(_03241_));
 sg13g2_nor2_1 _11947_ (.A(net5154),
    .B(_03201_),
    .Y(_03242_));
 sg13g2_nor2_1 _11948_ (.A(net3501),
    .B(net4765),
    .Y(_03243_));
 sg13g2_a21oi_1 _11949_ (.A1(net5428),
    .A2(net4765),
    .Y(_00243_),
    .B1(_03243_));
 sg13g2_nor2_1 _11950_ (.A(net3680),
    .B(net4765),
    .Y(_03244_));
 sg13g2_a21oi_1 _11951_ (.A1(net5473),
    .A2(net4765),
    .Y(_00244_),
    .B1(_03244_));
 sg13g2_nor2_1 _11952_ (.A(net3745),
    .B(net4764),
    .Y(_03245_));
 sg13g2_a21oi_1 _11953_ (.A1(net5520),
    .A2(net4764),
    .Y(_00245_),
    .B1(_03245_));
 sg13g2_nor2_1 _11954_ (.A(net3700),
    .B(net4764),
    .Y(_03246_));
 sg13g2_a21oi_1 _11955_ (.A1(net5562),
    .A2(net4764),
    .Y(_00246_),
    .B1(_03246_));
 sg13g2_nor2_1 _11956_ (.A(net4132),
    .B(net4764),
    .Y(_03247_));
 sg13g2_a21oi_1 _11957_ (.A1(net5609),
    .A2(net4764),
    .Y(_00247_),
    .B1(_03247_));
 sg13g2_nor2_1 _11958_ (.A(net3887),
    .B(net4765),
    .Y(_03248_));
 sg13g2_a21oi_1 _11959_ (.A1(net5654),
    .A2(net4765),
    .Y(_00248_),
    .B1(_03248_));
 sg13g2_nor2_1 _11960_ (.A(net3907),
    .B(net4765),
    .Y(_03249_));
 sg13g2_a21oi_1 _11961_ (.A1(net5700),
    .A2(_03242_),
    .Y(_00249_),
    .B1(_03249_));
 sg13g2_nor2_1 _11962_ (.A(net3605),
    .B(net4764),
    .Y(_03250_));
 sg13g2_a21oi_1 _11963_ (.A1(net5746),
    .A2(net4764),
    .Y(_00250_),
    .B1(_03250_));
 sg13g2_nand2_1 _11964_ (.Y(_03251_),
    .A(net5253),
    .B(net5216));
 sg13g2_nand2_1 _11965_ (.Y(_03252_),
    .A(net2489),
    .B(net5125));
 sg13g2_o21ai_1 _11966_ (.B1(_03252_),
    .Y(_00251_),
    .A1(net5437),
    .A2(net5125));
 sg13g2_nand2_1 _11967_ (.Y(_03253_),
    .A(net3122),
    .B(net5125));
 sg13g2_o21ai_1 _11968_ (.B1(_03253_),
    .Y(_00252_),
    .A1(net5482),
    .A2(net5125));
 sg13g2_nand2_1 _11969_ (.Y(_03254_),
    .A(net2757),
    .B(net5125));
 sg13g2_o21ai_1 _11970_ (.B1(_03254_),
    .Y(_00253_),
    .A1(net5528),
    .A2(net5125));
 sg13g2_nand2_1 _11971_ (.Y(_03255_),
    .A(net2960),
    .B(net5124));
 sg13g2_o21ai_1 _11972_ (.B1(_03255_),
    .Y(_00254_),
    .A1(net5569),
    .A2(net5124));
 sg13g2_nand2_1 _11973_ (.Y(_03256_),
    .A(net2824),
    .B(net5125));
 sg13g2_o21ai_1 _11974_ (.B1(_03256_),
    .Y(_00255_),
    .A1(net5617),
    .A2(net5125));
 sg13g2_nand2_1 _11975_ (.Y(_03257_),
    .A(net2456),
    .B(net5124));
 sg13g2_o21ai_1 _11976_ (.B1(_03257_),
    .Y(_00256_),
    .A1(net5662),
    .A2(net5124));
 sg13g2_nand2_1 _11977_ (.Y(_03258_),
    .A(net3163),
    .B(net5124));
 sg13g2_o21ai_1 _11978_ (.B1(_03258_),
    .Y(_00257_),
    .A1(net5706),
    .A2(net5124));
 sg13g2_nand2_1 _11979_ (.Y(_03259_),
    .A(net2668),
    .B(net5124));
 sg13g2_o21ai_1 _11980_ (.B1(_03259_),
    .Y(_00258_),
    .A1(net5752),
    .A2(net5124));
 sg13g2_nor2_1 _11981_ (.A(_02968_),
    .B(_03120_),
    .Y(_03260_));
 sg13g2_nor2_1 _11982_ (.A(net3918),
    .B(net5123),
    .Y(_03261_));
 sg13g2_a21oi_1 _11983_ (.A1(net5464),
    .A2(net5123),
    .Y(_00259_),
    .B1(_03261_));
 sg13g2_nor2_1 _11984_ (.A(net3460),
    .B(net5123),
    .Y(_03262_));
 sg13g2_a21oi_1 _11985_ (.A1(net5508),
    .A2(net5123),
    .Y(_00260_),
    .B1(_03262_));
 sg13g2_nor2_1 _11986_ (.A(net3465),
    .B(net5122),
    .Y(_03263_));
 sg13g2_a21oi_1 _11987_ (.A1(net5552),
    .A2(net5122),
    .Y(_00261_),
    .B1(_03263_));
 sg13g2_nor2_1 _11988_ (.A(net3817),
    .B(net5122),
    .Y(_03264_));
 sg13g2_a21oi_1 _11989_ (.A1(net5597),
    .A2(net5122),
    .Y(_00262_),
    .B1(_03264_));
 sg13g2_nor2_1 _11990_ (.A(net3679),
    .B(net5122),
    .Y(_03265_));
 sg13g2_a21oi_1 _11991_ (.A1(net5646),
    .A2(net5122),
    .Y(_00263_),
    .B1(_03265_));
 sg13g2_nor2_1 _11992_ (.A(net4066),
    .B(net5122),
    .Y(_03266_));
 sg13g2_a21oi_1 _11993_ (.A1(net5690),
    .A2(net5122),
    .Y(_00264_),
    .B1(_03266_));
 sg13g2_nor2_1 _11994_ (.A(net3866),
    .B(net5123),
    .Y(_03267_));
 sg13g2_a21oi_1 _11995_ (.A1(net5736),
    .A2(net5123),
    .Y(_00265_),
    .B1(_03267_));
 sg13g2_nor2_1 _11996_ (.A(net4139),
    .B(net5123),
    .Y(_03268_));
 sg13g2_a21oi_1 _11997_ (.A1(net5780),
    .A2(net5123),
    .Y(_00266_),
    .B1(_03268_));
 sg13g2_and2_1 _11998_ (.A(net6190),
    .B(net10),
    .X(_00267_));
 sg13g2_nor2_1 _11999_ (.A(_02968_),
    .B(_03080_),
    .Y(_03269_));
 sg13g2_nor2_1 _12000_ (.A(net3961),
    .B(net5121),
    .Y(_03270_));
 sg13g2_a21oi_1 _12001_ (.A1(net5463),
    .A2(net5121),
    .Y(_00268_),
    .B1(_03270_));
 sg13g2_nor2_1 _12002_ (.A(net3644),
    .B(net5121),
    .Y(_03271_));
 sg13g2_a21oi_1 _12003_ (.A1(net5508),
    .A2(net5121),
    .Y(_00269_),
    .B1(_03271_));
 sg13g2_nor2_1 _12004_ (.A(net3911),
    .B(net5120),
    .Y(_03272_));
 sg13g2_a21oi_1 _12005_ (.A1(net5551),
    .A2(net5120),
    .Y(_00270_),
    .B1(_03272_));
 sg13g2_nor2_1 _12006_ (.A(net4072),
    .B(net5120),
    .Y(_03273_));
 sg13g2_a21oi_1 _12007_ (.A1(net5598),
    .A2(net5120),
    .Y(_00271_),
    .B1(_03273_));
 sg13g2_nor2_1 _12008_ (.A(net3494),
    .B(net5120),
    .Y(_03274_));
 sg13g2_a21oi_1 _12009_ (.A1(net5646),
    .A2(net5120),
    .Y(_00272_),
    .B1(_03274_));
 sg13g2_nor2_1 _12010_ (.A(net3832),
    .B(net5120),
    .Y(_03275_));
 sg13g2_a21oi_1 _12011_ (.A1(net5690),
    .A2(net5120),
    .Y(_00273_),
    .B1(_03275_));
 sg13g2_nor2_1 _12012_ (.A(net3568),
    .B(net5121),
    .Y(_03276_));
 sg13g2_a21oi_1 _12013_ (.A1(net5736),
    .A2(net5121),
    .Y(_00274_),
    .B1(_03276_));
 sg13g2_nor2_1 _12014_ (.A(net3946),
    .B(net5121),
    .Y(_03277_));
 sg13g2_a21oi_1 _12015_ (.A1(net5780),
    .A2(net5121),
    .Y(_00275_),
    .B1(_03277_));
 sg13g2_nor2_1 _12016_ (.A(net5230),
    .B(net5258),
    .Y(_03278_));
 sg13g2_nand2_1 _12017_ (.Y(_03279_),
    .A(_03200_),
    .B(net5211));
 sg13g2_nand2_1 _12018_ (.Y(_03280_),
    .A(net2861),
    .B(net5118));
 sg13g2_o21ai_1 _12019_ (.B1(_03280_),
    .Y(_00276_),
    .A1(net5447),
    .A2(net5118));
 sg13g2_nand2_1 _12020_ (.Y(_03281_),
    .A(net2572),
    .B(net5118));
 sg13g2_o21ai_1 _12021_ (.B1(_03281_),
    .Y(_00277_),
    .A1(net5494),
    .A2(net5118));
 sg13g2_nand2_1 _12022_ (.Y(_03282_),
    .A(net2321),
    .B(net5118));
 sg13g2_o21ai_1 _12023_ (.B1(_03282_),
    .Y(_00278_),
    .A1(net5539),
    .A2(net5118));
 sg13g2_nand2_1 _12024_ (.Y(_03283_),
    .A(net3013),
    .B(net5118));
 sg13g2_o21ai_1 _12025_ (.B1(_03283_),
    .Y(_00279_),
    .A1(net5583),
    .A2(net5118));
 sg13g2_nand2_1 _12026_ (.Y(_03284_),
    .A(net3050),
    .B(net5119));
 sg13g2_o21ai_1 _12027_ (.B1(_03284_),
    .Y(_00280_),
    .A1(net5630),
    .A2(net5119));
 sg13g2_nand2_1 _12028_ (.Y(_03285_),
    .A(net2813),
    .B(net5119));
 sg13g2_o21ai_1 _12029_ (.B1(_03285_),
    .Y(_00281_),
    .A1(net5674),
    .A2(net5119));
 sg13g2_nand2_1 _12030_ (.Y(_03286_),
    .A(net2906),
    .B(net5119));
 sg13g2_o21ai_1 _12031_ (.B1(_03286_),
    .Y(_00282_),
    .A1(net5719),
    .A2(net5119));
 sg13g2_nand2_1 _12032_ (.Y(_03287_),
    .A(net3249),
    .B(net5119));
 sg13g2_o21ai_1 _12033_ (.B1(_03287_),
    .Y(_00283_),
    .A1(net5763),
    .A2(net5119));
 sg13g2_nor2_2 _12034_ (.A(net5795),
    .B(net5788),
    .Y(_03288_));
 sg13g2_or2_2 _12035_ (.X(_03289_),
    .B(net5788),
    .A(net5795));
 sg13g2_or2_1 _12036_ (.X(_03290_),
    .B(\state[5] ),
    .A(\state[6] ));
 sg13g2_nor4_2 _12037_ (.A(net5799),
    .B(net5791),
    .C(_03289_),
    .Y(_03291_),
    .D(net5257));
 sg13g2_inv_1 _12038_ (.Y(_03292_),
    .A(net5250));
 sg13g2_nor2_2 _12039_ (.A(net11),
    .B(_02884_),
    .Y(_03293_));
 sg13g2_nand2_1 _12040_ (.Y(_03294_),
    .A(_02930_),
    .B(_03293_));
 sg13g2_a22oi_1 _12041_ (.Y(_03295_),
    .B1(_03293_),
    .B2(_02930_),
    .A2(net5250),
    .A1(_02884_));
 sg13g2_o21ai_1 _12042_ (.B1(_03294_),
    .Y(_03296_),
    .A1(halted),
    .A2(_03292_));
 sg13g2_a22oi_1 _12043_ (.Y(_03297_),
    .B1(net4255),
    .B2(net5257),
    .A2(\B[0] ),
    .A1(net5799));
 sg13g2_o21ai_1 _12044_ (.B1(_03297_),
    .Y(_03298_),
    .A1(net5806),
    .A2(_03288_));
 sg13g2_a221oi_1 _12045_ (.B2(net4223),
    .C1(_03298_),
    .B1(net5250),
    .A1(net5791),
    .Y(_03299_),
    .A2(_02906_));
 sg13g2_o21ai_1 _12046_ (.B1(net6185),
    .Y(_03300_),
    .A1(net5806),
    .A2(net5116));
 sg13g2_a21oi_1 _12047_ (.A1(net5116),
    .A2(_03299_),
    .Y(_00284_),
    .B1(_03300_));
 sg13g2_nand3_1 _12048_ (.B(_02962_),
    .C(_03289_),
    .A(_02935_),
    .Y(_03301_));
 sg13g2_a22oi_1 _12049_ (.Y(_03302_),
    .B1(\A[1] ),
    .B2(net5257),
    .A2(\B[1] ),
    .A1(net5799));
 sg13g2_nand2_1 _12050_ (.Y(_03303_),
    .A(_03301_),
    .B(_03302_));
 sg13g2_a221oi_1 _12051_ (.B2(net4230),
    .C1(_03303_),
    .B1(net5250),
    .A1(net5791),
    .Y(_03304_),
    .A2(_02911_));
 sg13g2_o21ai_1 _12052_ (.B1(net6185),
    .Y(_03305_),
    .A1(net5805),
    .A2(net5116));
 sg13g2_a21oi_1 _12053_ (.A1(net5116),
    .A2(_03304_),
    .Y(_00285_),
    .B1(_03305_));
 sg13g2_nand2_1 _12054_ (.Y(_03306_),
    .A(net5791),
    .B(_02918_));
 sg13g2_a21oi_1 _12055_ (.A1(_02830_),
    .A2(_02962_),
    .Y(_03307_),
    .B1(_03288_));
 sg13g2_a22oi_1 _12056_ (.Y(_03308_),
    .B1(net4197),
    .B2(net5257),
    .A2(net4202),
    .A1(net5799));
 sg13g2_a22oi_1 _12057_ (.Y(_03309_),
    .B1(_03307_),
    .B2(_03002_),
    .A2(net5250),
    .A1(\PC[2] ));
 sg13g2_and3_1 _12058_ (.X(_03310_),
    .A(net5116),
    .B(_03308_),
    .C(_03309_));
 sg13g2_a221oi_1 _12059_ (.B2(_03310_),
    .C1(net6177),
    .B1(net4237),
    .A1(_02830_),
    .Y(_00286_),
    .A2(_03296_));
 sg13g2_and2_1 _12060_ (.A(net5790),
    .B(_02915_),
    .X(_03311_));
 sg13g2_xnor2_1 _12061_ (.Y(_03312_),
    .A(\mem.addr[3] ),
    .B(_03002_));
 sg13g2_a22oi_1 _12062_ (.Y(_03313_),
    .B1(net5250),
    .B2(\PC[3] ),
    .A2(\B[3] ),
    .A1(net5799));
 sg13g2_a22oi_1 _12063_ (.Y(_03314_),
    .B1(_03312_),
    .B2(_03289_),
    .A2(net5257),
    .A1(\A[3] ));
 sg13g2_nand3_1 _12064_ (.B(_03313_),
    .C(_03314_),
    .A(net5116),
    .Y(_03315_));
 sg13g2_o21ai_1 _12065_ (.B1(net6187),
    .Y(_03316_),
    .A1(_03311_),
    .A2(_03315_));
 sg13g2_a21oi_1 _12066_ (.A1(_02829_),
    .A2(_03296_),
    .Y(_00287_),
    .B1(_03316_));
 sg13g2_nand2_1 _12067_ (.Y(_03317_),
    .A(net5790),
    .B(_02905_));
 sg13g2_a22oi_1 _12068_ (.Y(_03318_),
    .B1(net5250),
    .B2(\PC[4] ),
    .A2(\B[4] ),
    .A1(net5800));
 sg13g2_xnor2_1 _12069_ (.Y(_03319_),
    .A(net5804),
    .B(net5241));
 sg13g2_a22oi_1 _12070_ (.Y(_03320_),
    .B1(_03319_),
    .B2(_03289_),
    .A2(_03290_),
    .A1(net4187));
 sg13g2_nand4_1 _12071_ (.B(_03317_),
    .C(_03318_),
    .A(net5117),
    .Y(_03321_),
    .D(_03320_));
 sg13g2_o21ai_1 _12072_ (.B1(_03321_),
    .Y(_03322_),
    .A1(net5804),
    .A2(net5117));
 sg13g2_nor2_1 _12073_ (.A(net6177),
    .B(_03322_),
    .Y(_00288_));
 sg13g2_nand2_1 _12074_ (.Y(_03323_),
    .A(net5792),
    .B(_02922_));
 sg13g2_a21oi_1 _12075_ (.A1(net5804),
    .A2(_03004_),
    .Y(_03324_),
    .B1(\mem.addr[5] ));
 sg13g2_and3_1 _12076_ (.X(_03325_),
    .A(\mem.addr[5] ),
    .B(net5804),
    .C(_03004_));
 sg13g2_nor3_1 _12077_ (.A(_03288_),
    .B(_03324_),
    .C(_03325_),
    .Y(_03326_));
 sg13g2_a221oi_1 _12078_ (.B2(net5257),
    .C1(_03326_),
    .B1(\A[5] ),
    .A1(net5799),
    .Y(_03327_),
    .A2(\B[5] ));
 sg13g2_a21oi_1 _12079_ (.A1(\PC[5] ),
    .A2(_03291_),
    .Y(_03328_),
    .B1(_03296_));
 sg13g2_nand3_1 _12080_ (.B(_03327_),
    .C(_03328_),
    .A(_03323_),
    .Y(_03329_));
 sg13g2_o21ai_1 _12081_ (.B1(_03329_),
    .Y(_03330_),
    .A1(net4252),
    .A2(net5117));
 sg13g2_nor2_1 _12082_ (.A(net6178),
    .B(_03330_),
    .Y(_00289_));
 sg13g2_nand2_1 _12083_ (.Y(_03331_),
    .A(net5802),
    .B(_03325_));
 sg13g2_a21o_1 _12084_ (.A2(_03331_),
    .A1(_03289_),
    .B1(_03296_),
    .X(_03332_));
 sg13g2_o21ai_1 _12085_ (.B1(_03332_),
    .Y(_03333_),
    .A1(net5802),
    .A2(_03325_));
 sg13g2_a22oi_1 _12086_ (.Y(_03334_),
    .B1(net4188),
    .B2(net5257),
    .A2(net4189),
    .A1(net5799));
 sg13g2_inv_1 _12087_ (.Y(_03335_),
    .A(_03334_));
 sg13g2_a221oi_1 _12088_ (.B2(net4221),
    .C1(_03335_),
    .B1(_03291_),
    .A1(net5793),
    .Y(_03336_),
    .A2(_02925_));
 sg13g2_o21ai_1 _12089_ (.B1(net6187),
    .Y(_03337_),
    .A1(net5802),
    .A2(net5117));
 sg13g2_a21oi_1 _12090_ (.A1(_03333_),
    .A2(_03336_),
    .Y(_00290_),
    .B1(_03337_));
 sg13g2_a21oi_1 _12091_ (.A1(_02831_),
    .A2(net5250),
    .Y(_03338_),
    .B1(_03296_));
 sg13g2_nand2b_1 _12092_ (.Y(_03339_),
    .B(net5792),
    .A_N(_02901_));
 sg13g2_a22oi_1 _12093_ (.Y(_03340_),
    .B1(net4257),
    .B2(net5257),
    .A2(\B[7] ),
    .A1(net5799));
 sg13g2_nand3_1 _12094_ (.B(_03289_),
    .C(_03325_),
    .A(_02949_),
    .Y(_03341_));
 sg13g2_nand4_1 _12095_ (.B(_03339_),
    .C(_03340_),
    .A(_03292_),
    .Y(_03342_),
    .D(_03341_));
 sg13g2_a22oi_1 _12096_ (.Y(_03343_),
    .B1(_03338_),
    .B2(_03342_),
    .A2(_03332_),
    .A1(net5801));
 sg13g2_nor2_1 _12097_ (.A(net6177),
    .B(_03343_),
    .Y(_00291_));
 sg13g2_nor2_1 _12098_ (.A(_02968_),
    .B(net5252),
    .Y(_03344_));
 sg13g2_nor2_1 _12099_ (.A(net3885),
    .B(_03344_),
    .Y(_03345_));
 sg13g2_a21oi_1 _12100_ (.A1(net5463),
    .A2(net5115),
    .Y(_00292_),
    .B1(_03345_));
 sg13g2_nor2_1 _12101_ (.A(net3429),
    .B(net5114),
    .Y(_03346_));
 sg13g2_a21oi_1 _12102_ (.A1(net5508),
    .A2(net5114),
    .Y(_00293_),
    .B1(_03346_));
 sg13g2_nor2_1 _12103_ (.A(net4155),
    .B(net5115),
    .Y(_03347_));
 sg13g2_a21oi_1 _12104_ (.A1(net5551),
    .A2(net5115),
    .Y(_00294_),
    .B1(_03347_));
 sg13g2_nor2_1 _12105_ (.A(net3390),
    .B(net5115),
    .Y(_03348_));
 sg13g2_a21oi_1 _12106_ (.A1(net5597),
    .A2(net5115),
    .Y(_00295_),
    .B1(_03348_));
 sg13g2_nor2_1 _12107_ (.A(net4137),
    .B(net5115),
    .Y(_03349_));
 sg13g2_a21oi_1 _12108_ (.A1(net5641),
    .A2(net5115),
    .Y(_00296_),
    .B1(_03349_));
 sg13g2_nor2_1 _12109_ (.A(net3461),
    .B(net5114),
    .Y(_03350_));
 sg13g2_a21oi_1 _12110_ (.A1(net5690),
    .A2(net5114),
    .Y(_00297_),
    .B1(_03350_));
 sg13g2_nor2_1 _12111_ (.A(net3580),
    .B(net5114),
    .Y(_03351_));
 sg13g2_a21oi_1 _12112_ (.A1(net5735),
    .A2(net5114),
    .Y(_00298_),
    .B1(_03351_));
 sg13g2_nor2_1 _12113_ (.A(net4082),
    .B(net5114),
    .Y(_03352_));
 sg13g2_a21oi_1 _12114_ (.A1(net5780),
    .A2(net5114),
    .Y(_00299_),
    .B1(_03352_));
 sg13g2_and2_2 _12115_ (.A(_02934_),
    .B(_03078_),
    .X(_03353_));
 sg13g2_nand2_1 _12116_ (.Y(_03354_),
    .A(_02967_),
    .B(net5249));
 sg13g2_nand2_1 _12117_ (.Y(_03355_),
    .A(net2235),
    .B(net5113));
 sg13g2_o21ai_1 _12118_ (.B1(_03355_),
    .Y(_00300_),
    .A1(net5463),
    .A2(net5113));
 sg13g2_nand2_1 _12119_ (.Y(_03356_),
    .A(net2271),
    .B(net5113));
 sg13g2_o21ai_1 _12120_ (.B1(_03356_),
    .Y(_00301_),
    .A1(net5508),
    .A2(net5113));
 sg13g2_nand2_1 _12121_ (.Y(_03357_),
    .A(net2353),
    .B(net5112));
 sg13g2_o21ai_1 _12122_ (.B1(_03357_),
    .Y(_00302_),
    .A1(net5551),
    .A2(net5112));
 sg13g2_nand2_1 _12123_ (.Y(_03358_),
    .A(net2883),
    .B(net5112));
 sg13g2_o21ai_1 _12124_ (.B1(_03358_),
    .Y(_00303_),
    .A1(net5597),
    .A2(net5112));
 sg13g2_nand2_1 _12125_ (.Y(_03359_),
    .A(net2341),
    .B(net5112));
 sg13g2_o21ai_1 _12126_ (.B1(_03359_),
    .Y(_00304_),
    .A1(net5641),
    .A2(net5112));
 sg13g2_nand2_1 _12127_ (.Y(_03360_),
    .A(net2253),
    .B(net5112));
 sg13g2_o21ai_1 _12128_ (.B1(_03360_),
    .Y(_00305_),
    .A1(net5690),
    .A2(net5112));
 sg13g2_nand2_1 _12129_ (.Y(_03361_),
    .A(net2461),
    .B(net5113));
 sg13g2_o21ai_1 _12130_ (.B1(_03361_),
    .Y(_00306_),
    .A1(net5735),
    .A2(net5113));
 sg13g2_nand2_1 _12131_ (.Y(_03362_),
    .A(net2982),
    .B(net5113));
 sg13g2_o21ai_1 _12132_ (.B1(_03362_),
    .Y(_00307_),
    .A1(net5780),
    .A2(net5113));
 sg13g2_nor2b_2 _12133_ (.A(net5230),
    .B_N(_02966_),
    .Y(_03363_));
 sg13g2_nand2b_2 _12134_ (.Y(_03364_),
    .B(_02966_),
    .A_N(net5230));
 sg13g2_nor2_1 _12135_ (.A(net5240),
    .B(_03364_),
    .Y(_03365_));
 sg13g2_nor2_1 _12136_ (.A(net3895),
    .B(net5111),
    .Y(_03366_));
 sg13g2_a21oi_1 _12137_ (.A1(net5459),
    .A2(net5111),
    .Y(_00308_),
    .B1(_03366_));
 sg13g2_nor2_1 _12138_ (.A(net3515),
    .B(net5110),
    .Y(_03367_));
 sg13g2_a21oi_1 _12139_ (.A1(net5510),
    .A2(net5110),
    .Y(_00309_),
    .B1(_03367_));
 sg13g2_nor2_1 _12140_ (.A(net3415),
    .B(net5111),
    .Y(_03368_));
 sg13g2_a21oi_1 _12141_ (.A1(net5551),
    .A2(net5111),
    .Y(_00310_),
    .B1(_03368_));
 sg13g2_nor2_1 _12142_ (.A(net3773),
    .B(_03365_),
    .Y(_03369_));
 sg13g2_a21oi_1 _12143_ (.A1(net5597),
    .A2(net5111),
    .Y(_00311_),
    .B1(_03369_));
 sg13g2_nor2_1 _12144_ (.A(net3795),
    .B(net5111),
    .Y(_03370_));
 sg13g2_a21oi_1 _12145_ (.A1(net5640),
    .A2(net5111),
    .Y(_00312_),
    .B1(_03370_));
 sg13g2_nor2_1 _12146_ (.A(net3688),
    .B(net5110),
    .Y(_03371_));
 sg13g2_a21oi_1 _12147_ (.A1(net5689),
    .A2(net5110),
    .Y(_00313_),
    .B1(_03371_));
 sg13g2_nor2_1 _12148_ (.A(net4024),
    .B(net5110),
    .Y(_03372_));
 sg13g2_a21oi_1 _12149_ (.A1(net5730),
    .A2(net5110),
    .Y(_00314_),
    .B1(_03372_));
 sg13g2_nor2_1 _12150_ (.A(net4021),
    .B(net5110),
    .Y(_03373_));
 sg13g2_a21oi_1 _12151_ (.A1(net5778),
    .A2(net5110),
    .Y(_00315_),
    .B1(_03373_));
 sg13g2_nor2_2 _12152_ (.A(_02943_),
    .B(_02979_),
    .Y(_03374_));
 sg13g2_nand2_2 _12153_ (.Y(_03375_),
    .A(_02942_),
    .B(_02978_));
 sg13g2_nand2_2 _12154_ (.Y(_03376_),
    .A(_02967_),
    .B(net5247));
 sg13g2_nand2_1 _12155_ (.Y(_03377_),
    .A(net2175),
    .B(net5108));
 sg13g2_o21ai_1 _12156_ (.B1(_03377_),
    .Y(_00316_),
    .A1(net5461),
    .A2(net5108));
 sg13g2_nand2_1 _12157_ (.Y(_03378_),
    .A(net2838),
    .B(net5108));
 sg13g2_o21ai_1 _12158_ (.B1(_03378_),
    .Y(_00317_),
    .A1(net5507),
    .A2(net5108));
 sg13g2_nand2_1 _12159_ (.Y(_03379_),
    .A(net2182),
    .B(net5109));
 sg13g2_o21ai_1 _12160_ (.B1(_03379_),
    .Y(_00318_),
    .A1(net5554),
    .A2(net5109));
 sg13g2_nand2_1 _12161_ (.Y(_03380_),
    .A(net2173),
    .B(net5109));
 sg13g2_o21ai_1 _12162_ (.B1(_03380_),
    .Y(_00319_),
    .A1(net5601),
    .A2(net5109));
 sg13g2_nand2_1 _12163_ (.Y(_03381_),
    .A(net2663),
    .B(net5109));
 sg13g2_o21ai_1 _12164_ (.B1(_03381_),
    .Y(_00320_),
    .A1(net5644),
    .A2(net5109));
 sg13g2_nand2_1 _12165_ (.Y(_03382_),
    .A(net2966),
    .B(net5108));
 sg13g2_o21ai_1 _12166_ (.B1(_03382_),
    .Y(_00321_),
    .A1(net5688),
    .A2(net5108));
 sg13g2_nand2_1 _12167_ (.Y(_03383_),
    .A(net2357),
    .B(net5108));
 sg13g2_o21ai_1 _12168_ (.B1(_03383_),
    .Y(_00322_),
    .A1(net5733),
    .A2(net5108));
 sg13g2_nand2_1 _12169_ (.Y(_03384_),
    .A(net2770),
    .B(net5109));
 sg13g2_o21ai_1 _12170_ (.B1(_03384_),
    .Y(_00323_),
    .A1(net5779),
    .A2(net5109));
 sg13g2_nand2_1 _12171_ (.Y(_03385_),
    .A(_03363_),
    .B(net5247));
 sg13g2_nand2_1 _12172_ (.Y(_03386_),
    .A(net2164),
    .B(net5107));
 sg13g2_o21ai_1 _12173_ (.B1(_03386_),
    .Y(_00324_),
    .A1(net5459),
    .A2(net5107));
 sg13g2_nand2_1 _12174_ (.Y(_03387_),
    .A(net2337),
    .B(net5106));
 sg13g2_o21ai_1 _12175_ (.B1(_03387_),
    .Y(_00325_),
    .A1(net5510),
    .A2(net5106));
 sg13g2_nand2_1 _12176_ (.Y(_03388_),
    .A(net2956),
    .B(net5107));
 sg13g2_o21ai_1 _12177_ (.B1(_03388_),
    .Y(_00326_),
    .A1(net5551),
    .A2(_03385_));
 sg13g2_nand2_1 _12178_ (.Y(_03389_),
    .A(net2689),
    .B(net5107));
 sg13g2_o21ai_1 _12179_ (.B1(_03389_),
    .Y(_00327_),
    .A1(net5595),
    .A2(net5107));
 sg13g2_nand2_1 _12180_ (.Y(_03390_),
    .A(net2915),
    .B(net5107));
 sg13g2_o21ai_1 _12181_ (.B1(_03390_),
    .Y(_00328_),
    .A1(net5641),
    .A2(net5107));
 sg13g2_nand2_1 _12182_ (.Y(_03391_),
    .A(net3017),
    .B(net5106));
 sg13g2_o21ai_1 _12183_ (.B1(_03391_),
    .Y(_00329_),
    .A1(net5689),
    .A2(net5106));
 sg13g2_nand2_1 _12184_ (.Y(_03392_),
    .A(net2462),
    .B(net5106));
 sg13g2_o21ai_1 _12185_ (.B1(_03392_),
    .Y(_00330_),
    .A1(net5730),
    .A2(net5106));
 sg13g2_nand2_1 _12186_ (.Y(_03393_),
    .A(net3079),
    .B(net5106));
 sg13g2_o21ai_1 _12187_ (.B1(_03393_),
    .Y(_00331_),
    .A1(net5778),
    .A2(net5106));
 sg13g2_nand2_2 _12188_ (.Y(_03394_),
    .A(_02967_),
    .B(_03211_));
 sg13g2_nand2_1 _12189_ (.Y(_03395_),
    .A(net2238),
    .B(net5105));
 sg13g2_o21ai_1 _12190_ (.B1(_03395_),
    .Y(_00332_),
    .A1(net5461),
    .A2(net5105));
 sg13g2_nand2_1 _12191_ (.Y(_03396_),
    .A(net2299),
    .B(net5105));
 sg13g2_o21ai_1 _12192_ (.B1(_03396_),
    .Y(_00333_),
    .A1(net5507),
    .A2(net5105));
 sg13g2_nand2_1 _12193_ (.Y(_03397_),
    .A(net2989),
    .B(_03394_));
 sg13g2_o21ai_1 _12194_ (.B1(_03397_),
    .Y(_00334_),
    .A1(net5554),
    .A2(net5105));
 sg13g2_nand2_1 _12195_ (.Y(_03398_),
    .A(net2660),
    .B(net5104));
 sg13g2_o21ai_1 _12196_ (.B1(_03398_),
    .Y(_00335_),
    .A1(net5600),
    .A2(net5104));
 sg13g2_nand2_1 _12197_ (.Y(_03399_),
    .A(net2935),
    .B(net5104));
 sg13g2_o21ai_1 _12198_ (.B1(_03399_),
    .Y(_00336_),
    .A1(net5644),
    .A2(net5104));
 sg13g2_nand2_1 _12199_ (.Y(_03400_),
    .A(net2741),
    .B(net5105));
 sg13g2_o21ai_1 _12200_ (.B1(_03400_),
    .Y(_00337_),
    .A1(net5689),
    .A2(net5105));
 sg13g2_nand2_1 _12201_ (.Y(_03401_),
    .A(net3218),
    .B(net5104));
 sg13g2_o21ai_1 _12202_ (.B1(_03401_),
    .Y(_00338_),
    .A1(net5734),
    .A2(net5104));
 sg13g2_nand2_1 _12203_ (.Y(_03402_),
    .A(net3241),
    .B(net5104));
 sg13g2_o21ai_1 _12204_ (.B1(_03402_),
    .Y(_00339_),
    .A1(net5782),
    .A2(net5104));
 sg13g2_nand2_1 _12205_ (.Y(_03403_),
    .A(net5223),
    .B(net5234));
 sg13g2_nand2_1 _12206_ (.Y(_03404_),
    .A(net2844),
    .B(net5103));
 sg13g2_o21ai_1 _12207_ (.B1(_03404_),
    .Y(_00340_),
    .A1(net5423),
    .A2(net5103));
 sg13g2_nand2_1 _12208_ (.Y(_03405_),
    .A(net2768),
    .B(net5102));
 sg13g2_o21ai_1 _12209_ (.B1(_03405_),
    .Y(_00341_),
    .A1(net5468),
    .A2(net5102));
 sg13g2_nand2_1 _12210_ (.Y(_03406_),
    .A(net2550),
    .B(net5102));
 sg13g2_o21ai_1 _12211_ (.B1(_03406_),
    .Y(_00342_),
    .A1(net5513),
    .A2(net5102));
 sg13g2_nand2_1 _12212_ (.Y(_03407_),
    .A(net2914),
    .B(net5102));
 sg13g2_o21ai_1 _12213_ (.B1(_03407_),
    .Y(_00343_),
    .A1(net5559),
    .A2(net5102));
 sg13g2_nand2_1 _12214_ (.Y(_03408_),
    .A(net2358),
    .B(net5103));
 sg13g2_o21ai_1 _12215_ (.B1(_03408_),
    .Y(_00344_),
    .A1(net5605),
    .A2(net5103));
 sg13g2_nand2_1 _12216_ (.Y(_03409_),
    .A(net2641),
    .B(net5102));
 sg13g2_o21ai_1 _12217_ (.B1(_03409_),
    .Y(_00345_),
    .A1(net5649),
    .A2(net5102));
 sg13g2_nand2_1 _12218_ (.Y(_03410_),
    .A(net2986),
    .B(net5103));
 sg13g2_o21ai_1 _12219_ (.B1(_03410_),
    .Y(_00346_),
    .A1(net5694),
    .A2(net5103));
 sg13g2_nand2_1 _12220_ (.Y(_03411_),
    .A(net2193),
    .B(net5103));
 sg13g2_o21ai_1 _12221_ (.B1(_03411_),
    .Y(_00347_),
    .A1(net5741),
    .A2(net5103));
 sg13g2_nand3_1 _12222_ (.B(net5221),
    .C(net5248),
    .A(_02949_),
    .Y(_03412_));
 sg13g2_nand2_1 _12223_ (.Y(_03413_),
    .A(net2187),
    .B(net5101));
 sg13g2_o21ai_1 _12224_ (.B1(_03413_),
    .Y(_00348_),
    .A1(net5429),
    .A2(net5101));
 sg13g2_nand2_1 _12225_ (.Y(_03414_),
    .A(net2896),
    .B(net5101));
 sg13g2_o21ai_1 _12226_ (.B1(_03414_),
    .Y(_00349_),
    .A1(net5473),
    .A2(net5101));
 sg13g2_nand2_1 _12227_ (.Y(_03415_),
    .A(net3007),
    .B(net5100));
 sg13g2_o21ai_1 _12228_ (.B1(_03415_),
    .Y(_00350_),
    .A1(net5514),
    .A2(net5100));
 sg13g2_nand2_1 _12229_ (.Y(_03416_),
    .A(net3609),
    .B(net5101));
 sg13g2_o21ai_1 _12230_ (.B1(_03416_),
    .Y(_00351_),
    .A1(net5562),
    .A2(_03412_));
 sg13g2_nand2_1 _12231_ (.Y(_03417_),
    .A(net3595),
    .B(net5101));
 sg13g2_o21ai_1 _12232_ (.B1(_03417_),
    .Y(_00352_),
    .A1(net5604),
    .A2(net5101));
 sg13g2_nand2_1 _12233_ (.Y(_03418_),
    .A(net2292),
    .B(net5100));
 sg13g2_o21ai_1 _12234_ (.B1(_03418_),
    .Y(_00353_),
    .A1(net5651),
    .A2(net5100));
 sg13g2_nand2_1 _12235_ (.Y(_03419_),
    .A(net2633),
    .B(net5100));
 sg13g2_o21ai_1 _12236_ (.B1(_03419_),
    .Y(_00354_),
    .A1(net5694),
    .A2(net5100));
 sg13g2_nand2_1 _12237_ (.Y(_03420_),
    .A(net2840),
    .B(net5100));
 sg13g2_o21ai_1 _12238_ (.B1(_03420_),
    .Y(_00355_),
    .A1(net5740),
    .A2(net5100));
 sg13g2_and2_2 _12239_ (.A(_03004_),
    .B(net5219),
    .X(_03421_));
 sg13g2_nor2_1 _12240_ (.A(net3586),
    .B(net5098),
    .Y(_03422_));
 sg13g2_a21oi_1 _12241_ (.A1(net5427),
    .A2(net5098),
    .Y(_00356_),
    .B1(_03422_));
 sg13g2_nor2_1 _12242_ (.A(net3629),
    .B(net5098),
    .Y(_03423_));
 sg13g2_a21oi_1 _12243_ (.A1(net5471),
    .A2(net5098),
    .Y(_00357_),
    .B1(_03423_));
 sg13g2_nor2_1 _12244_ (.A(net3716),
    .B(net5098),
    .Y(_03424_));
 sg13g2_a21oi_1 _12245_ (.A1(net5525),
    .A2(net5098),
    .Y(_00358_),
    .B1(_03424_));
 sg13g2_nor2_1 _12246_ (.A(net3809),
    .B(net5099),
    .Y(_03425_));
 sg13g2_a21oi_1 _12247_ (.A1(net5569),
    .A2(net5099),
    .Y(_00359_),
    .B1(_03425_));
 sg13g2_nor2_1 _12248_ (.A(net4126),
    .B(net5099),
    .Y(_03426_));
 sg13g2_a21oi_1 _12249_ (.A1(net5606),
    .A2(net5099),
    .Y(_00360_),
    .B1(_03426_));
 sg13g2_nor2_1 _12250_ (.A(net3844),
    .B(net5099),
    .Y(_03427_));
 sg13g2_a21oi_1 _12251_ (.A1(net5661),
    .A2(net5099),
    .Y(_00361_),
    .B1(_03427_));
 sg13g2_nor2_1 _12252_ (.A(net3715),
    .B(net5099),
    .Y(_03428_));
 sg13g2_a21oi_1 _12253_ (.A1(net5705),
    .A2(net5099),
    .Y(_00362_),
    .B1(_03428_));
 sg13g2_nor2_1 _12254_ (.A(net4087),
    .B(net5098),
    .Y(_03429_));
 sg13g2_a21oi_1 _12255_ (.A1(net5743),
    .A2(net5098),
    .Y(_00363_),
    .B1(_03429_));
 sg13g2_nand2_1 _12256_ (.Y(_03430_),
    .A(net5223),
    .B(net5235));
 sg13g2_nand2_1 _12257_ (.Y(_03431_),
    .A(net2152),
    .B(net5096));
 sg13g2_o21ai_1 _12258_ (.B1(_03431_),
    .Y(_00364_),
    .A1(net5423),
    .A2(net5096));
 sg13g2_nand2_1 _12259_ (.Y(_03432_),
    .A(net3300),
    .B(net5097));
 sg13g2_o21ai_1 _12260_ (.B1(_03432_),
    .Y(_00365_),
    .A1(net5468),
    .A2(net5097));
 sg13g2_nor2_1 _12261_ (.A(\mem.data_in[2] ),
    .B(net5097),
    .Y(_03433_));
 sg13g2_a21oi_1 _12262_ (.A1(_02847_),
    .A2(net5097),
    .Y(_00366_),
    .B1(_03433_));
 sg13g2_nand2_1 _12263_ (.Y(_03434_),
    .A(net3016),
    .B(net5096));
 sg13g2_o21ai_1 _12264_ (.B1(_03434_),
    .Y(_00367_),
    .A1(net5559),
    .A2(net5096));
 sg13g2_nand2_1 _12265_ (.Y(_03435_),
    .A(net2446),
    .B(net5096));
 sg13g2_o21ai_1 _12266_ (.B1(_03435_),
    .Y(_00368_),
    .A1(net5605),
    .A2(net5096));
 sg13g2_nand2_1 _12267_ (.Y(_03436_),
    .A(net2506),
    .B(net5097));
 sg13g2_o21ai_1 _12268_ (.B1(_03436_),
    .Y(_00369_),
    .A1(net5649),
    .A2(net5097));
 sg13g2_nand2_1 _12269_ (.Y(_03437_),
    .A(net2468),
    .B(net5096));
 sg13g2_o21ai_1 _12270_ (.B1(_03437_),
    .Y(_00370_),
    .A1(net5694),
    .A2(net5096));
 sg13g2_nand2_1 _12271_ (.Y(_03438_),
    .A(net3368),
    .B(net5097));
 sg13g2_o21ai_1 _12272_ (.B1(_03438_),
    .Y(_00371_),
    .A1(net5741),
    .A2(net5097));
 sg13g2_nand2_1 _12273_ (.Y(_03439_),
    .A(net5219),
    .B(net5246));
 sg13g2_nand2_1 _12274_ (.Y(_03440_),
    .A(net2951),
    .B(net5095));
 sg13g2_o21ai_1 _12275_ (.B1(_03440_),
    .Y(_00372_),
    .A1(net5427),
    .A2(net5095));
 sg13g2_nand2_1 _12276_ (.Y(_03441_),
    .A(net3210),
    .B(net5094));
 sg13g2_o21ai_1 _12277_ (.B1(_03441_),
    .Y(_00373_),
    .A1(net5471),
    .A2(net5094));
 sg13g2_nand2_1 _12278_ (.Y(_03442_),
    .A(net3155),
    .B(net5095));
 sg13g2_o21ai_1 _12279_ (.B1(_03442_),
    .Y(_00374_),
    .A1(net5524),
    .A2(net5095));
 sg13g2_nand2_1 _12280_ (.Y(_03443_),
    .A(net3222),
    .B(net5094));
 sg13g2_o21ai_1 _12281_ (.B1(_03443_),
    .Y(_00375_),
    .A1(net5570),
    .A2(net5094));
 sg13g2_nand2_1 _12282_ (.Y(_03444_),
    .A(net2801),
    .B(net5094));
 sg13g2_o21ai_1 _12283_ (.B1(_03444_),
    .Y(_00376_),
    .A1(net5607),
    .A2(net5094));
 sg13g2_nand2_1 _12284_ (.Y(_03445_),
    .A(net3930),
    .B(net5095));
 sg13g2_o21ai_1 _12285_ (.B1(_03445_),
    .Y(_00377_),
    .A1(net5661),
    .A2(_03439_));
 sg13g2_nand2_1 _12286_ (.Y(_03446_),
    .A(net2244),
    .B(net5094));
 sg13g2_o21ai_1 _12287_ (.B1(_03446_),
    .Y(_00378_),
    .A1(net5697),
    .A2(net5094));
 sg13g2_nor2_1 _12288_ (.A(\mem.data_in[7] ),
    .B(net5095),
    .Y(_03447_));
 sg13g2_a21oi_1 _12289_ (.A1(_02877_),
    .A2(net5095),
    .Y(_00379_),
    .B1(_03447_));
 sg13g2_nand2_1 _12290_ (.Y(_03448_),
    .A(net5219),
    .B(net5251));
 sg13g2_nand2_1 _12291_ (.Y(_03449_),
    .A(net2917),
    .B(net5092));
 sg13g2_o21ai_1 _12292_ (.B1(_03449_),
    .Y(_00380_),
    .A1(net5426),
    .A2(net5092));
 sg13g2_nand2_1 _12293_ (.Y(_03450_),
    .A(net2791),
    .B(net5092));
 sg13g2_o21ai_1 _12294_ (.B1(_03450_),
    .Y(_00381_),
    .A1(net5471),
    .A2(net5092));
 sg13g2_nand2_1 _12295_ (.Y(_03451_),
    .A(net2625),
    .B(net5093));
 sg13g2_o21ai_1 _12296_ (.B1(_03451_),
    .Y(_00382_),
    .A1(net5524),
    .A2(net5093));
 sg13g2_nand2_1 _12297_ (.Y(_03452_),
    .A(net2361),
    .B(net5093));
 sg13g2_o21ai_1 _12298_ (.B1(_03452_),
    .Y(_00383_),
    .A1(net5570),
    .A2(net5093));
 sg13g2_nand2_1 _12299_ (.Y(_03453_),
    .A(net2913),
    .B(net5092));
 sg13g2_o21ai_1 _12300_ (.B1(_03453_),
    .Y(_00384_),
    .A1(net5607),
    .A2(net5092));
 sg13g2_nand2_1 _12301_ (.Y(_03454_),
    .A(net2516),
    .B(net5093));
 sg13g2_o21ai_1 _12302_ (.B1(_03454_),
    .Y(_00385_),
    .A1(net5661),
    .A2(net5093));
 sg13g2_nand2_1 _12303_ (.Y(_03455_),
    .A(net3076),
    .B(net5092));
 sg13g2_o21ai_1 _12304_ (.B1(_03455_),
    .Y(_00386_),
    .A1(net5698),
    .A2(net5092));
 sg13g2_nand2_1 _12305_ (.Y(_03456_),
    .A(net2899),
    .B(net5093));
 sg13g2_o21ai_1 _12306_ (.B1(_03456_),
    .Y(_00387_),
    .A1(net5750),
    .A2(net5093));
 sg13g2_nand2_1 _12307_ (.Y(_03457_),
    .A(net5223),
    .B(net5253));
 sg13g2_nand2_1 _12308_ (.Y(_03458_),
    .A(net3237),
    .B(_03457_));
 sg13g2_o21ai_1 _12309_ (.B1(_03458_),
    .Y(_00388_),
    .A1(net5423),
    .A2(net5091));
 sg13g2_nand2_1 _12310_ (.Y(_03459_),
    .A(net2835),
    .B(net5091));
 sg13g2_o21ai_1 _12311_ (.B1(_03459_),
    .Y(_00389_),
    .A1(net5469),
    .A2(net5091));
 sg13g2_nand2_1 _12312_ (.Y(_03460_),
    .A(net2850),
    .B(net5090));
 sg13g2_o21ai_1 _12313_ (.B1(_03460_),
    .Y(_00390_),
    .A1(net5514),
    .A2(net5090));
 sg13g2_nand2_1 _12314_ (.Y(_03461_),
    .A(net2893),
    .B(net5090));
 sg13g2_o21ai_1 _12315_ (.B1(_03461_),
    .Y(_00391_),
    .A1(net5559),
    .A2(net5090));
 sg13g2_nand2_1 _12316_ (.Y(_03462_),
    .A(net2879),
    .B(net5091));
 sg13g2_o21ai_1 _12317_ (.B1(_03462_),
    .Y(_00392_),
    .A1(net5604),
    .A2(net5091));
 sg13g2_nand2_1 _12318_ (.Y(_03463_),
    .A(net2847),
    .B(net5090));
 sg13g2_o21ai_1 _12319_ (.B1(_03463_),
    .Y(_00393_),
    .A1(net5651),
    .A2(net5090));
 sg13g2_nand2_1 _12320_ (.Y(_03464_),
    .A(net3172),
    .B(net5091));
 sg13g2_o21ai_1 _12321_ (.B1(_03464_),
    .Y(_00394_),
    .A1(net5695),
    .A2(net5091));
 sg13g2_nand2_1 _12322_ (.Y(_03465_),
    .A(net2401),
    .B(net5090));
 sg13g2_o21ai_1 _12323_ (.B1(_03465_),
    .Y(_00395_),
    .A1(net5740),
    .A2(net5090));
 sg13g2_nor2_2 _12324_ (.A(_02935_),
    .B(_02943_),
    .Y(_03466_));
 sg13g2_nand2_2 _12325_ (.Y(_03467_),
    .A(_02934_),
    .B(_02942_));
 sg13g2_nand2_1 _12326_ (.Y(_03468_),
    .A(net5219),
    .B(net5245));
 sg13g2_nand2_1 _12327_ (.Y(_03469_),
    .A(net2192),
    .B(net5088));
 sg13g2_o21ai_1 _12328_ (.B1(_03469_),
    .Y(_00396_),
    .A1(net5426),
    .A2(net5088));
 sg13g2_nand2_1 _12329_ (.Y(_03470_),
    .A(net2185),
    .B(net5088));
 sg13g2_o21ai_1 _12330_ (.B1(_03470_),
    .Y(_00397_),
    .A1(net5472),
    .A2(net5088));
 sg13g2_nand2_1 _12331_ (.Y(_03471_),
    .A(net2924),
    .B(net5089));
 sg13g2_o21ai_1 _12332_ (.B1(_03471_),
    .Y(_00398_),
    .A1(net5524),
    .A2(net5089));
 sg13g2_nand2_1 _12333_ (.Y(_03472_),
    .A(net3052),
    .B(net5089));
 sg13g2_o21ai_1 _12334_ (.B1(_03472_),
    .Y(_00399_),
    .A1(net5570),
    .A2(net5089));
 sg13g2_nand2_1 _12335_ (.Y(_03473_),
    .A(net3015),
    .B(net5088));
 sg13g2_o21ai_1 _12336_ (.B1(_03473_),
    .Y(_00400_),
    .A1(net5607),
    .A2(net5088));
 sg13g2_nand2_1 _12337_ (.Y(_03474_),
    .A(net2280),
    .B(net5089));
 sg13g2_o21ai_1 _12338_ (.B1(_03474_),
    .Y(_00401_),
    .A1(net5661),
    .A2(net5089));
 sg13g2_nand2_1 _12339_ (.Y(_03475_),
    .A(net3383),
    .B(net5088));
 sg13g2_o21ai_1 _12340_ (.B1(_03475_),
    .Y(_00402_),
    .A1(net5697),
    .A2(net5088));
 sg13g2_nand2_1 _12341_ (.Y(_03476_),
    .A(net3029),
    .B(net5089));
 sg13g2_o21ai_1 _12342_ (.B1(_03476_),
    .Y(_00403_),
    .A1(net5750),
    .A2(net5089));
 sg13g2_nor2_1 _12343_ (.A(net5142),
    .B(_03201_),
    .Y(_03477_));
 sg13g2_nor2_1 _12344_ (.A(net3753),
    .B(net4762),
    .Y(_03478_));
 sg13g2_a21oi_1 _12345_ (.A1(net5436),
    .A2(net4762),
    .Y(_00404_),
    .B1(_03478_));
 sg13g2_nor2_1 _12346_ (.A(net3983),
    .B(net4763),
    .Y(_03479_));
 sg13g2_a21oi_1 _12347_ (.A1(net5494),
    .A2(net4763),
    .Y(_00405_),
    .B1(_03479_));
 sg13g2_nor2_1 _12348_ (.A(net3993),
    .B(net4763),
    .Y(_03480_));
 sg13g2_a21oi_1 _12349_ (.A1(net5527),
    .A2(net4763),
    .Y(_00406_),
    .B1(_03480_));
 sg13g2_nor2_1 _12350_ (.A(net3504),
    .B(net4762),
    .Y(_03481_));
 sg13g2_a21oi_1 _12351_ (.A1(net5571),
    .A2(net4762),
    .Y(_00407_),
    .B1(_03481_));
 sg13g2_nor2_1 _12352_ (.A(net3910),
    .B(net4762),
    .Y(_03482_));
 sg13g2_a21oi_1 _12353_ (.A1(net5617),
    .A2(net4762),
    .Y(_00408_),
    .B1(_03482_));
 sg13g2_nor2_1 _12354_ (.A(net3398),
    .B(net4763),
    .Y(_03483_));
 sg13g2_a21oi_1 _12355_ (.A1(net5673),
    .A2(net4763),
    .Y(_00409_),
    .B1(_03483_));
 sg13g2_nor2_1 _12356_ (.A(net3908),
    .B(net4762),
    .Y(_03484_));
 sg13g2_a21oi_1 _12357_ (.A1(net5717),
    .A2(net4762),
    .Y(_00410_),
    .B1(_03484_));
 sg13g2_nor2_1 _12358_ (.A(net3655),
    .B(net4763),
    .Y(_03485_));
 sg13g2_a21oi_1 _12359_ (.A1(net5762),
    .A2(net4763),
    .Y(_00411_),
    .B1(_03485_));
 sg13g2_nor3_2 _12360_ (.A(net5229),
    .B(net5259),
    .C(net5254),
    .Y(_03486_));
 sg13g2_nor2_1 _12361_ (.A(net4160),
    .B(_03486_),
    .Y(_03487_));
 sg13g2_a21oi_1 _12362_ (.A1(net5423),
    .A2(net5209),
    .Y(_00412_),
    .B1(_03487_));
 sg13g2_nor2_1 _12363_ (.A(net4128),
    .B(net5209),
    .Y(_03488_));
 sg13g2_a21oi_1 _12364_ (.A1(net5469),
    .A2(net5209),
    .Y(_00413_),
    .B1(_03488_));
 sg13g2_nor2_1 _12365_ (.A(net3865),
    .B(net5208),
    .Y(_03489_));
 sg13g2_a21oi_1 _12366_ (.A1(net5514),
    .A2(net5208),
    .Y(_00414_),
    .B1(_03489_));
 sg13g2_nor2_1 _12367_ (.A(net3782),
    .B(net5208),
    .Y(_03490_));
 sg13g2_a21oi_1 _12368_ (.A1(net5559),
    .A2(net5208),
    .Y(_00415_),
    .B1(_03490_));
 sg13g2_nor2_1 _12369_ (.A(net3363),
    .B(net5209),
    .Y(_03491_));
 sg13g2_a21oi_1 _12370_ (.A1(net5604),
    .A2(net5209),
    .Y(_00416_),
    .B1(_03491_));
 sg13g2_nor2_1 _12371_ (.A(net3428),
    .B(net5208),
    .Y(_03492_));
 sg13g2_a21oi_1 _12372_ (.A1(net5651),
    .A2(net5208),
    .Y(_00417_),
    .B1(_03492_));
 sg13g2_nor2_1 _12373_ (.A(net3664),
    .B(net5209),
    .Y(_03493_));
 sg13g2_a21oi_1 _12374_ (.A1(net5695),
    .A2(net5209),
    .Y(_00418_),
    .B1(_03493_));
 sg13g2_nor2_1 _12375_ (.A(net3972),
    .B(net5208),
    .Y(_03494_));
 sg13g2_a21oi_1 _12376_ (.A1(net5740),
    .A2(net5208),
    .Y(_00419_),
    .B1(_03494_));
 sg13g2_nand2_1 _12377_ (.Y(_03495_),
    .A(net5242),
    .B(net5218));
 sg13g2_nand2_1 _12378_ (.Y(_03496_),
    .A(net2169),
    .B(net5086));
 sg13g2_o21ai_1 _12379_ (.B1(_03496_),
    .Y(_00420_),
    .A1(net5426),
    .A2(net5086));
 sg13g2_nand2_1 _12380_ (.Y(_03497_),
    .A(net2288),
    .B(net5086));
 sg13g2_o21ai_1 _12381_ (.B1(_03497_),
    .Y(_00421_),
    .A1(net5472),
    .A2(net5086));
 sg13g2_nand2_1 _12382_ (.Y(_03498_),
    .A(net3042),
    .B(net5086));
 sg13g2_o21ai_1 _12383_ (.B1(_03498_),
    .Y(_00422_),
    .A1(net5516),
    .A2(net5086));
 sg13g2_nand2_1 _12384_ (.Y(_03499_),
    .A(net2284),
    .B(net5087));
 sg13g2_o21ai_1 _12385_ (.B1(_03499_),
    .Y(_00423_),
    .A1(net5560),
    .A2(_03495_));
 sg13g2_nand2_1 _12386_ (.Y(_03500_),
    .A(net3083),
    .B(net5087));
 sg13g2_o21ai_1 _12387_ (.B1(_03500_),
    .Y(_00424_),
    .A1(net5607),
    .A2(net5087));
 sg13g2_nand2_1 _12388_ (.Y(_03501_),
    .A(net2242),
    .B(net5086));
 sg13g2_o21ai_1 _12389_ (.B1(_03501_),
    .Y(_00425_),
    .A1(net5652),
    .A2(net5086));
 sg13g2_nand2_1 _12390_ (.Y(_03502_),
    .A(net2452),
    .B(net5087));
 sg13g2_o21ai_1 _12391_ (.B1(_03502_),
    .Y(_00426_),
    .A1(net5698),
    .A2(net5087));
 sg13g2_nand2_1 _12392_ (.Y(_03503_),
    .A(net2698),
    .B(net5087));
 sg13g2_o21ai_1 _12393_ (.B1(_03503_),
    .Y(_00427_),
    .A1(net5743),
    .A2(net5087));
 sg13g2_nand2_1 _12394_ (.Y(_03504_),
    .A(net5239),
    .B(net5218));
 sg13g2_nand2_1 _12395_ (.Y(_03505_),
    .A(net3228),
    .B(net5085));
 sg13g2_o21ai_1 _12396_ (.B1(_03505_),
    .Y(_00428_),
    .A1(net5426),
    .A2(net5085));
 sg13g2_nand2_1 _12397_ (.Y(_03506_),
    .A(net2336),
    .B(_03504_));
 sg13g2_o21ai_1 _12398_ (.B1(_03506_),
    .Y(_00429_),
    .A1(net5471),
    .A2(net5085));
 sg13g2_nand2_1 _12399_ (.Y(_03507_),
    .A(net3307),
    .B(net5085));
 sg13g2_o21ai_1 _12400_ (.B1(_03507_),
    .Y(_00430_),
    .A1(net5516),
    .A2(net5085));
 sg13g2_nand2_1 _12401_ (.Y(_03508_),
    .A(net3344),
    .B(net5084));
 sg13g2_o21ai_1 _12402_ (.B1(_03508_),
    .Y(_00431_),
    .A1(net5560),
    .A2(net5084));
 sg13g2_nand2_1 _12403_ (.Y(_03509_),
    .A(net3278),
    .B(net5084));
 sg13g2_o21ai_1 _12404_ (.B1(_03509_),
    .Y(_00432_),
    .A1(net5607),
    .A2(net5084));
 sg13g2_nand2_1 _12405_ (.Y(_03510_),
    .A(net2350),
    .B(net5085));
 sg13g2_o21ai_1 _12406_ (.B1(_03510_),
    .Y(_00433_),
    .A1(net5652),
    .A2(net5085));
 sg13g2_nand2_1 _12407_ (.Y(_03511_),
    .A(net3319),
    .B(net5084));
 sg13g2_o21ai_1 _12408_ (.B1(_03511_),
    .Y(_00434_),
    .A1(net5698),
    .A2(net5084));
 sg13g2_nand2_1 _12409_ (.Y(_03512_),
    .A(net2738),
    .B(net5084));
 sg13g2_o21ai_1 _12410_ (.B1(_03512_),
    .Y(_00435_),
    .A1(net5743),
    .A2(net5084));
 sg13g2_nor3_2 _12411_ (.A(net5229),
    .B(net5259),
    .C(net5252),
    .Y(_03513_));
 sg13g2_nor2_1 _12412_ (.A(net3855),
    .B(_03513_),
    .Y(_03514_));
 sg13g2_a21oi_1 _12413_ (.A1(net5423),
    .A2(net5207),
    .Y(_00436_),
    .B1(_03514_));
 sg13g2_nor2_1 _12414_ (.A(net3778),
    .B(net5206),
    .Y(_03515_));
 sg13g2_a21oi_1 _12415_ (.A1(net5469),
    .A2(net5206),
    .Y(_00437_),
    .B1(_03515_));
 sg13g2_nor2_1 _12416_ (.A(net3815),
    .B(net5206),
    .Y(_03516_));
 sg13g2_a21oi_1 _12417_ (.A1(net5514),
    .A2(net5206),
    .Y(_00438_),
    .B1(_03516_));
 sg13g2_nor2_1 _12418_ (.A(net3620),
    .B(net5206),
    .Y(_03517_));
 sg13g2_a21oi_1 _12419_ (.A1(net5559),
    .A2(net5206),
    .Y(_00439_),
    .B1(_03517_));
 sg13g2_nor2_1 _12420_ (.A(net3996),
    .B(net5207),
    .Y(_03518_));
 sg13g2_a21oi_1 _12421_ (.A1(net5604),
    .A2(net5207),
    .Y(_00440_),
    .B1(_03518_));
 sg13g2_nor2_1 _12422_ (.A(net3329),
    .B(net5206),
    .Y(_03519_));
 sg13g2_a21oi_1 _12423_ (.A1(net5651),
    .A2(net5206),
    .Y(_00441_),
    .B1(_03519_));
 sg13g2_nor2_1 _12424_ (.A(net3662),
    .B(net5207),
    .Y(_03520_));
 sg13g2_a21oi_1 _12425_ (.A1(net5695),
    .A2(net5207),
    .Y(_00442_),
    .B1(_03520_));
 sg13g2_nor2_1 _12426_ (.A(net3945),
    .B(net5207),
    .Y(_03521_));
 sg13g2_a21oi_1 _12427_ (.A1(net5740),
    .A2(net5207),
    .Y(_00443_),
    .B1(_03521_));
 sg13g2_nand2_1 _12428_ (.Y(_03522_),
    .A(net5244),
    .B(net5218));
 sg13g2_nand2_1 _12429_ (.Y(_03523_),
    .A(net2157),
    .B(net5082));
 sg13g2_o21ai_1 _12430_ (.B1(_03523_),
    .Y(_00444_),
    .A1(net5426),
    .A2(net5082));
 sg13g2_nor2_1 _12431_ (.A(\mem.data_in[1] ),
    .B(net5082),
    .Y(_03524_));
 sg13g2_a21oi_1 _12432_ (.A1(_02889_),
    .A2(net5082),
    .Y(_00445_),
    .B1(_03524_));
 sg13g2_nand2_1 _12433_ (.Y(_03525_),
    .A(net2672),
    .B(net5082));
 sg13g2_o21ai_1 _12434_ (.B1(_03525_),
    .Y(_00446_),
    .A1(net5516),
    .A2(net5082));
 sg13g2_nand2_1 _12435_ (.Y(_03526_),
    .A(net2437),
    .B(net5083));
 sg13g2_o21ai_1 _12436_ (.B1(_03526_),
    .Y(_00447_),
    .A1(net5560),
    .A2(net5083));
 sg13g2_nand2_1 _12437_ (.Y(_03527_),
    .A(net3149),
    .B(net5083));
 sg13g2_o21ai_1 _12438_ (.B1(_03527_),
    .Y(_00448_),
    .A1(net5607),
    .A2(net5083));
 sg13g2_nand2_1 _12439_ (.Y(_03528_),
    .A(net3116),
    .B(net5083));
 sg13g2_o21ai_1 _12440_ (.B1(_03528_),
    .Y(_00449_),
    .A1(net5652),
    .A2(net5083));
 sg13g2_nand2_1 _12441_ (.Y(_03529_),
    .A(net3054),
    .B(net5083));
 sg13g2_o21ai_1 _12442_ (.B1(_03529_),
    .Y(_00450_),
    .A1(net5698),
    .A2(net5083));
 sg13g2_nand2_1 _12443_ (.Y(_03530_),
    .A(net3238),
    .B(net5082));
 sg13g2_o21ai_1 _12444_ (.B1(_03530_),
    .Y(_00451_),
    .A1(net5743),
    .A2(net5082));
 sg13g2_nand2_1 _12445_ (.Y(_03531_),
    .A(net5237),
    .B(net5217));
 sg13g2_nand2_1 _12446_ (.Y(_03532_),
    .A(net2849),
    .B(net5081));
 sg13g2_o21ai_1 _12447_ (.B1(_03532_),
    .Y(_00452_),
    .A1(net5427),
    .A2(net5081));
 sg13g2_nand2_1 _12448_ (.Y(_03533_),
    .A(net2195),
    .B(net5080));
 sg13g2_o21ai_1 _12449_ (.B1(_03533_),
    .Y(_00453_),
    .A1(net5471),
    .A2(net5080));
 sg13g2_nand2_1 _12450_ (.Y(_03534_),
    .A(net2324),
    .B(net5081));
 sg13g2_o21ai_1 _12451_ (.B1(_03534_),
    .Y(_00454_),
    .A1(net5516),
    .A2(net5081));
 sg13g2_nand2_1 _12452_ (.Y(_03535_),
    .A(net3221),
    .B(net5081));
 sg13g2_o21ai_1 _12453_ (.B1(_03535_),
    .Y(_00455_),
    .A1(net5561),
    .A2(net5081));
 sg13g2_nand2_1 _12454_ (.Y(_03536_),
    .A(net2370),
    .B(net5080));
 sg13g2_o21ai_1 _12455_ (.B1(_03536_),
    .Y(_00456_),
    .A1(net5606),
    .A2(net5080));
 sg13g2_nand2_1 _12456_ (.Y(_03537_),
    .A(net2318),
    .B(net5081));
 sg13g2_o21ai_1 _12457_ (.B1(_03537_),
    .Y(_00457_),
    .A1(net5652),
    .A2(net5081));
 sg13g2_nand2_1 _12458_ (.Y(_03538_),
    .A(net2262),
    .B(net5080));
 sg13g2_o21ai_1 _12459_ (.B1(_03538_),
    .Y(_00458_),
    .A1(net5697),
    .A2(net5080));
 sg13g2_nand2_1 _12460_ (.Y(_03539_),
    .A(net2600),
    .B(net5080));
 sg13g2_o21ai_1 _12461_ (.B1(_03539_),
    .Y(_00459_),
    .A1(net5743),
    .A2(net5080));
 sg13g2_nand2_1 _12462_ (.Y(_03540_),
    .A(net5223),
    .B(net5248));
 sg13g2_nand2_1 _12463_ (.Y(_03541_),
    .A(net3199),
    .B(_03540_));
 sg13g2_o21ai_1 _12464_ (.B1(_03541_),
    .Y(_00460_),
    .A1(net5423),
    .A2(net5079));
 sg13g2_nand2_1 _12465_ (.Y(_03542_),
    .A(net2977),
    .B(net5078));
 sg13g2_o21ai_1 _12466_ (.B1(_03542_),
    .Y(_00461_),
    .A1(net5469),
    .A2(net5078));
 sg13g2_nand2_1 _12467_ (.Y(_03543_),
    .A(net2865),
    .B(net5078));
 sg13g2_o21ai_1 _12468_ (.B1(_03543_),
    .Y(_00462_),
    .A1(net5514),
    .A2(net5078));
 sg13g2_nand2_1 _12469_ (.Y(_03544_),
    .A(net2199),
    .B(net5078));
 sg13g2_o21ai_1 _12470_ (.B1(_03544_),
    .Y(_00463_),
    .A1(net5559),
    .A2(net5078));
 sg13g2_nand2_1 _12471_ (.Y(_03545_),
    .A(net2513),
    .B(net5079));
 sg13g2_o21ai_1 _12472_ (.B1(_03545_),
    .Y(_00464_),
    .A1(net5604),
    .A2(net5079));
 sg13g2_nand2_1 _12473_ (.Y(_03546_),
    .A(net2857),
    .B(net5078));
 sg13g2_o21ai_1 _12474_ (.B1(_03546_),
    .Y(_00465_),
    .A1(net5651),
    .A2(net5078));
 sg13g2_nand2_1 _12475_ (.Y(_03547_),
    .A(net2243),
    .B(net5079));
 sg13g2_o21ai_1 _12476_ (.B1(_03547_),
    .Y(_00466_),
    .A1(net5695),
    .A2(net5079));
 sg13g2_nand2_1 _12477_ (.Y(_03548_),
    .A(net3250),
    .B(net5079));
 sg13g2_o21ai_1 _12478_ (.B1(_03548_),
    .Y(_00467_),
    .A1(net5740),
    .A2(net5079));
 sg13g2_nand2_1 _12479_ (.Y(_03549_),
    .A(net5236),
    .B(net5217));
 sg13g2_nand2_1 _12480_ (.Y(_03550_),
    .A(net2162),
    .B(net5077));
 sg13g2_o21ai_1 _12481_ (.B1(_03550_),
    .Y(_00468_),
    .A1(net5427),
    .A2(net5077));
 sg13g2_nand2_1 _12482_ (.Y(_03551_),
    .A(net3128),
    .B(net5076));
 sg13g2_o21ai_1 _12483_ (.B1(_03551_),
    .Y(_00469_),
    .A1(net5471),
    .A2(net5076));
 sg13g2_nand2_1 _12484_ (.Y(_03552_),
    .A(net2611),
    .B(net5077));
 sg13g2_o21ai_1 _12485_ (.B1(_03552_),
    .Y(_00470_),
    .A1(net5516),
    .A2(net5077));
 sg13g2_nand2_1 _12486_ (.Y(_03553_),
    .A(net2713),
    .B(net5077));
 sg13g2_o21ai_1 _12487_ (.B1(_03553_),
    .Y(_00471_),
    .A1(net5560),
    .A2(net5077));
 sg13g2_nand2_1 _12488_ (.Y(_03554_),
    .A(net2236),
    .B(net5076));
 sg13g2_o21ai_1 _12489_ (.B1(_03554_),
    .Y(_00472_),
    .A1(net5606),
    .A2(net5076));
 sg13g2_nand2_1 _12490_ (.Y(_03555_),
    .A(net2330),
    .B(net5077));
 sg13g2_o21ai_1 _12491_ (.B1(_03555_),
    .Y(_00473_),
    .A1(net5652),
    .A2(net5077));
 sg13g2_nand2_1 _12492_ (.Y(_03556_),
    .A(net3369),
    .B(net5076));
 sg13g2_o21ai_1 _12493_ (.B1(_03556_),
    .Y(_00474_),
    .A1(net5697),
    .A2(net5076));
 sg13g2_nand2_1 _12494_ (.Y(_03557_),
    .A(net2623),
    .B(net5076));
 sg13g2_o21ai_1 _12495_ (.B1(_03557_),
    .Y(_00475_),
    .A1(net5743),
    .A2(net5076));
 sg13g2_nand2_1 _12496_ (.Y(_03558_),
    .A(net5217),
    .B(net5234));
 sg13g2_nand2_1 _12497_ (.Y(_03559_),
    .A(net3230),
    .B(net5075));
 sg13g2_o21ai_1 _12498_ (.B1(_03559_),
    .Y(_00476_),
    .A1(net5426),
    .A2(net5075));
 sg13g2_nand2_1 _12499_ (.Y(_03560_),
    .A(net3136),
    .B(net5074));
 sg13g2_o21ai_1 _12500_ (.B1(_03560_),
    .Y(_00477_),
    .A1(net5471),
    .A2(net5074));
 sg13g2_nand2_1 _12501_ (.Y(_03561_),
    .A(net3280),
    .B(net5074));
 sg13g2_o21ai_1 _12502_ (.B1(_03561_),
    .Y(_00478_),
    .A1(net5517),
    .A2(net5074));
 sg13g2_nand2_1 _12503_ (.Y(_03562_),
    .A(net2404),
    .B(net5075));
 sg13g2_o21ai_1 _12504_ (.B1(_03562_),
    .Y(_00479_),
    .A1(net5560),
    .A2(net5075));
 sg13g2_nand2_1 _12505_ (.Y(_03563_),
    .A(net3110),
    .B(net5075));
 sg13g2_o21ai_1 _12506_ (.B1(_03563_),
    .Y(_00480_),
    .A1(net5606),
    .A2(net5075));
 sg13g2_nand2_1 _12507_ (.Y(_03564_),
    .A(net2905),
    .B(net5075));
 sg13g2_o21ai_1 _12508_ (.B1(_03564_),
    .Y(_00481_),
    .A1(net5652),
    .A2(net5075));
 sg13g2_nand2_1 _12509_ (.Y(_03565_),
    .A(net2657),
    .B(net5074));
 sg13g2_o21ai_1 _12510_ (.B1(_03565_),
    .Y(_00482_),
    .A1(net5697),
    .A2(net5074));
 sg13g2_nand2_1 _12511_ (.Y(_03566_),
    .A(net2339),
    .B(net5074));
 sg13g2_o21ai_1 _12512_ (.B1(_03566_),
    .Y(_00483_),
    .A1(net5743),
    .A2(net5074));
 sg13g2_nand3_1 _12513_ (.B(net5220),
    .C(net5237),
    .A(_02966_),
    .Y(_03567_));
 sg13g2_nand2_1 _12514_ (.Y(_03568_),
    .A(net3166),
    .B(net5073));
 sg13g2_o21ai_1 _12515_ (.B1(_03568_),
    .Y(_00484_),
    .A1(net5436),
    .A2(net5073));
 sg13g2_nand2_1 _12516_ (.Y(_03569_),
    .A(net2345),
    .B(net5073));
 sg13g2_o21ai_1 _12517_ (.B1(_03569_),
    .Y(_00485_),
    .A1(net5483),
    .A2(net5073));
 sg13g2_nand2_1 _12518_ (.Y(_03570_),
    .A(net2519),
    .B(net5073));
 sg13g2_o21ai_1 _12519_ (.B1(_03570_),
    .Y(_00486_),
    .A1(net5527),
    .A2(net5072));
 sg13g2_nand2_1 _12520_ (.Y(_03571_),
    .A(net2269),
    .B(net5072));
 sg13g2_o21ai_1 _12521_ (.B1(_03571_),
    .Y(_00487_),
    .A1(net5571),
    .A2(net5072));
 sg13g2_nand2_1 _12522_ (.Y(_03572_),
    .A(net2378),
    .B(net5072));
 sg13g2_o21ai_1 _12523_ (.B1(_03572_),
    .Y(_00488_),
    .A1(net5617),
    .A2(net5072));
 sg13g2_nand2_1 _12524_ (.Y(_03573_),
    .A(net2254),
    .B(_03567_));
 sg13g2_o21ai_1 _12525_ (.B1(_03573_),
    .Y(_00489_),
    .A1(net5670),
    .A2(net5072));
 sg13g2_nand2_1 _12526_ (.Y(_03574_),
    .A(net3261),
    .B(net5073));
 sg13g2_o21ai_1 _12527_ (.B1(_03574_),
    .Y(_00490_),
    .A1(net5717),
    .A2(net5073));
 sg13g2_nand2_1 _12528_ (.Y(_03575_),
    .A(net2812),
    .B(net5072));
 sg13g2_o21ai_1 _12529_ (.B1(_03575_),
    .Y(_00491_),
    .A1(net5762),
    .A2(net5072));
 sg13g2_nand2_1 _12530_ (.Y(_03576_),
    .A(net5235),
    .B(net5217));
 sg13g2_nand2_1 _12531_ (.Y(_03577_),
    .A(net2142),
    .B(_03576_));
 sg13g2_o21ai_1 _12532_ (.B1(_03577_),
    .Y(_00492_),
    .A1(net5426),
    .A2(net5071));
 sg13g2_nand2_1 _12533_ (.Y(_03578_),
    .A(net2183),
    .B(net5070));
 sg13g2_o21ai_1 _12534_ (.B1(_03578_),
    .Y(_00493_),
    .A1(net5471),
    .A2(net5070));
 sg13g2_nand2_1 _12535_ (.Y(_03579_),
    .A(net2881),
    .B(net5071));
 sg13g2_o21ai_1 _12536_ (.B1(_03579_),
    .Y(_00494_),
    .A1(net5517),
    .A2(net5071));
 sg13g2_nand2_1 _12537_ (.Y(_03580_),
    .A(net3352),
    .B(net5071));
 sg13g2_o21ai_1 _12538_ (.B1(_03580_),
    .Y(_00495_),
    .A1(net5560),
    .A2(net5071));
 sg13g2_nor2_1 _12539_ (.A(\mem.data_in[4] ),
    .B(net5070),
    .Y(_03581_));
 sg13g2_a21oi_1 _12540_ (.A1(_02860_),
    .A2(net5070),
    .Y(_00496_),
    .B1(_03581_));
 sg13g2_nand2_1 _12541_ (.Y(_03582_),
    .A(net3185),
    .B(net5071));
 sg13g2_o21ai_1 _12542_ (.B1(_03582_),
    .Y(_00497_),
    .A1(net5652),
    .A2(net5071));
 sg13g2_nor2_1 _12543_ (.A(\mem.data_in[6] ),
    .B(net5070),
    .Y(_03583_));
 sg13g2_a21oi_1 _12544_ (.A1(_02871_),
    .A2(net5070),
    .Y(_00498_),
    .B1(_03583_));
 sg13g2_nand2_1 _12545_ (.Y(_03584_),
    .A(net2793),
    .B(net5070));
 sg13g2_o21ai_1 _12546_ (.B1(_03584_),
    .Y(_00499_),
    .A1(net5743),
    .A2(net5070));
 sg13g2_nand2_1 _12547_ (.Y(_03585_),
    .A(net5253),
    .B(net5217));
 sg13g2_nand2_1 _12548_ (.Y(_03586_),
    .A(net2259),
    .B(net5068));
 sg13g2_o21ai_1 _12549_ (.B1(_03586_),
    .Y(_00500_),
    .A1(net5424),
    .A2(net5068));
 sg13g2_nand2_1 _12550_ (.Y(_03587_),
    .A(net3224),
    .B(net5068));
 sg13g2_o21ai_1 _12551_ (.B1(_03587_),
    .Y(_00501_),
    .A1(net5468),
    .A2(net5068));
 sg13g2_nand2_1 _12552_ (.Y(_03588_),
    .A(net2372),
    .B(net5069));
 sg13g2_o21ai_1 _12553_ (.B1(_03588_),
    .Y(_00502_),
    .A1(net5513),
    .A2(_03585_));
 sg13g2_nand2_1 _12554_ (.Y(_03589_),
    .A(net2426),
    .B(net5069));
 sg13g2_o21ai_1 _12555_ (.B1(_03589_),
    .Y(_00503_),
    .A1(net5558),
    .A2(net5069));
 sg13g2_nand2_1 _12556_ (.Y(_03590_),
    .A(net3493),
    .B(net5069));
 sg13g2_o21ai_1 _12557_ (.B1(_03590_),
    .Y(_00504_),
    .A1(net5606),
    .A2(net5069));
 sg13g2_nand2_1 _12558_ (.Y(_03591_),
    .A(net2520),
    .B(net5069));
 sg13g2_o21ai_1 _12559_ (.B1(_03591_),
    .Y(_00505_),
    .A1(net5649),
    .A2(net5069));
 sg13g2_nand2_1 _12560_ (.Y(_03592_),
    .A(net3125),
    .B(net5068));
 sg13g2_o21ai_1 _12561_ (.B1(_03592_),
    .Y(_00506_),
    .A1(net5696),
    .A2(net5068));
 sg13g2_nand2_1 _12562_ (.Y(_03593_),
    .A(net2480),
    .B(net5068));
 sg13g2_o21ai_1 _12563_ (.B1(_03593_),
    .Y(_00507_),
    .A1(net5741),
    .A2(net5068));
 sg13g2_nor2_1 _12564_ (.A(net5155),
    .B(_03375_),
    .Y(_03594_));
 sg13g2_nor2_1 _12565_ (.A(net3616),
    .B(net4760),
    .Y(_03595_));
 sg13g2_a21oi_1 _12566_ (.A1(net5424),
    .A2(net4760),
    .Y(_00508_),
    .B1(_03595_));
 sg13g2_nor2_1 _12567_ (.A(net3526),
    .B(net4761),
    .Y(_03596_));
 sg13g2_a21oi_1 _12568_ (.A1(net5469),
    .A2(net4761),
    .Y(_00509_),
    .B1(_03596_));
 sg13g2_nor2_1 _12569_ (.A(net3714),
    .B(net4761),
    .Y(_03597_));
 sg13g2_a21oi_1 _12570_ (.A1(net5515),
    .A2(net4761),
    .Y(_00510_),
    .B1(_03597_));
 sg13g2_nor2_1 _12571_ (.A(net4013),
    .B(net4761),
    .Y(_03598_));
 sg13g2_a21oi_1 _12572_ (.A1(net5559),
    .A2(net4761),
    .Y(_00511_),
    .B1(_03598_));
 sg13g2_nor2_1 _12573_ (.A(net3676),
    .B(net4761),
    .Y(_03599_));
 sg13g2_a21oi_1 _12574_ (.A1(net5605),
    .A2(net4761),
    .Y(_00512_),
    .B1(_03599_));
 sg13g2_nor2_1 _12575_ (.A(net2912),
    .B(net4760),
    .Y(_03600_));
 sg13g2_a21oi_1 _12576_ (.A1(net5650),
    .A2(net4760),
    .Y(_00513_),
    .B1(_03600_));
 sg13g2_nor2_1 _12577_ (.A(net3785),
    .B(net4760),
    .Y(_03601_));
 sg13g2_a21oi_1 _12578_ (.A1(net5696),
    .A2(net4760),
    .Y(_00514_),
    .B1(_03601_));
 sg13g2_nor2_1 _12579_ (.A(net2829),
    .B(net4760),
    .Y(_03602_));
 sg13g2_a21oi_1 _12580_ (.A1(net5741),
    .A2(net4760),
    .Y(_00515_),
    .B1(_03602_));
 sg13g2_nand2_1 _12581_ (.Y(_03603_),
    .A(_03079_),
    .B(net5217));
 sg13g2_nand2_1 _12582_ (.Y(_03604_),
    .A(net2786),
    .B(net5065));
 sg13g2_o21ai_1 _12583_ (.B1(_03604_),
    .Y(_00516_),
    .A1(net5425),
    .A2(net5065));
 sg13g2_nand2_1 _12584_ (.Y(_03605_),
    .A(net2455),
    .B(net5065));
 sg13g2_o21ai_1 _12585_ (.B1(_03605_),
    .Y(_00517_),
    .A1(net5470),
    .A2(net5065));
 sg13g2_nand2_1 _12586_ (.Y(_03606_),
    .A(net2322),
    .B(net5066));
 sg13g2_o21ai_1 _12587_ (.B1(_03606_),
    .Y(_00518_),
    .A1(net5513),
    .A2(net5065));
 sg13g2_nand2_1 _12588_ (.Y(_03607_),
    .A(net2207),
    .B(net5066));
 sg13g2_o21ai_1 _12589_ (.B1(_03607_),
    .Y(_00519_),
    .A1(net5558),
    .A2(net5066));
 sg13g2_nand2_1 _12590_ (.Y(_03608_),
    .A(net3066),
    .B(net5067));
 sg13g2_o21ai_1 _12591_ (.B1(_03608_),
    .Y(_00520_),
    .A1(net5606),
    .A2(net5067));
 sg13g2_nand2_1 _12592_ (.Y(_03609_),
    .A(net2556),
    .B(net5066));
 sg13g2_o21ai_1 _12593_ (.B1(_03609_),
    .Y(_00521_),
    .A1(net5649),
    .A2(net5065));
 sg13g2_nand2_1 _12594_ (.Y(_03610_),
    .A(net2245),
    .B(net5067));
 sg13g2_o21ai_1 _12595_ (.B1(_03610_),
    .Y(_00522_),
    .A1(net5697),
    .A2(net5067));
 sg13g2_nand2_1 _12596_ (.Y(_03611_),
    .A(net2848),
    .B(net5065));
 sg13g2_o21ai_1 _12597_ (.B1(_03611_),
    .Y(_00523_),
    .A1(net5741),
    .A2(net5065));
 sg13g2_nor2_1 _12598_ (.A(net5142),
    .B(_03109_),
    .Y(_03612_));
 sg13g2_nor2_1 _12599_ (.A(net2771),
    .B(net4758),
    .Y(_03613_));
 sg13g2_a21oi_1 _12600_ (.A1(net5436),
    .A2(net4758),
    .Y(_00524_),
    .B1(_03613_));
 sg13g2_nor2_1 _12601_ (.A(net4049),
    .B(net4759),
    .Y(_03614_));
 sg13g2_a21oi_1 _12602_ (.A1(net5483),
    .A2(net4759),
    .Y(_00525_),
    .B1(_03614_));
 sg13g2_nor2_1 _12603_ (.A(net4115),
    .B(net4759),
    .Y(_03615_));
 sg13g2_a21oi_1 _12604_ (.A1(net5527),
    .A2(net4759),
    .Y(_00526_),
    .B1(_03615_));
 sg13g2_nor2_1 _12605_ (.A(net3916),
    .B(net4758),
    .Y(_03616_));
 sg13g2_a21oi_1 _12606_ (.A1(net5571),
    .A2(net4758),
    .Y(_00527_),
    .B1(_03616_));
 sg13g2_nor2_1 _12607_ (.A(net3888),
    .B(net4758),
    .Y(_03617_));
 sg13g2_a21oi_1 _12608_ (.A1(net5617),
    .A2(net4758),
    .Y(_00528_),
    .B1(_03617_));
 sg13g2_nor2_1 _12609_ (.A(net3879),
    .B(net4759),
    .Y(_03618_));
 sg13g2_a21oi_1 _12610_ (.A1(net5670),
    .A2(net4759),
    .Y(_00529_),
    .B1(_03618_));
 sg13g2_nor2_1 _12611_ (.A(net3600),
    .B(net4758),
    .Y(_03619_));
 sg13g2_a21oi_1 _12612_ (.A1(net5717),
    .A2(net4758),
    .Y(_00530_),
    .B1(_03619_));
 sg13g2_nor2_1 _12613_ (.A(net3477),
    .B(net4759),
    .Y(_03620_));
 sg13g2_a21oi_1 _12614_ (.A1(net5762),
    .A2(net4759),
    .Y(_00531_),
    .B1(_03620_));
 sg13g2_nor2_1 _12615_ (.A(net5155),
    .B(_03212_),
    .Y(_03621_));
 sg13g2_nor2_1 _12616_ (.A(net3730),
    .B(net4756),
    .Y(_03622_));
 sg13g2_a21oi_1 _12617_ (.A1(net5424),
    .A2(net4756),
    .Y(_00532_),
    .B1(_03622_));
 sg13g2_nor2_1 _12618_ (.A(net3928),
    .B(net4757),
    .Y(_03623_));
 sg13g2_a21oi_1 _12619_ (.A1(net5468),
    .A2(net4757),
    .Y(_00533_),
    .B1(_03623_));
 sg13g2_nor2_1 _12620_ (.A(net3393),
    .B(net4757),
    .Y(_03624_));
 sg13g2_a21oi_1 _12621_ (.A1(net5513),
    .A2(net4757),
    .Y(_00534_),
    .B1(_03624_));
 sg13g2_nor2_1 _12622_ (.A(net3328),
    .B(net4757),
    .Y(_03625_));
 sg13g2_a21oi_1 _12623_ (.A1(net5561),
    .A2(net4757),
    .Y(_00535_),
    .B1(_03625_));
 sg13g2_nor2_1 _12624_ (.A(net3594),
    .B(net4757),
    .Y(_03626_));
 sg13g2_a21oi_1 _12625_ (.A1(net5605),
    .A2(net4757),
    .Y(_00536_),
    .B1(_03626_));
 sg13g2_nor2_1 _12626_ (.A(net3724),
    .B(net4756),
    .Y(_03627_));
 sg13g2_a21oi_1 _12627_ (.A1(net5650),
    .A2(net4756),
    .Y(_00537_),
    .B1(_03627_));
 sg13g2_nor2_1 _12628_ (.A(net4064),
    .B(net4756),
    .Y(_03628_));
 sg13g2_a21oi_1 _12629_ (.A1(net5696),
    .A2(net4756),
    .Y(_00538_),
    .B1(_03628_));
 sg13g2_nor2_1 _12630_ (.A(net3762),
    .B(net4756),
    .Y(_03629_));
 sg13g2_a21oi_1 _12631_ (.A1(net5745),
    .A2(net4756),
    .Y(_00539_),
    .B1(_03629_));
 sg13g2_nand2_1 _12632_ (.Y(_03630_),
    .A(net5217),
    .B(net5248));
 sg13g2_nand2_1 _12633_ (.Y(_03631_),
    .A(net3583),
    .B(net5063));
 sg13g2_o21ai_1 _12634_ (.B1(_03631_),
    .Y(_00540_),
    .A1(net5425),
    .A2(net5063));
 sg13g2_nand2_1 _12635_ (.Y(_03632_),
    .A(net2420),
    .B(net5063));
 sg13g2_o21ai_1 _12636_ (.B1(_03632_),
    .Y(_00541_),
    .A1(net5470),
    .A2(net5063));
 sg13g2_nand2_1 _12637_ (.Y(_03633_),
    .A(net2377),
    .B(net5064));
 sg13g2_o21ai_1 _12638_ (.B1(_03633_),
    .Y(_00542_),
    .A1(net5516),
    .A2(_03630_));
 sg13g2_nand2_1 _12639_ (.Y(_03634_),
    .A(net2351),
    .B(net5064));
 sg13g2_o21ai_1 _12640_ (.B1(_03634_),
    .Y(_00543_),
    .A1(net5558),
    .A2(net5064));
 sg13g2_nand2_1 _12641_ (.Y(_03635_),
    .A(net2387),
    .B(net5064));
 sg13g2_o21ai_1 _12642_ (.B1(_03635_),
    .Y(_00544_),
    .A1(net5606),
    .A2(net5063));
 sg13g2_nand2_1 _12643_ (.Y(_03636_),
    .A(net2788),
    .B(net5064));
 sg13g2_o21ai_1 _12644_ (.B1(_03636_),
    .Y(_00545_),
    .A1(net5649),
    .A2(net5064));
 sg13g2_nand2_1 _12645_ (.Y(_03637_),
    .A(net3056),
    .B(net5063));
 sg13g2_o21ai_1 _12646_ (.B1(_03637_),
    .Y(_00546_),
    .A1(net5697),
    .A2(net5063));
 sg13g2_nand2_1 _12647_ (.Y(_03638_),
    .A(net2534),
    .B(net5064));
 sg13g2_o21ai_1 _12648_ (.B1(_03638_),
    .Y(_00547_),
    .A1(net5741),
    .A2(net5063));
 sg13g2_nor2_2 _12649_ (.A(_02941_),
    .B(_03212_),
    .Y(_03639_));
 sg13g2_nor3_1 _12650_ (.A(_02880_),
    .B(_02941_),
    .C(_03212_),
    .Y(_03640_));
 sg13g2_mux4_1 _12651_ (.S0(net6080),
    .A0(\mem.mem[0][0] ),
    .A1(\mem.mem[1][0] ),
    .A2(\mem.mem[2][0] ),
    .A3(\mem.mem[3][0] ),
    .S1(net5937),
    .X(_03641_));
 sg13g2_mux2_1 _12652_ (.A0(\mem.mem[4][0] ),
    .A1(\mem.mem[5][0] ),
    .S(net6075),
    .X(_03642_));
 sg13g2_nand2_1 _12653_ (.Y(_03643_),
    .A(net5356),
    .B(_03642_));
 sg13g2_mux2_1 _12654_ (.A0(\mem.mem[6][0] ),
    .A1(\mem.mem[7][0] ),
    .S(net6074),
    .X(_03644_));
 sg13g2_a21oi_1 _12655_ (.A1(net5934),
    .A2(_03644_),
    .Y(_03645_),
    .B1(net5320));
 sg13g2_a21oi_1 _12656_ (.A1(_03643_),
    .A2(_03645_),
    .Y(_03646_),
    .B1(net5836));
 sg13g2_o21ai_1 _12657_ (.B1(_03646_),
    .Y(_03647_),
    .A1(net5862),
    .A2(_03641_));
 sg13g2_mux4_1 _12658_ (.S0(net6083),
    .A0(\mem.mem[8][0] ),
    .A1(\mem.mem[9][0] ),
    .A2(\mem.mem[10][0] ),
    .A3(\mem.mem[11][0] ),
    .S1(net5939),
    .X(_03648_));
 sg13g2_nand2b_1 _12659_ (.Y(_03649_),
    .B(net5319),
    .A_N(_03648_));
 sg13g2_mux2_1 _12660_ (.A0(\mem.mem[12][0] ),
    .A1(\mem.mem[13][0] ),
    .S(net6109),
    .X(_03650_));
 sg13g2_nand2_1 _12661_ (.Y(_03651_),
    .A(net5364),
    .B(_03650_));
 sg13g2_mux2_1 _12662_ (.A0(\mem.mem[14][0] ),
    .A1(\mem.mem[15][0] ),
    .S(net6109),
    .X(_03652_));
 sg13g2_a21oi_1 _12663_ (.A1(net5958),
    .A2(_03652_),
    .Y(_03653_),
    .B1(net5329));
 sg13g2_a21oi_1 _12664_ (.A1(_03651_),
    .A2(_03653_),
    .Y(_03654_),
    .B1(net5283));
 sg13g2_a21oi_1 _12665_ (.A1(_03649_),
    .A2(_03654_),
    .Y(_03655_),
    .B1(net5820));
 sg13g2_nor2b_1 _12666_ (.A(\mem.mem[23][0] ),
    .B_N(net6125),
    .Y(_03656_));
 sg13g2_o21ai_1 _12667_ (.B1(net5966),
    .Y(_03657_),
    .A1(net6125),
    .A2(\mem.mem[22][0] ));
 sg13g2_mux2_1 _12668_ (.A0(\mem.mem[20][0] ),
    .A1(\mem.mem[21][0] ),
    .S(net6125),
    .X(_03658_));
 sg13g2_o21ai_1 _12669_ (.B1(net5873),
    .Y(_03659_),
    .A1(_03656_),
    .A2(_03657_));
 sg13g2_a21oi_1 _12670_ (.A1(net5363),
    .A2(_03658_),
    .Y(_03660_),
    .B1(_03659_));
 sg13g2_mux2_1 _12671_ (.A0(\mem.mem[18][0] ),
    .A1(\mem.mem[19][0] ),
    .S(net6123),
    .X(_03661_));
 sg13g2_nand2b_1 _12672_ (.Y(_03662_),
    .B(net6121),
    .A_N(\mem.mem[17][0] ));
 sg13g2_a21oi_1 _12673_ (.A1(net5406),
    .A2(_02885_),
    .Y(_03663_),
    .B1(net5966));
 sg13g2_a221oi_1 _12674_ (.B2(_03663_),
    .C1(net5871),
    .B1(_03662_),
    .A1(net5966),
    .Y(_03664_),
    .A2(_03661_));
 sg13g2_or3_2 _12675_ (.A(net5840),
    .B(_03660_),
    .C(_03664_),
    .X(_03665_));
 sg13g2_mux4_1 _12676_ (.S0(net6125),
    .A0(\mem.mem[24][0] ),
    .A1(\mem.mem[25][0] ),
    .A2(\mem.mem[26][0] ),
    .A3(\mem.mem[27][0] ),
    .S1(net5968),
    .X(_03666_));
 sg13g2_nand2b_1 _12677_ (.Y(_03667_),
    .B(net5333),
    .A_N(_03666_));
 sg13g2_mux2_1 _12678_ (.A0(\mem.mem[28][0] ),
    .A1(\mem.mem[29][0] ),
    .S(net6151),
    .X(_03668_));
 sg13g2_nand2_1 _12679_ (.Y(_03669_),
    .A(net5367),
    .B(_03668_));
 sg13g2_mux2_1 _12680_ (.A0(\mem.mem[30][0] ),
    .A1(\mem.mem[31][0] ),
    .S(net6152),
    .X(_03670_));
 sg13g2_a21oi_1 _12681_ (.A1(net5987),
    .A2(_03670_),
    .Y(_03671_),
    .B1(net5340));
 sg13g2_a21oi_2 _12682_ (.B1(net5295),
    .Y(_03672_),
    .A2(_03671_),
    .A1(_03669_));
 sg13g2_a21oi_2 _12683_ (.B1(net5274),
    .Y(_03673_),
    .A2(_03672_),
    .A1(_03667_));
 sg13g2_a221oi_1 _12684_ (.B2(_03673_),
    .C1(net5815),
    .B1(_03665_),
    .A1(_03647_),
    .Y(_03674_),
    .A2(_03655_));
 sg13g2_nand2b_1 _12685_ (.Y(_03675_),
    .B(net6162),
    .A_N(\mem.mem[45][0] ));
 sg13g2_o21ai_1 _12686_ (.B1(_03675_),
    .Y(_03676_),
    .A1(net6165),
    .A2(\mem.mem[44][0] ));
 sg13g2_mux2_1 _12687_ (.A0(\mem.mem[46][0] ),
    .A1(\mem.mem[47][0] ),
    .S(net6165),
    .X(_03677_));
 sg13g2_a21oi_1 _12688_ (.A1(net5998),
    .A2(_03677_),
    .Y(_03678_),
    .B1(net5344));
 sg13g2_o21ai_1 _12689_ (.B1(_03678_),
    .Y(_03679_),
    .A1(net5998),
    .A2(_03676_));
 sg13g2_mux4_1 _12690_ (.S0(net6166),
    .A0(\mem.mem[40][0] ),
    .A1(\mem.mem[41][0] ),
    .A2(\mem.mem[42][0] ),
    .A3(\mem.mem[43][0] ),
    .S1(net5999),
    .X(_03680_));
 sg13g2_o21ai_1 _12691_ (.B1(net5847),
    .Y(_03681_),
    .A1(net5881),
    .A2(_03680_));
 sg13g2_inv_1 _12692_ (.Y(_03682_),
    .A(_03681_));
 sg13g2_mux4_1 _12693_ (.S0(net6167),
    .A0(\mem.mem[32][0] ),
    .A1(\mem.mem[33][0] ),
    .A2(\mem.mem[34][0] ),
    .A3(\mem.mem[35][0] ),
    .S1(net6000),
    .X(_03683_));
 sg13g2_nand2b_1 _12694_ (.Y(_03684_),
    .B(net5345),
    .A_N(_03683_));
 sg13g2_mux2_1 _12695_ (.A0(\mem.mem[36][0] ),
    .A1(\mem.mem[37][0] ),
    .S(net6152),
    .X(_03685_));
 sg13g2_nand2_1 _12696_ (.Y(_03686_),
    .A(net5367),
    .B(_03685_));
 sg13g2_mux2_1 _12697_ (.A0(\mem.mem[38][0] ),
    .A1(\mem.mem[39][0] ),
    .S(net6162),
    .X(_03687_));
 sg13g2_a21oi_1 _12698_ (.A1(net5995),
    .A2(_03687_),
    .Y(_03688_),
    .B1(net5344));
 sg13g2_a21oi_1 _12699_ (.A1(_03686_),
    .A2(_03688_),
    .Y(_03689_),
    .B1(net5847));
 sg13g2_a221oi_1 _12700_ (.B2(_03689_),
    .C1(net5824),
    .B1(_03684_),
    .A1(_03679_),
    .Y(_03690_),
    .A2(_03682_));
 sg13g2_mux2_1 _12701_ (.A0(\mem.mem[58][0] ),
    .A1(\mem.mem[59][0] ),
    .S(net6030),
    .X(_03691_));
 sg13g2_nand2_1 _12702_ (.Y(_03692_),
    .A(net5903),
    .B(_03691_));
 sg13g2_mux2_1 _12703_ (.A0(\mem.mem[56][0] ),
    .A1(\mem.mem[57][0] ),
    .S(net6030),
    .X(_03693_));
 sg13g2_a21oi_1 _12704_ (.A1(net5350),
    .A2(_03693_),
    .Y(_03694_),
    .B1(net5854));
 sg13g2_mux2_1 _12705_ (.A0(\mem.mem[60][0] ),
    .A1(\mem.mem[61][0] ),
    .S(net6033),
    .X(_03695_));
 sg13g2_nor2_1 _12706_ (.A(net6033),
    .B(\mem.mem[62][0] ),
    .Y(_03696_));
 sg13g2_o21ai_1 _12707_ (.B1(net5906),
    .Y(_03697_),
    .A1(net5378),
    .A2(\mem.mem[63][0] ));
 sg13g2_a21oi_1 _12708_ (.A1(net5350),
    .A2(_03695_),
    .Y(_03698_),
    .B1(net5309));
 sg13g2_o21ai_1 _12709_ (.B1(_03698_),
    .Y(_03699_),
    .A1(_03696_),
    .A2(_03697_));
 sg13g2_a21oi_1 _12710_ (.A1(_03692_),
    .A2(_03694_),
    .Y(_03700_),
    .B1(net5279));
 sg13g2_mux4_1 _12711_ (.S0(net6010),
    .A0(\mem.mem[48][0] ),
    .A1(\mem.mem[49][0] ),
    .A2(\mem.mem[50][0] ),
    .A3(\mem.mem[51][0] ),
    .S1(net5889),
    .X(_03701_));
 sg13g2_nand2b_2 _12712_ (.Y(_03702_),
    .B(net5299),
    .A_N(_03701_));
 sg13g2_mux2_1 _12713_ (.A0(\mem.mem[52][0] ),
    .A1(\mem.mem[53][0] ),
    .S(net6030),
    .X(_03703_));
 sg13g2_nand2_1 _12714_ (.Y(_03704_),
    .A(net5350),
    .B(_03703_));
 sg13g2_mux2_1 _12715_ (.A0(\mem.mem[54][0] ),
    .A1(\mem.mem[55][0] ),
    .S(net6030),
    .X(_03705_));
 sg13g2_a21oi_1 _12716_ (.A1(net5903),
    .A2(_03705_),
    .Y(_03706_),
    .B1(net5304));
 sg13g2_a21oi_1 _12717_ (.A1(_03704_),
    .A2(_03706_),
    .Y(_03707_),
    .B1(net5829));
 sg13g2_a221oi_1 _12718_ (.B2(_03707_),
    .C1(net5270),
    .B1(_03702_),
    .A1(_03699_),
    .Y(_03708_),
    .A2(_03700_));
 sg13g2_nor3_1 _12719_ (.A(net5264),
    .B(_03690_),
    .C(_03708_),
    .Y(_03709_));
 sg13g2_or3_1 _12720_ (.A(net5808),
    .B(_03674_),
    .C(_03709_),
    .X(_03710_));
 sg13g2_mux2_1 _12721_ (.A0(\mem.mem[74][0] ),
    .A1(\mem.mem[75][0] ),
    .S(net6017),
    .X(_03711_));
 sg13g2_nand2_1 _12722_ (.Y(_03712_),
    .A(net5894),
    .B(_03711_));
 sg13g2_mux2_1 _12723_ (.A0(\mem.mem[72][0] ),
    .A1(\mem.mem[73][0] ),
    .S(net6017),
    .X(_03713_));
 sg13g2_a21oi_1 _12724_ (.A1(net5348),
    .A2(_03713_),
    .Y(_03714_),
    .B1(net5852));
 sg13g2_mux2_1 _12725_ (.A0(\mem.mem[76][0] ),
    .A1(\mem.mem[77][0] ),
    .S(net6022),
    .X(_03715_));
 sg13g2_nor2_1 _12726_ (.A(net6022),
    .B(\mem.mem[78][0] ),
    .Y(_03716_));
 sg13g2_o21ai_1 _12727_ (.B1(net5897),
    .Y(_03717_),
    .A1(net5374),
    .A2(\mem.mem[79][0] ));
 sg13g2_a21oi_1 _12728_ (.A1(net5349),
    .A2(_03715_),
    .Y(_03718_),
    .B1(net5309));
 sg13g2_o21ai_1 _12729_ (.B1(_03718_),
    .Y(_03719_),
    .A1(_03716_),
    .A2(_03717_));
 sg13g2_a21oi_1 _12730_ (.A1(_03712_),
    .A2(_03714_),
    .Y(_03720_),
    .B1(net5276));
 sg13g2_nand2b_1 _12731_ (.Y(_03721_),
    .B(net6019),
    .A_N(\mem.mem[71][0] ));
 sg13g2_o21ai_1 _12732_ (.B1(_03721_),
    .Y(_03722_),
    .A1(net6019),
    .A2(\mem.mem[70][0] ));
 sg13g2_mux2_1 _12733_ (.A0(\mem.mem[68][0] ),
    .A1(\mem.mem[69][0] ),
    .S(net6017),
    .X(_03723_));
 sg13g2_a21oi_1 _12734_ (.A1(net5348),
    .A2(_03723_),
    .Y(_03724_),
    .B1(net5302));
 sg13g2_o21ai_1 _12735_ (.B1(_03724_),
    .Y(_03725_),
    .A1(net5348),
    .A2(_03722_));
 sg13g2_mux2_1 _12736_ (.A0(\mem.mem[66][0] ),
    .A1(\mem.mem[67][0] ),
    .S(net6018),
    .X(_03726_));
 sg13g2_nand2_1 _12737_ (.Y(_03727_),
    .A(net5895),
    .B(_03726_));
 sg13g2_mux2_1 _12738_ (.A0(\mem.mem[64][0] ),
    .A1(\mem.mem[65][0] ),
    .S(net6016),
    .X(_03728_));
 sg13g2_a21oi_1 _12739_ (.A1(net5348),
    .A2(_03728_),
    .Y(_03729_),
    .B1(net5852));
 sg13g2_a21oi_1 _12740_ (.A1(_03727_),
    .A2(_03729_),
    .Y(_03730_),
    .B1(net5828));
 sg13g2_a221oi_1 _12741_ (.B2(_03730_),
    .C1(net5816),
    .B1(_03725_),
    .A1(_03719_),
    .Y(_03731_),
    .A2(_03720_));
 sg13g2_mux4_1 _12742_ (.S0(net6005),
    .A0(\mem.mem[80][0] ),
    .A1(\mem.mem[81][0] ),
    .A2(\mem.mem[82][0] ),
    .A3(\mem.mem[83][0] ),
    .S1(net5885),
    .X(_03732_));
 sg13g2_nor2_1 _12743_ (.A(net5850),
    .B(_03732_),
    .Y(_03733_));
 sg13g2_mux2_1 _12744_ (.A0(\mem.mem[86][0] ),
    .A1(\mem.mem[87][0] ),
    .S(net6005),
    .X(_03734_));
 sg13g2_nand2_1 _12745_ (.Y(_03735_),
    .A(net5885),
    .B(_03734_));
 sg13g2_mux2_1 _12746_ (.A0(\mem.mem[84][0] ),
    .A1(\mem.mem[85][0] ),
    .S(net6005),
    .X(_03736_));
 sg13g2_a21oi_1 _12747_ (.A1(net5349),
    .A2(_03736_),
    .Y(_03737_),
    .B1(net5298));
 sg13g2_a21oi_2 _12748_ (.B1(_03733_),
    .Y(_03738_),
    .A2(_03737_),
    .A1(_03735_));
 sg13g2_mux4_1 _12749_ (.S0(net6018),
    .A0(\mem.mem[88][0] ),
    .A1(\mem.mem[89][0] ),
    .A2(\mem.mem[90][0] ),
    .A3(\mem.mem[91][0] ),
    .S1(net5895),
    .X(_03739_));
 sg13g2_nand2b_1 _12750_ (.Y(_03740_),
    .B(net5302),
    .A_N(_03739_));
 sg13g2_mux2_1 _12751_ (.A0(\mem.mem[92][0] ),
    .A1(\mem.mem[93][0] ),
    .S(net6019),
    .X(_03741_));
 sg13g2_nand2_1 _12752_ (.Y(_03742_),
    .A(net5348),
    .B(_03741_));
 sg13g2_mux2_1 _12753_ (.A0(\mem.mem[94][0] ),
    .A1(\mem.mem[95][0] ),
    .S(net6024),
    .X(_03743_));
 sg13g2_a21oi_1 _12754_ (.A1(net5899),
    .A2(_03743_),
    .Y(_03744_),
    .B1(net5302));
 sg13g2_a21oi_1 _12755_ (.A1(_03742_),
    .A2(_03744_),
    .Y(_03745_),
    .B1(net5276));
 sg13g2_a221oi_1 _12756_ (.B2(_03745_),
    .C1(net5270),
    .B1(_03740_),
    .A1(net5276),
    .Y(_03746_),
    .A2(_03738_));
 sg13g2_nor3_2 _12757_ (.A(net5810),
    .B(_03731_),
    .C(_03746_),
    .Y(_03747_));
 sg13g2_mux2_1 _12758_ (.A0(\mem.mem[108][0] ),
    .A1(\mem.mem[109][0] ),
    .S(net6065),
    .X(_03748_));
 sg13g2_nand2_1 _12759_ (.Y(_03749_),
    .A(net5355),
    .B(_03748_));
 sg13g2_mux2_1 _12760_ (.A0(\mem.mem[110][0] ),
    .A1(\mem.mem[111][0] ),
    .S(net6074),
    .X(_03750_));
 sg13g2_a21oi_1 _12761_ (.A1(net5925),
    .A2(_03750_),
    .Y(_03751_),
    .B1(net5315));
 sg13g2_mux4_1 _12762_ (.S0(net6065),
    .A0(\mem.mem[104][0] ),
    .A1(\mem.mem[105][0] ),
    .A2(\mem.mem[106][0] ),
    .A3(\mem.mem[107][0] ),
    .S1(net5925),
    .X(_03752_));
 sg13g2_o21ai_1 _12763_ (.B1(net5833),
    .Y(_03753_),
    .A1(net5861),
    .A2(_03752_));
 sg13g2_a21oi_2 _12764_ (.B1(_03753_),
    .Y(_03754_),
    .A2(_03751_),
    .A1(_03749_));
 sg13g2_a21oi_1 _12765_ (.A1(net5390),
    .A2(_02886_),
    .Y(_03755_),
    .B1(net5355));
 sg13g2_o21ai_1 _12766_ (.B1(_03755_),
    .Y(_03756_),
    .A1(net5390),
    .A2(\mem.mem[103][0] ));
 sg13g2_mux2_1 _12767_ (.A0(\mem.mem[100][0] ),
    .A1(\mem.mem[101][0] ),
    .S(net6072),
    .X(_03757_));
 sg13g2_a21oi_1 _12768_ (.A1(net5355),
    .A2(_03757_),
    .Y(_03758_),
    .B1(net5317));
 sg13g2_mux2_1 _12769_ (.A0(\mem.mem[98][0] ),
    .A1(\mem.mem[99][0] ),
    .S(net6072),
    .X(_03759_));
 sg13g2_nand2_1 _12770_ (.Y(_03760_),
    .A(net5930),
    .B(_03759_));
 sg13g2_mux2_1 _12771_ (.A0(\mem.mem[96][0] ),
    .A1(\mem.mem[97][0] ),
    .S(net6072),
    .X(_03761_));
 sg13g2_a21oi_1 _12772_ (.A1(net5355),
    .A2(_03761_),
    .Y(_03762_),
    .B1(net5861));
 sg13g2_a221oi_1 _12773_ (.B2(_03762_),
    .C1(net5834),
    .B1(_03760_),
    .A1(_03756_),
    .Y(_03763_),
    .A2(_03758_));
 sg13g2_nor3_1 _12774_ (.A(net5820),
    .B(_03754_),
    .C(_03763_),
    .Y(_03764_));
 sg13g2_a21oi_1 _12775_ (.A1(net5383),
    .A2(_02887_),
    .Y(_03765_),
    .B1(net5350));
 sg13g2_o21ai_1 _12776_ (.B1(_03765_),
    .Y(_03766_),
    .A1(net5380),
    .A2(\mem.mem[119][0] ));
 sg13g2_mux2_1 _12777_ (.A0(\mem.mem[116][0] ),
    .A1(\mem.mem[117][0] ),
    .S(net6064),
    .X(_03767_));
 sg13g2_a21oi_1 _12778_ (.A1(net5351),
    .A2(_03767_),
    .Y(_03768_),
    .B1(net5306));
 sg13g2_mux2_1 _12779_ (.A0(\mem.mem[114][0] ),
    .A1(\mem.mem[115][0] ),
    .S(net6064),
    .X(_03769_));
 sg13g2_nand2_1 _12780_ (.Y(_03770_),
    .A(net5927),
    .B(_03769_));
 sg13g2_mux2_1 _12781_ (.A0(\mem.mem[112][0] ),
    .A1(\mem.mem[113][0] ),
    .S(net6064),
    .X(_03771_));
 sg13g2_a21oi_1 _12782_ (.A1(net5350),
    .A2(_03771_),
    .Y(_03772_),
    .B1(net5861));
 sg13g2_a221oi_1 _12783_ (.B2(_03772_),
    .C1(net5833),
    .B1(_03770_),
    .A1(_03766_),
    .Y(_03773_),
    .A2(_03768_));
 sg13g2_mux4_1 _12784_ (.S0(net6068),
    .A0(\mem.mem[120][0] ),
    .A1(\mem.mem[121][0] ),
    .A2(\mem.mem[122][0] ),
    .A3(\mem.mem[123][0] ),
    .S1(net5928),
    .X(_03774_));
 sg13g2_nor2_1 _12785_ (.A(net5864),
    .B(_03774_),
    .Y(_03775_));
 sg13g2_nor2b_1 _12786_ (.A(\mem.mem[125][0] ),
    .B_N(net6038),
    .Y(_03776_));
 sg13g2_nor2_1 _12787_ (.A(net6039),
    .B(\mem.mem[124][0] ),
    .Y(_03777_));
 sg13g2_nor3_1 _12788_ (.A(net5912),
    .B(_03776_),
    .C(_03777_),
    .Y(_03778_));
 sg13g2_nor2b_1 _12789_ (.A(\mem.mem[127][0] ),
    .B_N(net6038),
    .Y(_03779_));
 sg13g2_o21ai_1 _12790_ (.B1(net5912),
    .Y(_03780_),
    .A1(net6039),
    .A2(\mem.mem[126][0] ));
 sg13g2_o21ai_1 _12791_ (.B1(net5856),
    .Y(_03781_),
    .A1(_03779_),
    .A2(_03780_));
 sg13g2_o21ai_1 _12792_ (.B1(net5830),
    .Y(_03782_),
    .A1(_03778_),
    .A2(_03781_));
 sg13g2_o21ai_1 _12793_ (.B1(net5818),
    .Y(_03783_),
    .A1(_03775_),
    .A2(_03782_));
 sg13g2_o21ai_1 _12794_ (.B1(net5809),
    .Y(_03784_),
    .A1(_03773_),
    .A2(_03783_));
 sg13g2_nor2_1 _12795_ (.A(_03764_),
    .B(_03784_),
    .Y(_03785_));
 sg13g2_nand2b_1 _12796_ (.Y(_03786_),
    .B(net5808),
    .A_N(_03747_));
 sg13g2_o21ai_1 _12797_ (.B1(_03710_),
    .Y(_03787_),
    .A1(_03785_),
    .A2(_03786_));
 sg13g2_nand2_1 _12798_ (.Y(_03788_),
    .A(net5407),
    .B(\mem.mem[132][0] ));
 sg13g2_a21oi_1 _12799_ (.A1(net6118),
    .A2(\mem.mem[133][0] ),
    .Y(_03789_),
    .B1(net5964));
 sg13g2_and2_1 _12800_ (.A(net6118),
    .B(\mem.mem[135][0] ),
    .X(_03790_));
 sg13g2_a21oi_1 _12801_ (.A1(net5405),
    .A2(\mem.mem[134][0] ),
    .Y(_03791_),
    .B1(_03790_));
 sg13g2_a221oi_1 _12802_ (.B2(net5964),
    .C1(net5332),
    .B1(_03791_),
    .A1(_03788_),
    .Y(_03792_),
    .A2(_03789_));
 sg13g2_nand2_1 _12803_ (.Y(_03793_),
    .A(net5405),
    .B(\mem.mem[128][0] ));
 sg13g2_a21oi_1 _12804_ (.A1(net6116),
    .A2(\mem.mem[129][0] ),
    .Y(_03794_),
    .B1(net5965));
 sg13g2_nor2b_1 _12805_ (.A(net6117),
    .B_N(\mem.mem[130][0] ),
    .Y(_03795_));
 sg13g2_a21oi_1 _12806_ (.A1(net6117),
    .A2(\mem.mem[131][0] ),
    .Y(_03796_),
    .B1(_03795_));
 sg13g2_a221oi_1 _12807_ (.B2(net5965),
    .C1(net5872),
    .B1(_03796_),
    .A1(_03793_),
    .Y(_03797_),
    .A2(_03794_));
 sg13g2_o21ai_1 _12808_ (.B1(net5291),
    .Y(_03798_),
    .A1(_03792_),
    .A2(_03797_));
 sg13g2_nor2b_1 _12809_ (.A(net6114),
    .B_N(\mem.mem[142][0] ),
    .Y(_03799_));
 sg13g2_a21oi_1 _12810_ (.A1(net6114),
    .A2(\mem.mem[143][0] ),
    .Y(_03800_),
    .B1(_03799_));
 sg13g2_nand2_1 _12811_ (.Y(_03801_),
    .A(net5404),
    .B(\mem.mem[140][0] ));
 sg13g2_a21oi_1 _12812_ (.A1(net6122),
    .A2(\mem.mem[141][0] ),
    .Y(_03802_),
    .B1(net5959));
 sg13g2_a221oi_1 _12813_ (.B2(_03802_),
    .C1(net5330),
    .B1(_03801_),
    .A1(net5959),
    .Y(_03803_),
    .A2(_03800_));
 sg13g2_nand2_1 _12814_ (.Y(_03804_),
    .A(net5406),
    .B(\mem.mem[136][0] ));
 sg13g2_a21oi_1 _12815_ (.A1(net6122),
    .A2(\mem.mem[137][0] ),
    .Y(_03805_),
    .B1(net5967));
 sg13g2_nor2b_1 _12816_ (.A(net6113),
    .B_N(\mem.mem[138][0] ),
    .Y(_03806_));
 sg13g2_a21oi_1 _12817_ (.A1(net6121),
    .A2(\mem.mem[139][0] ),
    .Y(_03807_),
    .B1(_03806_));
 sg13g2_a221oi_1 _12818_ (.B2(net5960),
    .C1(net5871),
    .B1(_03807_),
    .A1(_03804_),
    .Y(_03808_),
    .A2(_03805_));
 sg13g2_o21ai_1 _12819_ (.B1(net5842),
    .Y(_03809_),
    .A1(_03803_),
    .A2(_03808_));
 sg13g2_nand3_1 _12820_ (.B(_03798_),
    .C(_03809_),
    .A(net5271),
    .Y(_03810_));
 sg13g2_nor2b_1 _12821_ (.A(net6105),
    .B_N(\mem.mem[150][0] ),
    .Y(_03811_));
 sg13g2_a21oi_1 _12822_ (.A1(net6105),
    .A2(\mem.mem[151][0] ),
    .Y(_03812_),
    .B1(_03811_));
 sg13g2_nand2_1 _12823_ (.Y(_03813_),
    .A(net5392),
    .B(\mem.mem[148][0] ));
 sg13g2_a21oi_1 _12824_ (.A1(net6105),
    .A2(\mem.mem[149][0] ),
    .Y(_03814_),
    .B1(net5956));
 sg13g2_a221oi_1 _12825_ (.B2(_03814_),
    .C1(net5320),
    .B1(_03813_),
    .A1(net5956),
    .Y(_03815_),
    .A2(_03812_));
 sg13g2_nand2_1 _12826_ (.Y(_03816_),
    .A(net5392),
    .B(\mem.mem[144][0] ));
 sg13g2_a21oi_1 _12827_ (.A1(net6077),
    .A2(\mem.mem[145][0] ),
    .Y(_03817_),
    .B1(net5933));
 sg13g2_nor2b_1 _12828_ (.A(net6076),
    .B_N(\mem.mem[146][0] ),
    .Y(_03818_));
 sg13g2_a21oi_1 _12829_ (.A1(net6076),
    .A2(\mem.mem[147][0] ),
    .Y(_03819_),
    .B1(_03818_));
 sg13g2_a221oi_1 _12830_ (.B2(net5933),
    .C1(net5863),
    .B1(_03819_),
    .A1(_03816_),
    .Y(_03820_),
    .A2(_03817_));
 sg13g2_o21ai_1 _12831_ (.B1(net5283),
    .Y(_03821_),
    .A1(_03815_),
    .A2(_03820_));
 sg13g2_nand2_1 _12832_ (.Y(_03822_),
    .A(net6106),
    .B(\mem.mem[157][0] ));
 sg13g2_a21oi_1 _12833_ (.A1(net5402),
    .A2(\mem.mem[156][0] ),
    .Y(_03823_),
    .B1(net5955));
 sg13g2_and2_1 _12834_ (.A(net6106),
    .B(\mem.mem[159][0] ),
    .X(_03824_));
 sg13g2_a21oi_1 _12835_ (.A1(net5402),
    .A2(\mem.mem[158][0] ),
    .Y(_03825_),
    .B1(_03824_));
 sg13g2_a221oi_1 _12836_ (.B2(net5955),
    .C1(net5328),
    .B1(_03825_),
    .A1(_03822_),
    .Y(_03826_),
    .A2(_03823_));
 sg13g2_nand2_1 _12837_ (.Y(_03827_),
    .A(net5397),
    .B(\mem.mem[152][0] ));
 sg13g2_a21oi_1 _12838_ (.A1(net6092),
    .A2(\mem.mem[153][0] ),
    .Y(_03828_),
    .B1(net5955));
 sg13g2_nor2b_1 _12839_ (.A(net6091),
    .B_N(\mem.mem[154][0] ),
    .Y(_03829_));
 sg13g2_a21oi_1 _12840_ (.A1(net6091),
    .A2(\mem.mem[155][0] ),
    .Y(_03830_),
    .B1(_03829_));
 sg13g2_a221oi_1 _12841_ (.B2(net5946),
    .C1(net5866),
    .B1(_03830_),
    .A1(_03827_),
    .Y(_03831_),
    .A2(_03828_));
 sg13g2_o21ai_1 _12842_ (.B1(net5841),
    .Y(_03832_),
    .A1(_03826_),
    .A2(_03831_));
 sg13g2_nand3_1 _12843_ (.B(_03821_),
    .C(_03832_),
    .A(net5822),
    .Y(_03833_));
 sg13g2_nand3_1 _12844_ (.B(_03810_),
    .C(_03833_),
    .A(net5265),
    .Y(_03834_));
 sg13g2_mux4_1 _12845_ (.S0(net6056),
    .A0(\mem.mem[160][0] ),
    .A1(\mem.mem[161][0] ),
    .A2(\mem.mem[162][0] ),
    .A3(\mem.mem[163][0] ),
    .S1(net5920),
    .X(_03835_));
 sg13g2_a21o_1 _12846_ (.A2(\mem.mem[165][0] ),
    .A1(net6056),
    .B1(net5920),
    .X(_03836_));
 sg13g2_a21oi_1 _12847_ (.A1(net5387),
    .A2(\mem.mem[164][0] ),
    .Y(_03837_),
    .B1(_03836_));
 sg13g2_mux2_1 _12848_ (.A0(\mem.mem[166][0] ),
    .A1(\mem.mem[167][0] ),
    .S(net6060),
    .X(_03838_));
 sg13g2_o21ai_1 _12849_ (.B1(net5859),
    .Y(_03839_),
    .A1(net5353),
    .A2(_03838_));
 sg13g2_mux4_1 _12850_ (.S0(net6086),
    .A0(\mem.mem[168][0] ),
    .A1(\mem.mem[169][0] ),
    .A2(\mem.mem[170][0] ),
    .A3(\mem.mem[171][0] ),
    .S1(net5943),
    .X(_03840_));
 sg13g2_a21oi_1 _12851_ (.A1(net6090),
    .A2(\mem.mem[175][0] ),
    .Y(_03841_),
    .B1(net5360));
 sg13g2_o21ai_1 _12852_ (.B1(_03841_),
    .Y(_03842_),
    .A1(net6091),
    .A2(_02888_));
 sg13g2_nand2_1 _12853_ (.Y(_03843_),
    .A(net6090),
    .B(\mem.mem[173][0] ));
 sg13g2_a21oi_1 _12854_ (.A1(net5397),
    .A2(\mem.mem[172][0] ),
    .Y(_03844_),
    .B1(net5946));
 sg13g2_a21oi_1 _12855_ (.A1(_03843_),
    .A2(_03844_),
    .Y(_03845_),
    .B1(net5323));
 sg13g2_o21ai_1 _12856_ (.B1(net5285),
    .Y(_03846_),
    .A1(_03837_),
    .A2(_03839_));
 sg13g2_a21oi_2 _12857_ (.B1(_03846_),
    .Y(_03847_),
    .A2(_03835_),
    .A1(net5313));
 sg13g2_a221oi_1 _12858_ (.B2(_03845_),
    .C1(net5288),
    .B1(_03842_),
    .A1(net5323),
    .Y(_03848_),
    .A2(_03840_));
 sg13g2_o21ai_1 _12859_ (.B1(net5272),
    .Y(_03849_),
    .A1(_03847_),
    .A2(_03848_));
 sg13g2_mux4_1 _12860_ (.S0(net6132),
    .A0(\mem.mem[176][0] ),
    .A1(\mem.mem[177][0] ),
    .A2(\mem.mem[178][0] ),
    .A3(\mem.mem[179][0] ),
    .S1(net5973),
    .X(_03850_));
 sg13g2_and2_1 _12861_ (.A(net5335),
    .B(_03850_),
    .X(_03851_));
 sg13g2_nor2b_1 _12862_ (.A(net6135),
    .B_N(\mem.mem[182][0] ),
    .Y(_03852_));
 sg13g2_a21oi_1 _12863_ (.A1(net6135),
    .A2(\mem.mem[183][0] ),
    .Y(_03853_),
    .B1(_03852_));
 sg13g2_nand2_1 _12864_ (.Y(_03854_),
    .A(net5410),
    .B(\mem.mem[180][0] ));
 sg13g2_a21oi_1 _12865_ (.A1(net6135),
    .A2(\mem.mem[181][0] ),
    .Y(_03855_),
    .B1(net5976));
 sg13g2_a221oi_1 _12866_ (.B2(_03855_),
    .C1(net5336),
    .B1(_03854_),
    .A1(net5976),
    .Y(_03856_),
    .A2(_03853_));
 sg13g2_o21ai_1 _12867_ (.B1(net5292),
    .Y(_03857_),
    .A1(_03851_),
    .A2(_03856_));
 sg13g2_nand2_1 _12868_ (.Y(_03858_),
    .A(net6102),
    .B(\mem.mem[189][0] ));
 sg13g2_a21oi_1 _12869_ (.A1(net5400),
    .A2(\mem.mem[188][0] ),
    .Y(_03859_),
    .B1(net5954));
 sg13g2_and2_1 _12870_ (.A(net6102),
    .B(\mem.mem[191][0] ),
    .X(_03860_));
 sg13g2_a21oi_1 _12871_ (.A1(net5400),
    .A2(\mem.mem[190][0] ),
    .Y(_03861_),
    .B1(_03860_));
 sg13g2_a221oi_1 _12872_ (.B2(net5953),
    .C1(net5327),
    .B1(_03861_),
    .A1(_03858_),
    .Y(_03862_),
    .A2(_03859_));
 sg13g2_nand2_1 _12873_ (.Y(_03863_),
    .A(net5401),
    .B(\mem.mem[184][0] ));
 sg13g2_a21oi_1 _12874_ (.A1(net6097),
    .A2(\mem.mem[185][0] ),
    .Y(_03864_),
    .B1(net5950));
 sg13g2_nor2b_1 _12875_ (.A(net6096),
    .B_N(\mem.mem[186][0] ),
    .Y(_03865_));
 sg13g2_a21oi_1 _12876_ (.A1(net6097),
    .A2(\mem.mem[187][0] ),
    .Y(_03866_),
    .B1(_03865_));
 sg13g2_a221oi_1 _12877_ (.B2(net5950),
    .C1(net5868),
    .B1(_03866_),
    .A1(_03863_),
    .Y(_03867_),
    .A2(_03864_));
 sg13g2_o21ai_1 _12878_ (.B1(net5838),
    .Y(_03868_),
    .A1(_03862_),
    .A2(_03867_));
 sg13g2_nand3_1 _12879_ (.B(_03857_),
    .C(_03868_),
    .A(net5823),
    .Y(_03869_));
 sg13g2_nand3_1 _12880_ (.B(_03849_),
    .C(_03869_),
    .A(net5815),
    .Y(_03870_));
 sg13g2_mux4_1 _12881_ (.S0(net6053),
    .A0(\mem.mem[244][0] ),
    .A1(\mem.mem[245][0] ),
    .A2(\mem.mem[246][0] ),
    .A3(\mem.mem[247][0] ),
    .S1(net5918),
    .X(_03871_));
 sg13g2_mux4_1 _12882_ (.S0(net6048),
    .A0(\mem.mem[240][0] ),
    .A1(\mem.mem[241][0] ),
    .A2(\mem.mem[242][0] ),
    .A3(\mem.mem[243][0] ),
    .S1(net5915),
    .X(_03872_));
 sg13g2_mux4_1 _12883_ (.S0(net6053),
    .A0(\mem.mem[248][0] ),
    .A1(\mem.mem[249][0] ),
    .A2(\mem.mem[250][0] ),
    .A3(\mem.mem[251][0] ),
    .S1(net5918),
    .X(_03873_));
 sg13g2_a21o_2 _12884_ (.A2(_03870_),
    .A1(_03834_),
    .B1(net5807),
    .X(_03874_));
 sg13g2_nand2_1 _12885_ (.Y(_03875_),
    .A(net5399),
    .B(\mem.mem[198][0] ));
 sg13g2_a21oi_1 _12886_ (.A1(net6100),
    .A2(\mem.mem[199][0] ),
    .Y(_03876_),
    .B1(net5358));
 sg13g2_and2_1 _12887_ (.A(net6099),
    .B(\mem.mem[197][0] ),
    .X(_03877_));
 sg13g2_a21oi_1 _12888_ (.A1(net5399),
    .A2(\mem.mem[196][0] ),
    .Y(_03878_),
    .B1(_03877_));
 sg13g2_a221oi_1 _12889_ (.B2(net5358),
    .C1(net5325),
    .B1(_03878_),
    .A1(_03875_),
    .Y(_03879_),
    .A2(_03876_));
 sg13g2_nand2_1 _12890_ (.Y(_03880_),
    .A(net6099),
    .B(\mem.mem[193][0] ));
 sg13g2_nand2_1 _12891_ (.Y(_03881_),
    .A(net5399),
    .B(\mem.mem[192][0] ));
 sg13g2_nand3_1 _12892_ (.B(_03880_),
    .C(_03881_),
    .A(net5358),
    .Y(_03882_));
 sg13g2_and2_1 _12893_ (.A(net6100),
    .B(\mem.mem[195][0] ),
    .X(_03883_));
 sg13g2_a21oi_1 _12894_ (.A1(net5399),
    .A2(\mem.mem[194][0] ),
    .Y(_03884_),
    .B1(_03883_));
 sg13g2_a21oi_1 _12895_ (.A1(net5953),
    .A2(_03884_),
    .Y(_03885_),
    .B1(net5868));
 sg13g2_a21oi_1 _12896_ (.A1(_03882_),
    .A2(_03885_),
    .Y(_03886_),
    .B1(_03879_));
 sg13g2_mux4_1 _12897_ (.S0(net6087),
    .A0(\mem.mem[200][0] ),
    .A1(\mem.mem[201][0] ),
    .A2(\mem.mem[202][0] ),
    .A3(\mem.mem[203][0] ),
    .S1(net5944),
    .X(_03887_));
 sg13g2_nand2_1 _12898_ (.Y(_03888_),
    .A(net5324),
    .B(_03887_));
 sg13g2_nor2b_1 _12899_ (.A(net6099),
    .B_N(\mem.mem[206][0] ),
    .Y(_03889_));
 sg13g2_a21oi_1 _12900_ (.A1(net6099),
    .A2(\mem.mem[207][0] ),
    .Y(_03890_),
    .B1(_03889_));
 sg13g2_nand2_1 _12901_ (.Y(_03891_),
    .A(net6099),
    .B(\mem.mem[205][0] ));
 sg13g2_a21oi_1 _12902_ (.A1(net5399),
    .A2(\mem.mem[204][0] ),
    .Y(_03892_),
    .B1(net5947));
 sg13g2_a221oi_1 _12903_ (.B2(_03892_),
    .C1(net5323),
    .B1(_03891_),
    .A1(net5947),
    .Y(_03893_),
    .A2(_03890_));
 sg13g2_nor2_1 _12904_ (.A(net5287),
    .B(_03893_),
    .Y(_03894_));
 sg13g2_a221oi_1 _12905_ (.B2(_03894_),
    .C1(net5822),
    .B1(_03888_),
    .A1(net5287),
    .Y(_03895_),
    .A2(_03886_));
 sg13g2_nor2b_1 _12906_ (.A(net6161),
    .B_N(\mem.mem[222][0] ),
    .Y(_03896_));
 sg13g2_a21oi_1 _12907_ (.A1(net6161),
    .A2(\mem.mem[223][0] ),
    .Y(_03897_),
    .B1(_03896_));
 sg13g2_nand2_1 _12908_ (.Y(_03898_),
    .A(net6161),
    .B(\mem.mem[221][0] ));
 sg13g2_a21oi_1 _12909_ (.A1(net5419),
    .A2(\mem.mem[220][0] ),
    .Y(_03899_),
    .B1(net5995));
 sg13g2_a221oi_1 _12910_ (.B2(_03899_),
    .C1(net5344),
    .B1(_03898_),
    .A1(net5995),
    .Y(_03900_),
    .A2(_03897_));
 sg13g2_mux4_1 _12911_ (.S0(net6153),
    .A0(\mem.mem[216][0] ),
    .A1(\mem.mem[217][0] ),
    .A2(\mem.mem[218][0] ),
    .A3(\mem.mem[219][0] ),
    .S1(net5989),
    .X(_03901_));
 sg13g2_nand2_1 _12912_ (.Y(_03902_),
    .A(net5343),
    .B(_03901_));
 sg13g2_nor2_1 _12913_ (.A(net5296),
    .B(_03900_),
    .Y(_03903_));
 sg13g2_nor2b_1 _12914_ (.A(net6144),
    .B_N(\mem.mem[214][0] ),
    .Y(_03904_));
 sg13g2_a21oi_1 _12915_ (.A1(net6144),
    .A2(\mem.mem[215][0] ),
    .Y(_03905_),
    .B1(_03904_));
 sg13g2_mux2_1 _12916_ (.A0(\mem.mem[212][0] ),
    .A1(\mem.mem[213][0] ),
    .S(net6144),
    .X(_03906_));
 sg13g2_a21oi_1 _12917_ (.A1(net5982),
    .A2(_03905_),
    .Y(_03907_),
    .B1(net5338));
 sg13g2_o21ai_1 _12918_ (.B1(_03907_),
    .Y(_03908_),
    .A1(net5982),
    .A2(_03906_));
 sg13g2_nand2_1 _12919_ (.Y(_03909_),
    .A(net6162),
    .B(\mem.mem[209][0] ));
 sg13g2_nand2_1 _12920_ (.Y(_03910_),
    .A(net5419),
    .B(\mem.mem[208][0] ));
 sg13g2_nand3_1 _12921_ (.B(_03909_),
    .C(_03910_),
    .A(net5367),
    .Y(_03911_));
 sg13g2_and2_1 _12922_ (.A(net6162),
    .B(\mem.mem[211][0] ),
    .X(_03912_));
 sg13g2_a21oi_1 _12923_ (.A1(net5419),
    .A2(\mem.mem[210][0] ),
    .Y(_03913_),
    .B1(_03912_));
 sg13g2_a21oi_1 _12924_ (.A1(net5995),
    .A2(_03913_),
    .Y(_03914_),
    .B1(net5882));
 sg13g2_a21oi_1 _12925_ (.A1(_03911_),
    .A2(_03914_),
    .Y(_03915_),
    .B1(net5847));
 sg13g2_a221oi_1 _12926_ (.B2(_03915_),
    .C1(net5274),
    .B1(_03908_),
    .A1(_03902_),
    .Y(_03916_),
    .A2(_03903_));
 sg13g2_or3_2 _12927_ (.A(net5814),
    .B(_03895_),
    .C(_03916_),
    .X(_03917_));
 sg13g2_mux4_1 _12928_ (.S0(net6138),
    .A0(\mem.mem[224][0] ),
    .A1(\mem.mem[225][0] ),
    .A2(\mem.mem[226][0] ),
    .A3(\mem.mem[227][0] ),
    .S1(net5978),
    .X(_03918_));
 sg13g2_and2_1 _12929_ (.A(net5339),
    .B(_03918_),
    .X(_03919_));
 sg13g2_and2_1 _12930_ (.A(net6142),
    .B(\mem.mem[231][0] ),
    .X(_03920_));
 sg13g2_a21oi_1 _12931_ (.A1(net5413),
    .A2(\mem.mem[230][0] ),
    .Y(_03921_),
    .B1(_03920_));
 sg13g2_nand2_1 _12932_ (.Y(_03922_),
    .A(net6142),
    .B(\mem.mem[229][0] ));
 sg13g2_a21oi_1 _12933_ (.A1(net5413),
    .A2(\mem.mem[228][0] ),
    .Y(_03923_),
    .B1(net5981));
 sg13g2_a221oi_1 _12934_ (.B2(_03923_),
    .C1(net5338),
    .B1(_03922_),
    .A1(net5981),
    .Y(_03924_),
    .A2(_03921_));
 sg13g2_nor3_1 _12935_ (.A(net5843),
    .B(_03919_),
    .C(_03924_),
    .Y(_03925_));
 sg13g2_mux4_1 _12936_ (.S0(net6140),
    .A0(\mem.mem[232][0] ),
    .A1(\mem.mem[233][0] ),
    .A2(\mem.mem[234][0] ),
    .A3(\mem.mem[235][0] ),
    .S1(net5979),
    .X(_03926_));
 sg13g2_nand2_1 _12937_ (.Y(_03927_),
    .A(net6140),
    .B(\mem.mem[237][0] ));
 sg13g2_nand2_1 _12938_ (.Y(_03928_),
    .A(net5414),
    .B(\mem.mem[236][0] ));
 sg13g2_nand3_1 _12939_ (.B(_03927_),
    .C(_03928_),
    .A(net5365),
    .Y(_03929_));
 sg13g2_and2_1 _12940_ (.A(net6145),
    .B(\mem.mem[239][0] ),
    .X(_03930_));
 sg13g2_a21oi_1 _12941_ (.A1(net5412),
    .A2(\mem.mem[238][0] ),
    .Y(_03931_),
    .B1(_03930_));
 sg13g2_a21oi_1 _12942_ (.A1(net5983),
    .A2(_03931_),
    .Y(_03932_),
    .B1(net5337));
 sg13g2_a221oi_1 _12943_ (.B2(_03932_),
    .C1(net5293),
    .B1(_03929_),
    .A1(net5339),
    .Y(_03933_),
    .A2(_03926_));
 sg13g2_or3_2 _12944_ (.A(net5824),
    .B(_03925_),
    .C(_03933_),
    .X(_03934_));
 sg13g2_nand2_1 _12945_ (.Y(_03935_),
    .A(net5310),
    .B(_03872_));
 sg13g2_a21oi_1 _12946_ (.A1(net5860),
    .A2(_03871_),
    .Y(_03936_),
    .B1(net5831));
 sg13g2_nand2_1 _12947_ (.Y(_03937_),
    .A(net5860),
    .B(\mem.mem[252][0] ));
 sg13g2_a21oi_1 _12948_ (.A1(net5310),
    .A2(_03873_),
    .Y(_03938_),
    .B1(net5281));
 sg13g2_a221oi_1 _12949_ (.B2(_03938_),
    .C1(net5269),
    .B1(_03937_),
    .A1(_03935_),
    .Y(_03939_),
    .A2(_03936_));
 sg13g2_nor2_1 _12950_ (.A(net5264),
    .B(_03939_),
    .Y(_03940_));
 sg13g2_a21oi_1 _12951_ (.A1(_03934_),
    .A2(_03940_),
    .Y(_03941_),
    .B1(net5262));
 sg13g2_a21oi_1 _12952_ (.A1(_03917_),
    .A2(_03941_),
    .Y(_03942_),
    .B1(_02840_));
 sg13g2_a221oi_1 _12953_ (.B2(_03942_),
    .C1(_02944_),
    .B1(_03874_),
    .A1(_02840_),
    .Y(_03943_),
    .A2(_03787_));
 sg13g2_nor2_2 _12954_ (.A(_03640_),
    .B(_03943_),
    .Y(_03944_));
 sg13g2_o21ai_1 _12955_ (.B1(net6185),
    .Y(_03945_),
    .A1(net5787),
    .A2(net4183));
 sg13g2_a21oi_1 _12956_ (.A1(net5787),
    .A2(_03944_),
    .Y(_00548_),
    .B1(_03945_));
 sg13g2_o21ai_1 _12957_ (.B1(_02944_),
    .Y(_03946_),
    .A1(_02841_),
    .A2(_03015_));
 sg13g2_nand2b_1 _12958_ (.Y(_03947_),
    .B(net6032),
    .A_N(\mem.mem[57][1] ));
 sg13g2_a21oi_1 _12959_ (.A1(net5377),
    .A2(_02889_),
    .Y(_03948_),
    .B1(net5903));
 sg13g2_mux2_1 _12960_ (.A0(\mem.mem[58][1] ),
    .A1(\mem.mem[59][1] ),
    .S(net6029),
    .X(_03949_));
 sg13g2_a221oi_1 _12961_ (.B2(net5904),
    .C1(net5855),
    .B1(_03949_),
    .A1(_03947_),
    .Y(_03950_),
    .A2(_03948_));
 sg13g2_mux2_1 _12962_ (.A0(\mem.mem[60][1] ),
    .A1(\mem.mem[61][1] ),
    .S(net6031),
    .X(_03951_));
 sg13g2_nor2b_1 _12963_ (.A(\mem.mem[63][1] ),
    .B_N(net6031),
    .Y(_03952_));
 sg13g2_o21ai_1 _12964_ (.B1(net5905),
    .Y(_03953_),
    .A1(net6031),
    .A2(\mem.mem[62][1] ));
 sg13g2_o21ai_1 _12965_ (.B1(net5854),
    .Y(_03954_),
    .A1(_03952_),
    .A2(_03953_));
 sg13g2_a21oi_1 _12966_ (.A1(net5350),
    .A2(_03951_),
    .Y(_03955_),
    .B1(_03954_));
 sg13g2_mux2_1 _12967_ (.A0(\mem.mem[52][1] ),
    .A1(\mem.mem[53][1] ),
    .S(net6028),
    .X(_03956_));
 sg13g2_nor2b_1 _12968_ (.A(\mem.mem[55][1] ),
    .B_N(net6028),
    .Y(_03957_));
 sg13g2_o21ai_1 _12969_ (.B1(net5901),
    .Y(_03958_),
    .A1(net6028),
    .A2(\mem.mem[54][1] ));
 sg13g2_o21ai_1 _12970_ (.B1(net5854),
    .Y(_03959_),
    .A1(_03957_),
    .A2(_03958_));
 sg13g2_a21oi_1 _12971_ (.A1(net5350),
    .A2(_03956_),
    .Y(_03960_),
    .B1(_03959_));
 sg13g2_mux4_1 _12972_ (.S0(net6010),
    .A0(\mem.mem[48][1] ),
    .A1(\mem.mem[49][1] ),
    .A2(\mem.mem[50][1] ),
    .A3(\mem.mem[51][1] ),
    .S1(net5889),
    .X(_03961_));
 sg13g2_nor2_2 _12973_ (.A(net5851),
    .B(_03961_),
    .Y(_03962_));
 sg13g2_nor2b_1 _12974_ (.A(net6035),
    .B_N(\mem.mem[124][1] ),
    .Y(_03963_));
 sg13g2_a21oi_1 _12975_ (.A1(net6035),
    .A2(\mem.mem[125][1] ),
    .Y(_03964_),
    .B1(_03963_));
 sg13g2_mux2_1 _12976_ (.A0(\mem.mem[126][1] ),
    .A1(\mem.mem[127][1] ),
    .S(net6037),
    .X(_03965_));
 sg13g2_o21ai_1 _12977_ (.B1(net5855),
    .Y(_03966_),
    .A1(net5351),
    .A2(_03965_));
 sg13g2_a21o_1 _12978_ (.A2(_03964_),
    .A1(net5351),
    .B1(_03966_),
    .X(_03967_));
 sg13g2_mux4_1 _12979_ (.S0(net6040),
    .A0(\mem.mem[120][1] ),
    .A1(\mem.mem[121][1] ),
    .A2(\mem.mem[122][1] ),
    .A3(\mem.mem[123][1] ),
    .S1(net5910),
    .X(_03968_));
 sg13g2_a21oi_1 _12980_ (.A1(net5307),
    .A2(_03968_),
    .Y(_03969_),
    .B1(net5280));
 sg13g2_mux4_1 _12981_ (.S0(net6023),
    .A0(\mem.mem[112][1] ),
    .A1(\mem.mem[113][1] ),
    .A2(\mem.mem[114][1] ),
    .A3(\mem.mem[115][1] ),
    .S1(net5898),
    .X(_03970_));
 sg13g2_nand2_1 _12982_ (.Y(_03971_),
    .A(net5308),
    .B(_03970_));
 sg13g2_nand2_1 _12983_ (.Y(_03972_),
    .A(net6036),
    .B(\mem.mem[119][1] ));
 sg13g2_nand2b_1 _12984_ (.Y(_03973_),
    .B(\mem.mem[118][1] ),
    .A_N(net6036));
 sg13g2_nand3_1 _12985_ (.B(_03972_),
    .C(_03973_),
    .A(net5908),
    .Y(_03974_));
 sg13g2_nand2b_1 _12986_ (.Y(_03975_),
    .B(\mem.mem[116][1] ),
    .A_N(net6035));
 sg13g2_a21oi_1 _12987_ (.A1(net6035),
    .A2(\mem.mem[117][1] ),
    .Y(_03976_),
    .B1(net5909));
 sg13g2_a21oi_1 _12988_ (.A1(_03975_),
    .A2(_03976_),
    .Y(_03977_),
    .B1(net5306));
 sg13g2_a21oi_1 _12989_ (.A1(_03974_),
    .A2(_03977_),
    .Y(_03978_),
    .B1(net5830));
 sg13g2_a221oi_1 _12990_ (.B2(_03978_),
    .C1(net5270),
    .B1(_03971_),
    .A1(_03967_),
    .Y(_03979_),
    .A2(_03969_));
 sg13g2_mux4_1 _12991_ (.S0(net6072),
    .A0(\mem.mem[96][1] ),
    .A1(\mem.mem[97][1] ),
    .A2(\mem.mem[98][1] ),
    .A3(\mem.mem[99][1] ),
    .S1(net5930),
    .X(_03980_));
 sg13g2_nand2_1 _12992_ (.Y(_03981_),
    .A(net6066),
    .B(\mem.mem[103][1] ));
 sg13g2_nand2_1 _12993_ (.Y(_03982_),
    .A(net5388),
    .B(\mem.mem[102][1] ));
 sg13g2_nand3_1 _12994_ (.B(_03981_),
    .C(_03982_),
    .A(net5926),
    .Y(_03983_));
 sg13g2_nand2_1 _12995_ (.Y(_03984_),
    .A(net5388),
    .B(\mem.mem[100][1] ));
 sg13g2_a21oi_1 _12996_ (.A1(net6067),
    .A2(\mem.mem[101][1] ),
    .Y(_03985_),
    .B1(net5926));
 sg13g2_a21oi_1 _12997_ (.A1(_03984_),
    .A2(_03985_),
    .Y(_03986_),
    .B1(net5317));
 sg13g2_a221oi_1 _12998_ (.B2(_03986_),
    .C1(net5833),
    .B1(_03983_),
    .A1(net5315),
    .Y(_03987_),
    .A2(_03980_));
 sg13g2_nand2_1 _12999_ (.Y(_03988_),
    .A(net5385),
    .B(\mem.mem[108][1] ));
 sg13g2_a21oi_1 _13000_ (.A1(net6052),
    .A2(\mem.mem[109][1] ),
    .Y(_03989_),
    .B1(net5918));
 sg13g2_and2_1 _13001_ (.A(net6058),
    .B(\mem.mem[111][1] ),
    .X(_03990_));
 sg13g2_a21oi_1 _13002_ (.A1(net5387),
    .A2(\mem.mem[110][1] ),
    .Y(_03991_),
    .B1(_03990_));
 sg13g2_a221oi_1 _13003_ (.B2(net5918),
    .C1(net5311),
    .B1(_03991_),
    .A1(_03988_),
    .Y(_03992_),
    .A2(_03989_));
 sg13g2_nor2b_1 _13004_ (.A(net6052),
    .B_N(\mem.mem[104][1] ),
    .Y(_03993_));
 sg13g2_a21oi_1 _13005_ (.A1(net6052),
    .A2(\mem.mem[105][1] ),
    .Y(_03994_),
    .B1(_03993_));
 sg13g2_nand2_1 _13006_ (.Y(_03995_),
    .A(net5385),
    .B(\mem.mem[106][1] ));
 sg13g2_a21oi_1 _13007_ (.A1(net6052),
    .A2(\mem.mem[107][1] ),
    .Y(_03996_),
    .B1(net5354));
 sg13g2_a221oi_1 _13008_ (.B2(_03996_),
    .C1(net5857),
    .B1(_03995_),
    .A1(net5354),
    .Y(_03997_),
    .A2(_03994_));
 sg13g2_nor3_1 _13009_ (.A(net5281),
    .B(_03992_),
    .C(_03997_),
    .Y(_03998_));
 sg13g2_or3_1 _13010_ (.A(net5820),
    .B(_03987_),
    .C(_03998_),
    .X(_03999_));
 sg13g2_nor2_1 _13011_ (.A(net5264),
    .B(_03979_),
    .Y(_04000_));
 sg13g2_nand2_1 _13012_ (.Y(_04001_),
    .A(net5372),
    .B(\mem.mem[68][1] ));
 sg13g2_a21oi_1 _13013_ (.A1(net6018),
    .A2(\mem.mem[69][1] ),
    .Y(_04002_),
    .B1(net5895));
 sg13g2_and2_1 _13014_ (.A(net6018),
    .B(\mem.mem[71][1] ),
    .X(_04003_));
 sg13g2_a21oi_1 _13015_ (.A1(net5373),
    .A2(\mem.mem[70][1] ),
    .Y(_04004_),
    .B1(_04003_));
 sg13g2_a221oi_1 _13016_ (.B2(net5892),
    .C1(net5302),
    .B1(_04004_),
    .A1(_04001_),
    .Y(_04005_),
    .A2(_04002_));
 sg13g2_and2_1 _13017_ (.A(net6018),
    .B(\mem.mem[67][1] ),
    .X(_04006_));
 sg13g2_a21oi_1 _13018_ (.A1(net5373),
    .A2(\mem.mem[66][1] ),
    .Y(_04007_),
    .B1(_04006_));
 sg13g2_nand2_1 _13019_ (.Y(_04008_),
    .A(net5372),
    .B(\mem.mem[64][1] ));
 sg13g2_a21oi_1 _13020_ (.A1(net6018),
    .A2(\mem.mem[65][1] ),
    .Y(_04009_),
    .B1(net5893));
 sg13g2_a221oi_1 _13021_ (.B2(_04009_),
    .C1(net5852),
    .B1(_04008_),
    .A1(net5893),
    .Y(_04010_),
    .A2(_04007_));
 sg13g2_nor3_2 _13022_ (.A(net5828),
    .B(_04005_),
    .C(_04010_),
    .Y(_04011_));
 sg13g2_nand2_1 _13023_ (.Y(_04012_),
    .A(net5370),
    .B(\mem.mem[76][1] ));
 sg13g2_a21oi_1 _13024_ (.A1(net6013),
    .A2(\mem.mem[77][1] ),
    .Y(_04013_),
    .B1(net5890));
 sg13g2_and2_1 _13025_ (.A(net6013),
    .B(\mem.mem[79][1] ),
    .X(_04014_));
 sg13g2_a21oi_1 _13026_ (.A1(net5370),
    .A2(\mem.mem[78][1] ),
    .Y(_04015_),
    .B1(_04014_));
 sg13g2_a221oi_1 _13027_ (.B2(net5890),
    .C1(net5300),
    .B1(_04015_),
    .A1(_04012_),
    .Y(_04016_),
    .A2(_04013_));
 sg13g2_nor2b_1 _13028_ (.A(net6021),
    .B_N(\mem.mem[72][1] ),
    .Y(_04017_));
 sg13g2_a21oi_1 _13029_ (.A1(net6023),
    .A2(\mem.mem[73][1] ),
    .Y(_04018_),
    .B1(_04017_));
 sg13g2_nand2_1 _13030_ (.Y(_04019_),
    .A(net5374),
    .B(\mem.mem[74][1] ));
 sg13g2_a21oi_1 _13031_ (.A1(net6023),
    .A2(\mem.mem[75][1] ),
    .Y(_04020_),
    .B1(net5348));
 sg13g2_a221oi_1 _13032_ (.B2(_04020_),
    .C1(net5853),
    .B1(_04019_),
    .A1(net5348),
    .Y(_04021_),
    .A2(_04018_));
 sg13g2_nor3_1 _13033_ (.A(net5277),
    .B(_04016_),
    .C(_04021_),
    .Y(_04022_));
 sg13g2_or3_1 _13034_ (.A(net5816),
    .B(_04011_),
    .C(_04022_),
    .X(_04023_));
 sg13g2_nor2b_1 _13035_ (.A(net6047),
    .B_N(\mem.mem[88][1] ),
    .Y(_04024_));
 sg13g2_a21oi_1 _13036_ (.A1(net6047),
    .A2(\mem.mem[89][1] ),
    .Y(_04025_),
    .B1(_04024_));
 sg13g2_nand2_1 _13037_ (.Y(_04026_),
    .A(net5386),
    .B(\mem.mem[90][1] ));
 sg13g2_a21oi_1 _13038_ (.A1(net6047),
    .A2(\mem.mem[91][1] ),
    .Y(_04027_),
    .B1(net5348));
 sg13g2_a221oi_1 _13039_ (.B2(_04027_),
    .C1(net5857),
    .B1(_04026_),
    .A1(net5354),
    .Y(_04028_),
    .A2(_04025_));
 sg13g2_nand2_1 _13040_ (.Y(_04029_),
    .A(net5386),
    .B(\mem.mem[92][1] ));
 sg13g2_a21oi_1 _13041_ (.A1(net6046),
    .A2(\mem.mem[93][1] ),
    .Y(_04030_),
    .B1(net5916));
 sg13g2_and2_1 _13042_ (.A(net6051),
    .B(\mem.mem[95][1] ),
    .X(_04031_));
 sg13g2_a21oi_1 _13043_ (.A1(net5385),
    .A2(\mem.mem[94][1] ),
    .Y(_04032_),
    .B1(_04031_));
 sg13g2_a221oi_1 _13044_ (.B2(net5917),
    .C1(net5310),
    .B1(_04032_),
    .A1(_04029_),
    .Y(_04033_),
    .A2(_04030_));
 sg13g2_or3_1 _13045_ (.A(net5276),
    .B(_04028_),
    .C(_04033_),
    .X(_04034_));
 sg13g2_mux4_1 _13046_ (.S0(net6005),
    .A0(\mem.mem[80][1] ),
    .A1(\mem.mem[81][1] ),
    .A2(\mem.mem[82][1] ),
    .A3(\mem.mem[83][1] ),
    .S1(net5885),
    .X(_04035_));
 sg13g2_nand2_1 _13047_ (.Y(_04036_),
    .A(net6009),
    .B(\mem.mem[87][1] ));
 sg13g2_nand2b_1 _13048_ (.Y(_04037_),
    .B(\mem.mem[86][1] ),
    .A_N(net6009));
 sg13g2_nand3_1 _13049_ (.B(_04036_),
    .C(_04037_),
    .A(net5888),
    .Y(_04038_));
 sg13g2_nand2b_1 _13050_ (.Y(_04039_),
    .B(\mem.mem[84][1] ),
    .A_N(net6008));
 sg13g2_a21oi_1 _13051_ (.A1(net6009),
    .A2(\mem.mem[85][1] ),
    .Y(_04040_),
    .B1(net5888));
 sg13g2_a21oi_1 _13052_ (.A1(_04039_),
    .A2(_04040_),
    .Y(_04041_),
    .B1(net5299));
 sg13g2_a221oi_1 _13053_ (.B2(_04041_),
    .C1(net5827),
    .B1(_04038_),
    .A1(net5299),
    .Y(_04042_),
    .A2(_04035_));
 sg13g2_nor2_1 _13054_ (.A(net5270),
    .B(_04042_),
    .Y(_04043_));
 sg13g2_a21oi_1 _13055_ (.A1(_04034_),
    .A2(_04043_),
    .Y(_04044_),
    .B1(net5810));
 sg13g2_a221oi_1 _13056_ (.B2(_04044_),
    .C1(net5262),
    .B1(_04023_),
    .A1(_03999_),
    .Y(_04045_),
    .A2(_04000_));
 sg13g2_o21ai_1 _13057_ (.B1(net5279),
    .Y(_04046_),
    .A1(_03960_),
    .A2(_03962_));
 sg13g2_o21ai_1 _13058_ (.B1(net5829),
    .Y(_04047_),
    .A1(_03950_),
    .A2(_03955_));
 sg13g2_nand3_1 _13059_ (.B(_04046_),
    .C(_04047_),
    .A(net5817),
    .Y(_04048_));
 sg13g2_mux4_1 _13060_ (.S0(net6166),
    .A0(\mem.mem[36][1] ),
    .A1(\mem.mem[37][1] ),
    .A2(\mem.mem[38][1] ),
    .A3(\mem.mem[39][1] ),
    .S1(net5999),
    .X(_04049_));
 sg13g2_mux4_1 _13061_ (.S0(net6167),
    .A0(\mem.mem[32][1] ),
    .A1(\mem.mem[33][1] ),
    .A2(\mem.mem[34][1] ),
    .A3(\mem.mem[35][1] ),
    .S1(net6002),
    .X(_04050_));
 sg13g2_mux4_1 _13062_ (.S0(net6162),
    .A0(\mem.mem[44][1] ),
    .A1(\mem.mem[45][1] ),
    .A2(\mem.mem[46][1] ),
    .A3(\mem.mem[47][1] ),
    .S1(net5995),
    .X(_04051_));
 sg13g2_mux4_1 _13063_ (.S0(net6171),
    .A0(\mem.mem[40][1] ),
    .A1(\mem.mem[41][1] ),
    .A2(\mem.mem[42][1] ),
    .A3(\mem.mem[43][1] ),
    .S1(net6001),
    .X(_04052_));
 sg13g2_mux4_1 _13064_ (.S0(net5344),
    .A0(_04049_),
    .A1(_04050_),
    .A2(_04051_),
    .A3(_04052_),
    .S1(net5847),
    .X(_04053_));
 sg13g2_a21oi_2 _13065_ (.B1(net5265),
    .Y(_04054_),
    .A2(_04053_),
    .A1(net5271));
 sg13g2_mux4_1 _13066_ (.S0(net6080),
    .A0(\mem.mem[0][1] ),
    .A1(\mem.mem[1][1] ),
    .A2(\mem.mem[2][1] ),
    .A3(\mem.mem[3][1] ),
    .S1(net5937),
    .X(_04055_));
 sg13g2_nand2_1 _13067_ (.Y(_04056_),
    .A(net6074),
    .B(\mem.mem[7][1] ));
 sg13g2_nand2_1 _13068_ (.Y(_04057_),
    .A(net5391),
    .B(\mem.mem[6][1] ));
 sg13g2_nand3_1 _13069_ (.B(_04056_),
    .C(_04057_),
    .A(net5934),
    .Y(_04058_));
 sg13g2_nand2_1 _13070_ (.Y(_04059_),
    .A(net5392),
    .B(\mem.mem[4][1] ));
 sg13g2_a21oi_1 _13071_ (.A1(net6077),
    .A2(\mem.mem[5][1] ),
    .Y(_04060_),
    .B1(net5935));
 sg13g2_a21oi_1 _13072_ (.A1(_04059_),
    .A2(_04060_),
    .Y(_04061_),
    .B1(net5320));
 sg13g2_a221oi_1 _13073_ (.B2(_04061_),
    .C1(net5836),
    .B1(_04058_),
    .A1(net5318),
    .Y(_04062_),
    .A2(_04055_));
 sg13g2_nand2_1 _13074_ (.Y(_04063_),
    .A(net5394),
    .B(\mem.mem[12][1] ));
 sg13g2_a21oi_1 _13075_ (.A1(net6109),
    .A2(\mem.mem[13][1] ),
    .Y(_04064_),
    .B1(net5938));
 sg13g2_and2_1 _13076_ (.A(net6109),
    .B(\mem.mem[15][1] ),
    .X(_04065_));
 sg13g2_a21oi_1 _13077_ (.A1(net5403),
    .A2(\mem.mem[14][1] ),
    .Y(_04066_),
    .B1(_04065_));
 sg13g2_a221oi_1 _13078_ (.B2(net5938),
    .C1(net5318),
    .B1(_04066_),
    .A1(_04063_),
    .Y(_04067_),
    .A2(_04064_));
 sg13g2_nor2b_1 _13079_ (.A(net6081),
    .B_N(\mem.mem[8][1] ),
    .Y(_04068_));
 sg13g2_a21oi_1 _13080_ (.A1(net6081),
    .A2(\mem.mem[9][1] ),
    .Y(_04069_),
    .B1(_04068_));
 sg13g2_nand2_1 _13081_ (.Y(_04070_),
    .A(net5394),
    .B(\mem.mem[10][1] ));
 sg13g2_a21oi_1 _13082_ (.A1(net6081),
    .A2(\mem.mem[11][1] ),
    .Y(_04071_),
    .B1(net5356));
 sg13g2_a221oi_1 _13083_ (.B2(_04071_),
    .C1(net5862),
    .B1(_04070_),
    .A1(net5356),
    .Y(_04072_),
    .A2(_04069_));
 sg13g2_nor3_1 _13084_ (.A(net5284),
    .B(_04067_),
    .C(_04072_),
    .Y(_04073_));
 sg13g2_or3_1 _13085_ (.A(net5826),
    .B(_04062_),
    .C(_04073_),
    .X(_04074_));
 sg13g2_nor2b_1 _13086_ (.A(net6119),
    .B_N(\mem.mem[24][1] ),
    .Y(_04075_));
 sg13g2_a21oi_1 _13087_ (.A1(net6120),
    .A2(\mem.mem[25][1] ),
    .Y(_04076_),
    .B1(_04075_));
 sg13g2_nand2_1 _13088_ (.Y(_04077_),
    .A(net5405),
    .B(\mem.mem[26][1] ));
 sg13g2_a21oi_1 _13089_ (.A1(net6120),
    .A2(\mem.mem[27][1] ),
    .Y(_04078_),
    .B1(net5362));
 sg13g2_a221oi_1 _13090_ (.B2(_04078_),
    .C1(net5872),
    .B1(_04077_),
    .A1(net5362),
    .Y(_04079_),
    .A2(_04076_));
 sg13g2_nand2_1 _13091_ (.Y(_04080_),
    .A(net5415),
    .B(\mem.mem[28][1] ));
 sg13g2_a21oi_1 _13092_ (.A1(net6149),
    .A2(\mem.mem[29][1] ),
    .Y(_04081_),
    .B1(net5987));
 sg13g2_and2_1 _13093_ (.A(net6150),
    .B(\mem.mem[31][1] ),
    .X(_04082_));
 sg13g2_a21oi_1 _13094_ (.A1(net5415),
    .A2(\mem.mem[30][1] ),
    .Y(_04083_),
    .B1(_04082_));
 sg13g2_a221oi_1 _13095_ (.B2(net5987),
    .C1(net5340),
    .B1(_04083_),
    .A1(_04080_),
    .Y(_04084_),
    .A2(_04081_));
 sg13g2_or3_1 _13096_ (.A(net5290),
    .B(_04079_),
    .C(_04084_),
    .X(_04085_));
 sg13g2_nand2b_1 _13097_ (.Y(_04086_),
    .B(\mem.mem[20][1] ),
    .A_N(net6125));
 sg13g2_a21oi_1 _13098_ (.A1(net6125),
    .A2(\mem.mem[21][1] ),
    .Y(_04087_),
    .B1(net5968));
 sg13g2_mux2_1 _13099_ (.A0(\mem.mem[22][1] ),
    .A1(\mem.mem[23][1] ),
    .S(net6124),
    .X(_04088_));
 sg13g2_a21oi_1 _13100_ (.A1(_04086_),
    .A2(_04087_),
    .Y(_04089_),
    .B1(net5331));
 sg13g2_o21ai_1 _13101_ (.B1(_04089_),
    .Y(_04090_),
    .A1(net5363),
    .A2(_04088_));
 sg13g2_nand2_1 _13102_ (.Y(_04091_),
    .A(net6122),
    .B(\mem.mem[19][1] ));
 sg13g2_nand2b_1 _13103_ (.Y(_04092_),
    .B(\mem.mem[18][1] ),
    .A_N(net6123));
 sg13g2_nand3_1 _13104_ (.B(_04091_),
    .C(_04092_),
    .A(net5967),
    .Y(_04093_));
 sg13g2_nand2b_1 _13105_ (.Y(_04094_),
    .B(\mem.mem[16][1] ),
    .A_N(net6121));
 sg13g2_a21oi_1 _13106_ (.A1(net6123),
    .A2(\mem.mem[17][1] ),
    .Y(_04095_),
    .B1(net5966));
 sg13g2_a21oi_1 _13107_ (.A1(_04094_),
    .A2(_04095_),
    .Y(_04096_),
    .B1(net5871));
 sg13g2_a21oi_2 _13108_ (.B1(net5842),
    .Y(_04097_),
    .A2(_04096_),
    .A1(_04093_));
 sg13g2_a21oi_1 _13109_ (.A1(_04090_),
    .A2(_04097_),
    .Y(_04098_),
    .B1(net5271));
 sg13g2_a21oi_2 _13110_ (.B1(net5814),
    .Y(_04099_),
    .A2(_04098_),
    .A1(_04085_));
 sg13g2_a221oi_1 _13111_ (.B2(_04099_),
    .C1(net5807),
    .B1(_04074_),
    .A1(_04048_),
    .Y(_04100_),
    .A2(_04054_));
 sg13g2_o21ai_1 _13112_ (.B1(_02840_),
    .Y(_04101_),
    .A1(_04045_),
    .A2(_04100_));
 sg13g2_a21oi_1 _13113_ (.A1(net6113),
    .A2(\mem.mem[143][1] ),
    .Y(_04102_),
    .B1(net5364));
 sg13g2_o21ai_1 _13114_ (.B1(_04102_),
    .Y(_04103_),
    .A1(net6113),
    .A2(_02890_));
 sg13g2_nand2_1 _13115_ (.Y(_04104_),
    .A(net6112),
    .B(\mem.mem[141][1] ));
 sg13g2_a21oi_1 _13116_ (.A1(net5403),
    .A2(\mem.mem[140][1] ),
    .Y(_04105_),
    .B1(net5958));
 sg13g2_a21oi_1 _13117_ (.A1(_04104_),
    .A2(_04105_),
    .Y(_04106_),
    .B1(net5329));
 sg13g2_mux4_1 _13118_ (.S0(net6113),
    .A0(\mem.mem[136][1] ),
    .A1(\mem.mem[137][1] ),
    .A2(\mem.mem[138][1] ),
    .A3(\mem.mem[139][1] ),
    .S1(net5959),
    .X(_04107_));
 sg13g2_a221oi_1 _13119_ (.B2(net5330),
    .C1(net5290),
    .B1(_04107_),
    .A1(_04103_),
    .Y(_04108_),
    .A2(_04106_));
 sg13g2_nand2_1 _13120_ (.Y(_04109_),
    .A(net5405),
    .B(\mem.mem[128][1] ));
 sg13g2_a21oi_1 _13121_ (.A1(net6100),
    .A2(\mem.mem[129][1] ),
    .Y(_04110_),
    .B1(net5953));
 sg13g2_nor2b_1 _13122_ (.A(net6100),
    .B_N(\mem.mem[130][1] ),
    .Y(_04111_));
 sg13g2_a21oi_1 _13123_ (.A1(net6100),
    .A2(\mem.mem[131][1] ),
    .Y(_04112_),
    .B1(_04111_));
 sg13g2_a221oi_1 _13124_ (.B2(net5953),
    .C1(net5868),
    .B1(_04112_),
    .A1(_04109_),
    .Y(_04113_),
    .A2(_04110_));
 sg13g2_nand2_1 _13125_ (.Y(_04114_),
    .A(net5405),
    .B(\mem.mem[132][1] ));
 sg13g2_a21oi_1 _13126_ (.A1(net6102),
    .A2(\mem.mem[133][1] ),
    .Y(_04115_),
    .B1(net5963));
 sg13g2_nor2b_1 _13127_ (.A(net6102),
    .B_N(\mem.mem[134][1] ),
    .Y(_04116_));
 sg13g2_a21oi_1 _13128_ (.A1(net6102),
    .A2(\mem.mem[135][1] ),
    .Y(_04117_),
    .B1(_04116_));
 sg13g2_a221oi_1 _13129_ (.B2(net5953),
    .C1(net5325),
    .B1(_04117_),
    .A1(_04114_),
    .Y(_04118_),
    .A2(_04115_));
 sg13g2_nor3_2 _13130_ (.A(net5839),
    .B(_04113_),
    .C(_04118_),
    .Y(_04119_));
 sg13g2_o21ai_1 _13131_ (.B1(net5275),
    .Y(_04120_),
    .A1(_04108_),
    .A2(_04119_));
 sg13g2_and2_1 _13132_ (.A(net6092),
    .B(\mem.mem[157][1] ),
    .X(_04121_));
 sg13g2_a21oi_1 _13133_ (.A1(net5398),
    .A2(\mem.mem[156][1] ),
    .Y(_04122_),
    .B1(_04121_));
 sg13g2_mux2_1 _13134_ (.A0(\mem.mem[158][1] ),
    .A1(\mem.mem[159][1] ),
    .S(net6092),
    .X(_04123_));
 sg13g2_a21oi_1 _13135_ (.A1(net5948),
    .A2(_04123_),
    .Y(_04124_),
    .B1(net5323));
 sg13g2_o21ai_1 _13136_ (.B1(_04124_),
    .Y(_04125_),
    .A1(net5948),
    .A2(_04122_));
 sg13g2_mux4_1 _13137_ (.S0(net6093),
    .A0(\mem.mem[152][1] ),
    .A1(\mem.mem[153][1] ),
    .A2(\mem.mem[154][1] ),
    .A3(\mem.mem[155][1] ),
    .S1(net5947),
    .X(_04126_));
 sg13g2_o21ai_1 _13138_ (.B1(net5838),
    .Y(_04127_),
    .A1(net5866),
    .A2(_04126_));
 sg13g2_inv_1 _13139_ (.Y(_04128_),
    .A(_04127_));
 sg13g2_a21o_1 _13140_ (.A2(\mem.mem[149][1] ),
    .A1(net6106),
    .B1(net5956),
    .X(_04129_));
 sg13g2_a21oi_1 _13141_ (.A1(net5402),
    .A2(\mem.mem[148][1] ),
    .Y(_04130_),
    .B1(_04129_));
 sg13g2_mux2_1 _13142_ (.A0(\mem.mem[150][1] ),
    .A1(\mem.mem[151][1] ),
    .S(net6105),
    .X(_04131_));
 sg13g2_o21ai_1 _13143_ (.B1(net5869),
    .Y(_04132_),
    .A1(net5361),
    .A2(_04131_));
 sg13g2_mux4_1 _13144_ (.S0(net6076),
    .A0(\mem.mem[144][1] ),
    .A1(\mem.mem[145][1] ),
    .A2(\mem.mem[146][1] ),
    .A3(\mem.mem[147][1] ),
    .S1(net5933),
    .X(_04133_));
 sg13g2_nand2_1 _13145_ (.Y(_04134_),
    .A(net5320),
    .B(_04133_));
 sg13g2_o21ai_1 _13146_ (.B1(_04134_),
    .Y(_04135_),
    .A1(_04130_),
    .A2(_04132_));
 sg13g2_a22oi_1 _13147_ (.Y(_04136_),
    .B1(_04135_),
    .B2(net5287),
    .A2(_04128_),
    .A1(_04125_));
 sg13g2_a21oi_1 _13148_ (.A1(net5821),
    .A2(_04136_),
    .Y(_04137_),
    .B1(net5812));
 sg13g2_mux4_1 _13149_ (.S0(net6130),
    .A0(\mem.mem[184][1] ),
    .A1(\mem.mem[185][1] ),
    .A2(\mem.mem[186][1] ),
    .A3(\mem.mem[187][1] ),
    .S1(net5972),
    .X(_04138_));
 sg13g2_nand2_1 _13150_ (.Y(_04139_),
    .A(net5334),
    .B(_04138_));
 sg13g2_mux4_1 _13151_ (.S0(net6101),
    .A0(\mem.mem[188][1] ),
    .A1(\mem.mem[189][1] ),
    .A2(\mem.mem[190][1] ),
    .A3(\mem.mem[191][1] ),
    .S1(net5952),
    .X(_04140_));
 sg13g2_a21oi_1 _13152_ (.A1(net5876),
    .A2(_04140_),
    .Y(_04141_),
    .B1(net5292));
 sg13g2_mux4_1 _13153_ (.S0(net6130),
    .A0(\mem.mem[180][1] ),
    .A1(\mem.mem[181][1] ),
    .A2(\mem.mem[182][1] ),
    .A3(\mem.mem[183][1] ),
    .S1(net5974),
    .X(_04142_));
 sg13g2_nand2_1 _13154_ (.Y(_04143_),
    .A(net5875),
    .B(_04142_));
 sg13g2_mux4_1 _13155_ (.S0(net6130),
    .A0(\mem.mem[176][1] ),
    .A1(\mem.mem[177][1] ),
    .A2(\mem.mem[178][1] ),
    .A3(\mem.mem[179][1] ),
    .S1(net5972),
    .X(_04144_));
 sg13g2_a21oi_1 _13156_ (.A1(net5334),
    .A2(_04144_),
    .Y(_04145_),
    .B1(net5845));
 sg13g2_a221oi_1 _13157_ (.B2(_04145_),
    .C1(net5273),
    .B1(_04143_),
    .A1(_04139_),
    .Y(_04146_),
    .A2(_04141_));
 sg13g2_mux4_1 _13158_ (.S0(net6060),
    .A0(\mem.mem[172][1] ),
    .A1(\mem.mem[173][1] ),
    .A2(\mem.mem[174][1] ),
    .A3(\mem.mem[175][1] ),
    .S1(net5923),
    .X(_04147_));
 sg13g2_mux4_1 _13159_ (.S0(net6056),
    .A0(\mem.mem[168][1] ),
    .A1(\mem.mem[169][1] ),
    .A2(\mem.mem[170][1] ),
    .A3(\mem.mem[171][1] ),
    .S1(net5920),
    .X(_04148_));
 sg13g2_mux4_1 _13160_ (.S0(net6060),
    .A0(\mem.mem[164][1] ),
    .A1(\mem.mem[165][1] ),
    .A2(\mem.mem[166][1] ),
    .A3(\mem.mem[167][1] ),
    .S1(net5923),
    .X(_04149_));
 sg13g2_mux4_1 _13161_ (.S0(net6056),
    .A0(\mem.mem[160][1] ),
    .A1(\mem.mem[161][1] ),
    .A2(\mem.mem[162][1] ),
    .A3(\mem.mem[163][1] ),
    .S1(net5920),
    .X(_04150_));
 sg13g2_mux4_1 _13162_ (.S0(net5314),
    .A0(_04147_),
    .A1(_04148_),
    .A2(_04149_),
    .A3(_04150_),
    .S1(net5282),
    .X(_04151_));
 sg13g2_a21o_1 _13163_ (.A2(_04151_),
    .A1(net5272),
    .B1(_04146_),
    .X(_04152_));
 sg13g2_a221oi_1 _13164_ (.B2(net5812),
    .C1(net5807),
    .B1(_04152_),
    .A1(_04120_),
    .Y(_04153_),
    .A2(_04137_));
 sg13g2_nand2_1 _13165_ (.Y(_04154_),
    .A(net5396),
    .B(\mem.mem[202][1] ));
 sg13g2_a21oi_1 _13166_ (.A1(net6088),
    .A2(\mem.mem[203][1] ),
    .Y(_04155_),
    .B1(net5357));
 sg13g2_nand2_1 _13167_ (.Y(_04156_),
    .A(net5396),
    .B(\mem.mem[200][1] ));
 sg13g2_a21oi_1 _13168_ (.A1(net6088),
    .A2(\mem.mem[201][1] ),
    .Y(_04157_),
    .B1(net5945));
 sg13g2_a221oi_1 _13169_ (.B2(_04157_),
    .C1(net5865),
    .B1(_04156_),
    .A1(_04154_),
    .Y(_04158_),
    .A2(_04155_));
 sg13g2_nand2_1 _13170_ (.Y(_04159_),
    .A(net5398),
    .B(\mem.mem[204][1] ));
 sg13g2_a21oi_1 _13171_ (.A1(net6088),
    .A2(\mem.mem[205][1] ),
    .Y(_04160_),
    .B1(net5945));
 sg13g2_nand2_1 _13172_ (.Y(_04161_),
    .A(net5398),
    .B(\mem.mem[206][1] ));
 sg13g2_a21oi_1 _13173_ (.A1(net6088),
    .A2(\mem.mem[207][1] ),
    .Y(_04162_),
    .B1(net5357));
 sg13g2_a221oi_1 _13174_ (.B2(_04162_),
    .C1(net5324),
    .B1(_04161_),
    .A1(_04159_),
    .Y(_04163_),
    .A2(_04160_));
 sg13g2_o21ai_1 _13175_ (.B1(net5838),
    .Y(_04164_),
    .A1(_04158_),
    .A2(_04163_));
 sg13g2_mux4_1 _13176_ (.S0(net6101),
    .A0(\mem.mem[196][1] ),
    .A1(\mem.mem[197][1] ),
    .A2(\mem.mem[198][1] ),
    .A3(\mem.mem[199][1] ),
    .S1(net5952),
    .X(_04165_));
 sg13g2_mux4_1 _13177_ (.S0(net6095),
    .A0(\mem.mem[192][1] ),
    .A1(\mem.mem[193][1] ),
    .A2(\mem.mem[194][1] ),
    .A3(\mem.mem[195][1] ),
    .S1(net5951),
    .X(_04166_));
 sg13g2_nor2_1 _13178_ (.A(net5867),
    .B(_04166_),
    .Y(_04167_));
 sg13g2_nor2_1 _13179_ (.A(net5839),
    .B(_04167_),
    .Y(_04168_));
 sg13g2_o21ai_1 _13180_ (.B1(_04168_),
    .Y(_04169_),
    .A1(net5326),
    .A2(_04165_));
 sg13g2_nand3_1 _13181_ (.B(_04164_),
    .C(_04169_),
    .A(net5272),
    .Y(_04170_));
 sg13g2_mux4_1 _13182_ (.S0(net6146),
    .A0(\mem.mem[212][1] ),
    .A1(\mem.mem[213][1] ),
    .A2(\mem.mem[214][1] ),
    .A3(\mem.mem[215][1] ),
    .S1(net5984),
    .X(_04171_));
 sg13g2_mux4_1 _13183_ (.S0(net6163),
    .A0(\mem.mem[208][1] ),
    .A1(\mem.mem[209][1] ),
    .A2(\mem.mem[210][1] ),
    .A3(\mem.mem[211][1] ),
    .S1(net5996),
    .X(_04172_));
 sg13g2_mux2_2 _13184_ (.A0(_04171_),
    .A1(_04172_),
    .S(net5337),
    .X(_04173_));
 sg13g2_mux4_1 _13185_ (.S0(net6134),
    .A0(\mem.mem[216][1] ),
    .A1(\mem.mem[217][1] ),
    .A2(\mem.mem[218][1] ),
    .A3(\mem.mem[219][1] ),
    .S1(net5975),
    .X(_04174_));
 sg13g2_or2_1 _13186_ (.X(_04175_),
    .B(_04174_),
    .A(net5876));
 sg13g2_mux2_1 _13187_ (.A0(\mem.mem[222][1] ),
    .A1(\mem.mem[223][1] ),
    .S(net6154),
    .X(_04176_));
 sg13g2_nand2_2 _13188_ (.Y(_04177_),
    .A(net5989),
    .B(_04176_));
 sg13g2_mux2_1 _13189_ (.A0(\mem.mem[220][1] ),
    .A1(\mem.mem[221][1] ),
    .S(net6136),
    .X(_04178_));
 sg13g2_a21oi_1 _13190_ (.A1(net5366),
    .A2(_04178_),
    .Y(_04179_),
    .B1(net5335));
 sg13g2_a21oi_1 _13191_ (.A1(_04177_),
    .A2(_04179_),
    .Y(_04180_),
    .B1(net5294));
 sg13g2_a22oi_1 _13192_ (.Y(_04181_),
    .B1(_04175_),
    .B2(_04180_),
    .A2(_04173_),
    .A1(net5292));
 sg13g2_a21oi_1 _13193_ (.A1(net5821),
    .A2(_04181_),
    .Y(_04182_),
    .B1(net5813));
 sg13g2_nand2_1 _13194_ (.Y(_04183_),
    .A(net6140),
    .B(\mem.mem[233][1] ));
 sg13g2_a21oi_1 _13195_ (.A1(net5414),
    .A2(\mem.mem[232][1] ),
    .Y(_04184_),
    .B1(net5979));
 sg13g2_nor2b_1 _13196_ (.A(net6141),
    .B_N(\mem.mem[234][1] ),
    .Y(_04185_));
 sg13g2_a21oi_1 _13197_ (.A1(net6141),
    .A2(\mem.mem[235][1] ),
    .Y(_04186_),
    .B1(_04185_));
 sg13g2_a221oi_1 _13198_ (.B2(net5979),
    .C1(net5878),
    .B1(_04186_),
    .A1(_04183_),
    .Y(_04187_),
    .A2(_04184_));
 sg13g2_nand2_1 _13199_ (.Y(_04188_),
    .A(net6145),
    .B(\mem.mem[237][1] ));
 sg13g2_a21oi_1 _13200_ (.A1(net5412),
    .A2(\mem.mem[236][1] ),
    .Y(_04189_),
    .B1(net5983));
 sg13g2_nor2b_1 _13201_ (.A(net6145),
    .B_N(\mem.mem[238][1] ),
    .Y(_04190_));
 sg13g2_a21oi_1 _13202_ (.A1(net6145),
    .A2(\mem.mem[239][1] ),
    .Y(_04191_),
    .B1(_04190_));
 sg13g2_a221oi_1 _13203_ (.B2(net5983),
    .C1(net5337),
    .B1(_04191_),
    .A1(_04188_),
    .Y(_04192_),
    .A2(_04189_));
 sg13g2_nor3_2 _13204_ (.A(net5293),
    .B(_04187_),
    .C(_04192_),
    .Y(_04193_));
 sg13g2_mux4_1 _13205_ (.S0(net6133),
    .A0(\mem.mem[224][1] ),
    .A1(\mem.mem[225][1] ),
    .A2(\mem.mem[226][1] ),
    .A3(\mem.mem[227][1] ),
    .S1(net5973),
    .X(_04194_));
 sg13g2_mux4_1 _13206_ (.S0(net6139),
    .A0(\mem.mem[228][1] ),
    .A1(\mem.mem[229][1] ),
    .A2(\mem.mem[230][1] ),
    .A3(\mem.mem[231][1] ),
    .S1(net5980),
    .X(_04195_));
 sg13g2_a21o_1 _13207_ (.A2(_04195_),
    .A1(net5877),
    .B1(net5843),
    .X(_04196_));
 sg13g2_a21oi_1 _13208_ (.A1(net5335),
    .A2(_04194_),
    .Y(_04197_),
    .B1(_04196_));
 sg13g2_o21ai_1 _13209_ (.B1(net5273),
    .Y(_04198_),
    .A1(_04193_),
    .A2(_04197_));
 sg13g2_mux4_1 _13210_ (.S0(net6055),
    .A0(\mem.mem[240][1] ),
    .A1(\mem.mem[241][1] ),
    .A2(\mem.mem[242][1] ),
    .A3(\mem.mem[243][1] ),
    .S1(net5921),
    .X(_04199_));
 sg13g2_nor2_1 _13211_ (.A(net5859),
    .B(_04199_),
    .Y(_04200_));
 sg13g2_mux2_1 _13212_ (.A0(\mem.mem[244][1] ),
    .A1(\mem.mem[245][1] ),
    .S(net6058),
    .X(_04201_));
 sg13g2_nand2_1 _13213_ (.Y(_04202_),
    .A(net5354),
    .B(_04201_));
 sg13g2_mux2_1 _13214_ (.A0(\mem.mem[246][1] ),
    .A1(\mem.mem[247][1] ),
    .S(net6058),
    .X(_04203_));
 sg13g2_a21oi_1 _13215_ (.A1(net5922),
    .A2(_04203_),
    .Y(_04204_),
    .B1(net5314));
 sg13g2_a21oi_1 _13216_ (.A1(_04202_),
    .A2(_04204_),
    .Y(_04205_),
    .B1(_04200_));
 sg13g2_mux4_1 _13217_ (.S0(net6053),
    .A0(\mem.mem[248][1] ),
    .A1(\mem.mem[249][1] ),
    .A2(\mem.mem[250][1] ),
    .A3(\mem.mem[251][1] ),
    .S1(net5918),
    .X(_04206_));
 sg13g2_nor2_1 _13218_ (.A(net5858),
    .B(_04206_),
    .Y(_04207_));
 sg13g2_o21ai_1 _13219_ (.B1(net5832),
    .Y(_04208_),
    .A1(net5312),
    .A2(\mem.mem[252][1] ));
 sg13g2_o21ai_1 _13220_ (.B1(net5820),
    .Y(_04209_),
    .A1(_04207_),
    .A2(_04208_));
 sg13g2_a21oi_1 _13221_ (.A1(net5285),
    .A2(_04205_),
    .Y(_04210_),
    .B1(_04209_));
 sg13g2_nor2_2 _13222_ (.A(net5264),
    .B(_04210_),
    .Y(_04211_));
 sg13g2_a221oi_1 _13223_ (.B2(_04211_),
    .C1(net5263),
    .B1(_04198_),
    .A1(_04170_),
    .Y(_04212_),
    .A2(_04182_));
 sg13g2_or3_2 _13224_ (.A(_02840_),
    .B(_04153_),
    .C(_04212_),
    .X(_04213_));
 sg13g2_nand3_1 _13225_ (.B(_04101_),
    .C(_04213_),
    .A(_02945_),
    .Y(_04214_));
 sg13g2_nand2_2 _13226_ (.Y(_04215_),
    .A(_03946_),
    .B(_04214_));
 sg13g2_o21ai_1 _13227_ (.B1(net6183),
    .Y(_04216_),
    .A1(net5787),
    .A2(net4195));
 sg13g2_a21oi_1 _13228_ (.A1(net5787),
    .A2(_04215_),
    .Y(_00549_),
    .B1(_04216_));
 sg13g2_nand2_1 _13229_ (.Y(_04217_),
    .A(net5372),
    .B(\mem.mem[68][2] ));
 sg13g2_a21oi_1 _13230_ (.A1(net6016),
    .A2(\mem.mem[69][2] ),
    .Y(_04218_),
    .B1(net5892));
 sg13g2_and2_1 _13231_ (.A(net6020),
    .B(\mem.mem[71][2] ),
    .X(_04219_));
 sg13g2_a21oi_1 _13232_ (.A1(net5372),
    .A2(\mem.mem[70][2] ),
    .Y(_04220_),
    .B1(_04219_));
 sg13g2_a221oi_1 _13233_ (.B2(net5892),
    .C1(net5302),
    .B1(_04220_),
    .A1(_04217_),
    .Y(_04221_),
    .A2(_04218_));
 sg13g2_nand2_1 _13234_ (.Y(_04222_),
    .A(net5371),
    .B(\mem.mem[64][2] ));
 sg13g2_a21oi_1 _13235_ (.A1(net6007),
    .A2(\mem.mem[65][2] ),
    .Y(_04223_),
    .B1(net5887));
 sg13g2_nor2b_1 _13236_ (.A(net6006),
    .B_N(\mem.mem[66][2] ),
    .Y(_04224_));
 sg13g2_a21oi_1 _13237_ (.A1(net6006),
    .A2(\mem.mem[67][2] ),
    .Y(_04225_),
    .B1(_04224_));
 sg13g2_a221oi_1 _13238_ (.B2(net5886),
    .C1(net5850),
    .B1(_04225_),
    .A1(_04222_),
    .Y(_04226_),
    .A2(_04223_));
 sg13g2_nor3_2 _13239_ (.A(net5828),
    .B(_04221_),
    .C(_04226_),
    .Y(_04227_));
 sg13g2_nand2_1 _13240_ (.Y(_04228_),
    .A(net5374),
    .B(\mem.mem[72][2] ));
 sg13g2_a21oi_1 _13241_ (.A1(net6022),
    .A2(\mem.mem[73][2] ),
    .Y(_04229_),
    .B1(net5897));
 sg13g2_nor2b_1 _13242_ (.A(net6021),
    .B_N(\mem.mem[74][2] ),
    .Y(_04230_));
 sg13g2_a21oi_1 _13243_ (.A1(net6025),
    .A2(\mem.mem[75][2] ),
    .Y(_04231_),
    .B1(_04230_));
 sg13g2_a221oi_1 _13244_ (.B2(net5897),
    .C1(net5853),
    .B1(_04231_),
    .A1(_04228_),
    .Y(_04232_),
    .A2(_04229_));
 sg13g2_nor2b_1 _13245_ (.A(net6013),
    .B_N(\mem.mem[78][2] ),
    .Y(_04233_));
 sg13g2_a21oi_1 _13246_ (.A1(net6013),
    .A2(\mem.mem[79][2] ),
    .Y(_04234_),
    .B1(_04233_));
 sg13g2_nand2_1 _13247_ (.Y(_04235_),
    .A(net5371),
    .B(\mem.mem[76][2] ));
 sg13g2_a21oi_1 _13248_ (.A1(net6021),
    .A2(\mem.mem[77][2] ),
    .Y(_04236_),
    .B1(net5891));
 sg13g2_a221oi_1 _13249_ (.B2(_04236_),
    .C1(net5299),
    .B1(_04235_),
    .A1(net5890),
    .Y(_04237_),
    .A2(_04234_));
 sg13g2_nor3_1 _13250_ (.A(net5277),
    .B(_04232_),
    .C(_04237_),
    .Y(_04238_));
 sg13g2_o21ai_1 _13251_ (.B1(net5270),
    .Y(_04239_),
    .A1(_04227_),
    .A2(_04238_));
 sg13g2_nor2b_1 _13252_ (.A(net6008),
    .B_N(\mem.mem[86][2] ),
    .Y(_04240_));
 sg13g2_a21oi_1 _13253_ (.A1(net6008),
    .A2(\mem.mem[87][2] ),
    .Y(_04241_),
    .B1(_04240_));
 sg13g2_a21oi_1 _13254_ (.A1(net6008),
    .A2(\mem.mem[85][2] ),
    .Y(_04242_),
    .B1(net5888));
 sg13g2_o21ai_1 _13255_ (.B1(_04242_),
    .Y(_04243_),
    .A1(net6008),
    .A2(_02847_));
 sg13g2_a21oi_1 _13256_ (.A1(net5888),
    .A2(_04241_),
    .Y(_04244_),
    .B1(net5299));
 sg13g2_mux4_1 _13257_ (.S0(net6007),
    .A0(\mem.mem[80][2] ),
    .A1(\mem.mem[81][2] ),
    .A2(\mem.mem[82][2] ),
    .A3(\mem.mem[83][2] ),
    .S1(net5885),
    .X(_04245_));
 sg13g2_a221oi_1 _13258_ (.B2(net5299),
    .C1(net5827),
    .B1(_04245_),
    .A1(_04243_),
    .Y(_04246_),
    .A2(_04244_));
 sg13g2_nand2_1 _13259_ (.Y(_04247_),
    .A(net5373),
    .B(\mem.mem[88][2] ));
 sg13g2_a21oi_1 _13260_ (.A1(net6046),
    .A2(\mem.mem[89][2] ),
    .Y(_04248_),
    .B1(net5896));
 sg13g2_nor2b_1 _13261_ (.A(net6047),
    .B_N(\mem.mem[90][2] ),
    .Y(_04249_));
 sg13g2_a21oi_1 _13262_ (.A1(net6047),
    .A2(\mem.mem[91][2] ),
    .Y(_04250_),
    .B1(_04249_));
 sg13g2_a221oi_1 _13263_ (.B2(net5896),
    .C1(net5853),
    .B1(_04250_),
    .A1(_04247_),
    .Y(_04251_),
    .A2(_04248_));
 sg13g2_nand2_1 _13264_ (.Y(_04252_),
    .A(net6024),
    .B(\mem.mem[93][2] ));
 sg13g2_a21oi_1 _13265_ (.A1(net5375),
    .A2(\mem.mem[92][2] ),
    .Y(_04253_),
    .B1(net5899));
 sg13g2_and2_1 _13266_ (.A(net6024),
    .B(\mem.mem[95][2] ),
    .X(_04254_));
 sg13g2_a21oi_1 _13267_ (.A1(net5375),
    .A2(\mem.mem[94][2] ),
    .Y(_04255_),
    .B1(_04254_));
 sg13g2_a221oi_1 _13268_ (.B2(net5899),
    .C1(net5303),
    .B1(_04255_),
    .A1(_04252_),
    .Y(_04256_),
    .A2(_04253_));
 sg13g2_nor3_1 _13269_ (.A(net5277),
    .B(_04251_),
    .C(_04256_),
    .Y(_04257_));
 sg13g2_o21ai_1 _13270_ (.B1(net5819),
    .Y(_04258_),
    .A1(_04246_),
    .A2(_04257_));
 sg13g2_nand3_1 _13271_ (.B(_04239_),
    .C(_04258_),
    .A(net5264),
    .Y(_04259_));
 sg13g2_a21oi_1 _13272_ (.A1(net6071),
    .A2(\mem.mem[101][2] ),
    .Y(_04260_),
    .B1(net5930));
 sg13g2_o21ai_1 _13273_ (.B1(_04260_),
    .Y(_04261_),
    .A1(net6071),
    .A2(_02848_));
 sg13g2_and2_1 _13274_ (.A(net6071),
    .B(\mem.mem[103][2] ),
    .X(_04262_));
 sg13g2_a21oi_1 _13275_ (.A1(net5390),
    .A2(\mem.mem[102][2] ),
    .Y(_04263_),
    .B1(_04262_));
 sg13g2_a21oi_1 _13276_ (.A1(net5931),
    .A2(_04263_),
    .Y(_04264_),
    .B1(net5316));
 sg13g2_mux4_1 _13277_ (.S0(net6072),
    .A0(\mem.mem[96][2] ),
    .A1(\mem.mem[97][2] ),
    .A2(\mem.mem[98][2] ),
    .A3(\mem.mem[99][2] ),
    .S1(net5930),
    .X(_04265_));
 sg13g2_a221oi_1 _13278_ (.B2(net5317),
    .C1(net5834),
    .B1(_04265_),
    .A1(_04261_),
    .Y(_04266_),
    .A2(_04264_));
 sg13g2_nand2_1 _13279_ (.Y(_04267_),
    .A(net5388),
    .B(\mem.mem[104][2] ));
 sg13g2_a21oi_1 _13280_ (.A1(net6066),
    .A2(\mem.mem[105][2] ),
    .Y(_04268_),
    .B1(net5926));
 sg13g2_nor2b_1 _13281_ (.A(net6066),
    .B_N(\mem.mem[106][2] ),
    .Y(_04269_));
 sg13g2_a21oi_1 _13282_ (.A1(net6066),
    .A2(\mem.mem[107][2] ),
    .Y(_04270_),
    .B1(_04269_));
 sg13g2_a221oi_1 _13283_ (.B2(net5926),
    .C1(net5861),
    .B1(_04270_),
    .A1(_04267_),
    .Y(_04271_),
    .A2(_04268_));
 sg13g2_nor2b_1 _13284_ (.A(net6065),
    .B_N(\mem.mem[110][2] ),
    .Y(_04272_));
 sg13g2_a21oi_1 _13285_ (.A1(net6065),
    .A2(\mem.mem[111][2] ),
    .Y(_04273_),
    .B1(_04272_));
 sg13g2_nand2_1 _13286_ (.Y(_04274_),
    .A(net5388),
    .B(\mem.mem[108][2] ));
 sg13g2_a21oi_1 _13287_ (.A1(net6065),
    .A2(\mem.mem[109][2] ),
    .Y(_04275_),
    .B1(net5925));
 sg13g2_a221oi_1 _13288_ (.B2(_04275_),
    .C1(net5317),
    .B1(_04274_),
    .A1(net5925),
    .Y(_04276_),
    .A2(_04273_));
 sg13g2_nor3_1 _13289_ (.A(net5284),
    .B(_04271_),
    .C(_04276_),
    .Y(_04277_));
 sg13g2_o21ai_1 _13290_ (.B1(net5268),
    .Y(_04278_),
    .A1(_04266_),
    .A2(_04277_));
 sg13g2_nor2b_1 _13291_ (.A(net6023),
    .B_N(\mem.mem[118][2] ),
    .Y(_04279_));
 sg13g2_a21oi_1 _13292_ (.A1(net6023),
    .A2(\mem.mem[119][2] ),
    .Y(_04280_),
    .B1(_04279_));
 sg13g2_nand2_1 _13293_ (.Y(_04281_),
    .A(net5374),
    .B(\mem.mem[116][2] ));
 sg13g2_a21oi_1 _13294_ (.A1(net6023),
    .A2(\mem.mem[117][2] ),
    .Y(_04282_),
    .B1(net5898));
 sg13g2_a221oi_1 _13295_ (.B2(_04282_),
    .C1(net5303),
    .B1(_04281_),
    .A1(net5898),
    .Y(_04283_),
    .A2(_04280_));
 sg13g2_nand2_1 _13296_ (.Y(_04284_),
    .A(net5380),
    .B(\mem.mem[112][2] ));
 sg13g2_a21oi_1 _13297_ (.A1(net6036),
    .A2(\mem.mem[113][2] ),
    .Y(_04285_),
    .B1(net5908));
 sg13g2_nor2b_1 _13298_ (.A(net6063),
    .B_N(\mem.mem[114][2] ),
    .Y(_04286_));
 sg13g2_a21oi_1 _13299_ (.A1(net6063),
    .A2(\mem.mem[115][2] ),
    .Y(_04287_),
    .B1(_04286_));
 sg13g2_a221oi_1 _13300_ (.B2(net5908),
    .C1(net5855),
    .B1(_04287_),
    .A1(_04284_),
    .Y(_04288_),
    .A2(_04285_));
 sg13g2_nor3_1 _13301_ (.A(net5830),
    .B(_04283_),
    .C(_04288_),
    .Y(_04289_));
 sg13g2_mux4_1 _13302_ (.S0(net6041),
    .A0(\mem.mem[120][2] ),
    .A1(\mem.mem[121][2] ),
    .A2(\mem.mem[122][2] ),
    .A3(\mem.mem[123][2] ),
    .S1(net5911),
    .X(_04290_));
 sg13g2_nand2_1 _13303_ (.Y(_04291_),
    .A(net6040),
    .B(\mem.mem[125][2] ));
 sg13g2_a21oi_1 _13304_ (.A1(net5382),
    .A2(\mem.mem[124][2] ),
    .Y(_04292_),
    .B1(net5910));
 sg13g2_a21oi_1 _13305_ (.A1(net6039),
    .A2(\mem.mem[127][2] ),
    .Y(_04293_),
    .B1(net5351));
 sg13g2_o21ai_1 _13306_ (.B1(_04293_),
    .Y(_04294_),
    .A1(net6039),
    .A2(_02849_));
 sg13g2_a21oi_1 _13307_ (.A1(_04291_),
    .A2(_04292_),
    .Y(_04295_),
    .B1(net5308));
 sg13g2_a221oi_1 _13308_ (.B2(_04295_),
    .C1(net5280),
    .B1(_04294_),
    .A1(net5308),
    .Y(_04296_),
    .A2(_04290_));
 sg13g2_o21ai_1 _13309_ (.B1(net5817),
    .Y(_04297_),
    .A1(_04289_),
    .A2(_04296_));
 sg13g2_nand3_1 _13310_ (.B(_04278_),
    .C(_04297_),
    .A(net5809),
    .Y(_04298_));
 sg13g2_a21oi_1 _13311_ (.A1(net6158),
    .A2(\mem.mem[37][2] ),
    .Y(_04299_),
    .B1(net5992));
 sg13g2_o21ai_1 _13312_ (.B1(_04299_),
    .Y(_04300_),
    .A1(net6152),
    .A2(_02846_));
 sg13g2_and2_1 _13313_ (.A(net6152),
    .B(\mem.mem[39][2] ),
    .X(_04301_));
 sg13g2_a21oi_1 _13314_ (.A1(net5418),
    .A2(\mem.mem[38][2] ),
    .Y(_04302_),
    .B1(_04301_));
 sg13g2_a21oi_1 _13315_ (.A1(net5989),
    .A2(_04302_),
    .Y(_04303_),
    .B1(net5340));
 sg13g2_mux4_1 _13316_ (.S0(net6159),
    .A0(\mem.mem[32][2] ),
    .A1(\mem.mem[33][2] ),
    .A2(\mem.mem[34][2] ),
    .A3(\mem.mem[35][2] ),
    .S1(net5994),
    .X(_04304_));
 sg13g2_a221oi_1 _13317_ (.B2(net5342),
    .C1(net5846),
    .B1(_04304_),
    .A1(_04300_),
    .Y(_04305_),
    .A2(_04303_));
 sg13g2_nand2_1 _13318_ (.Y(_04306_),
    .A(net5421),
    .B(\mem.mem[40][2] ));
 sg13g2_a21oi_1 _13319_ (.A1(net6170),
    .A2(\mem.mem[41][2] ),
    .Y(_04307_),
    .B1(net6001));
 sg13g2_nor2b_1 _13320_ (.A(net6170),
    .B_N(\mem.mem[42][2] ),
    .Y(_04308_));
 sg13g2_a21oi_1 _13321_ (.A1(net6170),
    .A2(\mem.mem[43][2] ),
    .Y(_04309_),
    .B1(_04308_));
 sg13g2_a221oi_1 _13322_ (.B2(net6001),
    .C1(net5882),
    .B1(_04309_),
    .A1(_04306_),
    .Y(_04310_),
    .A2(_04307_));
 sg13g2_nor2b_1 _13323_ (.A(net6165),
    .B_N(\mem.mem[46][2] ),
    .Y(_04311_));
 sg13g2_a21oi_1 _13324_ (.A1(net6164),
    .A2(\mem.mem[47][2] ),
    .Y(_04312_),
    .B1(_04311_));
 sg13g2_nand2_1 _13325_ (.Y(_04313_),
    .A(net5421),
    .B(\mem.mem[44][2] ));
 sg13g2_a21oi_1 _13326_ (.A1(net6164),
    .A2(\mem.mem[45][2] ),
    .Y(_04314_),
    .B1(net5997));
 sg13g2_a221oi_1 _13327_ (.B2(_04314_),
    .C1(net5344),
    .B1(_04313_),
    .A1(net5997),
    .Y(_04315_),
    .A2(_04312_));
 sg13g2_nor3_2 _13328_ (.A(net5296),
    .B(_04310_),
    .C(_04315_),
    .Y(_04316_));
 sg13g2_o21ai_1 _13329_ (.B1(net5273),
    .Y(_04317_),
    .A1(_04305_),
    .A2(_04316_));
 sg13g2_nor2b_1 _13330_ (.A(net6026),
    .B_N(\mem.mem[54][2] ),
    .Y(_04318_));
 sg13g2_a21oi_1 _13331_ (.A1(net6026),
    .A2(\mem.mem[55][2] ),
    .Y(_04319_),
    .B1(_04318_));
 sg13g2_nand2_1 _13332_ (.Y(_04320_),
    .A(net5379),
    .B(\mem.mem[52][2] ));
 sg13g2_a21oi_1 _13333_ (.A1(net6027),
    .A2(\mem.mem[53][2] ),
    .Y(_04321_),
    .B1(net5902));
 sg13g2_a221oi_1 _13334_ (.B2(_04321_),
    .C1(net5305),
    .B1(_04320_),
    .A1(net5902),
    .Y(_04322_),
    .A2(_04319_));
 sg13g2_nand2_1 _13335_ (.Y(_04323_),
    .A(net5379),
    .B(\mem.mem[48][2] ));
 sg13g2_a21oi_1 _13336_ (.A1(net6028),
    .A2(\mem.mem[49][2] ),
    .Y(_04324_),
    .B1(net5901));
 sg13g2_nor2b_1 _13337_ (.A(net6011),
    .B_N(\mem.mem[50][2] ),
    .Y(_04325_));
 sg13g2_a21oi_1 _13338_ (.A1(net6011),
    .A2(\mem.mem[51][2] ),
    .Y(_04326_),
    .B1(_04325_));
 sg13g2_a221oi_1 _13339_ (.B2(net5901),
    .C1(net5854),
    .B1(_04326_),
    .A1(_04323_),
    .Y(_04327_),
    .A2(_04324_));
 sg13g2_nor3_1 _13340_ (.A(net5829),
    .B(_04322_),
    .C(_04327_),
    .Y(_04328_));
 sg13g2_nand2_1 _13341_ (.Y(_04329_),
    .A(net5377),
    .B(\mem.mem[56][2] ));
 sg13g2_a21oi_1 _13342_ (.A1(net6033),
    .A2(\mem.mem[57][2] ),
    .Y(_04330_),
    .B1(net5903));
 sg13g2_nor2b_1 _13343_ (.A(net6030),
    .B_N(\mem.mem[58][2] ),
    .Y(_04331_));
 sg13g2_a21oi_1 _13344_ (.A1(net6030),
    .A2(\mem.mem[59][2] ),
    .Y(_04332_),
    .B1(_04331_));
 sg13g2_a221oi_1 _13345_ (.B2(net5903),
    .C1(net5855),
    .B1(_04332_),
    .A1(_04329_),
    .Y(_04333_),
    .A2(_04330_));
 sg13g2_nand2_1 _13346_ (.Y(_04334_),
    .A(net6039),
    .B(\mem.mem[61][2] ));
 sg13g2_a21oi_1 _13347_ (.A1(net5381),
    .A2(\mem.mem[60][2] ),
    .Y(_04335_),
    .B1(net5912));
 sg13g2_and2_1 _13348_ (.A(net6038),
    .B(\mem.mem[63][2] ),
    .X(_04336_));
 sg13g2_a21oi_1 _13349_ (.A1(net5381),
    .A2(\mem.mem[62][2] ),
    .Y(_04337_),
    .B1(_04336_));
 sg13g2_a221oi_1 _13350_ (.B2(net5912),
    .C1(net5307),
    .B1(_04337_),
    .A1(_04334_),
    .Y(_04338_),
    .A2(_04335_));
 sg13g2_nor3_1 _13351_ (.A(net5279),
    .B(_04333_),
    .C(_04338_),
    .Y(_04339_));
 sg13g2_o21ai_1 _13352_ (.B1(net5817),
    .Y(_04340_),
    .A1(_04328_),
    .A2(_04339_));
 sg13g2_nand3_1 _13353_ (.B(_04317_),
    .C(_04340_),
    .A(net5810),
    .Y(_04341_));
 sg13g2_a21oi_1 _13354_ (.A1(net6080),
    .A2(\mem.mem[5][2] ),
    .Y(_04342_),
    .B1(net5937));
 sg13g2_o21ai_1 _13355_ (.B1(_04342_),
    .Y(_04343_),
    .A1(net6080),
    .A2(_02844_));
 sg13g2_and2_1 _13356_ (.A(net6075),
    .B(\mem.mem[7][2] ),
    .X(_04344_));
 sg13g2_a21oi_2 _13357_ (.B1(_04344_),
    .Y(_04345_),
    .A2(\mem.mem[6][2] ),
    .A1(net5391));
 sg13g2_a21oi_1 _13358_ (.A1(net5937),
    .A2(_04345_),
    .Y(_04346_),
    .B1(net5318));
 sg13g2_mux4_1 _13359_ (.S0(net6080),
    .A0(\mem.mem[0][2] ),
    .A1(\mem.mem[1][2] ),
    .A2(\mem.mem[2][2] ),
    .A3(\mem.mem[3][2] ),
    .S1(net5937),
    .X(_04347_));
 sg13g2_a221oi_1 _13360_ (.B2(net5318),
    .C1(net5835),
    .B1(_04347_),
    .A1(_04343_),
    .Y(_04348_),
    .A2(_04346_));
 sg13g2_nand2_1 _13361_ (.Y(_04349_),
    .A(net5393),
    .B(\mem.mem[8][2] ));
 sg13g2_a21oi_1 _13362_ (.A1(net6082),
    .A2(\mem.mem[9][2] ),
    .Y(_04350_),
    .B1(net5939));
 sg13g2_nor2b_1 _13363_ (.A(net6082),
    .B_N(\mem.mem[10][2] ),
    .Y(_04351_));
 sg13g2_a21oi_1 _13364_ (.A1(net6082),
    .A2(\mem.mem[11][2] ),
    .Y(_04352_),
    .B1(_04351_));
 sg13g2_a221oi_1 _13365_ (.B2(net5936),
    .C1(net5863),
    .B1(_04352_),
    .A1(_04349_),
    .Y(_04353_),
    .A2(_04350_));
 sg13g2_nor2b_1 _13366_ (.A(net6111),
    .B_N(\mem.mem[14][2] ),
    .Y(_04354_));
 sg13g2_a21oi_1 _13367_ (.A1(net6111),
    .A2(\mem.mem[15][2] ),
    .Y(_04355_),
    .B1(_04354_));
 sg13g2_nand2_1 _13368_ (.Y(_04356_),
    .A(net5403),
    .B(\mem.mem[12][2] ));
 sg13g2_a21oi_1 _13369_ (.A1(net6110),
    .A2(\mem.mem[13][2] ),
    .Y(_04357_),
    .B1(net5958));
 sg13g2_a221oi_1 _13370_ (.B2(_04357_),
    .C1(net5330),
    .B1(_04356_),
    .A1(net5958),
    .Y(_04358_),
    .A2(_04355_));
 sg13g2_nor3_2 _13371_ (.A(net5284),
    .B(_04353_),
    .C(_04358_),
    .Y(_04359_));
 sg13g2_o21ai_1 _13372_ (.B1(net5269),
    .Y(_04360_),
    .A1(_04348_),
    .A2(_04359_));
 sg13g2_a21oi_1 _13373_ (.A1(net6127),
    .A2(\mem.mem[23][2] ),
    .Y(_04361_),
    .B1(net5362));
 sg13g2_o21ai_1 _13374_ (.B1(_04361_),
    .Y(_04362_),
    .A1(net6127),
    .A2(_02845_));
 sg13g2_nand2_1 _13375_ (.Y(_04363_),
    .A(net5406),
    .B(\mem.mem[20][2] ));
 sg13g2_a21oi_1 _13376_ (.A1(net6126),
    .A2(\mem.mem[21][2] ),
    .Y(_04364_),
    .B1(net5969));
 sg13g2_a21oi_1 _13377_ (.A1(_04363_),
    .A2(_04364_),
    .Y(_04365_),
    .B1(net5331));
 sg13g2_mux4_1 _13378_ (.S0(net6127),
    .A0(\mem.mem[16][2] ),
    .A1(\mem.mem[17][2] ),
    .A2(\mem.mem[18][2] ),
    .A3(\mem.mem[19][2] ),
    .S1(net5968),
    .X(_04366_));
 sg13g2_a221oi_1 _13379_ (.B2(net5331),
    .C1(net5840),
    .B1(_04366_),
    .A1(_04362_),
    .Y(_04367_),
    .A2(_04365_));
 sg13g2_nand2_1 _13380_ (.Y(_04368_),
    .A(net5407),
    .B(\mem.mem[24][2] ));
 sg13g2_a21oi_1 _13381_ (.A1(net6128),
    .A2(\mem.mem[25][2] ),
    .Y(_04369_),
    .B1(net5968));
 sg13g2_nor2b_1 _13382_ (.A(net6128),
    .B_N(\mem.mem[26][2] ),
    .Y(_04370_));
 sg13g2_a21oi_1 _13383_ (.A1(net6128),
    .A2(\mem.mem[27][2] ),
    .Y(_04371_),
    .B1(_04370_));
 sg13g2_a221oi_1 _13384_ (.B2(net5968),
    .C1(net5873),
    .B1(_04371_),
    .A1(_04368_),
    .Y(_04372_),
    .A2(_04369_));
 sg13g2_nand2_1 _13385_ (.Y(_04373_),
    .A(net6157),
    .B(\mem.mem[29][2] ));
 sg13g2_a21oi_1 _13386_ (.A1(net5416),
    .A2(\mem.mem[28][2] ),
    .Y(_04374_),
    .B1(net5990));
 sg13g2_and2_1 _13387_ (.A(net6157),
    .B(\mem.mem[31][2] ),
    .X(_04375_));
 sg13g2_a21oi_1 _13388_ (.A1(net5416),
    .A2(\mem.mem[30][2] ),
    .Y(_04376_),
    .B1(_04375_));
 sg13g2_a221oi_1 _13389_ (.B2(net5990),
    .C1(net5341),
    .B1(_04376_),
    .A1(_04373_),
    .Y(_04377_),
    .A2(_04374_));
 sg13g2_nor3_1 _13390_ (.A(net5290),
    .B(_04372_),
    .C(_04377_),
    .Y(_04378_));
 sg13g2_o21ai_1 _13391_ (.B1(net5824),
    .Y(_04379_),
    .A1(_04367_),
    .A2(_04378_));
 sg13g2_nand3_1 _13392_ (.B(_04360_),
    .C(_04379_),
    .A(net5267),
    .Y(_04380_));
 sg13g2_nand3_1 _13393_ (.B(_04341_),
    .C(_04380_),
    .A(net5262),
    .Y(_04381_));
 sg13g2_nand3_1 _13394_ (.B(_04259_),
    .C(_04298_),
    .A(net5808),
    .Y(_04382_));
 sg13g2_a21o_1 _13395_ (.A2(_04382_),
    .A1(_04381_),
    .B1(_00007_),
    .X(_04383_));
 sg13g2_nor2b_1 _13396_ (.A(net6118),
    .B_N(\mem.mem[134][2] ),
    .Y(_04384_));
 sg13g2_a21oi_1 _13397_ (.A1(net6118),
    .A2(\mem.mem[135][2] ),
    .Y(_04385_),
    .B1(_04384_));
 sg13g2_nand2_1 _13398_ (.Y(_04386_),
    .A(net5407),
    .B(\mem.mem[132][2] ));
 sg13g2_a21oi_1 _13399_ (.A1(net6118),
    .A2(\mem.mem[133][2] ),
    .Y(_04387_),
    .B1(net5964));
 sg13g2_a221oi_1 _13400_ (.B2(_04387_),
    .C1(net5332),
    .B1(_04386_),
    .A1(net5964),
    .Y(_04388_),
    .A2(_04385_));
 sg13g2_nand2_1 _13401_ (.Y(_04389_),
    .A(net5405),
    .B(\mem.mem[128][2] ));
 sg13g2_a21oi_1 _13402_ (.A1(net6116),
    .A2(\mem.mem[129][2] ),
    .Y(_04390_),
    .B1(net5963));
 sg13g2_nor2b_1 _13403_ (.A(net6116),
    .B_N(\mem.mem[130][2] ),
    .Y(_04391_));
 sg13g2_a21oi_1 _13404_ (.A1(net6116),
    .A2(\mem.mem[131][2] ),
    .Y(_04392_),
    .B1(_04391_));
 sg13g2_a221oi_1 _13405_ (.B2(net5963),
    .C1(net5872),
    .B1(_04392_),
    .A1(_04389_),
    .Y(_04393_),
    .A2(_04390_));
 sg13g2_o21ai_1 _13406_ (.B1(net5291),
    .Y(_04394_),
    .A1(_04388_),
    .A2(_04393_));
 sg13g2_nand2_1 _13407_ (.Y(_04395_),
    .A(net6122),
    .B(\mem.mem[141][2] ));
 sg13g2_a21oi_1 _13408_ (.A1(net5403),
    .A2(\mem.mem[140][2] ),
    .Y(_04396_),
    .B1(net5960));
 sg13g2_and2_1 _13409_ (.A(net6114),
    .B(\mem.mem[143][2] ),
    .X(_04397_));
 sg13g2_a21oi_1 _13410_ (.A1(net5403),
    .A2(\mem.mem[142][2] ),
    .Y(_04398_),
    .B1(_04397_));
 sg13g2_a221oi_1 _13411_ (.B2(net5960),
    .C1(net5329),
    .B1(_04398_),
    .A1(_04395_),
    .Y(_04399_),
    .A2(_04396_));
 sg13g2_nand2_1 _13412_ (.Y(_04400_),
    .A(net5406),
    .B(\mem.mem[136][2] ));
 sg13g2_a21oi_1 _13413_ (.A1(net6122),
    .A2(\mem.mem[137][2] ),
    .Y(_04401_),
    .B1(net5967));
 sg13g2_nor2b_1 _13414_ (.A(net6121),
    .B_N(\mem.mem[138][2] ),
    .Y(_04402_));
 sg13g2_a21oi_1 _13415_ (.A1(net6122),
    .A2(\mem.mem[139][2] ),
    .Y(_04403_),
    .B1(_04402_));
 sg13g2_a221oi_1 _13416_ (.B2(net5967),
    .C1(net5871),
    .B1(_04403_),
    .A1(_04400_),
    .Y(_04404_),
    .A2(_04401_));
 sg13g2_o21ai_1 _13417_ (.B1(net5840),
    .Y(_04405_),
    .A1(_04399_),
    .A2(_04404_));
 sg13g2_nand3_1 _13418_ (.B(_04394_),
    .C(_04405_),
    .A(net5271),
    .Y(_04406_));
 sg13g2_nand2_1 _13419_ (.Y(_04407_),
    .A(net5402),
    .B(\mem.mem[148][2] ));
 sg13g2_a21oi_1 _13420_ (.A1(net6105),
    .A2(\mem.mem[149][2] ),
    .Y(_04408_),
    .B1(net5956));
 sg13g2_and2_1 _13421_ (.A(net6105),
    .B(\mem.mem[151][2] ),
    .X(_04409_));
 sg13g2_a21oi_1 _13422_ (.A1(net5402),
    .A2(\mem.mem[150][2] ),
    .Y(_04410_),
    .B1(_04409_));
 sg13g2_a221oi_1 _13423_ (.B2(net5956),
    .C1(net5320),
    .B1(_04410_),
    .A1(_04407_),
    .Y(_04411_),
    .A2(_04408_));
 sg13g2_nand2_1 _13424_ (.Y(_04412_),
    .A(net5392),
    .B(\mem.mem[144][2] ));
 sg13g2_a21oi_1 _13425_ (.A1(net6076),
    .A2(\mem.mem[145][2] ),
    .Y(_04413_),
    .B1(net5933));
 sg13g2_nor2b_1 _13426_ (.A(net6077),
    .B_N(\mem.mem[146][2] ),
    .Y(_04414_));
 sg13g2_a21oi_1 _13427_ (.A1(net6076),
    .A2(\mem.mem[147][2] ),
    .Y(_04415_),
    .B1(_04414_));
 sg13g2_a221oi_1 _13428_ (.B2(net5933),
    .C1(net5863),
    .B1(_04415_),
    .A1(_04412_),
    .Y(_04416_),
    .A2(_04413_));
 sg13g2_o21ai_1 _13429_ (.B1(net5283),
    .Y(_04417_),
    .A1(_04411_),
    .A2(_04416_));
 sg13g2_nor2b_1 _13430_ (.A(net6107),
    .B_N(\mem.mem[158][2] ),
    .Y(_04418_));
 sg13g2_a21oi_1 _13431_ (.A1(net6107),
    .A2(\mem.mem[159][2] ),
    .Y(_04419_),
    .B1(_04418_));
 sg13g2_nand2_1 _13432_ (.Y(_04420_),
    .A(net5404),
    .B(\mem.mem[156][2] ));
 sg13g2_a21oi_1 _13433_ (.A1(net6107),
    .A2(\mem.mem[157][2] ),
    .Y(_04421_),
    .B1(net5955));
 sg13g2_a221oi_1 _13434_ (.B2(_04421_),
    .C1(net5329),
    .B1(_04420_),
    .A1(net5962),
    .Y(_04422_),
    .A2(_04419_));
 sg13g2_nand2_1 _13435_ (.Y(_04423_),
    .A(net5402),
    .B(\mem.mem[152][2] ));
 sg13g2_a21oi_1 _13436_ (.A1(net6107),
    .A2(\mem.mem[153][2] ),
    .Y(_04424_),
    .B1(net5957));
 sg13g2_nor2b_1 _13437_ (.A(net6092),
    .B_N(\mem.mem[154][2] ),
    .Y(_04425_));
 sg13g2_a21oi_1 _13438_ (.A1(net6092),
    .A2(\mem.mem[155][2] ),
    .Y(_04426_),
    .B1(_04425_));
 sg13g2_a221oi_1 _13439_ (.B2(net5957),
    .C1(net5869),
    .B1(_04426_),
    .A1(_04423_),
    .Y(_04427_),
    .A2(_04424_));
 sg13g2_o21ai_1 _13440_ (.B1(net5841),
    .Y(_04428_),
    .A1(_04422_),
    .A2(_04427_));
 sg13g2_nand3_1 _13441_ (.B(_04417_),
    .C(_04428_),
    .A(net5822),
    .Y(_04429_));
 sg13g2_nand3_1 _13442_ (.B(_04406_),
    .C(_04429_),
    .A(net5265),
    .Y(_04430_));
 sg13g2_mux4_1 _13443_ (.S0(net6055),
    .A0(\mem.mem[160][2] ),
    .A1(\mem.mem[161][2] ),
    .A2(\mem.mem[162][2] ),
    .A3(\mem.mem[163][2] ),
    .S1(net5921),
    .X(_04431_));
 sg13g2_and2_1 _13444_ (.A(net5312),
    .B(_04431_),
    .X(_04432_));
 sg13g2_nor2b_1 _13445_ (.A(net6055),
    .B_N(\mem.mem[166][2] ),
    .Y(_04433_));
 sg13g2_a21oi_1 _13446_ (.A1(net6057),
    .A2(\mem.mem[167][2] ),
    .Y(_04434_),
    .B1(_04433_));
 sg13g2_nand2_1 _13447_ (.Y(_04435_),
    .A(net5387),
    .B(\mem.mem[164][2] ));
 sg13g2_a21oi_1 _13448_ (.A1(net6055),
    .A2(\mem.mem[165][2] ),
    .Y(_04436_),
    .B1(net5921));
 sg13g2_a221oi_1 _13449_ (.B2(_04436_),
    .C1(net5312),
    .B1(_04435_),
    .A1(net5921),
    .Y(_04437_),
    .A2(_04434_));
 sg13g2_o21ai_1 _13450_ (.B1(net5282),
    .Y(_04438_),
    .A1(_04432_),
    .A2(_04437_));
 sg13g2_nand2_1 _13451_ (.Y(_04439_),
    .A(net6090),
    .B(\mem.mem[173][2] ));
 sg13g2_a21oi_1 _13452_ (.A1(net5397),
    .A2(\mem.mem[172][2] ),
    .Y(_04440_),
    .B1(net5946));
 sg13g2_and2_1 _13453_ (.A(net6090),
    .B(\mem.mem[175][2] ),
    .X(_04441_));
 sg13g2_a21oi_1 _13454_ (.A1(net5397),
    .A2(\mem.mem[174][2] ),
    .Y(_04442_),
    .B1(_04441_));
 sg13g2_a221oi_1 _13455_ (.B2(net5946),
    .C1(net5323),
    .B1(_04442_),
    .A1(_04439_),
    .Y(_04443_),
    .A2(_04440_));
 sg13g2_nand2_1 _13456_ (.Y(_04444_),
    .A(net5396),
    .B(\mem.mem[168][2] ));
 sg13g2_a21oi_1 _13457_ (.A1(net6086),
    .A2(\mem.mem[169][2] ),
    .Y(_04445_),
    .B1(net5943));
 sg13g2_nor2b_1 _13458_ (.A(net6086),
    .B_N(\mem.mem[170][2] ),
    .Y(_04446_));
 sg13g2_a21oi_1 _13459_ (.A1(net6085),
    .A2(\mem.mem[171][2] ),
    .Y(_04447_),
    .B1(_04446_));
 sg13g2_a221oi_1 _13460_ (.B2(net5943),
    .C1(net5865),
    .B1(_04447_),
    .A1(_04444_),
    .Y(_04448_),
    .A2(_04445_));
 sg13g2_o21ai_1 _13461_ (.B1(net5838),
    .Y(_04449_),
    .A1(_04443_),
    .A2(_04448_));
 sg13g2_nand3_1 _13462_ (.B(_04438_),
    .C(_04449_),
    .A(net5272),
    .Y(_04450_));
 sg13g2_nand2_1 _13463_ (.Y(_04451_),
    .A(net5410),
    .B(\mem.mem[180][2] ));
 sg13g2_a21oi_1 _13464_ (.A1(net6135),
    .A2(\mem.mem[181][2] ),
    .Y(_04452_),
    .B1(net5975));
 sg13g2_and2_1 _13465_ (.A(net6135),
    .B(\mem.mem[183][2] ),
    .X(_04453_));
 sg13g2_a21oi_1 _13466_ (.A1(net5409),
    .A2(\mem.mem[182][2] ),
    .Y(_04454_),
    .B1(_04453_));
 sg13g2_a221oi_1 _13467_ (.B2(net5975),
    .C1(net5336),
    .B1(_04454_),
    .A1(_04451_),
    .Y(_04455_),
    .A2(_04452_));
 sg13g2_nand2_1 _13468_ (.Y(_04456_),
    .A(net5411),
    .B(\mem.mem[176][2] ));
 sg13g2_a21oi_1 _13469_ (.A1(net6133),
    .A2(\mem.mem[177][2] ),
    .Y(_04457_),
    .B1(net5973));
 sg13g2_nor2b_1 _13470_ (.A(net6132),
    .B_N(\mem.mem[178][2] ),
    .Y(_04458_));
 sg13g2_a21oi_1 _13471_ (.A1(net6132),
    .A2(\mem.mem[179][2] ),
    .Y(_04459_),
    .B1(_04458_));
 sg13g2_a221oi_1 _13472_ (.B2(net5974),
    .C1(net5875),
    .B1(_04459_),
    .A1(_04456_),
    .Y(_04460_),
    .A2(_04457_));
 sg13g2_o21ai_1 _13473_ (.B1(net5292),
    .Y(_04461_),
    .A1(_04455_),
    .A2(_04460_));
 sg13g2_nor2b_1 _13474_ (.A(net6103),
    .B_N(\mem.mem[190][2] ),
    .Y(_04462_));
 sg13g2_a21oi_1 _13475_ (.A1(net6101),
    .A2(\mem.mem[191][2] ),
    .Y(_04463_),
    .B1(_04462_));
 sg13g2_nand2_1 _13476_ (.Y(_04464_),
    .A(net5400),
    .B(\mem.mem[188][2] ));
 sg13g2_a21oi_1 _13477_ (.A1(net6101),
    .A2(\mem.mem[189][2] ),
    .Y(_04465_),
    .B1(net5952));
 sg13g2_a221oi_1 _13478_ (.B2(_04465_),
    .C1(net5325),
    .B1(_04464_),
    .A1(net5952),
    .Y(_04466_),
    .A2(_04463_));
 sg13g2_nand2_1 _13479_ (.Y(_04467_),
    .A(net5401),
    .B(\mem.mem[184][2] ));
 sg13g2_a21oi_1 _13480_ (.A1(net6097),
    .A2(\mem.mem[185][2] ),
    .Y(_04468_),
    .B1(net5950));
 sg13g2_nor2b_1 _13481_ (.A(net6097),
    .B_N(\mem.mem[186][2] ),
    .Y(_04469_));
 sg13g2_a21oi_1 _13482_ (.A1(net6097),
    .A2(\mem.mem[187][2] ),
    .Y(_04470_),
    .B1(_04469_));
 sg13g2_a221oi_1 _13483_ (.B2(net5950),
    .C1(net5867),
    .B1(_04470_),
    .A1(_04467_),
    .Y(_04471_),
    .A2(_04468_));
 sg13g2_o21ai_1 _13484_ (.B1(net5838),
    .Y(_04472_),
    .A1(_04466_),
    .A2(_04471_));
 sg13g2_nand3_1 _13485_ (.B(_04461_),
    .C(_04472_),
    .A(net5823),
    .Y(_04473_));
 sg13g2_nand3_1 _13486_ (.B(_04450_),
    .C(_04473_),
    .A(net5815),
    .Y(_04474_));
 sg13g2_nand2_1 _13487_ (.Y(_04475_),
    .A(net6059),
    .B(\mem.mem[247][2] ));
 sg13g2_nand2b_1 _13488_ (.Y(_04476_),
    .B(\mem.mem[246][2] ),
    .A_N(net6059));
 sg13g2_nand3_1 _13489_ (.B(_04475_),
    .C(_04476_),
    .A(net5922),
    .Y(_04477_));
 sg13g2_nand2b_1 _13490_ (.Y(_04478_),
    .B(\mem.mem[244][2] ),
    .A_N(net6059));
 sg13g2_a21oi_1 _13491_ (.A1(net6059),
    .A2(\mem.mem[245][2] ),
    .Y(_04479_),
    .B1(net5922));
 sg13g2_mux4_1 _13492_ (.S0(net6057),
    .A0(\mem.mem[240][2] ),
    .A1(\mem.mem[241][2] ),
    .A2(\mem.mem[242][2] ),
    .A3(\mem.mem[243][2] ),
    .S1(net5921),
    .X(_04480_));
 sg13g2_a21o_1 _13493_ (.A2(_04474_),
    .A1(_04430_),
    .B1(_00006_),
    .X(_04481_));
 sg13g2_nand2_1 _13494_ (.Y(_04482_),
    .A(net5400),
    .B(\mem.mem[198][2] ));
 sg13g2_a21oi_1 _13495_ (.A1(net6101),
    .A2(\mem.mem[199][2] ),
    .Y(_04483_),
    .B1(net5360));
 sg13g2_and2_1 _13496_ (.A(net6101),
    .B(\mem.mem[197][2] ),
    .X(_04484_));
 sg13g2_a21oi_1 _13497_ (.A1(net5400),
    .A2(\mem.mem[196][2] ),
    .Y(_04485_),
    .B1(_04484_));
 sg13g2_a221oi_1 _13498_ (.B2(net5358),
    .C1(net5325),
    .B1(_04485_),
    .A1(_04482_),
    .Y(_04486_),
    .A2(_04483_));
 sg13g2_nand2_1 _13499_ (.Y(_04487_),
    .A(net6099),
    .B(\mem.mem[193][2] ));
 sg13g2_nand2_1 _13500_ (.Y(_04488_),
    .A(net5399),
    .B(\mem.mem[192][2] ));
 sg13g2_nand3_1 _13501_ (.B(_04487_),
    .C(_04488_),
    .A(net5358),
    .Y(_04489_));
 sg13g2_and2_1 _13502_ (.A(net6099),
    .B(\mem.mem[195][2] ),
    .X(_04490_));
 sg13g2_a21oi_1 _13503_ (.A1(net5399),
    .A2(\mem.mem[194][2] ),
    .Y(_04491_),
    .B1(_04490_));
 sg13g2_a21oi_1 _13504_ (.A1(net5953),
    .A2(_04491_),
    .Y(_04492_),
    .B1(net5868));
 sg13g2_a21oi_1 _13505_ (.A1(_04489_),
    .A2(_04492_),
    .Y(_04493_),
    .B1(_04486_));
 sg13g2_mux2_1 _13506_ (.A0(\mem.mem[204][2] ),
    .A1(\mem.mem[205][2] ),
    .S(net6093),
    .X(_04494_));
 sg13g2_nor2b_1 _13507_ (.A(net6093),
    .B_N(\mem.mem[206][2] ),
    .Y(_04495_));
 sg13g2_a21oi_1 _13508_ (.A1(net6093),
    .A2(\mem.mem[207][2] ),
    .Y(_04496_),
    .B1(_04495_));
 sg13g2_a21oi_1 _13509_ (.A1(net5947),
    .A2(_04496_),
    .Y(_04497_),
    .B1(net5323));
 sg13g2_o21ai_1 _13510_ (.B1(_04497_),
    .Y(_04498_),
    .A1(net5947),
    .A2(_04494_));
 sg13g2_nand2_1 _13511_ (.Y(_04499_),
    .A(net6085),
    .B(\mem.mem[201][2] ));
 sg13g2_nand2_1 _13512_ (.Y(_04500_),
    .A(net5396),
    .B(\mem.mem[200][2] ));
 sg13g2_nand3_1 _13513_ (.B(_04499_),
    .C(_04500_),
    .A(net5357),
    .Y(_04501_));
 sg13g2_and2_1 _13514_ (.A(net6087),
    .B(\mem.mem[203][2] ),
    .X(_04502_));
 sg13g2_a21oi_1 _13515_ (.A1(net5396),
    .A2(\mem.mem[202][2] ),
    .Y(_04503_),
    .B1(_04502_));
 sg13g2_a21oi_1 _13516_ (.A1(net5943),
    .A2(_04503_),
    .Y(_04504_),
    .B1(net5865));
 sg13g2_a21oi_2 _13517_ (.B1(net5288),
    .Y(_04505_),
    .A2(_04504_),
    .A1(_04501_));
 sg13g2_a221oi_1 _13518_ (.B2(_04505_),
    .C1(net5821),
    .B1(_04498_),
    .A1(net5289),
    .Y(_04506_),
    .A2(_04493_));
 sg13g2_nand2_1 _13519_ (.Y(_04507_),
    .A(net6136),
    .B(\mem.mem[217][2] ));
 sg13g2_nand2_1 _13520_ (.Y(_04508_),
    .A(net5410),
    .B(\mem.mem[216][2] ));
 sg13g2_nand3_1 _13521_ (.B(_04507_),
    .C(_04508_),
    .A(net5366),
    .Y(_04509_));
 sg13g2_and2_1 _13522_ (.A(net6136),
    .B(\mem.mem[219][2] ),
    .X(_04510_));
 sg13g2_a21oi_1 _13523_ (.A1(net5409),
    .A2(\mem.mem[218][2] ),
    .Y(_04511_),
    .B1(_04510_));
 sg13g2_a21oi_1 _13524_ (.A1(net5976),
    .A2(_04511_),
    .Y(_04512_),
    .B1(net5876));
 sg13g2_a21oi_1 _13525_ (.A1(net5409),
    .A2(\mem.mem[220][2] ),
    .Y(_04513_),
    .B1(net5977));
 sg13g2_o21ai_1 _13526_ (.B1(_04513_),
    .Y(_04514_),
    .A1(net5409),
    .A2(_02850_));
 sg13g2_nor2b_1 _13527_ (.A(net6153),
    .B_N(\mem.mem[222][2] ),
    .Y(_04515_));
 sg13g2_a21oi_1 _13528_ (.A1(net6153),
    .A2(\mem.mem[223][2] ),
    .Y(_04516_),
    .B1(_04515_));
 sg13g2_a21oi_2 _13529_ (.B1(net5343),
    .Y(_04517_),
    .A2(_04516_),
    .A1(net5989));
 sg13g2_a221oi_1 _13530_ (.B2(_04517_),
    .C1(net5294),
    .B1(_04514_),
    .A1(_04509_),
    .Y(_04518_),
    .A2(_04512_));
 sg13g2_mux4_1 _13531_ (.S0(net6163),
    .A0(\mem.mem[208][2] ),
    .A1(\mem.mem[209][2] ),
    .A2(\mem.mem[210][2] ),
    .A3(\mem.mem[211][2] ),
    .S1(net5996),
    .X(_04519_));
 sg13g2_nand2_1 _13532_ (.Y(_04520_),
    .A(net6146),
    .B(\mem.mem[213][2] ));
 sg13g2_nand2_1 _13533_ (.Y(_04521_),
    .A(net5412),
    .B(\mem.mem[212][2] ));
 sg13g2_nand3_1 _13534_ (.B(_04520_),
    .C(_04521_),
    .A(net5368),
    .Y(_04522_));
 sg13g2_nor2b_1 _13535_ (.A(net6146),
    .B_N(\mem.mem[214][2] ),
    .Y(_04523_));
 sg13g2_a21oi_1 _13536_ (.A1(net6146),
    .A2(\mem.mem[215][2] ),
    .Y(_04524_),
    .B1(_04523_));
 sg13g2_a21oi_1 _13537_ (.A1(net5984),
    .A2(_04524_),
    .Y(_04525_),
    .B1(net5339));
 sg13g2_a221oi_1 _13538_ (.B2(_04525_),
    .C1(net5844),
    .B1(_04522_),
    .A1(net5337),
    .Y(_04526_),
    .A2(_04519_));
 sg13g2_nor3_2 _13539_ (.A(net5274),
    .B(_04518_),
    .C(_04526_),
    .Y(_04527_));
 sg13g2_or3_1 _13540_ (.A(net5812),
    .B(_04506_),
    .C(_04527_),
    .X(_04528_));
 sg13g2_mux4_1 _13541_ (.S0(net6135),
    .A0(\mem.mem[224][2] ),
    .A1(\mem.mem[225][2] ),
    .A2(\mem.mem[226][2] ),
    .A3(\mem.mem[227][2] ),
    .S1(net5976),
    .X(_04529_));
 sg13g2_nand2_1 _13542_ (.Y(_04530_),
    .A(net6135),
    .B(\mem.mem[229][2] ));
 sg13g2_nand2_1 _13543_ (.Y(_04531_),
    .A(net5410),
    .B(\mem.mem[228][2] ));
 sg13g2_nand3_1 _13544_ (.B(_04530_),
    .C(_04531_),
    .A(net5366),
    .Y(_04532_));
 sg13g2_nor2b_1 _13545_ (.A(net6142),
    .B_N(\mem.mem[230][2] ),
    .Y(_04533_));
 sg13g2_a21oi_1 _13546_ (.A1(net6142),
    .A2(\mem.mem[231][2] ),
    .Y(_04534_),
    .B1(_04533_));
 sg13g2_a21oi_1 _13547_ (.A1(net5976),
    .A2(_04534_),
    .Y(_04535_),
    .B1(net5335));
 sg13g2_a221oi_1 _13548_ (.B2(_04535_),
    .C1(net5844),
    .B1(_04532_),
    .A1(net5336),
    .Y(_04536_),
    .A2(_04529_));
 sg13g2_a21oi_1 _13549_ (.A1(net5414),
    .A2(\mem.mem[236][2] ),
    .Y(_04537_),
    .B1(net5983));
 sg13g2_o21ai_1 _13550_ (.B1(_04537_),
    .Y(_04538_),
    .A1(net5412),
    .A2(_02851_));
 sg13g2_nand2_1 _13551_ (.Y(_04539_),
    .A(net5412),
    .B(\mem.mem[238][2] ));
 sg13g2_a21oi_1 _13552_ (.A1(net6147),
    .A2(\mem.mem[239][2] ),
    .Y(_04540_),
    .B1(net5368));
 sg13g2_a21oi_1 _13553_ (.A1(_04539_),
    .A2(_04540_),
    .Y(_04541_),
    .B1(net5337));
 sg13g2_nand2_1 _13554_ (.Y(_04542_),
    .A(net6140),
    .B(\mem.mem[233][2] ));
 sg13g2_nand2_1 _13555_ (.Y(_04543_),
    .A(net5414),
    .B(\mem.mem[232][2] ));
 sg13g2_nand3_1 _13556_ (.B(_04542_),
    .C(_04543_),
    .A(net5365),
    .Y(_04544_));
 sg13g2_and2_1 _13557_ (.A(net6140),
    .B(\mem.mem[235][2] ),
    .X(_04545_));
 sg13g2_a21oi_1 _13558_ (.A1(net5414),
    .A2(\mem.mem[234][2] ),
    .Y(_04546_),
    .B1(_04545_));
 sg13g2_a21oi_1 _13559_ (.A1(net5979),
    .A2(_04546_),
    .Y(_04547_),
    .B1(net5878));
 sg13g2_a221oi_1 _13560_ (.B2(_04547_),
    .C1(net5293),
    .B1(_04544_),
    .A1(_04538_),
    .Y(_04548_),
    .A2(_04541_));
 sg13g2_or3_2 _13561_ (.A(net5823),
    .B(_04536_),
    .C(_04548_),
    .X(_04549_));
 sg13g2_nand2_1 _13562_ (.Y(_04550_),
    .A(net5312),
    .B(_04480_));
 sg13g2_a21oi_1 _13563_ (.A1(_04478_),
    .A2(_04479_),
    .Y(_04551_),
    .B1(net5314));
 sg13g2_a21oi_1 _13564_ (.A1(_04477_),
    .A2(_04551_),
    .Y(_04552_),
    .B1(net5832));
 sg13g2_nand2_1 _13565_ (.Y(_04553_),
    .A(net5858),
    .B(\mem.mem[252][2] ));
 sg13g2_mux4_1 _13566_ (.S0(net6048),
    .A0(\mem.mem[248][2] ),
    .A1(\mem.mem[249][2] ),
    .A2(\mem.mem[250][2] ),
    .A3(\mem.mem[251][2] ),
    .S1(net5915),
    .X(_04554_));
 sg13g2_a21oi_1 _13567_ (.A1(net5312),
    .A2(_04554_),
    .Y(_04555_),
    .B1(net5281));
 sg13g2_a221oi_1 _13568_ (.B2(_04555_),
    .C1(net5269),
    .B1(_04553_),
    .A1(_04550_),
    .Y(_04556_),
    .A2(_04552_));
 sg13g2_nor2_1 _13569_ (.A(net5265),
    .B(_04556_),
    .Y(_04557_));
 sg13g2_a21oi_1 _13570_ (.A1(_04549_),
    .A2(_04557_),
    .Y(_04558_),
    .B1(net5263));
 sg13g2_a21oi_1 _13571_ (.A1(_04528_),
    .A2(_04558_),
    .Y(_04559_),
    .B1(_02840_));
 sg13g2_a21oi_2 _13572_ (.B1(_02944_),
    .Y(_04560_),
    .A2(_04559_),
    .A1(_04481_));
 sg13g2_a22oi_1 _13573_ (.Y(_04561_),
    .B1(_04383_),
    .B2(_04560_),
    .A2(_03639_),
    .A1(net4));
 sg13g2_o21ai_1 _13574_ (.B1(net6185),
    .Y(_04562_),
    .A1(net5787),
    .A2(net4197));
 sg13g2_a21oi_1 _13575_ (.A1(net5787),
    .A2(_04561_),
    .Y(_00550_),
    .B1(_04562_));
 sg13g2_nand2_1 _13576_ (.Y(_04563_),
    .A(net5372),
    .B(\mem.mem[68][3] ));
 sg13g2_a21oi_1 _13577_ (.A1(net6015),
    .A2(\mem.mem[69][3] ),
    .Y(_04564_),
    .B1(net5892));
 sg13g2_and2_1 _13578_ (.A(net6015),
    .B(\mem.mem[71][3] ),
    .X(_04565_));
 sg13g2_a21oi_1 _13579_ (.A1(net5372),
    .A2(\mem.mem[70][3] ),
    .Y(_04566_),
    .B1(_04565_));
 sg13g2_a221oi_1 _13580_ (.B2(net5892),
    .C1(net5302),
    .B1(_04566_),
    .A1(_04563_),
    .Y(_04567_),
    .A2(_04564_));
 sg13g2_nand2_1 _13581_ (.Y(_04568_),
    .A(net5372),
    .B(\mem.mem[64][3] ));
 sg13g2_a21oi_1 _13582_ (.A1(net6015),
    .A2(\mem.mem[65][3] ),
    .Y(_04569_),
    .B1(net5893));
 sg13g2_nor2b_1 _13583_ (.A(net6016),
    .B_N(\mem.mem[66][3] ),
    .Y(_04570_));
 sg13g2_a21oi_1 _13584_ (.A1(net6016),
    .A2(\mem.mem[67][3] ),
    .Y(_04571_),
    .B1(_04570_));
 sg13g2_a221oi_1 _13585_ (.B2(net5893),
    .C1(net5852),
    .B1(_04571_),
    .A1(_04568_),
    .Y(_04572_),
    .A2(_04569_));
 sg13g2_nor3_2 _13586_ (.A(net5828),
    .B(_04567_),
    .C(_04572_),
    .Y(_04573_));
 sg13g2_mux4_1 _13587_ (.S0(net6021),
    .A0(\mem.mem[72][3] ),
    .A1(\mem.mem[73][3] ),
    .A2(\mem.mem[74][3] ),
    .A3(\mem.mem[75][3] ),
    .S1(net5897),
    .X(_04574_));
 sg13g2_a21oi_1 _13588_ (.A1(net6021),
    .A2(\mem.mem[79][3] ),
    .Y(_04575_),
    .B1(net5349));
 sg13g2_o21ai_1 _13589_ (.B1(_04575_),
    .Y(_04576_),
    .A1(net6021),
    .A2(_02854_));
 sg13g2_nand2_1 _13590_ (.Y(_04577_),
    .A(net6021),
    .B(\mem.mem[77][3] ));
 sg13g2_a21oi_1 _13591_ (.A1(net5374),
    .A2(\mem.mem[76][3] ),
    .Y(_04578_),
    .B1(net5900));
 sg13g2_a21oi_1 _13592_ (.A1(_04577_),
    .A2(_04578_),
    .Y(_04579_),
    .B1(net5303));
 sg13g2_a221oi_1 _13593_ (.B2(_04579_),
    .C1(net5278),
    .B1(_04576_),
    .A1(net5303),
    .Y(_04580_),
    .A2(_04574_));
 sg13g2_nor2_2 _13594_ (.A(_04573_),
    .B(_04580_),
    .Y(_04581_));
 sg13g2_nor2b_1 _13595_ (.A(net6005),
    .B_N(\mem.mem[86][3] ),
    .Y(_04582_));
 sg13g2_a21oi_1 _13596_ (.A1(net6007),
    .A2(\mem.mem[87][3] ),
    .Y(_04583_),
    .B1(_04582_));
 sg13g2_nand2_1 _13597_ (.Y(_04584_),
    .A(net5371),
    .B(\mem.mem[84][3] ));
 sg13g2_a21oi_1 _13598_ (.A1(net6007),
    .A2(\mem.mem[85][3] ),
    .Y(_04585_),
    .B1(net5885));
 sg13g2_a221oi_1 _13599_ (.B2(_04585_),
    .C1(net5298),
    .B1(_04584_),
    .A1(net5885),
    .Y(_04586_),
    .A2(_04583_));
 sg13g2_mux4_1 _13600_ (.S0(net6005),
    .A0(\mem.mem[80][3] ),
    .A1(\mem.mem[81][3] ),
    .A2(\mem.mem[82][3] ),
    .A3(\mem.mem[83][3] ),
    .S1(net5885),
    .X(_04587_));
 sg13g2_a21oi_2 _13601_ (.B1(_04586_),
    .Y(_04588_),
    .A2(_04587_),
    .A1(net5298));
 sg13g2_mux4_1 _13602_ (.S0(net6046),
    .A0(\mem.mem[88][3] ),
    .A1(\mem.mem[89][3] ),
    .A2(\mem.mem[90][3] ),
    .A3(\mem.mem[91][3] ),
    .S1(net5916),
    .X(_04589_));
 sg13g2_nand2_1 _13603_ (.Y(_04590_),
    .A(net5310),
    .B(_04589_));
 sg13g2_nand2_1 _13604_ (.Y(_04591_),
    .A(net6046),
    .B(\mem.mem[93][3] ));
 sg13g2_a21oi_1 _13605_ (.A1(net5386),
    .A2(\mem.mem[92][3] ),
    .Y(_04592_),
    .B1(net5916));
 sg13g2_a21oi_1 _13606_ (.A1(net6051),
    .A2(\mem.mem[95][3] ),
    .Y(_04593_),
    .B1(net5352));
 sg13g2_o21ai_1 _13607_ (.B1(_04593_),
    .Y(_04594_),
    .A1(net6051),
    .A2(_02855_));
 sg13g2_a21oi_1 _13608_ (.A1(_04591_),
    .A2(_04592_),
    .Y(_04595_),
    .B1(net5310));
 sg13g2_a21oi_1 _13609_ (.A1(_04594_),
    .A2(_04595_),
    .Y(_04596_),
    .B1(net5276));
 sg13g2_a22oi_1 _13610_ (.Y(_04597_),
    .B1(_04590_),
    .B2(_04596_),
    .A2(_04588_),
    .A1(net5276));
 sg13g2_nand2_1 _13611_ (.Y(_04598_),
    .A(net5389),
    .B(\mem.mem[100][3] ));
 sg13g2_a21oi_1 _13612_ (.A1(net6071),
    .A2(\mem.mem[101][3] ),
    .Y(_04599_),
    .B1(net5930));
 sg13g2_and2_1 _13613_ (.A(net6071),
    .B(\mem.mem[103][3] ),
    .X(_04600_));
 sg13g2_a21oi_1 _13614_ (.A1(net5389),
    .A2(\mem.mem[102][3] ),
    .Y(_04601_),
    .B1(_04600_));
 sg13g2_a221oi_1 _13615_ (.B2(net5930),
    .C1(net5316),
    .B1(_04601_),
    .A1(_04598_),
    .Y(_04602_),
    .A2(_04599_));
 sg13g2_mux4_1 _13616_ (.S0(net6064),
    .A0(\mem.mem[96][3] ),
    .A1(\mem.mem[97][3] ),
    .A2(\mem.mem[98][3] ),
    .A3(\mem.mem[99][3] ),
    .S1(net5927),
    .X(_04603_));
 sg13g2_nand2_1 _13617_ (.Y(_04604_),
    .A(net5315),
    .B(_04603_));
 sg13g2_nor2_1 _13618_ (.A(net5834),
    .B(_04602_),
    .Y(_04605_));
 sg13g2_nand2_1 _13619_ (.Y(_04606_),
    .A(net5388),
    .B(\mem.mem[104][3] ));
 sg13g2_a21oi_1 _13620_ (.A1(net6063),
    .A2(\mem.mem[105][3] ),
    .Y(_04607_),
    .B1(net5927));
 sg13g2_nor2b_1 _13621_ (.A(net6054),
    .B_N(\mem.mem[106][3] ),
    .Y(_04608_));
 sg13g2_a21oi_1 _13622_ (.A1(net6063),
    .A2(\mem.mem[107][3] ),
    .Y(_04609_),
    .B1(_04608_));
 sg13g2_a221oi_1 _13623_ (.B2(net5927),
    .C1(net5861),
    .B1(_04609_),
    .A1(_04606_),
    .Y(_04610_),
    .A2(_04607_));
 sg13g2_nor2b_1 _13624_ (.A(net6074),
    .B_N(\mem.mem[110][3] ),
    .Y(_04611_));
 sg13g2_a21oi_1 _13625_ (.A1(net6074),
    .A2(\mem.mem[111][3] ),
    .Y(_04612_),
    .B1(_04611_));
 sg13g2_nand2_1 _13626_ (.Y(_04613_),
    .A(net5390),
    .B(\mem.mem[108][3] ));
 sg13g2_a21oi_1 _13627_ (.A1(net6067),
    .A2(\mem.mem[109][3] ),
    .Y(_04614_),
    .B1(net5925));
 sg13g2_a221oi_1 _13628_ (.B2(_04614_),
    .C1(net5315),
    .B1(_04613_),
    .A1(net5925),
    .Y(_04615_),
    .A2(_04612_));
 sg13g2_nor3_2 _13629_ (.A(net5284),
    .B(_04610_),
    .C(_04615_),
    .Y(_04616_));
 sg13g2_a21oi_1 _13630_ (.A1(_04604_),
    .A2(_04605_),
    .Y(_04617_),
    .B1(_04616_));
 sg13g2_nor2b_1 _13631_ (.A(net6024),
    .B_N(\mem.mem[118][3] ),
    .Y(_04618_));
 sg13g2_a21oi_1 _13632_ (.A1(net6024),
    .A2(\mem.mem[119][3] ),
    .Y(_04619_),
    .B1(_04618_));
 sg13g2_nand2_1 _13633_ (.Y(_04620_),
    .A(net5375),
    .B(\mem.mem[116][3] ));
 sg13g2_a21oi_1 _13634_ (.A1(net6023),
    .A2(\mem.mem[117][3] ),
    .Y(_04621_),
    .B1(net5898));
 sg13g2_a221oi_1 _13635_ (.B2(_04621_),
    .C1(net5303),
    .B1(_04620_),
    .A1(net5898),
    .Y(_04622_),
    .A2(_04619_));
 sg13g2_nand2_1 _13636_ (.Y(_04623_),
    .A(net5374),
    .B(\mem.mem[112][3] ));
 sg13g2_a21oi_1 _13637_ (.A1(net6050),
    .A2(\mem.mem[113][3] ),
    .Y(_04624_),
    .B1(net5898));
 sg13g2_nor2b_1 _13638_ (.A(net6051),
    .B_N(\mem.mem[114][3] ),
    .Y(_04625_));
 sg13g2_a21oi_1 _13639_ (.A1(net6050),
    .A2(\mem.mem[115][3] ),
    .Y(_04626_),
    .B1(_04625_));
 sg13g2_a221oi_1 _13640_ (.B2(net5898),
    .C1(net5853),
    .B1(_04626_),
    .A1(_04623_),
    .Y(_04627_),
    .A2(_04624_));
 sg13g2_nor3_2 _13641_ (.A(net5828),
    .B(_04622_),
    .C(_04627_),
    .Y(_04628_));
 sg13g2_nand2_1 _13642_ (.Y(_04629_),
    .A(net5381),
    .B(\mem.mem[120][3] ));
 sg13g2_a21oi_1 _13643_ (.A1(net6043),
    .A2(\mem.mem[121][3] ),
    .Y(_04630_),
    .B1(net5910));
 sg13g2_nor2b_1 _13644_ (.A(net6068),
    .B_N(\mem.mem[122][3] ),
    .Y(_04631_));
 sg13g2_a21oi_1 _13645_ (.A1(net6069),
    .A2(\mem.mem[123][3] ),
    .Y(_04632_),
    .B1(_04631_));
 sg13g2_a221oi_1 _13646_ (.B2(net5910),
    .C1(net5856),
    .B1(_04632_),
    .A1(_04629_),
    .Y(_04633_),
    .A2(_04630_));
 sg13g2_nand2_1 _13647_ (.Y(_04634_),
    .A(net6036),
    .B(\mem.mem[125][3] ));
 sg13g2_a21oi_1 _13648_ (.A1(net5380),
    .A2(\mem.mem[124][3] ),
    .Y(_04635_),
    .B1(net5908));
 sg13g2_and2_1 _13649_ (.A(net6036),
    .B(\mem.mem[127][3] ),
    .X(_04636_));
 sg13g2_a21oi_1 _13650_ (.A1(net5380),
    .A2(\mem.mem[126][3] ),
    .Y(_04637_),
    .B1(_04636_));
 sg13g2_a221oi_1 _13651_ (.B2(net5908),
    .C1(net5306),
    .B1(_04637_),
    .A1(_04634_),
    .Y(_04638_),
    .A2(_04635_));
 sg13g2_nor3_1 _13652_ (.A(net5280),
    .B(_04633_),
    .C(_04638_),
    .Y(_04639_));
 sg13g2_nor2_1 _13653_ (.A(_04628_),
    .B(_04639_),
    .Y(_04640_));
 sg13g2_mux4_1 _13654_ (.S0(net5818),
    .A0(_04581_),
    .A1(_04597_),
    .A2(_04617_),
    .A3(_04640_),
    .S1(net5809),
    .X(_04641_));
 sg13g2_nand2_1 _13655_ (.Y(_04642_),
    .A(net5808),
    .B(_04641_));
 sg13g2_a21oi_1 _13656_ (.A1(net6158),
    .A2(\mem.mem[37][3] ),
    .Y(_04643_),
    .B1(net5992));
 sg13g2_o21ai_1 _13657_ (.B1(_04643_),
    .Y(_04644_),
    .A1(net6158),
    .A2(_02853_));
 sg13g2_and2_1 _13658_ (.A(net6158),
    .B(\mem.mem[39][3] ),
    .X(_04645_));
 sg13g2_a21oi_1 _13659_ (.A1(net5417),
    .A2(\mem.mem[38][3] ),
    .Y(_04646_),
    .B1(_04645_));
 sg13g2_a21oi_1 _13660_ (.A1(net5992),
    .A2(_04646_),
    .Y(_04647_),
    .B1(net5341));
 sg13g2_mux4_1 _13661_ (.S0(net6159),
    .A0(\mem.mem[32][3] ),
    .A1(\mem.mem[33][3] ),
    .A2(\mem.mem[34][3] ),
    .A3(\mem.mem[35][3] ),
    .S1(net5993),
    .X(_04648_));
 sg13g2_a221oi_1 _13662_ (.B2(net5342),
    .C1(net5846),
    .B1(_04648_),
    .A1(_04644_),
    .Y(_04649_),
    .A2(_04647_));
 sg13g2_nand2_1 _13663_ (.Y(_04650_),
    .A(net5420),
    .B(\mem.mem[40][3] ));
 sg13g2_a21oi_1 _13664_ (.A1(net6171),
    .A2(\mem.mem[41][3] ),
    .Y(_04651_),
    .B1(net6002));
 sg13g2_nor2b_1 _13665_ (.A(net6171),
    .B_N(\mem.mem[42][3] ),
    .Y(_04652_));
 sg13g2_a21oi_1 _13666_ (.A1(net6171),
    .A2(\mem.mem[43][3] ),
    .Y(_04653_),
    .B1(_04652_));
 sg13g2_a221oi_1 _13667_ (.B2(net6002),
    .C1(net5882),
    .B1(_04653_),
    .A1(_04650_),
    .Y(_04654_),
    .A2(_04651_));
 sg13g2_nor2b_1 _13668_ (.A(net6164),
    .B_N(\mem.mem[46][3] ),
    .Y(_04655_));
 sg13g2_a21oi_1 _13669_ (.A1(net6171),
    .A2(\mem.mem[47][3] ),
    .Y(_04656_),
    .B1(_04655_));
 sg13g2_nand2_1 _13670_ (.Y(_04657_),
    .A(net5421),
    .B(\mem.mem[44][3] ));
 sg13g2_a21oi_1 _13671_ (.A1(net6171),
    .A2(\mem.mem[45][3] ),
    .Y(_04658_),
    .B1(net6001));
 sg13g2_a221oi_1 _13672_ (.B2(_04658_),
    .C1(net5345),
    .B1(_04657_),
    .A1(net6001),
    .Y(_04659_),
    .A2(_04656_));
 sg13g2_nor3_2 _13673_ (.A(net5295),
    .B(_04654_),
    .C(_04659_),
    .Y(_04660_));
 sg13g2_o21ai_1 _13674_ (.B1(net5273),
    .Y(_04661_),
    .A1(_04649_),
    .A2(_04660_));
 sg13g2_nor2b_1 _13675_ (.A(net6027),
    .B_N(\mem.mem[54][3] ),
    .Y(_04662_));
 sg13g2_a21oi_1 _13676_ (.A1(net6026),
    .A2(\mem.mem[55][3] ),
    .Y(_04663_),
    .B1(_04662_));
 sg13g2_nand2_1 _13677_ (.Y(_04664_),
    .A(net5379),
    .B(\mem.mem[52][3] ));
 sg13g2_a21oi_1 _13678_ (.A1(net6027),
    .A2(\mem.mem[53][3] ),
    .Y(_04665_),
    .B1(net5902));
 sg13g2_a221oi_1 _13679_ (.B2(_04665_),
    .C1(net5304),
    .B1(_04664_),
    .A1(net5901),
    .Y(_04666_),
    .A2(_04663_));
 sg13g2_nand2_1 _13680_ (.Y(_04667_),
    .A(net5370),
    .B(\mem.mem[48][3] ));
 sg13g2_a21oi_1 _13681_ (.A1(net6011),
    .A2(\mem.mem[49][3] ),
    .Y(_04668_),
    .B1(net5889));
 sg13g2_nor2b_1 _13682_ (.A(net6010),
    .B_N(\mem.mem[50][3] ),
    .Y(_04669_));
 sg13g2_a21oi_1 _13683_ (.A1(net6010),
    .A2(\mem.mem[51][3] ),
    .Y(_04670_),
    .B1(_04669_));
 sg13g2_a221oi_1 _13684_ (.B2(net5889),
    .C1(net5851),
    .B1(_04670_),
    .A1(_04667_),
    .Y(_04671_),
    .A2(_04668_));
 sg13g2_nor3_1 _13685_ (.A(net5829),
    .B(_04666_),
    .C(_04671_),
    .Y(_04672_));
 sg13g2_nand2_1 _13686_ (.Y(_04673_),
    .A(net5378),
    .B(\mem.mem[56][3] ));
 sg13g2_a21oi_1 _13687_ (.A1(net6032),
    .A2(\mem.mem[57][3] ),
    .Y(_04674_),
    .B1(net5905));
 sg13g2_nor2b_1 _13688_ (.A(net6032),
    .B_N(\mem.mem[58][3] ),
    .Y(_04675_));
 sg13g2_a21oi_1 _13689_ (.A1(net6032),
    .A2(\mem.mem[59][3] ),
    .Y(_04676_),
    .B1(_04675_));
 sg13g2_a221oi_1 _13690_ (.B2(net5905),
    .C1(net5854),
    .B1(_04676_),
    .A1(_04673_),
    .Y(_04677_),
    .A2(_04674_));
 sg13g2_nand2_1 _13691_ (.Y(_04678_),
    .A(net6038),
    .B(\mem.mem[61][3] ));
 sg13g2_a21oi_1 _13692_ (.A1(net5381),
    .A2(\mem.mem[60][3] ),
    .Y(_04679_),
    .B1(net5912));
 sg13g2_and2_1 _13693_ (.A(net6038),
    .B(\mem.mem[63][3] ),
    .X(_04680_));
 sg13g2_a21oi_1 _13694_ (.A1(net5381),
    .A2(\mem.mem[62][3] ),
    .Y(_04681_),
    .B1(_04680_));
 sg13g2_a221oi_1 _13695_ (.B2(net5912),
    .C1(net5307),
    .B1(_04681_),
    .A1(_04678_),
    .Y(_04682_),
    .A2(_04679_));
 sg13g2_nor3_2 _13696_ (.A(net5279),
    .B(_04677_),
    .C(_04682_),
    .Y(_04683_));
 sg13g2_o21ai_1 _13697_ (.B1(net5817),
    .Y(_04684_),
    .A1(_04672_),
    .A2(_04683_));
 sg13g2_nand3_1 _13698_ (.B(_04661_),
    .C(_04684_),
    .A(net5811),
    .Y(_04685_));
 sg13g2_nand2_1 _13699_ (.Y(_04686_),
    .A(net5391),
    .B(\mem.mem[4][3] ));
 sg13g2_a21oi_1 _13700_ (.A1(net6078),
    .A2(\mem.mem[5][3] ),
    .Y(_04687_),
    .B1(net5934));
 sg13g2_and2_1 _13701_ (.A(net6075),
    .B(\mem.mem[7][3] ),
    .X(_04688_));
 sg13g2_a21oi_1 _13702_ (.A1(net5391),
    .A2(\mem.mem[6][3] ),
    .Y(_04689_),
    .B1(_04688_));
 sg13g2_a221oi_1 _13703_ (.B2(net5934),
    .C1(net5320),
    .B1(_04689_),
    .A1(_04686_),
    .Y(_04690_),
    .A2(_04687_));
 sg13g2_nand2_1 _13704_ (.Y(_04691_),
    .A(net5393),
    .B(\mem.mem[0][3] ));
 sg13g2_a21oi_1 _13705_ (.A1(net6079),
    .A2(\mem.mem[1][3] ),
    .Y(_04692_),
    .B1(net5936));
 sg13g2_nor2b_1 _13706_ (.A(net6079),
    .B_N(\mem.mem[2][3] ),
    .Y(_04693_));
 sg13g2_a21oi_1 _13707_ (.A1(net6079),
    .A2(\mem.mem[3][3] ),
    .Y(_04694_),
    .B1(_04693_));
 sg13g2_a221oi_1 _13708_ (.B2(net5936),
    .C1(net5862),
    .B1(_04694_),
    .A1(_04691_),
    .Y(_04695_),
    .A2(_04692_));
 sg13g2_nor3_1 _13709_ (.A(net5835),
    .B(_04690_),
    .C(_04695_),
    .Y(_04696_));
 sg13g2_nand2_1 _13710_ (.Y(_04697_),
    .A(net5393),
    .B(\mem.mem[8][3] ));
 sg13g2_a21oi_1 _13711_ (.A1(net6081),
    .A2(\mem.mem[9][3] ),
    .Y(_04698_),
    .B1(net5938));
 sg13g2_nor2b_1 _13712_ (.A(net6082),
    .B_N(\mem.mem[10][3] ),
    .Y(_04699_));
 sg13g2_a21oi_1 _13713_ (.A1(net6081),
    .A2(\mem.mem[11][3] ),
    .Y(_04700_),
    .B1(_04699_));
 sg13g2_a221oi_1 _13714_ (.B2(net5938),
    .C1(net5862),
    .B1(_04700_),
    .A1(_04697_),
    .Y(_04701_),
    .A2(_04698_));
 sg13g2_nor2b_1 _13715_ (.A(net6111),
    .B_N(\mem.mem[14][3] ),
    .Y(_04702_));
 sg13g2_a21oi_1 _13716_ (.A1(net6111),
    .A2(\mem.mem[15][3] ),
    .Y(_04703_),
    .B1(_04702_));
 sg13g2_nand2_1 _13717_ (.Y(_04704_),
    .A(net5403),
    .B(\mem.mem[12][3] ));
 sg13g2_a21oi_1 _13718_ (.A1(net6110),
    .A2(\mem.mem[13][3] ),
    .Y(_04705_),
    .B1(net5961));
 sg13g2_a221oi_1 _13719_ (.B2(_04705_),
    .C1(net5330),
    .B1(_04704_),
    .A1(net5958),
    .Y(_04706_),
    .A2(_04703_));
 sg13g2_nor3_1 _13720_ (.A(net5283),
    .B(_04701_),
    .C(_04706_),
    .Y(_04707_));
 sg13g2_o21ai_1 _13721_ (.B1(net5268),
    .Y(_04708_),
    .A1(_04696_),
    .A2(_04707_));
 sg13g2_nor2b_1 _13722_ (.A(net6126),
    .B_N(\mem.mem[22][3] ),
    .Y(_04709_));
 sg13g2_a21oi_1 _13723_ (.A1(net6126),
    .A2(\mem.mem[23][3] ),
    .Y(_04710_),
    .B1(_04709_));
 sg13g2_nand2_1 _13724_ (.Y(_04711_),
    .A(net5406),
    .B(\mem.mem[20][3] ));
 sg13g2_a21oi_1 _13725_ (.A1(net6126),
    .A2(\mem.mem[21][3] ),
    .Y(_04712_),
    .B1(net5969));
 sg13g2_a221oi_1 _13726_ (.B2(_04712_),
    .C1(net5331),
    .B1(_04711_),
    .A1(net5969),
    .Y(_04713_),
    .A2(_04710_));
 sg13g2_nand2_1 _13727_ (.Y(_04714_),
    .A(net5417),
    .B(\mem.mem[16][3] ));
 sg13g2_a21oi_1 _13728_ (.A1(net6156),
    .A2(\mem.mem[17][3] ),
    .Y(_04715_),
    .B1(net5991));
 sg13g2_nor2b_1 _13729_ (.A(net6156),
    .B_N(\mem.mem[18][3] ),
    .Y(_04716_));
 sg13g2_a21oi_1 _13730_ (.A1(net6157),
    .A2(\mem.mem[19][3] ),
    .Y(_04717_),
    .B1(_04716_));
 sg13g2_a221oi_1 _13731_ (.B2(net5991),
    .C1(net5880),
    .B1(_04717_),
    .A1(_04714_),
    .Y(_04718_),
    .A2(_04715_));
 sg13g2_nor3_2 _13732_ (.A(net5848),
    .B(_04713_),
    .C(_04718_),
    .Y(_04719_));
 sg13g2_nand2_1 _13733_ (.Y(_04720_),
    .A(net5416),
    .B(\mem.mem[24][3] ));
 sg13g2_a21oi_1 _13734_ (.A1(net6155),
    .A2(\mem.mem[25][3] ),
    .Y(_04721_),
    .B1(net5990));
 sg13g2_nor2b_1 _13735_ (.A(net6155),
    .B_N(\mem.mem[26][3] ),
    .Y(_04722_));
 sg13g2_a21oi_1 _13736_ (.A1(net6155),
    .A2(\mem.mem[27][3] ),
    .Y(_04723_),
    .B1(_04722_));
 sg13g2_a221oi_1 _13737_ (.B2(net5990),
    .C1(net5880),
    .B1(_04723_),
    .A1(_04720_),
    .Y(_04724_),
    .A2(_04721_));
 sg13g2_nand2_1 _13738_ (.Y(_04725_),
    .A(net6155),
    .B(\mem.mem[29][3] ));
 sg13g2_a21oi_1 _13739_ (.A1(net5416),
    .A2(\mem.mem[28][3] ),
    .Y(_04726_),
    .B1(net5990));
 sg13g2_and2_1 _13740_ (.A(net6155),
    .B(\mem.mem[31][3] ),
    .X(_04727_));
 sg13g2_a21oi_1 _13741_ (.A1(net5416),
    .A2(\mem.mem[30][3] ),
    .Y(_04728_),
    .B1(_04727_));
 sg13g2_a221oi_1 _13742_ (.B2(net5990),
    .C1(net5341),
    .B1(_04728_),
    .A1(_04725_),
    .Y(_04729_),
    .A2(_04726_));
 sg13g2_nor3_1 _13743_ (.A(net5295),
    .B(_04724_),
    .C(_04729_),
    .Y(_04730_));
 sg13g2_o21ai_1 _13744_ (.B1(net5824),
    .Y(_04731_),
    .A1(_04719_),
    .A2(_04730_));
 sg13g2_nand3_1 _13745_ (.B(_04708_),
    .C(_04731_),
    .A(net5267),
    .Y(_04732_));
 sg13g2_a21o_2 _13746_ (.A2(_04732_),
    .A1(_04685_),
    .B1(net5807),
    .X(_04733_));
 sg13g2_nand3_1 _13747_ (.B(_04642_),
    .C(_04733_),
    .A(_02840_),
    .Y(_04734_));
 sg13g2_mux2_1 _13748_ (.A0(\mem.mem[140][3] ),
    .A1(\mem.mem[141][3] ),
    .S(net6110),
    .X(_04735_));
 sg13g2_nand2_1 _13749_ (.Y(_04736_),
    .A(net5361),
    .B(_04735_));
 sg13g2_mux2_1 _13750_ (.A0(\mem.mem[142][3] ),
    .A1(\mem.mem[143][3] ),
    .S(net6110),
    .X(_04737_));
 sg13g2_a21oi_1 _13751_ (.A1(net5958),
    .A2(_04737_),
    .Y(_04738_),
    .B1(net5329));
 sg13g2_mux4_1 _13752_ (.S0(net6114),
    .A0(\mem.mem[136][3] ),
    .A1(\mem.mem[137][3] ),
    .A2(\mem.mem[138][3] ),
    .A3(\mem.mem[139][3] ),
    .S1(net5960),
    .X(_04739_));
 sg13g2_a21oi_1 _13753_ (.A1(_04736_),
    .A2(_04738_),
    .Y(_04740_),
    .B1(net5290));
 sg13g2_o21ai_1 _13754_ (.B1(_04740_),
    .Y(_04741_),
    .A1(net5870),
    .A2(_04739_));
 sg13g2_mux4_1 _13755_ (.S0(net6117),
    .A0(\mem.mem[128][3] ),
    .A1(\mem.mem[129][3] ),
    .A2(\mem.mem[130][3] ),
    .A3(\mem.mem[131][3] ),
    .S1(net5965),
    .X(_04742_));
 sg13g2_nand2b_1 _13756_ (.Y(_04743_),
    .B(net5332),
    .A_N(_04742_));
 sg13g2_mux2_1 _13757_ (.A0(\mem.mem[132][3] ),
    .A1(\mem.mem[133][3] ),
    .S(net6116),
    .X(_04744_));
 sg13g2_nand2_1 _13758_ (.Y(_04745_),
    .A(net5362),
    .B(_04744_));
 sg13g2_mux2_1 _13759_ (.A0(\mem.mem[134][3] ),
    .A1(\mem.mem[135][3] ),
    .S(net6116),
    .X(_04746_));
 sg13g2_a21oi_1 _13760_ (.A1(net5963),
    .A2(_04746_),
    .Y(_04747_),
    .B1(net5332));
 sg13g2_a21oi_1 _13761_ (.A1(_04745_),
    .A2(_04747_),
    .Y(_04748_),
    .B1(net5840));
 sg13g2_a21oi_1 _13762_ (.A1(_04743_),
    .A2(_04748_),
    .Y(_04749_),
    .B1(net5822));
 sg13g2_nor2b_1 _13763_ (.A(\mem.mem[151][3] ),
    .B_N(net6112),
    .Y(_04750_));
 sg13g2_o21ai_1 _13764_ (.B1(net5955),
    .Y(_04751_),
    .A1(net6105),
    .A2(\mem.mem[150][3] ));
 sg13g2_mux2_1 _13765_ (.A0(\mem.mem[148][3] ),
    .A1(\mem.mem[149][3] ),
    .S(net6106),
    .X(_04752_));
 sg13g2_o21ai_1 _13766_ (.B1(net5870),
    .Y(_04753_),
    .A1(_04750_),
    .A2(_04751_));
 sg13g2_a21oi_1 _13767_ (.A1(net5361),
    .A2(_04752_),
    .Y(_04754_),
    .B1(_04753_));
 sg13g2_mux2_1 _13768_ (.A0(\mem.mem[146][3] ),
    .A1(\mem.mem[147][3] ),
    .S(net6076),
    .X(_04755_));
 sg13g2_nand2b_1 _13769_ (.Y(_04756_),
    .B(net6076),
    .A_N(\mem.mem[145][3] ));
 sg13g2_a21oi_1 _13770_ (.A1(net5392),
    .A2(_02856_),
    .Y(_04757_),
    .B1(net5934));
 sg13g2_a221oi_1 _13771_ (.B2(_04757_),
    .C1(net5863),
    .B1(_04756_),
    .A1(net5933),
    .Y(_04758_),
    .A2(_04755_));
 sg13g2_or3_1 _13772_ (.A(net5841),
    .B(_04754_),
    .C(_04758_),
    .X(_04759_));
 sg13g2_mux4_1 _13773_ (.S0(net6093),
    .A0(\mem.mem[152][3] ),
    .A1(\mem.mem[153][3] ),
    .A2(\mem.mem[154][3] ),
    .A3(\mem.mem[155][3] ),
    .S1(net5948),
    .X(_04760_));
 sg13g2_nand2b_1 _13774_ (.Y(_04761_),
    .B(net5328),
    .A_N(_04760_));
 sg13g2_mux2_1 _13775_ (.A0(\mem.mem[156][3] ),
    .A1(\mem.mem[157][3] ),
    .S(net6107),
    .X(_04762_));
 sg13g2_nand2_1 _13776_ (.Y(_04763_),
    .A(net5361),
    .B(_04762_));
 sg13g2_mux2_1 _13777_ (.A0(\mem.mem[158][3] ),
    .A1(\mem.mem[159][3] ),
    .S(net6107),
    .X(_04764_));
 sg13g2_a21oi_1 _13778_ (.A1(net5957),
    .A2(_04764_),
    .Y(_04765_),
    .B1(net5328));
 sg13g2_a21oi_1 _13779_ (.A1(_04763_),
    .A2(_04765_),
    .Y(_04766_),
    .B1(net5290));
 sg13g2_a21oi_1 _13780_ (.A1(_04761_),
    .A2(_04766_),
    .Y(_04767_),
    .B1(net5271));
 sg13g2_a221oi_1 _13781_ (.B2(_04767_),
    .C1(net5814),
    .B1(_04759_),
    .A1(_04741_),
    .Y(_04768_),
    .A2(_04749_));
 sg13g2_mux2_1 _13782_ (.A0(\mem.mem[170][3] ),
    .A1(\mem.mem[171][3] ),
    .S(net6085),
    .X(_04769_));
 sg13g2_nand2_1 _13783_ (.Y(_04770_),
    .A(net5945),
    .B(_04769_));
 sg13g2_mux2_1 _13784_ (.A0(\mem.mem[168][3] ),
    .A1(\mem.mem[169][3] ),
    .S(net6085),
    .X(_04771_));
 sg13g2_a21oi_1 _13785_ (.A1(net5357),
    .A2(_04771_),
    .Y(_04772_),
    .B1(net5865));
 sg13g2_mux2_1 _13786_ (.A0(\mem.mem[172][3] ),
    .A1(\mem.mem[173][3] ),
    .S(net6094),
    .X(_04773_));
 sg13g2_nor2_1 _13787_ (.A(net6090),
    .B(\mem.mem[174][3] ),
    .Y(_04774_));
 sg13g2_o21ai_1 _13788_ (.B1(net5946),
    .Y(_04775_),
    .A1(net5397),
    .A2(\mem.mem[175][3] ));
 sg13g2_a21oi_1 _13789_ (.A1(net5360),
    .A2(_04773_),
    .Y(_04776_),
    .B1(net5323));
 sg13g2_o21ai_1 _13790_ (.B1(_04776_),
    .Y(_04777_),
    .A1(_04774_),
    .A2(_04775_));
 sg13g2_a21oi_1 _13791_ (.A1(_04770_),
    .A2(_04772_),
    .Y(_04778_),
    .B1(net5288));
 sg13g2_mux4_1 _13792_ (.S0(net6085),
    .A0(\mem.mem[160][3] ),
    .A1(\mem.mem[161][3] ),
    .A2(\mem.mem[162][3] ),
    .A3(\mem.mem[163][3] ),
    .S1(net5943),
    .X(_04779_));
 sg13g2_nand2b_1 _13793_ (.Y(_04780_),
    .B(net5324),
    .A_N(_04779_));
 sg13g2_mux2_1 _13794_ (.A0(\mem.mem[166][3] ),
    .A1(\mem.mem[167][3] ),
    .S(net6060),
    .X(_04781_));
 sg13g2_nand2_1 _13795_ (.Y(_04782_),
    .A(net5920),
    .B(_04781_));
 sg13g2_mux2_1 _13796_ (.A0(\mem.mem[164][3] ),
    .A1(\mem.mem[165][3] ),
    .S(net6056),
    .X(_04783_));
 sg13g2_a21oi_1 _13797_ (.A1(net5353),
    .A2(_04783_),
    .Y(_04784_),
    .B1(net5313));
 sg13g2_a21oi_2 _13798_ (.B1(net5832),
    .Y(_04785_),
    .A2(_04784_),
    .A1(_04782_));
 sg13g2_a221oi_1 _13799_ (.B2(_04785_),
    .C1(net5821),
    .B1(_04780_),
    .A1(_04777_),
    .Y(_04786_),
    .A2(_04778_));
 sg13g2_mux4_1 _13800_ (.S0(net6132),
    .A0(\mem.mem[176][3] ),
    .A1(\mem.mem[177][3] ),
    .A2(\mem.mem[178][3] ),
    .A3(\mem.mem[179][3] ),
    .S1(net5973),
    .X(_04787_));
 sg13g2_nor2_2 _13801_ (.A(net5875),
    .B(_04787_),
    .Y(_04788_));
 sg13g2_mux2_1 _13802_ (.A0(\mem.mem[182][3] ),
    .A1(\mem.mem[183][3] ),
    .S(net6135),
    .X(_04789_));
 sg13g2_nand2_1 _13803_ (.Y(_04790_),
    .A(net5976),
    .B(_04789_));
 sg13g2_mux2_1 _13804_ (.A0(\mem.mem[180][3] ),
    .A1(\mem.mem[181][3] ),
    .S(net6132),
    .X(_04791_));
 sg13g2_a21oi_1 _13805_ (.A1(net5366),
    .A2(_04791_),
    .Y(_04792_),
    .B1(net5335));
 sg13g2_a21oi_2 _13806_ (.B1(_04788_),
    .Y(_04793_),
    .A2(_04792_),
    .A1(_04790_));
 sg13g2_mux2_1 _13807_ (.A0(\mem.mem[188][3] ),
    .A1(\mem.mem[189][3] ),
    .S(net6102),
    .X(_04794_));
 sg13g2_nor2_1 _13808_ (.A(net6103),
    .B(\mem.mem[190][3] ),
    .Y(_04795_));
 sg13g2_o21ai_1 _13809_ (.B1(net5954),
    .Y(_04796_),
    .A1(net5400),
    .A2(\mem.mem[191][3] ));
 sg13g2_a21oi_1 _13810_ (.A1(net5358),
    .A2(_04794_),
    .Y(_04797_),
    .B1(net5325));
 sg13g2_o21ai_1 _13811_ (.B1(_04797_),
    .Y(_04798_),
    .A1(_04795_),
    .A2(_04796_));
 sg13g2_mux2_1 _13812_ (.A0(\mem.mem[186][3] ),
    .A1(\mem.mem[187][3] ),
    .S(net6097),
    .X(_04799_));
 sg13g2_nand2_1 _13813_ (.Y(_04800_),
    .A(net5950),
    .B(_04799_));
 sg13g2_mux2_1 _13814_ (.A0(\mem.mem[184][3] ),
    .A1(\mem.mem[185][3] ),
    .S(net6096),
    .X(_04801_));
 sg13g2_a21oi_1 _13815_ (.A1(net5359),
    .A2(_04801_),
    .Y(_04802_),
    .B1(net5875));
 sg13g2_a21oi_1 _13816_ (.A1(_04800_),
    .A2(_04802_),
    .Y(_04803_),
    .B1(net5289));
 sg13g2_a221oi_1 _13817_ (.B2(_04803_),
    .C1(net5273),
    .B1(_04798_),
    .A1(net5289),
    .Y(_04804_),
    .A2(_04793_));
 sg13g2_nor3_2 _13818_ (.A(net5265),
    .B(_04786_),
    .C(_04804_),
    .Y(_04805_));
 sg13g2_nor3_1 _13819_ (.A(net5807),
    .B(_04768_),
    .C(_04805_),
    .Y(_04806_));
 sg13g2_mux4_1 _13820_ (.S0(net6153),
    .A0(\mem.mem[220][3] ),
    .A1(\mem.mem[221][3] ),
    .A2(\mem.mem[222][3] ),
    .A3(\mem.mem[223][3] ),
    .S1(net5989),
    .X(_04807_));
 sg13g2_nor2_1 _13821_ (.A(net5343),
    .B(_04807_),
    .Y(_04808_));
 sg13g2_mux4_1 _13822_ (.S0(net6134),
    .A0(\mem.mem[216][3] ),
    .A1(\mem.mem[217][3] ),
    .A2(\mem.mem[218][3] ),
    .A3(\mem.mem[219][3] ),
    .S1(net5977),
    .X(_04809_));
 sg13g2_o21ai_1 _13823_ (.B1(net5845),
    .Y(_04810_),
    .A1(net5876),
    .A2(_04809_));
 sg13g2_mux4_1 _13824_ (.S0(net6147),
    .A0(\mem.mem[212][3] ),
    .A1(\mem.mem[213][3] ),
    .A2(\mem.mem[214][3] ),
    .A3(\mem.mem[215][3] ),
    .S1(net5983),
    .X(_04811_));
 sg13g2_mux4_1 _13825_ (.S0(net6163),
    .A0(\mem.mem[208][3] ),
    .A1(\mem.mem[209][3] ),
    .A2(\mem.mem[210][3] ),
    .A3(\mem.mem[211][3] ),
    .S1(net5996),
    .X(_04812_));
 sg13g2_mux2_1 _13826_ (.A0(_04811_),
    .A1(_04812_),
    .S(net5337),
    .X(_04813_));
 sg13g2_a21oi_2 _13827_ (.B1(net5274),
    .Y(_04814_),
    .A2(_04813_),
    .A1(net5293));
 sg13g2_o21ai_1 _13828_ (.B1(_04814_),
    .Y(_04815_),
    .A1(_04808_),
    .A2(_04810_));
 sg13g2_mux4_1 _13829_ (.S0(net6096),
    .A0(\mem.mem[196][3] ),
    .A1(\mem.mem[197][3] ),
    .A2(\mem.mem[198][3] ),
    .A3(\mem.mem[199][3] ),
    .S1(net5950),
    .X(_04816_));
 sg13g2_nor2_1 _13830_ (.A(net5326),
    .B(_04816_),
    .Y(_04817_));
 sg13g2_mux4_1 _13831_ (.S0(net6095),
    .A0(\mem.mem[192][3] ),
    .A1(\mem.mem[193][3] ),
    .A2(\mem.mem[194][3] ),
    .A3(\mem.mem[195][3] ),
    .S1(net5951),
    .X(_04818_));
 sg13g2_o21ai_1 _13832_ (.B1(net5289),
    .Y(_04819_),
    .A1(net5867),
    .A2(_04818_));
 sg13g2_mux2_1 _13833_ (.A0(\mem.mem[204][3] ),
    .A1(\mem.mem[205][3] ),
    .S(net6087),
    .X(_04820_));
 sg13g2_nand2_1 _13834_ (.Y(_04821_),
    .A(net5357),
    .B(_04820_));
 sg13g2_mux2_1 _13835_ (.A0(\mem.mem[206][3] ),
    .A1(\mem.mem[207][3] ),
    .S(net6088),
    .X(_04822_));
 sg13g2_a21oi_1 _13836_ (.A1(net5945),
    .A2(_04822_),
    .Y(_04823_),
    .B1(net5324));
 sg13g2_mux4_1 _13837_ (.S0(net6085),
    .A0(\mem.mem[200][3] ),
    .A1(\mem.mem[201][3] ),
    .A2(\mem.mem[202][3] ),
    .A3(\mem.mem[203][3] ),
    .S1(net5943),
    .X(_04824_));
 sg13g2_o21ai_1 _13838_ (.B1(net5838),
    .Y(_04825_),
    .A1(net5865),
    .A2(_04824_));
 sg13g2_a21oi_1 _13839_ (.A1(_04821_),
    .A2(_04823_),
    .Y(_04826_),
    .B1(_04825_));
 sg13g2_o21ai_1 _13840_ (.B1(net5272),
    .Y(_04827_),
    .A1(_04817_),
    .A2(_04819_));
 sg13g2_nor2_1 _13841_ (.A(_04826_),
    .B(_04827_),
    .Y(_04828_));
 sg13g2_nor2_1 _13842_ (.A(net5812),
    .B(_04828_),
    .Y(_04829_));
 sg13g2_nand2b_1 _13843_ (.Y(_04830_),
    .B(net6143),
    .A_N(\mem.mem[237][3] ));
 sg13g2_o21ai_1 _13844_ (.B1(_04830_),
    .Y(_04831_),
    .A1(net6142),
    .A2(\mem.mem[236][3] ));
 sg13g2_mux2_1 _13845_ (.A0(\mem.mem[238][3] ),
    .A1(\mem.mem[239][3] ),
    .S(net6143),
    .X(_04832_));
 sg13g2_a21oi_1 _13846_ (.A1(net5981),
    .A2(_04832_),
    .Y(_04833_),
    .B1(net5338));
 sg13g2_o21ai_1 _13847_ (.B1(_04833_),
    .Y(_04834_),
    .A1(net5981),
    .A2(_04831_));
 sg13g2_mux4_1 _13848_ (.S0(net6141),
    .A0(\mem.mem[232][3] ),
    .A1(\mem.mem[233][3] ),
    .A2(\mem.mem[234][3] ),
    .A3(\mem.mem[235][3] ),
    .S1(net5979),
    .X(_04835_));
 sg13g2_o21ai_1 _13849_ (.B1(net5843),
    .Y(_04836_),
    .A1(net5877),
    .A2(_04835_));
 sg13g2_inv_1 _13850_ (.Y(_04837_),
    .A(_04836_));
 sg13g2_nand2b_1 _13851_ (.Y(_04838_),
    .B(net6142),
    .A_N(\mem.mem[231][3] ));
 sg13g2_o21ai_1 _13852_ (.B1(_04838_),
    .Y(_04839_),
    .A1(net6142),
    .A2(\mem.mem[230][3] ));
 sg13g2_mux2_1 _13853_ (.A0(\mem.mem[228][3] ),
    .A1(\mem.mem[229][3] ),
    .S(net6143),
    .X(_04840_));
 sg13g2_a21oi_1 _13854_ (.A1(net5366),
    .A2(_04840_),
    .Y(_04841_),
    .B1(net5338));
 sg13g2_o21ai_1 _13855_ (.B1(_04841_),
    .Y(_04842_),
    .A1(net5366),
    .A2(_04839_));
 sg13g2_mux2_1 _13856_ (.A0(\mem.mem[226][3] ),
    .A1(\mem.mem[227][3] ),
    .S(net6139),
    .X(_04843_));
 sg13g2_nand2_1 _13857_ (.Y(_04844_),
    .A(net5981),
    .B(_04843_));
 sg13g2_mux2_1 _13858_ (.A0(\mem.mem[224][3] ),
    .A1(\mem.mem[225][3] ),
    .S(net6142),
    .X(_04845_));
 sg13g2_a21oi_1 _13859_ (.A1(net5365),
    .A2(_04845_),
    .Y(_04846_),
    .B1(net5879));
 sg13g2_a21oi_1 _13860_ (.A1(_04844_),
    .A2(_04846_),
    .Y(_04847_),
    .B1(net5843));
 sg13g2_a221oi_1 _13861_ (.B2(_04847_),
    .C1(net5823),
    .B1(_04842_),
    .A1(_04834_),
    .Y(_04848_),
    .A2(_04837_));
 sg13g2_mux4_1 _13862_ (.S0(net6048),
    .A0(\mem.mem[248][3] ),
    .A1(\mem.mem[249][3] ),
    .A2(\mem.mem[250][3] ),
    .A3(\mem.mem[251][3] ),
    .S1(net5915),
    .X(_04849_));
 sg13g2_nand2_1 _13863_ (.Y(_04850_),
    .A(net5831),
    .B(_04849_));
 sg13g2_mux4_1 _13864_ (.S0(net6048),
    .A0(\mem.mem[240][3] ),
    .A1(\mem.mem[241][3] ),
    .A2(\mem.mem[242][3] ),
    .A3(\mem.mem[243][3] ),
    .S1(net5915),
    .X(_04851_));
 sg13g2_nand2_1 _13865_ (.Y(_04852_),
    .A(net5281),
    .B(_04851_));
 sg13g2_a21oi_1 _13866_ (.A1(_04850_),
    .A2(_04852_),
    .Y(_04853_),
    .B1(net5859));
 sg13g2_nor2_1 _13867_ (.A(net5282),
    .B(\mem.mem[252][3] ),
    .Y(_04854_));
 sg13g2_mux4_1 _13868_ (.S0(net6052),
    .A0(\mem.mem[244][3] ),
    .A1(\mem.mem[245][3] ),
    .A2(\mem.mem[246][3] ),
    .A3(\mem.mem[247][3] ),
    .S1(net5922),
    .X(_04855_));
 sg13g2_o21ai_1 _13869_ (.B1(net5858),
    .Y(_04856_),
    .A1(net5832),
    .A2(_04855_));
 sg13g2_o21ai_1 _13870_ (.B1(net5820),
    .Y(_04857_),
    .A1(_04854_),
    .A2(_04856_));
 sg13g2_o21ai_1 _13871_ (.B1(net5811),
    .Y(_04858_),
    .A1(_04853_),
    .A2(_04857_));
 sg13g2_o21ai_1 _13872_ (.B1(net5807),
    .Y(_04859_),
    .A1(_04848_),
    .A2(_04858_));
 sg13g2_a21oi_2 _13873_ (.B1(_04859_),
    .Y(_04860_),
    .A2(_04829_),
    .A1(_04815_));
 sg13g2_o21ai_1 _13874_ (.B1(_00007_),
    .Y(_04861_),
    .A1(_04806_),
    .A2(_04860_));
 sg13g2_and2_1 _13875_ (.A(_02945_),
    .B(_04861_),
    .X(_04862_));
 sg13g2_a22oi_1 _13876_ (.Y(_04863_),
    .B1(_04734_),
    .B2(_04862_),
    .A2(_03639_),
    .A1(net5));
 sg13g2_o21ai_1 _13877_ (.B1(net6185),
    .Y(_04864_),
    .A1(net5787),
    .A2(net4181));
 sg13g2_a21oi_1 _13878_ (.A1(net5789),
    .A2(_04863_),
    .Y(_00551_),
    .B1(_04864_));
 sg13g2_nand2_1 _13879_ (.Y(_04865_),
    .A(net6015),
    .B(\mem.mem[69][4] ));
 sg13g2_nand2_1 _13880_ (.Y(_04866_),
    .A(net5371),
    .B(\mem.mem[68][4] ));
 sg13g2_nand3_1 _13881_ (.B(_04865_),
    .C(_04866_),
    .A(net5349),
    .Y(_04867_));
 sg13g2_and2_1 _13882_ (.A(net6015),
    .B(\mem.mem[71][4] ),
    .X(_04868_));
 sg13g2_a21oi_1 _13883_ (.A1(net5372),
    .A2(\mem.mem[70][4] ),
    .Y(_04869_),
    .B1(_04868_));
 sg13g2_a21oi_1 _13884_ (.A1(net5892),
    .A2(_04869_),
    .Y(_04870_),
    .B1(net5298));
 sg13g2_mux4_1 _13885_ (.S0(net6006),
    .A0(\mem.mem[64][4] ),
    .A1(\mem.mem[65][4] ),
    .A2(\mem.mem[66][4] ),
    .A3(\mem.mem[67][4] ),
    .S1(net5886),
    .X(_04871_));
 sg13g2_a221oi_1 _13886_ (.B2(net5298),
    .C1(net5827),
    .B1(_04871_),
    .A1(_04867_),
    .Y(_04872_),
    .A2(_04870_));
 sg13g2_mux4_1 _13887_ (.S0(net6021),
    .A0(\mem.mem[72][4] ),
    .A1(\mem.mem[73][4] ),
    .A2(\mem.mem[74][4] ),
    .A3(\mem.mem[75][4] ),
    .S1(net5897),
    .X(_04873_));
 sg13g2_mux4_1 _13888_ (.S0(net6013),
    .A0(\mem.mem[76][4] ),
    .A1(\mem.mem[77][4] ),
    .A2(\mem.mem[78][4] ),
    .A3(\mem.mem[79][4] ),
    .S1(net5890),
    .X(_04874_));
 sg13g2_a21o_1 _13889_ (.A2(_04874_),
    .A1(net5851),
    .B1(net5278),
    .X(_04875_));
 sg13g2_a21oi_1 _13890_ (.A1(net5300),
    .A2(_04873_),
    .Y(_04876_),
    .B1(_04875_));
 sg13g2_o21ai_1 _13891_ (.B1(net5270),
    .Y(_04877_),
    .A1(_04872_),
    .A2(_04876_));
 sg13g2_mux4_1 _13892_ (.S0(net6019),
    .A0(\mem.mem[88][4] ),
    .A1(\mem.mem[89][4] ),
    .A2(\mem.mem[90][4] ),
    .A3(\mem.mem[91][4] ),
    .S1(net5895),
    .X(_04878_));
 sg13g2_mux4_1 _13893_ (.S0(net6019),
    .A0(\mem.mem[92][4] ),
    .A1(\mem.mem[93][4] ),
    .A2(\mem.mem[94][4] ),
    .A3(\mem.mem[95][4] ),
    .S1(net5895),
    .X(_04879_));
 sg13g2_a21o_1 _13894_ (.A2(_04879_),
    .A1(net5852),
    .B1(net5276),
    .X(_04880_));
 sg13g2_a21oi_1 _13895_ (.A1(net5302),
    .A2(_04878_),
    .Y(_04881_),
    .B1(_04880_));
 sg13g2_mux4_1 _13896_ (.S0(net6006),
    .A0(\mem.mem[80][4] ),
    .A1(\mem.mem[81][4] ),
    .A2(\mem.mem[82][4] ),
    .A3(\mem.mem[83][4] ),
    .S1(net5887),
    .X(_04882_));
 sg13g2_and2_1 _13897_ (.A(net6012),
    .B(\mem.mem[87][4] ),
    .X(_04883_));
 sg13g2_a21oi_1 _13898_ (.A1(net5370),
    .A2(\mem.mem[86][4] ),
    .Y(_04884_),
    .B1(_04883_));
 sg13g2_nand2_1 _13899_ (.Y(_04885_),
    .A(net6012),
    .B(\mem.mem[85][4] ));
 sg13g2_nand2_1 _13900_ (.Y(_04886_),
    .A(net5370),
    .B(\mem.mem[84][4] ));
 sg13g2_nand3_1 _13901_ (.B(_04885_),
    .C(_04886_),
    .A(net5349),
    .Y(_04887_));
 sg13g2_a21oi_1 _13902_ (.A1(net5890),
    .A2(_04884_),
    .Y(_04888_),
    .B1(net5300));
 sg13g2_a221oi_1 _13903_ (.B2(_04888_),
    .C1(net5827),
    .B1(_04887_),
    .A1(net5300),
    .Y(_04889_),
    .A2(_04882_));
 sg13g2_o21ai_1 _13904_ (.B1(net5816),
    .Y(_04890_),
    .A1(_04881_),
    .A2(_04889_));
 sg13g2_nand3_1 _13905_ (.B(_04877_),
    .C(_04890_),
    .A(net5264),
    .Y(_04891_));
 sg13g2_nor2b_1 _13906_ (.A(net6071),
    .B_N(\mem.mem[102][4] ),
    .Y(_04892_));
 sg13g2_a21oi_1 _13907_ (.A1(net6072),
    .A2(\mem.mem[103][4] ),
    .Y(_04893_),
    .B1(_04892_));
 sg13g2_nand2_1 _13908_ (.Y(_04894_),
    .A(net5389),
    .B(\mem.mem[100][4] ));
 sg13g2_a21oi_1 _13909_ (.A1(net6072),
    .A2(\mem.mem[101][4] ),
    .Y(_04895_),
    .B1(net5930));
 sg13g2_a221oi_1 _13910_ (.B2(_04895_),
    .C1(net5316),
    .B1(_04894_),
    .A1(net5930),
    .Y(_04896_),
    .A2(_04893_));
 sg13g2_nand2_1 _13911_ (.Y(_04897_),
    .A(net5388),
    .B(\mem.mem[96][4] ));
 sg13g2_a21oi_1 _13912_ (.A1(net6066),
    .A2(\mem.mem[97][4] ),
    .Y(_04898_),
    .B1(net5926));
 sg13g2_nor2b_1 _13913_ (.A(net6066),
    .B_N(\mem.mem[98][4] ),
    .Y(_04899_));
 sg13g2_a21oi_1 _13914_ (.A1(net6066),
    .A2(\mem.mem[99][4] ),
    .Y(_04900_),
    .B1(_04899_));
 sg13g2_a221oi_1 _13915_ (.B2(net5926),
    .C1(net5861),
    .B1(_04900_),
    .A1(_04897_),
    .Y(_04901_),
    .A2(_04898_));
 sg13g2_nor3_1 _13916_ (.A(net5833),
    .B(_04896_),
    .C(_04901_),
    .Y(_04902_));
 sg13g2_mux4_1 _13917_ (.S0(net6063),
    .A0(\mem.mem[104][4] ),
    .A1(\mem.mem[105][4] ),
    .A2(\mem.mem[106][4] ),
    .A3(\mem.mem[107][4] ),
    .S1(net5927),
    .X(_04903_));
 sg13g2_nand2_1 _13918_ (.Y(_04904_),
    .A(net6065),
    .B(\mem.mem[109][4] ));
 sg13g2_a21oi_1 _13919_ (.A1(net5388),
    .A2(\mem.mem[108][4] ),
    .Y(_04905_),
    .B1(net5925));
 sg13g2_a21oi_1 _13920_ (.A1(net6074),
    .A2(\mem.mem[111][4] ),
    .Y(_04906_),
    .B1(net5355));
 sg13g2_o21ai_1 _13921_ (.B1(_04906_),
    .Y(_04907_),
    .A1(net6065),
    .A2(_02861_));
 sg13g2_a21oi_1 _13922_ (.A1(_04904_),
    .A2(_04905_),
    .Y(_04908_),
    .B1(net5315));
 sg13g2_a221oi_1 _13923_ (.B2(_04908_),
    .C1(net5284),
    .B1(_04907_),
    .A1(net5315),
    .Y(_04909_),
    .A2(_04903_));
 sg13g2_o21ai_1 _13924_ (.B1(net5268),
    .Y(_04910_),
    .A1(_04902_),
    .A2(_04909_));
 sg13g2_a21oi_1 _13925_ (.A1(net6035),
    .A2(\mem.mem[117][4] ),
    .Y(_04911_),
    .B1(net5908));
 sg13g2_o21ai_1 _13926_ (.B1(_04911_),
    .Y(_04912_),
    .A1(net6035),
    .A2(_02862_));
 sg13g2_and2_1 _13927_ (.A(net6036),
    .B(\mem.mem[119][4] ),
    .X(_04913_));
 sg13g2_a21oi_1 _13928_ (.A1(net5380),
    .A2(\mem.mem[118][4] ),
    .Y(_04914_),
    .B1(_04913_));
 sg13g2_a21oi_1 _13929_ (.A1(net5908),
    .A2(_04914_),
    .Y(_04915_),
    .B1(net5306));
 sg13g2_mux4_1 _13930_ (.S0(net6063),
    .A0(\mem.mem[112][4] ),
    .A1(\mem.mem[113][4] ),
    .A2(\mem.mem[114][4] ),
    .A3(\mem.mem[115][4] ),
    .S1(net5927),
    .X(_04916_));
 sg13g2_a221oi_1 _13931_ (.B2(net5306),
    .C1(net5830),
    .B1(_04916_),
    .A1(_04912_),
    .Y(_04917_),
    .A2(_04915_));
 sg13g2_nand2_1 _13932_ (.Y(_04918_),
    .A(net5381),
    .B(\mem.mem[120][4] ));
 sg13g2_a21oi_1 _13933_ (.A1(net6042),
    .A2(\mem.mem[121][4] ),
    .Y(_04919_),
    .B1(net5911));
 sg13g2_nor2b_1 _13934_ (.A(net6042),
    .B_N(\mem.mem[122][4] ),
    .Y(_04920_));
 sg13g2_a21oi_1 _13935_ (.A1(net6042),
    .A2(\mem.mem[123][4] ),
    .Y(_04921_),
    .B1(_04920_));
 sg13g2_a221oi_1 _13936_ (.B2(net5911),
    .C1(net5855),
    .B1(_04921_),
    .A1(_04918_),
    .Y(_04922_),
    .A2(_04919_));
 sg13g2_nor2b_1 _13937_ (.A(net6041),
    .B_N(\mem.mem[126][4] ),
    .Y(_04923_));
 sg13g2_a21oi_1 _13938_ (.A1(net6041),
    .A2(\mem.mem[127][4] ),
    .Y(_04924_),
    .B1(_04923_));
 sg13g2_nand2_1 _13939_ (.Y(_04925_),
    .A(net5382),
    .B(\mem.mem[124][4] ));
 sg13g2_a21oi_1 _13940_ (.A1(net6041),
    .A2(\mem.mem[125][4] ),
    .Y(_04926_),
    .B1(net5911));
 sg13g2_a221oi_1 _13941_ (.B2(_04926_),
    .C1(net5307),
    .B1(_04925_),
    .A1(net5911),
    .Y(_04927_),
    .A2(_04924_));
 sg13g2_nor3_2 _13942_ (.A(net5280),
    .B(_04922_),
    .C(_04927_),
    .Y(_04928_));
 sg13g2_o21ai_1 _13943_ (.B1(net5817),
    .Y(_04929_),
    .A1(_04917_),
    .A2(_04928_));
 sg13g2_nand3_1 _13944_ (.B(_04910_),
    .C(_04929_),
    .A(net5809),
    .Y(_04930_));
 sg13g2_a21oi_1 _13945_ (.A1(_04891_),
    .A2(_04930_),
    .Y(_04931_),
    .B1(net5262));
 sg13g2_nor2b_1 _13946_ (.A(net6159),
    .B_N(\mem.mem[38][4] ),
    .Y(_04932_));
 sg13g2_a21oi_1 _13947_ (.A1(net6158),
    .A2(\mem.mem[39][4] ),
    .Y(_04933_),
    .B1(_04932_));
 sg13g2_a21oi_1 _13948_ (.A1(net6158),
    .A2(\mem.mem[37][4] ),
    .Y(_04934_),
    .B1(net5992));
 sg13g2_o21ai_1 _13949_ (.B1(_04934_),
    .Y(_04935_),
    .A1(net6158),
    .A2(_02859_));
 sg13g2_a21oi_1 _13950_ (.A1(net5992),
    .A2(_04933_),
    .Y(_04936_),
    .B1(net5341));
 sg13g2_mux4_1 _13951_ (.S0(net6159),
    .A0(\mem.mem[32][4] ),
    .A1(\mem.mem[33][4] ),
    .A2(\mem.mem[34][4] ),
    .A3(\mem.mem[35][4] ),
    .S1(net5993),
    .X(_04937_));
 sg13g2_a221oi_1 _13952_ (.B2(net5341),
    .C1(net5846),
    .B1(_04937_),
    .A1(_04935_),
    .Y(_04938_),
    .A2(_04936_));
 sg13g2_nand2_1 _13953_ (.Y(_04939_),
    .A(net5420),
    .B(\mem.mem[40][4] ));
 sg13g2_a21oi_1 _13954_ (.A1(net6170),
    .A2(\mem.mem[41][4] ),
    .Y(_04940_),
    .B1(net6001));
 sg13g2_nor2b_1 _13955_ (.A(net6170),
    .B_N(\mem.mem[42][4] ),
    .Y(_04941_));
 sg13g2_a21oi_1 _13956_ (.A1(net6170),
    .A2(\mem.mem[43][4] ),
    .Y(_04942_),
    .B1(_04941_));
 sg13g2_a221oi_1 _13957_ (.B2(net5999),
    .C1(net5881),
    .B1(_04942_),
    .A1(_04939_),
    .Y(_04943_),
    .A2(_04940_));
 sg13g2_nand2_1 _13958_ (.Y(_04944_),
    .A(net6164),
    .B(\mem.mem[45][4] ));
 sg13g2_a21oi_1 _13959_ (.A1(net5421),
    .A2(\mem.mem[44][4] ),
    .Y(_04945_),
    .B1(net5997));
 sg13g2_and2_1 _13960_ (.A(net6165),
    .B(\mem.mem[47][4] ),
    .X(_04946_));
 sg13g2_a21oi_1 _13961_ (.A1(net5419),
    .A2(\mem.mem[46][4] ),
    .Y(_04947_),
    .B1(_04946_));
 sg13g2_a221oi_1 _13962_ (.B2(net5997),
    .C1(net5344),
    .B1(_04947_),
    .A1(_04944_),
    .Y(_04948_),
    .A2(_04945_));
 sg13g2_nor3_2 _13963_ (.A(net5295),
    .B(_04943_),
    .C(_04948_),
    .Y(_04949_));
 sg13g2_o21ai_1 _13964_ (.B1(net5273),
    .Y(_04950_),
    .A1(_04938_),
    .A2(_04949_));
 sg13g2_a21oi_1 _13965_ (.A1(net6027),
    .A2(\mem.mem[53][4] ),
    .Y(_04951_),
    .B1(net5902));
 sg13g2_o21ai_1 _13966_ (.B1(_04951_),
    .Y(_04952_),
    .A1(net6026),
    .A2(_02860_));
 sg13g2_and2_1 _13967_ (.A(net6028),
    .B(\mem.mem[55][4] ),
    .X(_04953_));
 sg13g2_a21oi_1 _13968_ (.A1(net5379),
    .A2(\mem.mem[54][4] ),
    .Y(_04954_),
    .B1(_04953_));
 sg13g2_a21oi_1 _13969_ (.A1(net5901),
    .A2(_04954_),
    .Y(_04955_),
    .B1(net5305));
 sg13g2_mux4_1 _13970_ (.S0(net6028),
    .A0(\mem.mem[48][4] ),
    .A1(\mem.mem[49][4] ),
    .A2(\mem.mem[50][4] ),
    .A3(\mem.mem[51][4] ),
    .S1(net5901),
    .X(_04956_));
 sg13g2_a221oi_1 _13971_ (.B2(net5305),
    .C1(net5829),
    .B1(_04956_),
    .A1(_04952_),
    .Y(_04957_),
    .A2(_04955_));
 sg13g2_nand2_1 _13972_ (.Y(_04958_),
    .A(net5377),
    .B(\mem.mem[56][4] ));
 sg13g2_a21oi_1 _13973_ (.A1(net6029),
    .A2(\mem.mem[57][4] ),
    .Y(_04959_),
    .B1(net5904));
 sg13g2_nor2b_1 _13974_ (.A(net6029),
    .B_N(\mem.mem[58][4] ),
    .Y(_04960_));
 sg13g2_a21oi_1 _13975_ (.A1(net6029),
    .A2(\mem.mem[59][4] ),
    .Y(_04961_),
    .B1(_04960_));
 sg13g2_a221oi_1 _13976_ (.B2(net5904),
    .C1(net5854),
    .B1(_04961_),
    .A1(_04958_),
    .Y(_04962_),
    .A2(_04959_));
 sg13g2_nor2b_1 _13977_ (.A(net6032),
    .B_N(\mem.mem[62][4] ),
    .Y(_04963_));
 sg13g2_a21oi_1 _13978_ (.A1(net6031),
    .A2(\mem.mem[63][4] ),
    .Y(_04964_),
    .B1(_04963_));
 sg13g2_nand2_1 _13979_ (.Y(_04965_),
    .A(net5378),
    .B(\mem.mem[60][4] ));
 sg13g2_a21oi_1 _13980_ (.A1(net6031),
    .A2(\mem.mem[61][4] ),
    .Y(_04966_),
    .B1(net5905));
 sg13g2_a221oi_1 _13981_ (.B2(_04966_),
    .C1(net5304),
    .B1(_04965_),
    .A1(net5906),
    .Y(_04967_),
    .A2(_04964_));
 sg13g2_nor3_2 _13982_ (.A(net5279),
    .B(_04962_),
    .C(_04967_),
    .Y(_04968_));
 sg13g2_o21ai_1 _13983_ (.B1(net5817),
    .Y(_04969_),
    .A1(_04957_),
    .A2(_04968_));
 sg13g2_nand3_1 _13984_ (.B(_04950_),
    .C(_04969_),
    .A(net5809),
    .Y(_04970_));
 sg13g2_nand2_1 _13985_ (.Y(_04971_),
    .A(net5393),
    .B(\mem.mem[4][4] ));
 sg13g2_a21oi_1 _13986_ (.A1(net6075),
    .A2(\mem.mem[5][4] ),
    .Y(_04972_),
    .B1(net5937));
 sg13g2_and2_1 _13987_ (.A(net6074),
    .B(\mem.mem[7][4] ),
    .X(_04973_));
 sg13g2_a21oi_1 _13988_ (.A1(net5391),
    .A2(\mem.mem[6][4] ),
    .Y(_04974_),
    .B1(_04973_));
 sg13g2_a221oi_1 _13989_ (.B2(net5937),
    .C1(net5318),
    .B1(_04974_),
    .A1(_04971_),
    .Y(_04975_),
    .A2(_04972_));
 sg13g2_nand2_1 _13990_ (.Y(_04976_),
    .A(net5393),
    .B(\mem.mem[0][4] ));
 sg13g2_a21oi_1 _13991_ (.A1(net6080),
    .A2(\mem.mem[1][4] ),
    .Y(_04977_),
    .B1(net5936));
 sg13g2_nor2b_1 _13992_ (.A(net6079),
    .B_N(\mem.mem[2][4] ),
    .Y(_04978_));
 sg13g2_a21oi_1 _13993_ (.A1(net6079),
    .A2(\mem.mem[3][4] ),
    .Y(_04979_),
    .B1(_04978_));
 sg13g2_a221oi_1 _13994_ (.B2(net5936),
    .C1(net5862),
    .B1(_04979_),
    .A1(_04976_),
    .Y(_04980_),
    .A2(_04977_));
 sg13g2_nor3_1 _13995_ (.A(net5835),
    .B(_04975_),
    .C(_04980_),
    .Y(_04981_));
 sg13g2_nand2_1 _13996_ (.Y(_04982_),
    .A(net5393),
    .B(\mem.mem[8][4] ));
 sg13g2_a21oi_1 _13997_ (.A1(net6082),
    .A2(\mem.mem[9][4] ),
    .Y(_04983_),
    .B1(net5939));
 sg13g2_nor2b_1 _13998_ (.A(net6082),
    .B_N(\mem.mem[10][4] ),
    .Y(_04984_));
 sg13g2_a21oi_1 _13999_ (.A1(net6082),
    .A2(\mem.mem[11][4] ),
    .Y(_04985_),
    .B1(_04984_));
 sg13g2_a221oi_1 _14000_ (.B2(net5936),
    .C1(net5862),
    .B1(_04985_),
    .A1(_04982_),
    .Y(_04986_),
    .A2(_04983_));
 sg13g2_nor2b_1 _14001_ (.A(net6110),
    .B_N(\mem.mem[14][4] ),
    .Y(_04987_));
 sg13g2_a21oi_1 _14002_ (.A1(net6110),
    .A2(\mem.mem[15][4] ),
    .Y(_04988_),
    .B1(_04987_));
 sg13g2_nand2_1 _14003_ (.Y(_04989_),
    .A(net5393),
    .B(\mem.mem[12][4] ));
 sg13g2_a21oi_1 _14004_ (.A1(net6110),
    .A2(\mem.mem[13][4] ),
    .Y(_04990_),
    .B1(net5939));
 sg13g2_a221oi_1 _14005_ (.B2(_04990_),
    .C1(net5319),
    .B1(_04989_),
    .A1(net5939),
    .Y(_04991_),
    .A2(_04988_));
 sg13g2_nor3_2 _14006_ (.A(net5283),
    .B(_04986_),
    .C(_04991_),
    .Y(_04992_));
 sg13g2_o21ai_1 _14007_ (.B1(net5268),
    .Y(_04993_),
    .A1(_04981_),
    .A2(_04992_));
 sg13g2_nor2b_1 _14008_ (.A(net6127),
    .B_N(\mem.mem[22][4] ),
    .Y(_04994_));
 sg13g2_a21oi_1 _14009_ (.A1(net6127),
    .A2(\mem.mem[23][4] ),
    .Y(_04995_),
    .B1(_04994_));
 sg13g2_a21oi_1 _14010_ (.A1(net6126),
    .A2(\mem.mem[21][4] ),
    .Y(_04996_),
    .B1(net5969));
 sg13g2_o21ai_1 _14011_ (.B1(_04996_),
    .Y(_04997_),
    .A1(net6126),
    .A2(_02858_));
 sg13g2_a21oi_1 _14012_ (.A1(net5969),
    .A2(_04995_),
    .Y(_04998_),
    .B1(net5331));
 sg13g2_mux4_1 _14013_ (.S0(net6156),
    .A0(\mem.mem[16][4] ),
    .A1(\mem.mem[17][4] ),
    .A2(\mem.mem[18][4] ),
    .A3(\mem.mem[19][4] ),
    .S1(net5991),
    .X(_04999_));
 sg13g2_a221oi_1 _14014_ (.B2(net5331),
    .C1(net5846),
    .B1(_04999_),
    .A1(_04997_),
    .Y(_05000_),
    .A2(_04998_));
 sg13g2_nand2_1 _14015_ (.Y(_05001_),
    .A(net5406),
    .B(\mem.mem[24][4] ));
 sg13g2_a21oi_1 _14016_ (.A1(net6125),
    .A2(\mem.mem[25][4] ),
    .Y(_05002_),
    .B1(net5968));
 sg13g2_nor2b_1 _14017_ (.A(net6119),
    .B_N(\mem.mem[26][4] ),
    .Y(_05003_));
 sg13g2_a21oi_1 _14018_ (.A1(net6119),
    .A2(\mem.mem[27][4] ),
    .Y(_05004_),
    .B1(_05003_));
 sg13g2_a221oi_1 _14019_ (.B2(net5968),
    .C1(net5873),
    .B1(_05004_),
    .A1(_05001_),
    .Y(_05005_),
    .A2(_05002_));
 sg13g2_nand2_1 _14020_ (.Y(_05006_),
    .A(net6155),
    .B(\mem.mem[29][4] ));
 sg13g2_a21oi_1 _14021_ (.A1(net5416),
    .A2(\mem.mem[28][4] ),
    .Y(_05007_),
    .B1(net5990));
 sg13g2_and2_1 _14022_ (.A(net6155),
    .B(\mem.mem[31][4] ),
    .X(_05008_));
 sg13g2_a21oi_1 _14023_ (.A1(net5416),
    .A2(\mem.mem[30][4] ),
    .Y(_05009_),
    .B1(_05008_));
 sg13g2_a221oi_1 _14024_ (.B2(net5990),
    .C1(net5341),
    .B1(_05009_),
    .A1(_05006_),
    .Y(_05010_),
    .A2(_05007_));
 sg13g2_nor3_1 _14025_ (.A(net5291),
    .B(_05005_),
    .C(_05010_),
    .Y(_05011_));
 sg13g2_o21ai_1 _14026_ (.B1(net5824),
    .Y(_05012_),
    .A1(_05000_),
    .A2(_05011_));
 sg13g2_nand3_1 _14027_ (.B(_04993_),
    .C(_05012_),
    .A(net5267),
    .Y(_05013_));
 sg13g2_a21oi_1 _14028_ (.A1(_04970_),
    .A2(_05013_),
    .Y(_05014_),
    .B1(net5808));
 sg13g2_nor3_1 _14029_ (.A(_00007_),
    .B(_04931_),
    .C(_05014_),
    .Y(_05015_));
 sg13g2_mux4_1 _14030_ (.S0(net6133),
    .A0(\mem.mem[224][4] ),
    .A1(\mem.mem[225][4] ),
    .A2(\mem.mem[226][4] ),
    .A3(\mem.mem[227][4] ),
    .S1(net5973),
    .X(_05016_));
 sg13g2_mux4_1 _14031_ (.S0(net6139),
    .A0(\mem.mem[228][4] ),
    .A1(\mem.mem[229][4] ),
    .A2(\mem.mem[230][4] ),
    .A3(\mem.mem[231][4] ),
    .S1(net5980),
    .X(_05017_));
 sg13g2_nand2_1 _14032_ (.Y(_05018_),
    .A(net5877),
    .B(_05017_));
 sg13g2_a21oi_1 _14033_ (.A1(net5334),
    .A2(_05016_),
    .Y(_05019_),
    .B1(net5843));
 sg13g2_nor2b_1 _14034_ (.A(net6139),
    .B_N(\mem.mem[234][4] ),
    .Y(_05020_));
 sg13g2_a21oi_1 _14035_ (.A1(net6139),
    .A2(\mem.mem[235][4] ),
    .Y(_05021_),
    .B1(_05020_));
 sg13g2_mux2_1 _14036_ (.A0(\mem.mem[232][4] ),
    .A1(\mem.mem[233][4] ),
    .S(net6138),
    .X(_05022_));
 sg13g2_a21oi_1 _14037_ (.A1(net5980),
    .A2(_05021_),
    .Y(_05023_),
    .B1(net5877));
 sg13g2_o21ai_1 _14038_ (.B1(_05023_),
    .Y(_05024_),
    .A1(net5978),
    .A2(_05022_));
 sg13g2_mux4_1 _14039_ (.S0(net6143),
    .A0(\mem.mem[236][4] ),
    .A1(\mem.mem[237][4] ),
    .A2(\mem.mem[238][4] ),
    .A3(\mem.mem[239][4] ),
    .S1(net5981),
    .X(_05025_));
 sg13g2_a21oi_1 _14040_ (.A1(net5879),
    .A2(_05025_),
    .Y(_05026_),
    .B1(net5294));
 sg13g2_mux4_1 _14041_ (.S0(net6053),
    .A0(\mem.mem[244][4] ),
    .A1(\mem.mem[245][4] ),
    .A2(\mem.mem[246][4] ),
    .A3(\mem.mem[247][4] ),
    .S1(net5919),
    .X(_05027_));
 sg13g2_nand2_1 _14042_ (.Y(_05028_),
    .A(net5859),
    .B(_05027_));
 sg13g2_mux4_1 _14043_ (.S0(net6055),
    .A0(\mem.mem[240][4] ),
    .A1(\mem.mem[241][4] ),
    .A2(\mem.mem[242][4] ),
    .A3(\mem.mem[243][4] ),
    .S1(net5921),
    .X(_05029_));
 sg13g2_a21oi_1 _14044_ (.A1(net5312),
    .A2(_05029_),
    .Y(_05030_),
    .B1(net5831));
 sg13g2_mux4_1 _14045_ (.S0(net6049),
    .A0(\mem.mem[248][4] ),
    .A1(\mem.mem[249][4] ),
    .A2(\mem.mem[250][4] ),
    .A3(\mem.mem[251][4] ),
    .S1(net5916),
    .X(_05031_));
 sg13g2_nand2_1 _14046_ (.Y(_05032_),
    .A(net5859),
    .B(\mem.mem[252][4] ));
 sg13g2_a21oi_1 _14047_ (.A1(net5310),
    .A2(_05031_),
    .Y(_05033_),
    .B1(net5281));
 sg13g2_a221oi_1 _14048_ (.B2(_05026_),
    .C1(net5823),
    .B1(_05024_),
    .A1(_05018_),
    .Y(_05034_),
    .A2(_05019_));
 sg13g2_a221oi_1 _14049_ (.B2(_05033_),
    .C1(net5269),
    .B1(_05032_),
    .A1(_05028_),
    .Y(_05035_),
    .A2(_05030_));
 sg13g2_o21ai_1 _14050_ (.B1(net5813),
    .Y(_05036_),
    .A1(_05034_),
    .A2(_05035_));
 sg13g2_mux2_1 _14051_ (.A0(\mem.mem[202][4] ),
    .A1(\mem.mem[203][4] ),
    .S(net6087),
    .X(_05037_));
 sg13g2_nand2_1 _14052_ (.Y(_05038_),
    .A(net5944),
    .B(_05037_));
 sg13g2_mux2_1 _14053_ (.A0(\mem.mem[200][4] ),
    .A1(\mem.mem[201][4] ),
    .S(net6088),
    .X(_05039_));
 sg13g2_a21oi_1 _14054_ (.A1(net5357),
    .A2(_05039_),
    .Y(_05040_),
    .B1(net5865));
 sg13g2_a21oi_1 _14055_ (.A1(net5396),
    .A2(_02863_),
    .Y(_05041_),
    .B1(net5944));
 sg13g2_o21ai_1 _14056_ (.B1(_05041_),
    .Y(_05042_),
    .A1(net5396),
    .A2(\mem.mem[205][4] ));
 sg13g2_mux2_1 _14057_ (.A0(\mem.mem[206][4] ),
    .A1(\mem.mem[207][4] ),
    .S(net6087),
    .X(_05043_));
 sg13g2_a21oi_1 _14058_ (.A1(net5944),
    .A2(_05043_),
    .Y(_05044_),
    .B1(net5324));
 sg13g2_a221oi_1 _14059_ (.B2(_05044_),
    .C1(net5288),
    .B1(_05042_),
    .A1(_05038_),
    .Y(_05045_),
    .A2(_05040_));
 sg13g2_mux2_1 _14060_ (.A0(\mem.mem[198][4] ),
    .A1(\mem.mem[199][4] ),
    .S(net6098),
    .X(_05046_));
 sg13g2_mux2_1 _14061_ (.A0(\mem.mem[196][4] ),
    .A1(\mem.mem[197][4] ),
    .S(net6095),
    .X(_05047_));
 sg13g2_nand2_1 _14062_ (.Y(_05048_),
    .A(net5359),
    .B(_05047_));
 sg13g2_a21oi_1 _14063_ (.A1(net5951),
    .A2(_05046_),
    .Y(_05049_),
    .B1(net5326));
 sg13g2_mux2_1 _14064_ (.A0(\mem.mem[194][4] ),
    .A1(\mem.mem[195][4] ),
    .S(net6095),
    .X(_05050_));
 sg13g2_nand2_1 _14065_ (.Y(_05051_),
    .A(net5951),
    .B(_05050_));
 sg13g2_mux2_1 _14066_ (.A0(\mem.mem[192][4] ),
    .A1(\mem.mem[193][4] ),
    .S(net6099),
    .X(_05052_));
 sg13g2_a21oi_1 _14067_ (.A1(net5359),
    .A2(_05052_),
    .Y(_05053_),
    .B1(net5868));
 sg13g2_a221oi_1 _14068_ (.B2(_05053_),
    .C1(net5839),
    .B1(_05051_),
    .A1(_05048_),
    .Y(_05054_),
    .A2(_05049_));
 sg13g2_nor3_1 _14069_ (.A(net5821),
    .B(_05045_),
    .C(_05054_),
    .Y(_05055_));
 sg13g2_nand2_1 _14070_ (.Y(_05056_),
    .A(net5413),
    .B(\mem.mem[212][4] ));
 sg13g2_a21oi_1 _14071_ (.A1(net6146),
    .A2(\mem.mem[213][4] ),
    .Y(_05057_),
    .B1(net5996));
 sg13g2_and2_1 _14072_ (.A(net6146),
    .B(\mem.mem[215][4] ),
    .X(_05058_));
 sg13g2_a21oi_1 _14073_ (.A1(net5413),
    .A2(\mem.mem[214][4] ),
    .Y(_05059_),
    .B1(_05058_));
 sg13g2_a221oi_1 _14074_ (.B2(net5984),
    .C1(net5337),
    .B1(_05059_),
    .A1(_05056_),
    .Y(_05060_),
    .A2(_05057_));
 sg13g2_nand2_1 _14075_ (.Y(_05061_),
    .A(net5419),
    .B(\mem.mem[208][4] ));
 sg13g2_a21oi_1 _14076_ (.A1(net6164),
    .A2(\mem.mem[209][4] ),
    .Y(_05062_),
    .B1(net5996));
 sg13g2_nor2b_1 _14077_ (.A(net6163),
    .B_N(\mem.mem[210][4] ),
    .Y(_05063_));
 sg13g2_a21oi_1 _14078_ (.A1(net6163),
    .A2(\mem.mem[211][4] ),
    .Y(_05064_),
    .B1(_05063_));
 sg13g2_a221oi_1 _14079_ (.B2(net5996),
    .C1(net5882),
    .B1(_05064_),
    .A1(_05061_),
    .Y(_05065_),
    .A2(_05062_));
 sg13g2_nor3_2 _14080_ (.A(net5847),
    .B(_05060_),
    .C(_05065_),
    .Y(_05066_));
 sg13g2_mux4_1 _14081_ (.S0(net6151),
    .A0(\mem.mem[216][4] ),
    .A1(\mem.mem[217][4] ),
    .A2(\mem.mem[218][4] ),
    .A3(\mem.mem[219][4] ),
    .S1(net5988),
    .X(_05067_));
 sg13g2_a21oi_1 _14082_ (.A1(net6152),
    .A2(\mem.mem[223][4] ),
    .Y(_05068_),
    .B1(net5367));
 sg13g2_o21ai_1 _14083_ (.B1(_05068_),
    .Y(_05069_),
    .A1(net6152),
    .A2(_02864_));
 sg13g2_nand2_1 _14084_ (.Y(_05070_),
    .A(net6153),
    .B(\mem.mem[221][4] ));
 sg13g2_a21oi_1 _14085_ (.A1(net5415),
    .A2(\mem.mem[220][4] ),
    .Y(_05071_),
    .B1(net5989));
 sg13g2_a21oi_1 _14086_ (.A1(_05070_),
    .A2(_05071_),
    .Y(_05072_),
    .B1(net5340));
 sg13g2_a221oi_1 _14087_ (.B2(_05072_),
    .C1(net5295),
    .B1(_05069_),
    .A1(net5340),
    .Y(_05073_),
    .A2(_05067_));
 sg13g2_o21ai_1 _14088_ (.B1(net5824),
    .Y(_05074_),
    .A1(_05066_),
    .A2(_05073_));
 sg13g2_nand2_2 _14089_ (.Y(_05075_),
    .A(net5266),
    .B(_05074_));
 sg13g2_o21ai_1 _14090_ (.B1(_05036_),
    .Y(_05076_),
    .A1(_05055_),
    .A2(_05075_));
 sg13g2_nand2_1 _14091_ (.Y(_05077_),
    .A(_00006_),
    .B(_05076_));
 sg13g2_mux4_1 _14092_ (.S0(net6056),
    .A0(\mem.mem[160][4] ),
    .A1(\mem.mem[161][4] ),
    .A2(\mem.mem[162][4] ),
    .A3(\mem.mem[163][4] ),
    .S1(net5920),
    .X(_05078_));
 sg13g2_nand2_1 _14093_ (.Y(_05079_),
    .A(net5387),
    .B(\mem.mem[166][4] ));
 sg13g2_a21oi_1 _14094_ (.A1(net6058),
    .A2(\mem.mem[167][4] ),
    .Y(_05080_),
    .B1(net5353));
 sg13g2_nand2b_1 _14095_ (.Y(_05081_),
    .B(net6058),
    .A_N(\mem.mem[165][4] ));
 sg13g2_o21ai_1 _14096_ (.B1(_05081_),
    .Y(_05082_),
    .A1(net6058),
    .A2(\mem.mem[164][4] ));
 sg13g2_a221oi_1 _14097_ (.B2(net5353),
    .C1(net5314),
    .B1(_05082_),
    .A1(_05079_),
    .Y(_05083_),
    .A2(_05080_));
 sg13g2_a21oi_2 _14098_ (.B1(_05083_),
    .Y(_05084_),
    .A2(_05078_),
    .A1(net5314));
 sg13g2_mux4_1 _14099_ (.S0(net6091),
    .A0(\mem.mem[172][4] ),
    .A1(\mem.mem[173][4] ),
    .A2(\mem.mem[174][4] ),
    .A3(\mem.mem[175][4] ),
    .S1(net5949),
    .X(_05085_));
 sg13g2_nor2b_1 _14100_ (.A(net6085),
    .B_N(\mem.mem[170][4] ),
    .Y(_05086_));
 sg13g2_a21oi_2 _14101_ (.B1(_05086_),
    .Y(_05087_),
    .A2(\mem.mem[171][4] ),
    .A1(net6090));
 sg13g2_nand2_1 _14102_ (.Y(_05088_),
    .A(net6090),
    .B(\mem.mem[169][4] ));
 sg13g2_nand2_1 _14103_ (.Y(_05089_),
    .A(net5397),
    .B(\mem.mem[168][4] ));
 sg13g2_nand3_1 _14104_ (.B(_05088_),
    .C(_05089_),
    .A(net5357),
    .Y(_05090_));
 sg13g2_a21oi_1 _14105_ (.A1(net5946),
    .A2(_05087_),
    .Y(_05091_),
    .B1(net5866));
 sg13g2_a221oi_1 _14106_ (.B2(_05091_),
    .C1(net5287),
    .B1(_05090_),
    .A1(net5866),
    .Y(_05092_),
    .A2(_05085_));
 sg13g2_a21oi_1 _14107_ (.A1(net5287),
    .A2(_05084_),
    .Y(_05093_),
    .B1(_05092_));
 sg13g2_mux4_1 _14108_ (.S0(net6137),
    .A0(\mem.mem[188][4] ),
    .A1(\mem.mem[189][4] ),
    .A2(\mem.mem[190][4] ),
    .A3(\mem.mem[191][4] ),
    .S1(net5977),
    .X(_05094_));
 sg13g2_nor2b_1 _14109_ (.A(net6131),
    .B_N(\mem.mem[186][4] ),
    .Y(_05095_));
 sg13g2_a21oi_1 _14110_ (.A1(net6131),
    .A2(\mem.mem[187][4] ),
    .Y(_05096_),
    .B1(_05095_));
 sg13g2_mux2_1 _14111_ (.A0(\mem.mem[184][4] ),
    .A1(\mem.mem[185][4] ),
    .S(net6130),
    .X(_05097_));
 sg13g2_a21oi_1 _14112_ (.A1(net5972),
    .A2(_05096_),
    .Y(_05098_),
    .B1(net5875));
 sg13g2_o21ai_1 _14113_ (.B1(_05098_),
    .Y(_05099_),
    .A1(net5972),
    .A2(_05097_));
 sg13g2_a21oi_1 _14114_ (.A1(net5876),
    .A2(_05094_),
    .Y(_05100_),
    .B1(net5292));
 sg13g2_mux2_1 _14115_ (.A0(\mem.mem[180][4] ),
    .A1(\mem.mem[181][4] ),
    .S(net6137),
    .X(_05101_));
 sg13g2_and2_1 _14116_ (.A(net6134),
    .B(\mem.mem[183][4] ),
    .X(_05102_));
 sg13g2_a21oi_1 _14117_ (.A1(net5409),
    .A2(\mem.mem[182][4] ),
    .Y(_05103_),
    .B1(_05102_));
 sg13g2_a21oi_1 _14118_ (.A1(net5975),
    .A2(_05103_),
    .Y(_05104_),
    .B1(net5336));
 sg13g2_o21ai_1 _14119_ (.B1(_05104_),
    .Y(_05105_),
    .A1(net5977),
    .A2(_05101_));
 sg13g2_mux4_1 _14120_ (.S0(net6130),
    .A0(\mem.mem[176][4] ),
    .A1(\mem.mem[177][4] ),
    .A2(\mem.mem[178][4] ),
    .A3(\mem.mem[179][4] ),
    .S1(net5972),
    .X(_05106_));
 sg13g2_a21oi_2 _14121_ (.B1(net5845),
    .Y(_05107_),
    .A2(_05106_),
    .A1(net5334));
 sg13g2_a22oi_1 _14122_ (.Y(_05108_),
    .B1(_05105_),
    .B2(_05107_),
    .A2(_05100_),
    .A1(_05099_));
 sg13g2_nand2b_1 _14123_ (.Y(_05109_),
    .B(net6102),
    .A_N(\mem.mem[133][4] ));
 sg13g2_o21ai_1 _14124_ (.B1(_05109_),
    .Y(_05110_),
    .A1(net6119),
    .A2(\mem.mem[132][4] ));
 sg13g2_nand2_1 _14125_ (.Y(_05111_),
    .A(net5399),
    .B(\mem.mem[134][4] ));
 sg13g2_a21oi_1 _14126_ (.A1(net6102),
    .A2(\mem.mem[135][4] ),
    .Y(_05112_),
    .B1(net5360));
 sg13g2_a221oi_1 _14127_ (.B2(_05112_),
    .C1(net5325),
    .B1(_05111_),
    .A1(net5358),
    .Y(_05113_),
    .A2(_05110_));
 sg13g2_mux4_1 _14128_ (.S0(net6100),
    .A0(\mem.mem[128][4] ),
    .A1(\mem.mem[129][4] ),
    .A2(\mem.mem[130][4] ),
    .A3(\mem.mem[131][4] ),
    .S1(net5953),
    .X(_05114_));
 sg13g2_a21oi_2 _14129_ (.B1(_05113_),
    .Y(_05115_),
    .A2(_05114_),
    .A1(net5325));
 sg13g2_mux4_1 _14130_ (.S0(net6111),
    .A0(\mem.mem[140][4] ),
    .A1(\mem.mem[141][4] ),
    .A2(\mem.mem[142][4] ),
    .A3(\mem.mem[143][4] ),
    .S1(net5958),
    .X(_05116_));
 sg13g2_nor2b_1 _14131_ (.A(net6113),
    .B_N(\mem.mem[138][4] ),
    .Y(_05117_));
 sg13g2_a21oi_1 _14132_ (.A1(net6113),
    .A2(\mem.mem[139][4] ),
    .Y(_05118_),
    .B1(_05117_));
 sg13g2_nand2_1 _14133_ (.Y(_05119_),
    .A(net6113),
    .B(\mem.mem[137][4] ));
 sg13g2_nand2_1 _14134_ (.Y(_05120_),
    .A(net5403),
    .B(\mem.mem[136][4] ));
 sg13g2_nand3_1 _14135_ (.B(_05119_),
    .C(_05120_),
    .A(net5364),
    .Y(_05121_));
 sg13g2_a21oi_1 _14136_ (.A1(net5959),
    .A2(_05118_),
    .Y(_05122_),
    .B1(net5870));
 sg13g2_a221oi_1 _14137_ (.B2(_05122_),
    .C1(net5290),
    .B1(_05121_),
    .A1(net5870),
    .Y(_05123_),
    .A2(_05116_));
 sg13g2_a21oi_1 _14138_ (.A1(net5287),
    .A2(_05115_),
    .Y(_05124_),
    .B1(_05123_));
 sg13g2_mux4_1 _14139_ (.S0(net6091),
    .A0(\mem.mem[156][4] ),
    .A1(\mem.mem[157][4] ),
    .A2(\mem.mem[158][4] ),
    .A3(\mem.mem[159][4] ),
    .S1(net5949),
    .X(_05125_));
 sg13g2_mux4_1 _14140_ (.S0(net6093),
    .A0(\mem.mem[152][4] ),
    .A1(\mem.mem[153][4] ),
    .A2(\mem.mem[154][4] ),
    .A3(\mem.mem[155][4] ),
    .S1(net5947),
    .X(_05126_));
 sg13g2_nand2_1 _14141_ (.Y(_05127_),
    .A(net5327),
    .B(_05126_));
 sg13g2_a21oi_1 _14142_ (.A1(net5866),
    .A2(_05125_),
    .Y(_05128_),
    .B1(net5287));
 sg13g2_mux2_1 _14143_ (.A0(\mem.mem[148][4] ),
    .A1(\mem.mem[149][4] ),
    .S(net6108),
    .X(_05129_));
 sg13g2_and2_1 _14144_ (.A(net6108),
    .B(\mem.mem[151][4] ),
    .X(_05130_));
 sg13g2_a21oi_1 _14145_ (.A1(net5404),
    .A2(\mem.mem[150][4] ),
    .Y(_05131_),
    .B1(_05130_));
 sg13g2_a21oi_1 _14146_ (.A1(net5957),
    .A2(_05131_),
    .Y(_05132_),
    .B1(net5329));
 sg13g2_o21ai_1 _14147_ (.B1(_05132_),
    .Y(_05133_),
    .A1(net5962),
    .A2(_05129_));
 sg13g2_mux4_1 _14148_ (.S0(net6061),
    .A0(\mem.mem[144][4] ),
    .A1(\mem.mem[145][4] ),
    .A2(\mem.mem[146][4] ),
    .A3(\mem.mem[147][4] ),
    .S1(net5922),
    .X(_05134_));
 sg13g2_a21oi_1 _14149_ (.A1(net5323),
    .A2(_05134_),
    .Y(_05135_),
    .B1(net5838));
 sg13g2_a22oi_1 _14150_ (.Y(_05136_),
    .B1(_05133_),
    .B2(_05135_),
    .A2(_05128_),
    .A1(_05127_));
 sg13g2_mux4_1 _14151_ (.S0(net5821),
    .A0(_05093_),
    .A1(_05108_),
    .A2(_05124_),
    .A3(_05136_),
    .S1(net5266),
    .X(_05137_));
 sg13g2_a21oi_1 _14152_ (.A1(net5263),
    .A2(_05137_),
    .Y(_05138_),
    .B1(_02840_));
 sg13g2_nand2_2 _14153_ (.Y(_05139_),
    .A(_05077_),
    .B(_05138_));
 sg13g2_nor2_1 _14154_ (.A(_02944_),
    .B(_05015_),
    .Y(_05140_));
 sg13g2_a22oi_1 _14155_ (.Y(_05141_),
    .B1(_05139_),
    .B2(_05140_),
    .A2(_03639_),
    .A1(net6));
 sg13g2_o21ai_1 _14156_ (.B1(net6187),
    .Y(_05142_),
    .A1(net5788),
    .A2(net4187));
 sg13g2_a21oi_1 _14157_ (.A1(net5788),
    .A2(_05141_),
    .Y(_00552_),
    .B1(_05142_));
 sg13g2_nand2_1 _14158_ (.Y(_05143_),
    .A(net5371),
    .B(\mem.mem[68][5] ));
 sg13g2_a21oi_1 _14159_ (.A1(net6017),
    .A2(\mem.mem[69][5] ),
    .Y(_05144_),
    .B1(net5886));
 sg13g2_and2_1 _14160_ (.A(net6007),
    .B(\mem.mem[71][5] ),
    .X(_05145_));
 sg13g2_a21oi_1 _14161_ (.A1(net5371),
    .A2(\mem.mem[70][5] ),
    .Y(_05146_),
    .B1(_05145_));
 sg13g2_a221oi_1 _14162_ (.B2(net5887),
    .C1(net5301),
    .B1(_05146_),
    .A1(_05143_),
    .Y(_05147_),
    .A2(_05144_));
 sg13g2_mux4_1 _14163_ (.S0(net6007),
    .A0(\mem.mem[64][5] ),
    .A1(\mem.mem[65][5] ),
    .A2(\mem.mem[66][5] ),
    .A3(\mem.mem[67][5] ),
    .S1(net5886),
    .X(_05148_));
 sg13g2_nand2_1 _14164_ (.Y(_05149_),
    .A(net5298),
    .B(_05148_));
 sg13g2_nor2_1 _14165_ (.A(net5827),
    .B(_05147_),
    .Y(_05150_));
 sg13g2_nand2_1 _14166_ (.Y(_05151_),
    .A(net5374),
    .B(\mem.mem[72][5] ));
 sg13g2_a21oi_1 _14167_ (.A1(net6022),
    .A2(\mem.mem[73][5] ),
    .Y(_05152_),
    .B1(net5897));
 sg13g2_nor2b_1 _14168_ (.A(net6022),
    .B_N(\mem.mem[74][5] ),
    .Y(_05153_));
 sg13g2_a21oi_1 _14169_ (.A1(net6022),
    .A2(\mem.mem[75][5] ),
    .Y(_05154_),
    .B1(_05153_));
 sg13g2_a221oi_1 _14170_ (.B2(net5897),
    .C1(net5853),
    .B1(_05154_),
    .A1(_05151_),
    .Y(_05155_),
    .A2(_05152_));
 sg13g2_mux2_1 _14171_ (.A0(\mem.mem[78][5] ),
    .A1(\mem.mem[79][5] ),
    .S(net6012),
    .X(_05156_));
 sg13g2_nand2_1 _14172_ (.Y(_05157_),
    .A(net6012),
    .B(\mem.mem[77][5] ));
 sg13g2_a21oi_1 _14173_ (.A1(net5370),
    .A2(\mem.mem[76][5] ),
    .Y(_05158_),
    .B1(net5890));
 sg13g2_a21oi_1 _14174_ (.A1(_05157_),
    .A2(_05158_),
    .Y(_05159_),
    .B1(net5300));
 sg13g2_o21ai_1 _14175_ (.B1(_05159_),
    .Y(_05160_),
    .A1(net5349),
    .A2(_05156_));
 sg13g2_nor2_1 _14176_ (.A(net5278),
    .B(_05155_),
    .Y(_05161_));
 sg13g2_a22oi_1 _14177_ (.Y(_05162_),
    .B1(_05160_),
    .B2(_05161_),
    .A2(_05150_),
    .A1(_05149_));
 sg13g2_nor2b_1 _14178_ (.A(net6008),
    .B_N(\mem.mem[86][5] ),
    .Y(_05163_));
 sg13g2_a21oi_1 _14179_ (.A1(net6008),
    .A2(\mem.mem[87][5] ),
    .Y(_05164_),
    .B1(_05163_));
 sg13g2_nand2_1 _14180_ (.Y(_05165_),
    .A(net5370),
    .B(\mem.mem[84][5] ));
 sg13g2_a21oi_1 _14181_ (.A1(net6008),
    .A2(\mem.mem[85][5] ),
    .Y(_05166_),
    .B1(net5888));
 sg13g2_a221oi_1 _14182_ (.B2(_05166_),
    .C1(net5299),
    .B1(_05165_),
    .A1(net5888),
    .Y(_05167_),
    .A2(_05164_));
 sg13g2_mux4_1 _14183_ (.S0(net6005),
    .A0(\mem.mem[80][5] ),
    .A1(\mem.mem[81][5] ),
    .A2(\mem.mem[82][5] ),
    .A3(\mem.mem[83][5] ),
    .S1(net5887),
    .X(_05168_));
 sg13g2_a21oi_2 _14184_ (.B1(_05167_),
    .Y(_05169_),
    .A2(_05168_),
    .A1(net5299));
 sg13g2_nand2_1 _14185_ (.Y(_05170_),
    .A(net5386),
    .B(\mem.mem[88][5] ));
 sg13g2_a21oi_1 _14186_ (.A1(net6046),
    .A2(\mem.mem[89][5] ),
    .Y(_05171_),
    .B1(net5916));
 sg13g2_nor2b_1 _14187_ (.A(net6046),
    .B_N(\mem.mem[90][5] ),
    .Y(_05172_));
 sg13g2_a21oi_1 _14188_ (.A1(net6046),
    .A2(\mem.mem[91][5] ),
    .Y(_05173_),
    .B1(_05172_));
 sg13g2_a221oi_1 _14189_ (.B2(net5916),
    .C1(net5857),
    .B1(_05173_),
    .A1(_05170_),
    .Y(_05174_),
    .A2(_05171_));
 sg13g2_nand2_1 _14190_ (.Y(_05175_),
    .A(net6051),
    .B(\mem.mem[93][5] ));
 sg13g2_a21oi_1 _14191_ (.A1(net5385),
    .A2(\mem.mem[92][5] ),
    .Y(_05176_),
    .B1(net5917));
 sg13g2_and2_1 _14192_ (.A(net6051),
    .B(\mem.mem[95][5] ),
    .X(_05177_));
 sg13g2_a21oi_1 _14193_ (.A1(net5385),
    .A2(\mem.mem[94][5] ),
    .Y(_05178_),
    .B1(_05177_));
 sg13g2_a221oi_1 _14194_ (.B2(net5917),
    .C1(net5311),
    .B1(_05178_),
    .A1(_05175_),
    .Y(_05179_),
    .A2(_05176_));
 sg13g2_nor3_1 _14195_ (.A(net5282),
    .B(_05174_),
    .C(_05179_),
    .Y(_05180_));
 sg13g2_a21oi_1 _14196_ (.A1(net5277),
    .A2(_05169_),
    .Y(_05181_),
    .B1(_05180_));
 sg13g2_nor2b_1 _14197_ (.A(net6071),
    .B_N(\mem.mem[102][5] ),
    .Y(_05182_));
 sg13g2_a21oi_1 _14198_ (.A1(net6071),
    .A2(\mem.mem[103][5] ),
    .Y(_05183_),
    .B1(_05182_));
 sg13g2_nand2_1 _14199_ (.Y(_05184_),
    .A(net5389),
    .B(\mem.mem[100][5] ));
 sg13g2_a21oi_1 _14200_ (.A1(net6068),
    .A2(\mem.mem[101][5] ),
    .Y(_05185_),
    .B1(net5928));
 sg13g2_a221oi_1 _14201_ (.B2(_05185_),
    .C1(net5316),
    .B1(_05184_),
    .A1(net5928),
    .Y(_05186_),
    .A2(_05183_));
 sg13g2_mux4_1 _14202_ (.S0(net6069),
    .A0(\mem.mem[96][5] ),
    .A1(\mem.mem[97][5] ),
    .A2(\mem.mem[98][5] ),
    .A3(\mem.mem[99][5] ),
    .S1(net5928),
    .X(_05187_));
 sg13g2_a21oi_2 _14203_ (.B1(_05186_),
    .Y(_05188_),
    .A2(_05187_),
    .A1(net5316));
 sg13g2_mux4_1 _14204_ (.S0(net6054),
    .A0(\mem.mem[104][5] ),
    .A1(\mem.mem[105][5] ),
    .A2(\mem.mem[106][5] ),
    .A3(\mem.mem[107][5] ),
    .S1(net5917),
    .X(_05189_));
 sg13g2_nand2_1 _14205_ (.Y(_05190_),
    .A(net6052),
    .B(\mem.mem[109][5] ));
 sg13g2_a21oi_1 _14206_ (.A1(net5386),
    .A2(\mem.mem[108][5] ),
    .Y(_05191_),
    .B1(net5919));
 sg13g2_a21oi_1 _14207_ (.A1(net6052),
    .A2(\mem.mem[111][5] ),
    .Y(_05192_),
    .B1(net5354));
 sg13g2_o21ai_1 _14208_ (.B1(_05192_),
    .Y(_05193_),
    .A1(net6052),
    .A2(_02867_));
 sg13g2_a21oi_1 _14209_ (.A1(_05190_),
    .A2(_05191_),
    .Y(_05194_),
    .B1(net5311));
 sg13g2_a221oi_1 _14210_ (.B2(_05194_),
    .C1(net5281),
    .B1(_05193_),
    .A1(net5311),
    .Y(_05195_),
    .A2(_05189_));
 sg13g2_a21oi_1 _14211_ (.A1(net5282),
    .A2(_05188_),
    .Y(_05196_),
    .B1(_05195_));
 sg13g2_nand2_1 _14212_ (.Y(_05197_),
    .A(net5374),
    .B(\mem.mem[116][5] ));
 sg13g2_a21oi_1 _14213_ (.A1(net6023),
    .A2(\mem.mem[117][5] ),
    .Y(_05198_),
    .B1(net5899));
 sg13g2_and2_1 _14214_ (.A(net6024),
    .B(\mem.mem[119][5] ),
    .X(_05199_));
 sg13g2_a21oi_1 _14215_ (.A1(net5375),
    .A2(\mem.mem[118][5] ),
    .Y(_05200_),
    .B1(_05199_));
 sg13g2_a221oi_1 _14216_ (.B2(net5898),
    .C1(net5303),
    .B1(_05200_),
    .A1(_05197_),
    .Y(_05201_),
    .A2(_05198_));
 sg13g2_nand2_1 _14217_ (.Y(_05202_),
    .A(net5385),
    .B(\mem.mem[112][5] ));
 sg13g2_a21oi_1 _14218_ (.A1(net6050),
    .A2(\mem.mem[113][5] ),
    .Y(_05203_),
    .B1(net5917));
 sg13g2_nor2b_1 _14219_ (.A(net6050),
    .B_N(\mem.mem[114][5] ),
    .Y(_05204_));
 sg13g2_a21oi_1 _14220_ (.A1(net6050),
    .A2(\mem.mem[115][5] ),
    .Y(_05205_),
    .B1(_05204_));
 sg13g2_a221oi_1 _14221_ (.B2(net5917),
    .C1(net5857),
    .B1(_05205_),
    .A1(_05202_),
    .Y(_05206_),
    .A2(_05203_));
 sg13g2_nor3_1 _14222_ (.A(net5831),
    .B(_05201_),
    .C(_05206_),
    .Y(_05207_));
 sg13g2_nand2_1 _14223_ (.Y(_05208_),
    .A(net5389),
    .B(\mem.mem[120][5] ));
 sg13g2_a21oi_1 _14224_ (.A1(net6069),
    .A2(\mem.mem[121][5] ),
    .Y(_05209_),
    .B1(net5928));
 sg13g2_nor2b_1 _14225_ (.A(net6069),
    .B_N(\mem.mem[122][5] ),
    .Y(_05210_));
 sg13g2_a21oi_1 _14226_ (.A1(net6069),
    .A2(\mem.mem[123][5] ),
    .Y(_05211_),
    .B1(_05210_));
 sg13g2_a221oi_1 _14227_ (.B2(net5928),
    .C1(net5855),
    .B1(_05211_),
    .A1(_05208_),
    .Y(_05212_),
    .A2(_05209_));
 sg13g2_nor2b_1 _14228_ (.A(net6040),
    .B_N(\mem.mem[126][5] ),
    .Y(_05213_));
 sg13g2_a21oi_1 _14229_ (.A1(net6040),
    .A2(\mem.mem[127][5] ),
    .Y(_05214_),
    .B1(_05213_));
 sg13g2_nand2_1 _14230_ (.Y(_05215_),
    .A(net5381),
    .B(\mem.mem[124][5] ));
 sg13g2_a21oi_1 _14231_ (.A1(net6040),
    .A2(\mem.mem[125][5] ),
    .Y(_05216_),
    .B1(net5910));
 sg13g2_a221oi_1 _14232_ (.B2(_05216_),
    .C1(net5307),
    .B1(_05215_),
    .A1(net5910),
    .Y(_05217_),
    .A2(_05214_));
 sg13g2_nor3_2 _14233_ (.A(net5280),
    .B(_05212_),
    .C(_05217_),
    .Y(_05218_));
 sg13g2_nor2_1 _14234_ (.A(_05207_),
    .B(_05218_),
    .Y(_05219_));
 sg13g2_mux4_1 _14235_ (.S0(net5816),
    .A0(_05162_),
    .A1(_05181_),
    .A2(_05196_),
    .A3(_05219_),
    .S1(net5810),
    .X(_05220_));
 sg13g2_nand2_1 _14236_ (.Y(_05221_),
    .A(net5418),
    .B(\mem.mem[36][5] ));
 sg13g2_a21oi_1 _14237_ (.A1(net6160),
    .A2(\mem.mem[37][5] ),
    .Y(_05222_),
    .B1(net5992));
 sg13g2_and2_1 _14238_ (.A(net6159),
    .B(\mem.mem[39][5] ),
    .X(_05223_));
 sg13g2_a21oi_1 _14239_ (.A1(net5417),
    .A2(\mem.mem[38][5] ),
    .Y(_05224_),
    .B1(_05223_));
 sg13g2_a221oi_1 _14240_ (.B2(net5992),
    .C1(net5342),
    .B1(_05224_),
    .A1(_05221_),
    .Y(_05225_),
    .A2(_05222_));
 sg13g2_nand2_1 _14241_ (.Y(_05226_),
    .A(net5417),
    .B(\mem.mem[32][5] ));
 sg13g2_a21oi_1 _14242_ (.A1(net6159),
    .A2(\mem.mem[33][5] ),
    .Y(_05227_),
    .B1(net5993));
 sg13g2_nor2b_1 _14243_ (.A(net6159),
    .B_N(\mem.mem[34][5] ),
    .Y(_05228_));
 sg13g2_a21oi_1 _14244_ (.A1(net6159),
    .A2(\mem.mem[35][5] ),
    .Y(_05229_),
    .B1(_05228_));
 sg13g2_a221oi_1 _14245_ (.B2(net5993),
    .C1(net5880),
    .B1(_05229_),
    .A1(_05226_),
    .Y(_05230_),
    .A2(_05227_));
 sg13g2_nor3_1 _14246_ (.A(net5846),
    .B(_05225_),
    .C(_05230_),
    .Y(_05231_));
 sg13g2_nand2_1 _14247_ (.Y(_05232_),
    .A(net5420),
    .B(\mem.mem[40][5] ));
 sg13g2_a21oi_1 _14248_ (.A1(net6168),
    .A2(\mem.mem[41][5] ),
    .Y(_05233_),
    .B1(net6000));
 sg13g2_nor2b_1 _14249_ (.A(net6167),
    .B_N(\mem.mem[42][5] ),
    .Y(_05234_));
 sg13g2_a21oi_1 _14250_ (.A1(net6167),
    .A2(\mem.mem[43][5] ),
    .Y(_05235_),
    .B1(_05234_));
 sg13g2_a221oi_1 _14251_ (.B2(net6000),
    .C1(net5881),
    .B1(_05235_),
    .A1(_05232_),
    .Y(_05236_),
    .A2(_05233_));
 sg13g2_nor2b_1 _14252_ (.A(net6162),
    .B_N(\mem.mem[46][5] ),
    .Y(_05237_));
 sg13g2_a21oi_1 _14253_ (.A1(net6162),
    .A2(\mem.mem[47][5] ),
    .Y(_05238_),
    .B1(_05237_));
 sg13g2_nand2_1 _14254_ (.Y(_05239_),
    .A(net5420),
    .B(\mem.mem[44][5] ));
 sg13g2_a21oi_1 _14255_ (.A1(net6169),
    .A2(\mem.mem[45][5] ),
    .Y(_05240_),
    .B1(net6000));
 sg13g2_a221oi_1 _14256_ (.B2(_05240_),
    .C1(net5345),
    .B1(_05239_),
    .A1(net5999),
    .Y(_05241_),
    .A2(_05238_));
 sg13g2_nor3_2 _14257_ (.A(net5295),
    .B(_05236_),
    .C(_05241_),
    .Y(_05242_));
 sg13g2_nor2_2 _14258_ (.A(_05231_),
    .B(_05242_),
    .Y(_05243_));
 sg13g2_nand2_1 _14259_ (.Y(_05244_),
    .A(net5377),
    .B(\mem.mem[52][5] ));
 sg13g2_a21oi_1 _14260_ (.A1(net6030),
    .A2(\mem.mem[53][5] ),
    .Y(_05245_),
    .B1(net5903));
 sg13g2_and2_1 _14261_ (.A(net6030),
    .B(\mem.mem[55][5] ),
    .X(_05246_));
 sg13g2_a21oi_1 _14262_ (.A1(net5377),
    .A2(\mem.mem[54][5] ),
    .Y(_05247_),
    .B1(_05246_));
 sg13g2_a221oi_1 _14263_ (.B2(net5903),
    .C1(net5304),
    .B1(_05247_),
    .A1(_05244_),
    .Y(_05248_),
    .A2(_05245_));
 sg13g2_mux4_1 _14264_ (.S0(net6010),
    .A0(\mem.mem[48][5] ),
    .A1(\mem.mem[49][5] ),
    .A2(\mem.mem[50][5] ),
    .A3(\mem.mem[51][5] ),
    .S1(net5889),
    .X(_05249_));
 sg13g2_nand2_1 _14265_ (.Y(_05250_),
    .A(net5304),
    .B(_05249_));
 sg13g2_nor2_1 _14266_ (.A(net5829),
    .B(_05248_),
    .Y(_05251_));
 sg13g2_nand2_1 _14267_ (.Y(_05252_),
    .A(net5377),
    .B(\mem.mem[56][5] ));
 sg13g2_a21oi_1 _14268_ (.A1(net6029),
    .A2(\mem.mem[57][5] ),
    .Y(_05253_),
    .B1(net5903));
 sg13g2_nor2b_1 _14269_ (.A(net6029),
    .B_N(\mem.mem[58][5] ),
    .Y(_05254_));
 sg13g2_a21oi_1 _14270_ (.A1(net6034),
    .A2(\mem.mem[59][5] ),
    .Y(_05255_),
    .B1(_05254_));
 sg13g2_a221oi_1 _14271_ (.B2(net5904),
    .C1(net5854),
    .B1(_05255_),
    .A1(_05252_),
    .Y(_05256_),
    .A2(_05253_));
 sg13g2_nor2b_1 _14272_ (.A(net6038),
    .B_N(\mem.mem[62][5] ),
    .Y(_05257_));
 sg13g2_a21oi_1 _14273_ (.A1(net6038),
    .A2(\mem.mem[63][5] ),
    .Y(_05258_),
    .B1(_05257_));
 sg13g2_nand2_1 _14274_ (.Y(_05259_),
    .A(net5378),
    .B(\mem.mem[60][5] ));
 sg13g2_a21oi_1 _14275_ (.A1(net6038),
    .A2(\mem.mem[61][5] ),
    .Y(_05260_),
    .B1(net5912));
 sg13g2_a221oi_1 _14276_ (.B2(_05260_),
    .C1(net5304),
    .B1(_05259_),
    .A1(net5905),
    .Y(_05261_),
    .A2(_05258_));
 sg13g2_nor3_2 _14277_ (.A(net5279),
    .B(_05256_),
    .C(_05261_),
    .Y(_05262_));
 sg13g2_a21oi_2 _14278_ (.B1(_05262_),
    .Y(_05263_),
    .A2(_05251_),
    .A1(_05250_));
 sg13g2_nand2_1 _14279_ (.Y(_05264_),
    .A(net5392),
    .B(\mem.mem[4][5] ));
 sg13g2_a21oi_1 _14280_ (.A1(net6077),
    .A2(\mem.mem[5][5] ),
    .Y(_05265_),
    .B1(net5935));
 sg13g2_and2_1 _14281_ (.A(net6077),
    .B(\mem.mem[7][5] ),
    .X(_05266_));
 sg13g2_a21oi_1 _14282_ (.A1(net5392),
    .A2(\mem.mem[6][5] ),
    .Y(_05267_),
    .B1(_05266_));
 sg13g2_a221oi_1 _14283_ (.B2(net5935),
    .C1(net5320),
    .B1(_05267_),
    .A1(_05264_),
    .Y(_05268_),
    .A2(_05265_));
 sg13g2_mux4_1 _14284_ (.S0(net6079),
    .A0(\mem.mem[0][5] ),
    .A1(\mem.mem[1][5] ),
    .A2(\mem.mem[2][5] ),
    .A3(\mem.mem[3][5] ),
    .S1(net5940),
    .X(_05269_));
 sg13g2_nand2_1 _14285_ (.Y(_05270_),
    .A(net5319),
    .B(_05269_));
 sg13g2_nor2_1 _14286_ (.A(net5835),
    .B(_05268_),
    .Y(_05271_));
 sg13g2_mux4_1 _14287_ (.S0(net6083),
    .A0(\mem.mem[8][5] ),
    .A1(\mem.mem[9][5] ),
    .A2(\mem.mem[10][5] ),
    .A3(\mem.mem[11][5] ),
    .S1(net5938),
    .X(_05272_));
 sg13g2_a21oi_1 _14288_ (.A1(net6109),
    .A2(\mem.mem[15][5] ),
    .Y(_05273_),
    .B1(net5356));
 sg13g2_o21ai_1 _14289_ (.B1(_05273_),
    .Y(_05274_),
    .A1(net6109),
    .A2(_02866_));
 sg13g2_nand2_1 _14290_ (.Y(_05275_),
    .A(net6081),
    .B(\mem.mem[13][5] ));
 sg13g2_a21oi_1 _14291_ (.A1(net5394),
    .A2(\mem.mem[12][5] ),
    .Y(_05276_),
    .B1(net5938));
 sg13g2_a21oi_1 _14292_ (.A1(_05275_),
    .A2(_05276_),
    .Y(_05277_),
    .B1(net5318));
 sg13g2_a221oi_1 _14293_ (.B2(_05277_),
    .C1(net5283),
    .B1(_05274_),
    .A1(net5319),
    .Y(_05278_),
    .A2(_05272_));
 sg13g2_a21oi_1 _14294_ (.A1(_05270_),
    .A2(_05271_),
    .Y(_05279_),
    .B1(_05278_));
 sg13g2_nor2b_1 _14295_ (.A(net6126),
    .B_N(\mem.mem[22][5] ),
    .Y(_05280_));
 sg13g2_a21oi_1 _14296_ (.A1(net6126),
    .A2(\mem.mem[23][5] ),
    .Y(_05281_),
    .B1(_05280_));
 sg13g2_nand2_1 _14297_ (.Y(_05282_),
    .A(net5417),
    .B(\mem.mem[20][5] ));
 sg13g2_a21oi_1 _14298_ (.A1(net6156),
    .A2(\mem.mem[21][5] ),
    .Y(_05283_),
    .B1(net5969));
 sg13g2_a221oi_1 _14299_ (.B2(_05283_),
    .C1(net5341),
    .B1(_05282_),
    .A1(net5991),
    .Y(_05284_),
    .A2(_05281_));
 sg13g2_nand2_1 _14300_ (.Y(_05285_),
    .A(net5417),
    .B(\mem.mem[16][5] ));
 sg13g2_a21oi_1 _14301_ (.A1(net6156),
    .A2(\mem.mem[17][5] ),
    .Y(_05286_),
    .B1(net5991));
 sg13g2_nor2b_1 _14302_ (.A(net6156),
    .B_N(\mem.mem[18][5] ),
    .Y(_05287_));
 sg13g2_a21oi_1 _14303_ (.A1(net6156),
    .A2(\mem.mem[19][5] ),
    .Y(_05288_),
    .B1(_05287_));
 sg13g2_a221oi_1 _14304_ (.B2(net5991),
    .C1(net5883),
    .B1(_05288_),
    .A1(_05285_),
    .Y(_05289_),
    .A2(_05286_));
 sg13g2_nor3_2 _14305_ (.A(net5848),
    .B(_05284_),
    .C(_05289_),
    .Y(_05290_));
 sg13g2_nand2_1 _14306_ (.Y(_05291_),
    .A(net5405),
    .B(\mem.mem[24][5] ));
 sg13g2_a21oi_1 _14307_ (.A1(net6149),
    .A2(\mem.mem[25][5] ),
    .Y(_05292_),
    .B1(net5964));
 sg13g2_nor2b_1 _14308_ (.A(net6149),
    .B_N(\mem.mem[26][5] ),
    .Y(_05293_));
 sg13g2_a21oi_1 _14309_ (.A1(net6149),
    .A2(\mem.mem[27][5] ),
    .Y(_05294_),
    .B1(_05293_));
 sg13g2_a221oi_1 _14310_ (.B2(net5965),
    .C1(net5880),
    .B1(_05294_),
    .A1(_05291_),
    .Y(_05295_),
    .A2(_05292_));
 sg13g2_nand2_1 _14311_ (.Y(_05296_),
    .A(net6150),
    .B(\mem.mem[29][5] ));
 sg13g2_a21oi_1 _14312_ (.A1(net5415),
    .A2(\mem.mem[28][5] ),
    .Y(_05297_),
    .B1(net5987));
 sg13g2_and2_1 _14313_ (.A(net6152),
    .B(\mem.mem[31][5] ),
    .X(_05298_));
 sg13g2_a21oi_1 _14314_ (.A1(net5418),
    .A2(\mem.mem[30][5] ),
    .Y(_05299_),
    .B1(_05298_));
 sg13g2_a221oi_1 _14315_ (.B2(net5987),
    .C1(net5340),
    .B1(_05299_),
    .A1(_05296_),
    .Y(_05300_),
    .A2(_05297_));
 sg13g2_nor3_1 _14316_ (.A(net5295),
    .B(_05295_),
    .C(_05300_),
    .Y(_05301_));
 sg13g2_nor2_2 _14317_ (.A(_05290_),
    .B(_05301_),
    .Y(_05302_));
 sg13g2_mux4_1 _14318_ (.S0(net5825),
    .A0(_05243_),
    .A1(_05263_),
    .A2(_05279_),
    .A3(_05302_),
    .S1(net5265),
    .X(_05303_));
 sg13g2_mux2_1 _14319_ (.A0(\mem.mem[194][5] ),
    .A1(\mem.mem[195][5] ),
    .S(net6095),
    .X(_05304_));
 sg13g2_mux2_1 _14320_ (.A0(\mem.mem[192][5] ),
    .A1(\mem.mem[193][5] ),
    .S(net6098),
    .X(_05305_));
 sg13g2_nor2_1 _14321_ (.A(net5951),
    .B(_05305_),
    .Y(_05306_));
 sg13g2_o21ai_1 _14322_ (.B1(net5326),
    .Y(_05307_),
    .A1(net5359),
    .A2(_05304_));
 sg13g2_mux4_1 _14323_ (.S0(net6096),
    .A0(\mem.mem[196][5] ),
    .A1(\mem.mem[197][5] ),
    .A2(\mem.mem[198][5] ),
    .A3(\mem.mem[199][5] ),
    .S1(net5950),
    .X(_05308_));
 sg13g2_a21oi_1 _14324_ (.A1(net5868),
    .A2(_05308_),
    .Y(_05309_),
    .B1(net5839));
 sg13g2_o21ai_1 _14325_ (.B1(_05309_),
    .Y(_05310_),
    .A1(_05306_),
    .A2(_05307_));
 sg13g2_mux4_1 _14326_ (.S0(net6086),
    .A0(\mem.mem[200][5] ),
    .A1(\mem.mem[201][5] ),
    .A2(\mem.mem[202][5] ),
    .A3(\mem.mem[203][5] ),
    .S1(net5943),
    .X(_05311_));
 sg13g2_nand2_1 _14327_ (.Y(_05312_),
    .A(net5324),
    .B(_05311_));
 sg13g2_mux4_1 _14328_ (.S0(net6087),
    .A0(\mem.mem[204][5] ),
    .A1(\mem.mem[205][5] ),
    .A2(\mem.mem[206][5] ),
    .A3(\mem.mem[207][5] ),
    .S1(net5944),
    .X(_05313_));
 sg13g2_a21oi_1 _14329_ (.A1(net5865),
    .A2(_05313_),
    .Y(_05314_),
    .B1(net5288));
 sg13g2_and2_1 _14330_ (.A(net6161),
    .B(\mem.mem[223][5] ),
    .X(_05315_));
 sg13g2_a21oi_1 _14331_ (.A1(net5419),
    .A2(\mem.mem[222][5] ),
    .Y(_05316_),
    .B1(_05315_));
 sg13g2_mux2_1 _14332_ (.A0(\mem.mem[220][5] ),
    .A1(\mem.mem[221][5] ),
    .S(net6144),
    .X(_05317_));
 sg13g2_o21ai_1 _14333_ (.B1(net5879),
    .Y(_05318_),
    .A1(net5982),
    .A2(_05317_));
 sg13g2_a21o_1 _14334_ (.A2(_05316_),
    .A1(net5982),
    .B1(_05318_),
    .X(_05319_));
 sg13g2_mux4_1 _14335_ (.S0(net6136),
    .A0(\mem.mem[216][5] ),
    .A1(\mem.mem[217][5] ),
    .A2(\mem.mem[218][5] ),
    .A3(\mem.mem[219][5] ),
    .S1(net5976),
    .X(_05320_));
 sg13g2_a21oi_1 _14336_ (.A1(net5335),
    .A2(_05320_),
    .Y(_05321_),
    .B1(net5292));
 sg13g2_mux2_1 _14337_ (.A0(\mem.mem[210][5] ),
    .A1(\mem.mem[211][5] ),
    .S(net6161),
    .X(_05322_));
 sg13g2_mux2_1 _14338_ (.A0(\mem.mem[208][5] ),
    .A1(\mem.mem[209][5] ),
    .S(net6161),
    .X(_05323_));
 sg13g2_nor2_1 _14339_ (.A(net5995),
    .B(_05323_),
    .Y(_05324_));
 sg13g2_o21ai_1 _14340_ (.B1(net5344),
    .Y(_05325_),
    .A1(net5368),
    .A2(_05322_));
 sg13g2_nand2_1 _14341_ (.Y(_05326_),
    .A(net5413),
    .B(\mem.mem[214][5] ));
 sg13g2_a21oi_1 _14342_ (.A1(net6148),
    .A2(\mem.mem[215][5] ),
    .Y(_05327_),
    .B1(net5365));
 sg13g2_nand2b_1 _14343_ (.Y(_05328_),
    .B(net6144),
    .A_N(\mem.mem[213][5] ));
 sg13g2_o21ai_1 _14344_ (.B1(_05328_),
    .Y(_05329_),
    .A1(net6144),
    .A2(\mem.mem[212][5] ));
 sg13g2_a221oi_1 _14345_ (.B2(net5365),
    .C1(net5338),
    .B1(_05329_),
    .A1(_05326_),
    .Y(_05330_),
    .A2(_05327_));
 sg13g2_o21ai_1 _14346_ (.B1(net5293),
    .Y(_05331_),
    .A1(_05324_),
    .A2(_05325_));
 sg13g2_a21oi_1 _14347_ (.A1(_05312_),
    .A2(_05314_),
    .Y(_05332_),
    .B1(net5821));
 sg13g2_nand2_1 _14348_ (.Y(_05333_),
    .A(_05310_),
    .B(_05332_));
 sg13g2_a21oi_1 _14349_ (.A1(_05319_),
    .A2(_05321_),
    .Y(_05334_),
    .B1(net5273));
 sg13g2_o21ai_1 _14350_ (.B1(_05334_),
    .Y(_05335_),
    .A1(_05330_),
    .A2(_05331_));
 sg13g2_a21oi_1 _14351_ (.A1(_05333_),
    .A2(_05335_),
    .Y(_05336_),
    .B1(net5812));
 sg13g2_and2_1 _14352_ (.A(net6132),
    .B(\mem.mem[227][5] ),
    .X(_05337_));
 sg13g2_a21oi_1 _14353_ (.A1(net5411),
    .A2(\mem.mem[226][5] ),
    .Y(_05338_),
    .B1(_05337_));
 sg13g2_nand2_1 _14354_ (.Y(_05339_),
    .A(net6132),
    .B(\mem.mem[225][5] ));
 sg13g2_a21oi_1 _14355_ (.A1(net5411),
    .A2(\mem.mem[224][5] ),
    .Y(_05340_),
    .B1(net5973));
 sg13g2_a221oi_1 _14356_ (.B2(_05340_),
    .C1(net5875),
    .B1(_05339_),
    .A1(net5973),
    .Y(_05341_),
    .A2(_05338_));
 sg13g2_mux4_1 _14357_ (.S0(net6138),
    .A0(\mem.mem[228][5] ),
    .A1(\mem.mem[229][5] ),
    .A2(\mem.mem[230][5] ),
    .A3(\mem.mem[231][5] ),
    .S1(net5978),
    .X(_05342_));
 sg13g2_a21oi_2 _14358_ (.B1(_05341_),
    .Y(_05343_),
    .A2(_05342_),
    .A1(net5877));
 sg13g2_mux4_1 _14359_ (.S0(net6139),
    .A0(\mem.mem[232][5] ),
    .A1(\mem.mem[233][5] ),
    .A2(\mem.mem[234][5] ),
    .A3(\mem.mem[235][5] ),
    .S1(net5978),
    .X(_05344_));
 sg13g2_nand2_1 _14360_ (.Y(_05345_),
    .A(net5339),
    .B(_05344_));
 sg13g2_mux4_1 _14361_ (.S0(net6145),
    .A0(\mem.mem[236][5] ),
    .A1(\mem.mem[237][5] ),
    .A2(\mem.mem[238][5] ),
    .A3(\mem.mem[239][5] ),
    .S1(net5983),
    .X(_05346_));
 sg13g2_a21oi_1 _14362_ (.A1(net5877),
    .A2(_05346_),
    .Y(_05347_),
    .B1(net5293));
 sg13g2_mux4_1 _14363_ (.S0(net6048),
    .A0(\mem.mem[248][5] ),
    .A1(\mem.mem[249][5] ),
    .A2(\mem.mem[250][5] ),
    .A3(\mem.mem[251][5] ),
    .S1(net5915),
    .X(_05348_));
 sg13g2_nand2_1 _14364_ (.Y(_05349_),
    .A(net5857),
    .B(\mem.mem[252][5] ));
 sg13g2_a21oi_1 _14365_ (.A1(net5310),
    .A2(_05348_),
    .Y(_05350_),
    .B1(net5281));
 sg13g2_mux4_1 _14366_ (.S0(net6055),
    .A0(\mem.mem[240][5] ),
    .A1(\mem.mem[241][5] ),
    .A2(\mem.mem[242][5] ),
    .A3(\mem.mem[243][5] ),
    .S1(net5921),
    .X(_05351_));
 sg13g2_mux4_1 _14367_ (.S0(net6053),
    .A0(\mem.mem[244][5] ),
    .A1(\mem.mem[245][5] ),
    .A2(\mem.mem[246][5] ),
    .A3(\mem.mem[247][5] ),
    .S1(net5918),
    .X(_05352_));
 sg13g2_nand2_1 _14368_ (.Y(_05353_),
    .A(net5857),
    .B(_05352_));
 sg13g2_a21oi_1 _14369_ (.A1(net5311),
    .A2(_05351_),
    .Y(_05354_),
    .B1(net5831));
 sg13g2_a22oi_1 _14370_ (.Y(_05355_),
    .B1(_05353_),
    .B2(_05354_),
    .A2(_05350_),
    .A1(_05349_));
 sg13g2_a221oi_1 _14371_ (.B2(_05347_),
    .C1(net5823),
    .B1(_05345_),
    .A1(net5293),
    .Y(_05356_),
    .A2(_05343_));
 sg13g2_a21o_1 _14372_ (.A2(_05355_),
    .A1(net5821),
    .B1(_05356_),
    .X(_05357_));
 sg13g2_a21o_2 _14373_ (.A2(_05357_),
    .A1(net5812),
    .B1(_05336_),
    .X(_05358_));
 sg13g2_mux4_1 _14374_ (.S0(net6061),
    .A0(\mem.mem[164][5] ),
    .A1(\mem.mem[165][5] ),
    .A2(\mem.mem[166][5] ),
    .A3(\mem.mem[167][5] ),
    .S1(net5922),
    .X(_05359_));
 sg13g2_mux4_1 _14375_ (.S0(net6056),
    .A0(\mem.mem[160][5] ),
    .A1(\mem.mem[161][5] ),
    .A2(\mem.mem[162][5] ),
    .A3(\mem.mem[163][5] ),
    .S1(net5920),
    .X(_05360_));
 sg13g2_nand2_1 _14376_ (.Y(_05361_),
    .A(net5313),
    .B(_05360_));
 sg13g2_a21oi_1 _14377_ (.A1(net5858),
    .A2(_05359_),
    .Y(_05362_),
    .B1(net5831));
 sg13g2_nor2b_1 _14378_ (.A(net6060),
    .B_N(\mem.mem[170][5] ),
    .Y(_05363_));
 sg13g2_a21oi_1 _14379_ (.A1(net6060),
    .A2(\mem.mem[171][5] ),
    .Y(_05364_),
    .B1(_05363_));
 sg13g2_nand2_1 _14380_ (.Y(_05365_),
    .A(net6060),
    .B(\mem.mem[169][5] ));
 sg13g2_nand2_1 _14381_ (.Y(_05366_),
    .A(net5387),
    .B(\mem.mem[168][5] ));
 sg13g2_nand3_1 _14382_ (.B(_05365_),
    .C(_05366_),
    .A(net5353),
    .Y(_05367_));
 sg13g2_a21oi_1 _14383_ (.A1(net5923),
    .A2(_05364_),
    .Y(_05368_),
    .B1(net5858));
 sg13g2_mux4_1 _14384_ (.S0(net6061),
    .A0(\mem.mem[172][5] ),
    .A1(\mem.mem[173][5] ),
    .A2(\mem.mem[174][5] ),
    .A3(\mem.mem[175][5] ),
    .S1(net5923),
    .X(_05369_));
 sg13g2_a221oi_1 _14385_ (.B2(net5858),
    .C1(net5282),
    .B1(_05369_),
    .A1(_05367_),
    .Y(_05370_),
    .A2(_05368_));
 sg13g2_a21oi_2 _14386_ (.B1(_05370_),
    .Y(_05371_),
    .A2(_05362_),
    .A1(_05361_));
 sg13g2_and2_1 _14387_ (.A(net6137),
    .B(\mem.mem[191][5] ),
    .X(_05372_));
 sg13g2_a21oi_1 _14388_ (.A1(net5409),
    .A2(\mem.mem[190][5] ),
    .Y(_05373_),
    .B1(_05372_));
 sg13g2_mux2_1 _14389_ (.A0(\mem.mem[188][5] ),
    .A1(\mem.mem[189][5] ),
    .S(net6101),
    .X(_05374_));
 sg13g2_o21ai_1 _14390_ (.B1(net5876),
    .Y(_05375_),
    .A1(net5952),
    .A2(_05374_));
 sg13g2_a21o_1 _14391_ (.A2(_05373_),
    .A1(net5975),
    .B1(_05375_),
    .X(_05376_));
 sg13g2_mux4_1 _14392_ (.S0(net6131),
    .A0(\mem.mem[184][5] ),
    .A1(\mem.mem[185][5] ),
    .A2(\mem.mem[186][5] ),
    .A3(\mem.mem[187][5] ),
    .S1(net5972),
    .X(_05377_));
 sg13g2_a21oi_1 _14393_ (.A1(net5334),
    .A2(_05377_),
    .Y(_05378_),
    .B1(net5292));
 sg13g2_mux4_1 _14394_ (.S0(net6131),
    .A0(\mem.mem[176][5] ),
    .A1(\mem.mem[177][5] ),
    .A2(\mem.mem[178][5] ),
    .A3(\mem.mem[179][5] ),
    .S1(net5974),
    .X(_05379_));
 sg13g2_nand2_1 _14395_ (.Y(_05380_),
    .A(net5334),
    .B(_05379_));
 sg13g2_mux4_1 _14396_ (.S0(net6134),
    .A0(\mem.mem[180][5] ),
    .A1(\mem.mem[181][5] ),
    .A2(\mem.mem[182][5] ),
    .A3(\mem.mem[183][5] ),
    .S1(net5975),
    .X(_05381_));
 sg13g2_a21oi_1 _14397_ (.A1(net5876),
    .A2(_05381_),
    .Y(_05382_),
    .B1(net5845));
 sg13g2_a22oi_1 _14398_ (.Y(_05383_),
    .B1(_05380_),
    .B2(_05382_),
    .A2(_05378_),
    .A1(_05376_));
 sg13g2_mux4_1 _14399_ (.S0(net6116),
    .A0(\mem.mem[128][5] ),
    .A1(\mem.mem[129][5] ),
    .A2(\mem.mem[130][5] ),
    .A3(\mem.mem[131][5] ),
    .S1(net5963),
    .X(_05384_));
 sg13g2_nand2_1 _14400_ (.Y(_05385_),
    .A(net5332),
    .B(_05384_));
 sg13g2_mux4_1 _14401_ (.S0(net6119),
    .A0(\mem.mem[132][5] ),
    .A1(\mem.mem[133][5] ),
    .A2(\mem.mem[134][5] ),
    .A3(\mem.mem[135][5] ),
    .S1(net5964),
    .X(_05386_));
 sg13g2_a21oi_1 _14402_ (.A1(net5872),
    .A2(_05386_),
    .Y(_05387_),
    .B1(net5840));
 sg13g2_nor2b_1 _14403_ (.A(net6121),
    .B_N(\mem.mem[138][5] ),
    .Y(_05388_));
 sg13g2_a21oi_1 _14404_ (.A1(net6121),
    .A2(\mem.mem[139][5] ),
    .Y(_05389_),
    .B1(_05388_));
 sg13g2_nand2_1 _14405_ (.Y(_05390_),
    .A(net6121),
    .B(\mem.mem[137][5] ));
 sg13g2_nand2_1 _14406_ (.Y(_05391_),
    .A(net5406),
    .B(\mem.mem[136][5] ));
 sg13g2_nand3_1 _14407_ (.B(_05390_),
    .C(_05391_),
    .A(net5363),
    .Y(_05392_));
 sg13g2_a21oi_1 _14408_ (.A1(net5966),
    .A2(_05389_),
    .Y(_05393_),
    .B1(net5871));
 sg13g2_mux4_1 _14409_ (.S0(net6113),
    .A0(\mem.mem[140][5] ),
    .A1(\mem.mem[141][5] ),
    .A2(\mem.mem[142][5] ),
    .A3(\mem.mem[143][5] ),
    .S1(net5959),
    .X(_05394_));
 sg13g2_a221oi_1 _14410_ (.B2(net5871),
    .C1(net5291),
    .B1(_05394_),
    .A1(_05392_),
    .Y(_05395_),
    .A2(_05393_));
 sg13g2_a21oi_2 _14411_ (.B1(_05395_),
    .Y(_05396_),
    .A2(_05387_),
    .A1(_05385_));
 sg13g2_mux4_1 _14412_ (.S0(net6090),
    .A0(\mem.mem[152][5] ),
    .A1(\mem.mem[153][5] ),
    .A2(\mem.mem[154][5] ),
    .A3(\mem.mem[155][5] ),
    .S1(net5946),
    .X(_05397_));
 sg13g2_nand2_1 _14413_ (.Y(_05398_),
    .A(net5328),
    .B(_05397_));
 sg13g2_mux4_1 _14414_ (.S0(net6106),
    .A0(\mem.mem[156][5] ),
    .A1(\mem.mem[157][5] ),
    .A2(\mem.mem[158][5] ),
    .A3(\mem.mem[159][5] ),
    .S1(net5955),
    .X(_05399_));
 sg13g2_a21oi_1 _14415_ (.A1(net5869),
    .A2(_05399_),
    .Y(_05400_),
    .B1(net5290));
 sg13g2_mux4_1 _14416_ (.S0(net6106),
    .A0(\mem.mem[144][5] ),
    .A1(\mem.mem[145][5] ),
    .A2(\mem.mem[146][5] ),
    .A3(\mem.mem[147][5] ),
    .S1(net5955),
    .X(_05401_));
 sg13g2_nand2_1 _14417_ (.Y(_05402_),
    .A(net5328),
    .B(_05401_));
 sg13g2_nand2_1 _14418_ (.Y(_05403_),
    .A(net5402),
    .B(\mem.mem[150][5] ));
 sg13g2_a21oi_1 _14419_ (.A1(net6108),
    .A2(\mem.mem[151][5] ),
    .Y(_05404_),
    .B1(net5361));
 sg13g2_nand2b_1 _14420_ (.Y(_05405_),
    .B(net6108),
    .A_N(\mem.mem[149][5] ));
 sg13g2_o21ai_1 _14421_ (.B1(_05405_),
    .Y(_05406_),
    .A1(net6108),
    .A2(\mem.mem[148][5] ));
 sg13g2_a221oi_1 _14422_ (.B2(net5361),
    .C1(net5328),
    .B1(_05406_),
    .A1(_05403_),
    .Y(_05407_),
    .A2(_05404_));
 sg13g2_nor2_1 _14423_ (.A(net5841),
    .B(_05407_),
    .Y(_05408_));
 sg13g2_a22oi_1 _14424_ (.Y(_05409_),
    .B1(_05402_),
    .B2(_05408_),
    .A2(_05400_),
    .A1(_05398_));
 sg13g2_mux4_1 _14425_ (.S0(net5825),
    .A0(_05371_),
    .A1(_05383_),
    .A2(_05396_),
    .A3(_05409_),
    .S1(net5265),
    .X(_05410_));
 sg13g2_mux4_1 _14426_ (.S0(net5263),
    .A0(_05220_),
    .A1(_05303_),
    .A2(_05358_),
    .A3(_05410_),
    .S1(_00007_),
    .X(_05411_));
 sg13g2_a22oi_1 _14427_ (.Y(_05412_),
    .B1(_05411_),
    .B2(_02945_),
    .A2(_03639_),
    .A1(net7));
 sg13g2_o21ai_1 _14428_ (.B1(net6187),
    .Y(_05413_),
    .A1(net5788),
    .A2(net4178));
 sg13g2_a21oi_1 _14429_ (.A1(net5789),
    .A2(_05412_),
    .Y(_00553_),
    .B1(_05413_));
 sg13g2_a21oi_1 _14430_ (.A1(net6078),
    .A2(\mem.mem[5][6] ),
    .Y(_05414_),
    .B1(net5934));
 sg13g2_o21ai_1 _14431_ (.B1(_05414_),
    .Y(_05415_),
    .A1(net6075),
    .A2(_02869_));
 sg13g2_and2_1 _14432_ (.A(net6075),
    .B(\mem.mem[7][6] ),
    .X(_05416_));
 sg13g2_a21oi_1 _14433_ (.A1(net5391),
    .A2(\mem.mem[6][6] ),
    .Y(_05417_),
    .B1(_05416_));
 sg13g2_a21oi_1 _14434_ (.A1(net5934),
    .A2(_05417_),
    .Y(_05418_),
    .B1(net5320));
 sg13g2_mux4_1 _14435_ (.S0(net6079),
    .A0(\mem.mem[0][6] ),
    .A1(\mem.mem[1][6] ),
    .A2(\mem.mem[2][6] ),
    .A3(\mem.mem[3][6] ),
    .S1(net5936),
    .X(_05419_));
 sg13g2_a221oi_1 _14436_ (.B2(net5318),
    .C1(net5835),
    .B1(_05419_),
    .A1(_05415_),
    .Y(_05420_),
    .A2(_05418_));
 sg13g2_mux4_1 _14437_ (.S0(net6081),
    .A0(\mem.mem[8][6] ),
    .A1(\mem.mem[9][6] ),
    .A2(\mem.mem[10][6] ),
    .A3(\mem.mem[11][6] ),
    .S1(net5938),
    .X(_05421_));
 sg13g2_a21oi_1 _14438_ (.A1(net6109),
    .A2(\mem.mem[15][6] ),
    .Y(_05422_),
    .B1(net5356));
 sg13g2_o21ai_1 _14439_ (.B1(_05422_),
    .Y(_05423_),
    .A1(net6109),
    .A2(_02870_));
 sg13g2_nand2_1 _14440_ (.Y(_05424_),
    .A(net6081),
    .B(\mem.mem[13][6] ));
 sg13g2_a21oi_1 _14441_ (.A1(net5393),
    .A2(\mem.mem[12][6] ),
    .Y(_05425_),
    .B1(net5938));
 sg13g2_a21oi_1 _14442_ (.A1(_05424_),
    .A2(_05425_),
    .Y(_05426_),
    .B1(net5319));
 sg13g2_a221oi_1 _14443_ (.B2(_05426_),
    .C1(net5283),
    .B1(_05423_),
    .A1(net5318),
    .Y(_05427_),
    .A2(_05421_));
 sg13g2_o21ai_1 _14444_ (.B1(net5268),
    .Y(_05428_),
    .A1(_05420_),
    .A2(_05427_));
 sg13g2_mux2_1 _14445_ (.A0(\mem.mem[22][6] ),
    .A1(\mem.mem[23][6] ),
    .S(net6125),
    .X(_05429_));
 sg13g2_a21o_1 _14446_ (.A2(\mem.mem[21][6] ),
    .A1(net6155),
    .B1(net5968),
    .X(_05430_));
 sg13g2_a21oi_1 _14447_ (.A1(net5416),
    .A2(\mem.mem[20][6] ),
    .Y(_05431_),
    .B1(_05430_));
 sg13g2_o21ai_1 _14448_ (.B1(net5880),
    .Y(_05432_),
    .A1(net5363),
    .A2(_05429_));
 sg13g2_mux4_1 _14449_ (.S0(net6156),
    .A0(\mem.mem[16][6] ),
    .A1(\mem.mem[17][6] ),
    .A2(\mem.mem[18][6] ),
    .A3(\mem.mem[19][6] ),
    .S1(net5991),
    .X(_05433_));
 sg13g2_a21oi_1 _14450_ (.A1(net5341),
    .A2(_05433_),
    .Y(_05434_),
    .B1(net5846));
 sg13g2_o21ai_1 _14451_ (.B1(_05434_),
    .Y(_05435_),
    .A1(_05431_),
    .A2(_05432_));
 sg13g2_nand2_1 _14452_ (.Y(_05436_),
    .A(net5415),
    .B(\mem.mem[24][6] ));
 sg13g2_a21oi_1 _14453_ (.A1(net6149),
    .A2(\mem.mem[25][6] ),
    .Y(_05437_),
    .B1(net5987));
 sg13g2_nor2b_1 _14454_ (.A(net6149),
    .B_N(\mem.mem[26][6] ),
    .Y(_05438_));
 sg13g2_a21oi_1 _14455_ (.A1(net6149),
    .A2(\mem.mem[27][6] ),
    .Y(_05439_),
    .B1(_05438_));
 sg13g2_a221oi_1 _14456_ (.B2(net5987),
    .C1(net5880),
    .B1(_05439_),
    .A1(_05436_),
    .Y(_05440_),
    .A2(_05437_));
 sg13g2_mux2_1 _14457_ (.A0(\mem.mem[28][6] ),
    .A1(\mem.mem[29][6] ),
    .S(net6149),
    .X(_05441_));
 sg13g2_a21o_1 _14458_ (.A2(\mem.mem[30][6] ),
    .A1(net5415),
    .B1(net5367),
    .X(_05442_));
 sg13g2_a21oi_1 _14459_ (.A1(net6150),
    .A2(\mem.mem[31][6] ),
    .Y(_05443_),
    .B1(_05442_));
 sg13g2_o21ai_1 _14460_ (.B1(net5880),
    .Y(_05444_),
    .A1(net5987),
    .A2(_05441_));
 sg13g2_o21ai_1 _14461_ (.B1(net5846),
    .Y(_05445_),
    .A1(_05443_),
    .A2(_05444_));
 sg13g2_o21ai_1 _14462_ (.B1(_05435_),
    .Y(_05446_),
    .A1(_05440_),
    .A2(_05445_));
 sg13g2_a21oi_1 _14463_ (.A1(net5820),
    .A2(_05446_),
    .Y(_05447_),
    .B1(net5815));
 sg13g2_nor2b_1 _14464_ (.A(net6166),
    .B_N(\mem.mem[38][6] ),
    .Y(_05448_));
 sg13g2_a21oi_1 _14465_ (.A1(net6166),
    .A2(\mem.mem[39][6] ),
    .Y(_05449_),
    .B1(_05448_));
 sg13g2_nand2_1 _14466_ (.Y(_05450_),
    .A(net5420),
    .B(\mem.mem[36][6] ));
 sg13g2_a21oi_1 _14467_ (.A1(net6166),
    .A2(\mem.mem[37][6] ),
    .Y(_05451_),
    .B1(net5999));
 sg13g2_a221oi_1 _14468_ (.B2(_05451_),
    .C1(net5344),
    .B1(_05450_),
    .A1(net5999),
    .Y(_05452_),
    .A2(_05449_));
 sg13g2_nand2_1 _14469_ (.Y(_05453_),
    .A(net5420),
    .B(\mem.mem[32][6] ));
 sg13g2_a21oi_1 _14470_ (.A1(net6166),
    .A2(\mem.mem[33][6] ),
    .Y(_05454_),
    .B1(net6000));
 sg13g2_nor2b_1 _14471_ (.A(net6167),
    .B_N(\mem.mem[34][6] ),
    .Y(_05455_));
 sg13g2_a21oi_1 _14472_ (.A1(net6167),
    .A2(\mem.mem[35][6] ),
    .Y(_05456_),
    .B1(_05455_));
 sg13g2_a221oi_1 _14473_ (.B2(net5999),
    .C1(net5881),
    .B1(_05456_),
    .A1(_05453_),
    .Y(_05457_),
    .A2(_05454_));
 sg13g2_or3_1 _14474_ (.A(net5847),
    .B(_05452_),
    .C(_05457_),
    .X(_05458_));
 sg13g2_nand2_1 _14475_ (.Y(_05459_),
    .A(net5420),
    .B(\mem.mem[40][6] ));
 sg13g2_a21oi_1 _14476_ (.A1(net6168),
    .A2(\mem.mem[41][6] ),
    .Y(_05460_),
    .B1(net6000));
 sg13g2_nor2b_1 _14477_ (.A(net6168),
    .B_N(\mem.mem[42][6] ),
    .Y(_05461_));
 sg13g2_a21oi_1 _14478_ (.A1(net6168),
    .A2(\mem.mem[43][6] ),
    .Y(_05462_),
    .B1(_05461_));
 sg13g2_a221oi_1 _14479_ (.B2(net6000),
    .C1(net5881),
    .B1(_05462_),
    .A1(_05459_),
    .Y(_05463_),
    .A2(_05460_));
 sg13g2_mux2_1 _14480_ (.A0(\mem.mem[44][6] ),
    .A1(\mem.mem[45][6] ),
    .S(net6164),
    .X(_05464_));
 sg13g2_a21o_1 _14481_ (.A2(\mem.mem[46][6] ),
    .A1(net5419),
    .B1(net5367),
    .X(_05465_));
 sg13g2_a21oi_1 _14482_ (.A1(net6164),
    .A2(\mem.mem[47][6] ),
    .Y(_05466_),
    .B1(_05465_));
 sg13g2_o21ai_1 _14483_ (.B1(net5881),
    .Y(_05467_),
    .A1(net5999),
    .A2(_05464_));
 sg13g2_o21ai_1 _14484_ (.B1(net5847),
    .Y(_05468_),
    .A1(_05466_),
    .A2(_05467_));
 sg13g2_o21ai_1 _14485_ (.B1(_05458_),
    .Y(_05469_),
    .A1(_05463_),
    .A2(_05468_));
 sg13g2_a21oi_1 _14486_ (.A1(net6026),
    .A2(\mem.mem[53][6] ),
    .Y(_05470_),
    .B1(net5902));
 sg13g2_o21ai_1 _14487_ (.B1(_05470_),
    .Y(_05471_),
    .A1(net6026),
    .A2(_02871_));
 sg13g2_and2_1 _14488_ (.A(net6028),
    .B(\mem.mem[55][6] ),
    .X(_05472_));
 sg13g2_a21oi_1 _14489_ (.A1(net5379),
    .A2(\mem.mem[54][6] ),
    .Y(_05473_),
    .B1(_05472_));
 sg13g2_a21oi_1 _14490_ (.A1(net5901),
    .A2(_05473_),
    .Y(_05474_),
    .B1(net5305));
 sg13g2_mux4_1 _14491_ (.S0(net6028),
    .A0(\mem.mem[48][6] ),
    .A1(\mem.mem[49][6] ),
    .A2(\mem.mem[50][6] ),
    .A3(\mem.mem[51][6] ),
    .S1(net5901),
    .X(_05475_));
 sg13g2_a221oi_1 _14492_ (.B2(net5305),
    .C1(net5829),
    .B1(_05475_),
    .A1(_05471_),
    .Y(_05476_),
    .A2(_05474_));
 sg13g2_nand2_1 _14493_ (.Y(_05477_),
    .A(net5377),
    .B(\mem.mem[56][6] ));
 sg13g2_a21oi_1 _14494_ (.A1(net6029),
    .A2(\mem.mem[57][6] ),
    .Y(_05478_),
    .B1(net5904));
 sg13g2_nor2b_1 _14495_ (.A(net6029),
    .B_N(\mem.mem[58][6] ),
    .Y(_05479_));
 sg13g2_a21oi_1 _14496_ (.A1(net6034),
    .A2(\mem.mem[59][6] ),
    .Y(_05480_),
    .B1(_05479_));
 sg13g2_a221oi_1 _14497_ (.B2(net5904),
    .C1(net5854),
    .B1(_05480_),
    .A1(_05477_),
    .Y(_05481_),
    .A2(_05478_));
 sg13g2_nor2b_1 _14498_ (.A(net6031),
    .B_N(\mem.mem[62][6] ),
    .Y(_05482_));
 sg13g2_a21oi_1 _14499_ (.A1(net6031),
    .A2(\mem.mem[63][6] ),
    .Y(_05483_),
    .B1(_05482_));
 sg13g2_nand2_1 _14500_ (.Y(_05484_),
    .A(net5377),
    .B(\mem.mem[60][6] ));
 sg13g2_a21oi_1 _14501_ (.A1(net6031),
    .A2(\mem.mem[61][6] ),
    .Y(_05485_),
    .B1(net5905));
 sg13g2_a221oi_1 _14502_ (.B2(_05485_),
    .C1(net5304),
    .B1(_05484_),
    .A1(net5905),
    .Y(_05486_),
    .A2(_05483_));
 sg13g2_nor3_2 _14503_ (.A(net5279),
    .B(_05481_),
    .C(_05486_),
    .Y(_05487_));
 sg13g2_o21ai_1 _14504_ (.B1(net5817),
    .Y(_05488_),
    .A1(_05476_),
    .A2(_05487_));
 sg13g2_a21oi_2 _14505_ (.B1(net5265),
    .Y(_05489_),
    .A2(_05469_),
    .A1(net5271));
 sg13g2_a221oi_1 _14506_ (.B2(_05489_),
    .C1(net5807),
    .B1(_05488_),
    .A1(_05428_),
    .Y(_05490_),
    .A2(_05447_));
 sg13g2_mux4_1 _14507_ (.S0(net6012),
    .A0(\mem.mem[76][6] ),
    .A1(\mem.mem[77][6] ),
    .A2(\mem.mem[78][6] ),
    .A3(\mem.mem[79][6] ),
    .S1(net5890),
    .X(_05491_));
 sg13g2_nand2_1 _14508_ (.Y(_05492_),
    .A(net5850),
    .B(_05491_));
 sg13g2_mux4_1 _14509_ (.S0(net6017),
    .A0(\mem.mem[72][6] ),
    .A1(\mem.mem[73][6] ),
    .A2(\mem.mem[74][6] ),
    .A3(\mem.mem[75][6] ),
    .S1(net5894),
    .X(_05493_));
 sg13g2_mux4_1 _14510_ (.S0(net6017),
    .A0(\mem.mem[68][6] ),
    .A1(\mem.mem[69][6] ),
    .A2(\mem.mem[70][6] ),
    .A3(\mem.mem[71][6] ),
    .S1(net5894),
    .X(_05494_));
 sg13g2_nand2_1 _14511_ (.Y(_05495_),
    .A(net5852),
    .B(_05494_));
 sg13g2_mux4_1 _14512_ (.S0(net6006),
    .A0(\mem.mem[64][6] ),
    .A1(\mem.mem[65][6] ),
    .A2(\mem.mem[66][6] ),
    .A3(\mem.mem[67][6] ),
    .S1(net5886),
    .X(_05496_));
 sg13g2_and2_1 _14513_ (.A(net6024),
    .B(\mem.mem[95][6] ),
    .X(_05497_));
 sg13g2_a21oi_1 _14514_ (.A1(net5373),
    .A2(\mem.mem[94][6] ),
    .Y(_05498_),
    .B1(_05497_));
 sg13g2_mux2_1 _14515_ (.A0(\mem.mem[92][6] ),
    .A1(\mem.mem[93][6] ),
    .S(net6019),
    .X(_05499_));
 sg13g2_o21ai_1 _14516_ (.B1(net5852),
    .Y(_05500_),
    .A1(net5895),
    .A2(_05499_));
 sg13g2_a21o_1 _14517_ (.A2(_05498_),
    .A1(net5895),
    .B1(_05500_),
    .X(_05501_));
 sg13g2_mux4_1 _14518_ (.S0(net6018),
    .A0(\mem.mem[88][6] ),
    .A1(\mem.mem[89][6] ),
    .A2(\mem.mem[90][6] ),
    .A3(\mem.mem[91][6] ),
    .S1(net5895),
    .X(_05502_));
 sg13g2_a21oi_1 _14519_ (.A1(net5303),
    .A2(_05502_),
    .Y(_05503_),
    .B1(net5276));
 sg13g2_mux4_1 _14520_ (.S0(net6006),
    .A0(\mem.mem[80][6] ),
    .A1(\mem.mem[81][6] ),
    .A2(\mem.mem[82][6] ),
    .A3(\mem.mem[83][6] ),
    .S1(net5886),
    .X(_05504_));
 sg13g2_nand2_2 _14521_ (.Y(_05505_),
    .A(net5298),
    .B(_05504_));
 sg13g2_mux4_1 _14522_ (.S0(net6006),
    .A0(\mem.mem[84][6] ),
    .A1(\mem.mem[85][6] ),
    .A2(\mem.mem[86][6] ),
    .A3(\mem.mem[87][6] ),
    .S1(net5886),
    .X(_05506_));
 sg13g2_a21oi_2 _14523_ (.B1(net5827),
    .Y(_05507_),
    .A2(_05506_),
    .A1(net5850));
 sg13g2_a21oi_1 _14524_ (.A1(net5298),
    .A2(_05496_),
    .Y(_05508_),
    .B1(net5827));
 sg13g2_a21oi_1 _14525_ (.A1(net5302),
    .A2(_05493_),
    .Y(_05509_),
    .B1(net5278));
 sg13g2_a221oi_1 _14526_ (.B2(_05492_),
    .C1(net5816),
    .B1(_05509_),
    .A1(_05495_),
    .Y(_05510_),
    .A2(_05508_));
 sg13g2_a221oi_1 _14527_ (.B2(_05507_),
    .C1(net5270),
    .B1(_05505_),
    .A1(_05501_),
    .Y(_05511_),
    .A2(_05503_));
 sg13g2_or2_2 _14528_ (.X(_05512_),
    .B(_05511_),
    .A(_05510_));
 sg13g2_a21oi_1 _14529_ (.A1(net6068),
    .A2(\mem.mem[103][6] ),
    .Y(_05513_),
    .B1(net5355));
 sg13g2_o21ai_1 _14530_ (.B1(_05513_),
    .Y(_05514_),
    .A1(net6068),
    .A2(_02872_));
 sg13g2_nand2_1 _14531_ (.Y(_05515_),
    .A(net5389),
    .B(\mem.mem[100][6] ));
 sg13g2_a21oi_1 _14532_ (.A1(net6070),
    .A2(\mem.mem[101][6] ),
    .Y(_05516_),
    .B1(net5929));
 sg13g2_a21oi_1 _14533_ (.A1(_05515_),
    .A2(_05516_),
    .Y(_05517_),
    .B1(net5316));
 sg13g2_mux4_1 _14534_ (.S0(net6069),
    .A0(\mem.mem[96][6] ),
    .A1(\mem.mem[97][6] ),
    .A2(\mem.mem[98][6] ),
    .A3(\mem.mem[99][6] ),
    .S1(net5928),
    .X(_05518_));
 sg13g2_a221oi_1 _14535_ (.B2(net5316),
    .C1(net5834),
    .B1(_05518_),
    .A1(_05514_),
    .Y(_05519_),
    .A2(_05517_));
 sg13g2_mux4_1 _14536_ (.S0(net6063),
    .A0(\mem.mem[104][6] ),
    .A1(\mem.mem[105][6] ),
    .A2(\mem.mem[106][6] ),
    .A3(\mem.mem[107][6] ),
    .S1(net5927),
    .X(_05520_));
 sg13g2_mux2_1 _14537_ (.A0(\mem.mem[108][6] ),
    .A1(\mem.mem[109][6] ),
    .S(net6066),
    .X(_05521_));
 sg13g2_a21o_1 _14538_ (.A2(\mem.mem[110][6] ),
    .A1(net5391),
    .B1(net5355),
    .X(_05522_));
 sg13g2_a21oi_1 _14539_ (.A1(net6074),
    .A2(\mem.mem[111][6] ),
    .Y(_05523_),
    .B1(_05522_));
 sg13g2_o21ai_1 _14540_ (.B1(net5861),
    .Y(_05524_),
    .A1(net5925),
    .A2(_05521_));
 sg13g2_o21ai_1 _14541_ (.B1(net5833),
    .Y(_05525_),
    .A1(_05523_),
    .A2(_05524_));
 sg13g2_a21oi_1 _14542_ (.A1(net5315),
    .A2(_05520_),
    .Y(_05526_),
    .B1(_05525_));
 sg13g2_o21ai_1 _14543_ (.B1(net5268),
    .Y(_05527_),
    .A1(_05519_),
    .A2(_05526_));
 sg13g2_a21oi_1 _14544_ (.A1(net6035),
    .A2(\mem.mem[117][6] ),
    .Y(_05528_),
    .B1(net5908));
 sg13g2_o21ai_1 _14545_ (.B1(_05528_),
    .Y(_05529_),
    .A1(net6037),
    .A2(_02873_));
 sg13g2_and2_1 _14546_ (.A(net6036),
    .B(\mem.mem[119][6] ),
    .X(_05530_));
 sg13g2_a21oi_1 _14547_ (.A1(net5380),
    .A2(\mem.mem[118][6] ),
    .Y(_05531_),
    .B1(_05530_));
 sg13g2_a21oi_1 _14548_ (.A1(net5909),
    .A2(_05531_),
    .Y(_05532_),
    .B1(net5306));
 sg13g2_mux4_1 _14549_ (.S0(net6037),
    .A0(\mem.mem[112][6] ),
    .A1(\mem.mem[113][6] ),
    .A2(\mem.mem[114][6] ),
    .A3(\mem.mem[115][6] ),
    .S1(net5909),
    .X(_05533_));
 sg13g2_a221oi_1 _14550_ (.B2(net5306),
    .C1(net5830),
    .B1(_05533_),
    .A1(_05529_),
    .Y(_05534_),
    .A2(_05532_));
 sg13g2_nand2_1 _14551_ (.Y(_05535_),
    .A(net5382),
    .B(\mem.mem[120][6] ));
 sg13g2_a21oi_1 _14552_ (.A1(net6068),
    .A2(\mem.mem[121][6] ),
    .Y(_05536_),
    .B1(net5911));
 sg13g2_nor2b_1 _14553_ (.A(net6042),
    .B_N(\mem.mem[122][6] ),
    .Y(_05537_));
 sg13g2_a21oi_1 _14554_ (.A1(net6042),
    .A2(\mem.mem[123][6] ),
    .Y(_05538_),
    .B1(_05537_));
 sg13g2_a221oi_1 _14555_ (.B2(net5911),
    .C1(net5855),
    .B1(_05538_),
    .A1(_05535_),
    .Y(_05539_),
    .A2(_05536_));
 sg13g2_nor2b_1 _14556_ (.A(net6040),
    .B_N(\mem.mem[126][6] ),
    .Y(_05540_));
 sg13g2_a21oi_1 _14557_ (.A1(net6040),
    .A2(\mem.mem[127][6] ),
    .Y(_05541_),
    .B1(_05540_));
 sg13g2_nand2_1 _14558_ (.Y(_05542_),
    .A(net5382),
    .B(\mem.mem[124][6] ));
 sg13g2_a21oi_1 _14559_ (.A1(net6040),
    .A2(\mem.mem[125][6] ),
    .Y(_05543_),
    .B1(net5910));
 sg13g2_a221oi_1 _14560_ (.B2(_05543_),
    .C1(net5307),
    .B1(_05542_),
    .A1(net5910),
    .Y(_05544_),
    .A2(_05541_));
 sg13g2_nor3_1 _14561_ (.A(net5280),
    .B(_05539_),
    .C(_05544_),
    .Y(_05545_));
 sg13g2_o21ai_1 _14562_ (.B1(net5818),
    .Y(_05546_),
    .A1(_05534_),
    .A2(_05545_));
 sg13g2_and2_1 _14563_ (.A(net5809),
    .B(_05546_),
    .X(_05547_));
 sg13g2_a221oi_1 _14564_ (.B2(_05547_),
    .C1(net5262),
    .B1(_05527_),
    .A1(net5264),
    .Y(_05548_),
    .A2(_05512_));
 sg13g2_o21ai_1 _14565_ (.B1(_02840_),
    .Y(_05549_),
    .A1(_05490_),
    .A2(_05548_));
 sg13g2_mux4_1 _14566_ (.S0(net6085),
    .A0(\mem.mem[160][6] ),
    .A1(\mem.mem[161][6] ),
    .A2(\mem.mem[162][6] ),
    .A3(\mem.mem[163][6] ),
    .S1(net5943),
    .X(_05550_));
 sg13g2_nand2_1 _14567_ (.Y(_05551_),
    .A(net5313),
    .B(_05550_));
 sg13g2_mux4_1 _14568_ (.S0(net6058),
    .A0(\mem.mem[164][6] ),
    .A1(\mem.mem[165][6] ),
    .A2(\mem.mem[166][6] ),
    .A3(\mem.mem[167][6] ),
    .S1(net5922),
    .X(_05552_));
 sg13g2_a21oi_1 _14569_ (.A1(net5858),
    .A2(_05552_),
    .Y(_05553_),
    .B1(net5831));
 sg13g2_mux4_1 _14570_ (.S0(net6057),
    .A0(\mem.mem[168][6] ),
    .A1(\mem.mem[169][6] ),
    .A2(\mem.mem[170][6] ),
    .A3(\mem.mem[171][6] ),
    .S1(net5920),
    .X(_05554_));
 sg13g2_nand2_1 _14571_ (.Y(_05555_),
    .A(net5313),
    .B(_05554_));
 sg13g2_mux4_1 _14572_ (.S0(net6060),
    .A0(\mem.mem[172][6] ),
    .A1(\mem.mem[173][6] ),
    .A2(\mem.mem[174][6] ),
    .A3(\mem.mem[175][6] ),
    .S1(net5923),
    .X(_05556_));
 sg13g2_a21oi_1 _14573_ (.A1(net5858),
    .A2(_05556_),
    .Y(_05557_),
    .B1(net5282));
 sg13g2_nand2_1 _14574_ (.Y(_05558_),
    .A(net6134),
    .B(\mem.mem[189][6] ));
 sg13g2_a21oi_1 _14575_ (.A1(net5409),
    .A2(\mem.mem[188][6] ),
    .Y(_05559_),
    .B1(net5952));
 sg13g2_and2_1 _14576_ (.A(net6134),
    .B(\mem.mem[191][6] ),
    .X(_05560_));
 sg13g2_a21oi_1 _14577_ (.A1(net5409),
    .A2(\mem.mem[190][6] ),
    .Y(_05561_),
    .B1(_05560_));
 sg13g2_a221oi_1 _14578_ (.B2(net5952),
    .C1(net5325),
    .B1(_05561_),
    .A1(_05558_),
    .Y(_05562_),
    .A2(_05559_));
 sg13g2_mux4_1 _14579_ (.S0(net6130),
    .A0(\mem.mem[184][6] ),
    .A1(\mem.mem[185][6] ),
    .A2(\mem.mem[186][6] ),
    .A3(\mem.mem[187][6] ),
    .S1(net5972),
    .X(_05563_));
 sg13g2_nand2_1 _14580_ (.Y(_05564_),
    .A(net5334),
    .B(_05563_));
 sg13g2_nor2_1 _14581_ (.A(net5292),
    .B(_05562_),
    .Y(_05565_));
 sg13g2_mux4_1 _14582_ (.S0(net6134),
    .A0(\mem.mem[180][6] ),
    .A1(\mem.mem[181][6] ),
    .A2(\mem.mem[182][6] ),
    .A3(\mem.mem[183][6] ),
    .S1(net5975),
    .X(_05566_));
 sg13g2_nand2_1 _14583_ (.Y(_05567_),
    .A(net5876),
    .B(_05566_));
 sg13g2_mux4_1 _14584_ (.S0(net6130),
    .A0(\mem.mem[176][6] ),
    .A1(\mem.mem[177][6] ),
    .A2(\mem.mem[178][6] ),
    .A3(\mem.mem[179][6] ),
    .S1(net5972),
    .X(_05568_));
 sg13g2_a21oi_1 _14585_ (.A1(net5334),
    .A2(_05568_),
    .Y(_05569_),
    .B1(net5845));
 sg13g2_a221oi_1 _14586_ (.B2(_05557_),
    .C1(net5820),
    .B1(_05555_),
    .A1(_05551_),
    .Y(_05570_),
    .A2(_05553_));
 sg13g2_a221oi_1 _14587_ (.B2(_05569_),
    .C1(net5273),
    .B1(_05567_),
    .A1(_05564_),
    .Y(_05571_),
    .A2(_05565_));
 sg13g2_o21ai_1 _14588_ (.B1(net5812),
    .Y(_05572_),
    .A1(_05570_),
    .A2(_05571_));
 sg13g2_mux4_1 _14589_ (.S0(net6121),
    .A0(\mem.mem[136][6] ),
    .A1(\mem.mem[137][6] ),
    .A2(\mem.mem[138][6] ),
    .A3(\mem.mem[139][6] ),
    .S1(net5966),
    .X(_05573_));
 sg13g2_mux4_1 _14590_ (.S0(net6122),
    .A0(\mem.mem[140][6] ),
    .A1(\mem.mem[141][6] ),
    .A2(\mem.mem[142][6] ),
    .A3(\mem.mem[143][6] ),
    .S1(net5966),
    .X(_05574_));
 sg13g2_nand2_1 _14591_ (.Y(_05575_),
    .A(net5871),
    .B(_05574_));
 sg13g2_a21oi_1 _14592_ (.A1(net5331),
    .A2(_05573_),
    .Y(_05576_),
    .B1(net5291));
 sg13g2_nor2b_1 _14593_ (.A(net6117),
    .B_N(\mem.mem[130][6] ),
    .Y(_05577_));
 sg13g2_a21oi_1 _14594_ (.A1(net6117),
    .A2(\mem.mem[131][6] ),
    .Y(_05578_),
    .B1(_05577_));
 sg13g2_mux2_1 _14595_ (.A0(\mem.mem[128][6] ),
    .A1(\mem.mem[129][6] ),
    .S(net6116),
    .X(_05579_));
 sg13g2_a21oi_1 _14596_ (.A1(net5963),
    .A2(_05578_),
    .Y(_05580_),
    .B1(net5872));
 sg13g2_o21ai_1 _14597_ (.B1(_05580_),
    .Y(_05581_),
    .A1(net5963),
    .A2(_05579_));
 sg13g2_nand2_1 _14598_ (.Y(_05582_),
    .A(net5405),
    .B(\mem.mem[134][6] ));
 sg13g2_a21oi_1 _14599_ (.A1(net6119),
    .A2(\mem.mem[135][6] ),
    .Y(_05583_),
    .B1(net5362));
 sg13g2_nand2b_1 _14600_ (.Y(_05584_),
    .B(net6118),
    .A_N(\mem.mem[133][6] ));
 sg13g2_o21ai_1 _14601_ (.B1(_05584_),
    .Y(_05585_),
    .A1(net6118),
    .A2(\mem.mem[132][6] ));
 sg13g2_a221oi_1 _14602_ (.B2(net5362),
    .C1(net5332),
    .B1(_05585_),
    .A1(_05582_),
    .Y(_05586_),
    .A2(_05583_));
 sg13g2_nor2_1 _14603_ (.A(net5840),
    .B(_05586_),
    .Y(_05587_));
 sg13g2_mux4_1 _14604_ (.S0(net6092),
    .A0(\mem.mem[152][6] ),
    .A1(\mem.mem[153][6] ),
    .A2(\mem.mem[154][6] ),
    .A3(\mem.mem[155][6] ),
    .S1(net5947),
    .X(_05588_));
 sg13g2_nand2_1 _14605_ (.Y(_05589_),
    .A(net5328),
    .B(_05588_));
 sg13g2_mux4_1 _14606_ (.S0(net6107),
    .A0(\mem.mem[156][6] ),
    .A1(\mem.mem[157][6] ),
    .A2(\mem.mem[158][6] ),
    .A3(\mem.mem[159][6] ),
    .S1(net5957),
    .X(_05590_));
 sg13g2_mux4_1 _14607_ (.S0(net6076),
    .A0(\mem.mem[144][6] ),
    .A1(\mem.mem[145][6] ),
    .A2(\mem.mem[146][6] ),
    .A3(\mem.mem[147][6] ),
    .S1(net5933),
    .X(_05591_));
 sg13g2_nand2_1 _14608_ (.Y(_05592_),
    .A(net5328),
    .B(_05591_));
 sg13g2_mux4_1 _14609_ (.S0(net6108),
    .A0(\mem.mem[148][6] ),
    .A1(\mem.mem[149][6] ),
    .A2(\mem.mem[150][6] ),
    .A3(\mem.mem[151][6] ),
    .S1(net5957),
    .X(_05593_));
 sg13g2_a221oi_1 _14610_ (.B2(_05587_),
    .C1(net5825),
    .B1(_05581_),
    .A1(_05575_),
    .Y(_05594_),
    .A2(_05576_));
 sg13g2_a21oi_1 _14611_ (.A1(net5869),
    .A2(_05593_),
    .Y(_05595_),
    .B1(net5841));
 sg13g2_a21oi_1 _14612_ (.A1(net5869),
    .A2(_05590_),
    .Y(_05596_),
    .B1(net5290));
 sg13g2_a221oi_1 _14613_ (.B2(_05589_),
    .C1(net5271),
    .B1(_05596_),
    .A1(_05592_),
    .Y(_05597_),
    .A2(_05595_));
 sg13g2_nor2_1 _14614_ (.A(_05594_),
    .B(_05597_),
    .Y(_05598_));
 sg13g2_nor2_1 _14615_ (.A(net5813),
    .B(_05598_),
    .Y(_05599_));
 sg13g2_nor2_1 _14616_ (.A(net5807),
    .B(_05599_),
    .Y(_05600_));
 sg13g2_mux2_1 _14617_ (.A0(\mem.mem[204][6] ),
    .A1(\mem.mem[205][6] ),
    .S(net6098),
    .X(_05601_));
 sg13g2_nor2_1 _14618_ (.A(net5396),
    .B(\mem.mem[207][6] ),
    .Y(_05602_));
 sg13g2_o21ai_1 _14619_ (.B1(net5944),
    .Y(_05603_),
    .A1(net6098),
    .A2(\mem.mem[206][6] ));
 sg13g2_o21ai_1 _14620_ (.B1(net5867),
    .Y(_05604_),
    .A1(_05602_),
    .A2(_05603_));
 sg13g2_a21oi_1 _14621_ (.A1(net5357),
    .A2(_05601_),
    .Y(_05605_),
    .B1(_05604_));
 sg13g2_mux4_1 _14622_ (.S0(net6087),
    .A0(\mem.mem[200][6] ),
    .A1(\mem.mem[201][6] ),
    .A2(\mem.mem[202][6] ),
    .A3(\mem.mem[203][6] ),
    .S1(net5944),
    .X(_05606_));
 sg13g2_nor2_1 _14623_ (.A(net5289),
    .B(_05605_),
    .Y(_05607_));
 sg13g2_o21ai_1 _14624_ (.B1(_05607_),
    .Y(_05608_),
    .A1(net5867),
    .A2(_05606_));
 sg13g2_mux4_1 _14625_ (.S0(net6095),
    .A0(\mem.mem[192][6] ),
    .A1(\mem.mem[193][6] ),
    .A2(\mem.mem[194][6] ),
    .A3(\mem.mem[195][6] ),
    .S1(net5951),
    .X(_05609_));
 sg13g2_mux2_1 _14626_ (.A0(\mem.mem[198][6] ),
    .A1(\mem.mem[199][6] ),
    .S(net6098),
    .X(_05610_));
 sg13g2_nand2_1 _14627_ (.Y(_05611_),
    .A(net5954),
    .B(_05610_));
 sg13g2_mux2_1 _14628_ (.A0(\mem.mem[196][6] ),
    .A1(\mem.mem[197][6] ),
    .S(net6097),
    .X(_05612_));
 sg13g2_a21oi_1 _14629_ (.A1(net5359),
    .A2(_05612_),
    .Y(_05613_),
    .B1(net5326));
 sg13g2_a21oi_1 _14630_ (.A1(_05611_),
    .A2(_05613_),
    .Y(_05614_),
    .B1(net5839));
 sg13g2_o21ai_1 _14631_ (.B1(_05614_),
    .Y(_05615_),
    .A1(net5867),
    .A2(_05609_));
 sg13g2_nand3_1 _14632_ (.B(_05608_),
    .C(_05615_),
    .A(net5272),
    .Y(_05616_));
 sg13g2_nand2_1 _14633_ (.Y(_05617_),
    .A(net5413),
    .B(\mem.mem[212][6] ));
 sg13g2_a21oi_1 _14634_ (.A1(net6146),
    .A2(\mem.mem[213][6] ),
    .Y(_05618_),
    .B1(net5981));
 sg13g2_and2_1 _14635_ (.A(net6146),
    .B(\mem.mem[215][6] ),
    .X(_05619_));
 sg13g2_a21oi_1 _14636_ (.A1(net5412),
    .A2(\mem.mem[214][6] ),
    .Y(_05620_),
    .B1(_05619_));
 sg13g2_a221oi_1 _14637_ (.B2(net5981),
    .C1(net5338),
    .B1(_05620_),
    .A1(_05617_),
    .Y(_05621_),
    .A2(_05618_));
 sg13g2_nand2_1 _14638_ (.Y(_05622_),
    .A(net5419),
    .B(\mem.mem[208][6] ));
 sg13g2_a21oi_1 _14639_ (.A1(net6163),
    .A2(\mem.mem[209][6] ),
    .Y(_05623_),
    .B1(net5996));
 sg13g2_nor2b_1 _14640_ (.A(net6163),
    .B_N(\mem.mem[210][6] ),
    .Y(_05624_));
 sg13g2_a21oi_1 _14641_ (.A1(net6163),
    .A2(\mem.mem[211][6] ),
    .Y(_05625_),
    .B1(_05624_));
 sg13g2_a221oi_1 _14642_ (.B2(net5996),
    .C1(net5882),
    .B1(_05625_),
    .A1(_05622_),
    .Y(_05626_),
    .A2(_05623_));
 sg13g2_nor3_2 _14643_ (.A(net5844),
    .B(_05621_),
    .C(_05626_),
    .Y(_05627_));
 sg13g2_mux4_1 _14644_ (.S0(net6153),
    .A0(\mem.mem[216][6] ),
    .A1(\mem.mem[217][6] ),
    .A2(\mem.mem[218][6] ),
    .A3(\mem.mem[219][6] ),
    .S1(net6003),
    .X(_05628_));
 sg13g2_a21oi_1 _14645_ (.A1(net6154),
    .A2(\mem.mem[223][6] ),
    .Y(_05629_),
    .B1(net5367));
 sg13g2_o21ai_1 _14646_ (.B1(_05629_),
    .Y(_05630_),
    .A1(net6152),
    .A2(_02874_));
 sg13g2_nand2_1 _14647_ (.Y(_05631_),
    .A(net6153),
    .B(\mem.mem[221][6] ));
 sg13g2_a21oi_1 _14648_ (.A1(net5418),
    .A2(\mem.mem[220][6] ),
    .Y(_05632_),
    .B1(net5989));
 sg13g2_a21oi_1 _14649_ (.A1(_05631_),
    .A2(_05632_),
    .Y(_05633_),
    .B1(net5340));
 sg13g2_a221oi_1 _14650_ (.B2(_05633_),
    .C1(net5295),
    .B1(_05630_),
    .A1(net5340),
    .Y(_05634_),
    .A2(_05628_));
 sg13g2_o21ai_1 _14651_ (.B1(net5823),
    .Y(_05635_),
    .A1(_05627_),
    .A2(_05634_));
 sg13g2_nand3_1 _14652_ (.B(_05616_),
    .C(_05635_),
    .A(net5266),
    .Y(_05636_));
 sg13g2_a21o_1 _14653_ (.A2(\mem.mem[231][6] ),
    .A1(net6138),
    .B1(net5365),
    .X(_05637_));
 sg13g2_a21oi_1 _14654_ (.A1(net5414),
    .A2(\mem.mem[230][6] ),
    .Y(_05638_),
    .B1(_05637_));
 sg13g2_mux2_1 _14655_ (.A0(\mem.mem[228][6] ),
    .A1(\mem.mem[229][6] ),
    .S(net6138),
    .X(_05639_));
 sg13g2_o21ai_1 _14656_ (.B1(net5877),
    .Y(_05640_),
    .A1(net5978),
    .A2(_05639_));
 sg13g2_mux4_1 _14657_ (.S0(net6138),
    .A0(\mem.mem[224][6] ),
    .A1(\mem.mem[225][6] ),
    .A2(\mem.mem[226][6] ),
    .A3(\mem.mem[227][6] ),
    .S1(net5978),
    .X(_05641_));
 sg13g2_a21oi_1 _14658_ (.A1(net5339),
    .A2(_05641_),
    .Y(_05642_),
    .B1(net5843));
 sg13g2_o21ai_1 _14659_ (.B1(_05642_),
    .Y(_05643_),
    .A1(_05638_),
    .A2(_05640_));
 sg13g2_nand2_1 _14660_ (.Y(_05644_),
    .A(net5414),
    .B(\mem.mem[232][6] ));
 sg13g2_a21oi_1 _14661_ (.A1(net6140),
    .A2(\mem.mem[233][6] ),
    .Y(_05645_),
    .B1(net5979));
 sg13g2_nor2b_1 _14662_ (.A(net6141),
    .B_N(\mem.mem[234][6] ),
    .Y(_05646_));
 sg13g2_a21oi_1 _14663_ (.A1(net6140),
    .A2(\mem.mem[235][6] ),
    .Y(_05647_),
    .B1(_05646_));
 sg13g2_a221oi_1 _14664_ (.B2(net5980),
    .C1(net5878),
    .B1(_05647_),
    .A1(_05644_),
    .Y(_05648_),
    .A2(_05645_));
 sg13g2_mux2_1 _14665_ (.A0(\mem.mem[236][6] ),
    .A1(\mem.mem[237][6] ),
    .S(net6140),
    .X(_05649_));
 sg13g2_a21o_1 _14666_ (.A2(\mem.mem[238][6] ),
    .A1(net5412),
    .B1(net5365),
    .X(_05650_));
 sg13g2_a21oi_1 _14667_ (.A1(net6145),
    .A2(\mem.mem[239][6] ),
    .Y(_05651_),
    .B1(_05650_));
 sg13g2_o21ai_1 _14668_ (.B1(net5877),
    .Y(_05652_),
    .A1(net5979),
    .A2(_05649_));
 sg13g2_o21ai_1 _14669_ (.B1(net5843),
    .Y(_05653_),
    .A1(_05651_),
    .A2(_05652_));
 sg13g2_o21ai_1 _14670_ (.B1(_05643_),
    .Y(_05654_),
    .A1(_05648_),
    .A2(_05653_));
 sg13g2_mux4_1 _14671_ (.S0(net6048),
    .A0(\mem.mem[248][6] ),
    .A1(\mem.mem[249][6] ),
    .A2(\mem.mem[250][6] ),
    .A3(\mem.mem[251][6] ),
    .S1(net5915),
    .X(_05655_));
 sg13g2_mux4_1 _14672_ (.S0(net6058),
    .A0(\mem.mem[244][6] ),
    .A1(\mem.mem[245][6] ),
    .A2(\mem.mem[246][6] ),
    .A3(\mem.mem[247][6] ),
    .S1(net5922),
    .X(_05656_));
 sg13g2_mux4_1 _14673_ (.S0(net6057),
    .A0(\mem.mem[240][6] ),
    .A1(\mem.mem[241][6] ),
    .A2(\mem.mem[242][6] ),
    .A3(\mem.mem[243][6] ),
    .S1(net5921),
    .X(_05657_));
 sg13g2_mux4_1 _14674_ (.S0(net5312),
    .A0(\mem.mem[252][6] ),
    .A1(_05655_),
    .A2(_05656_),
    .A3(_05657_),
    .S1(net5285),
    .X(_05658_));
 sg13g2_o21ai_1 _14675_ (.B1(net5811),
    .Y(_05659_),
    .A1(net5269),
    .A2(_05658_));
 sg13g2_a21oi_2 _14676_ (.B1(_05659_),
    .Y(_05660_),
    .A2(_05654_),
    .A1(net5272));
 sg13g2_nor2_1 _14677_ (.A(net5263),
    .B(_05660_),
    .Y(_05661_));
 sg13g2_a22oi_1 _14678_ (.Y(_05662_),
    .B1(_05636_),
    .B2(_05661_),
    .A2(_05600_),
    .A1(_05572_));
 sg13g2_nand2b_2 _14679_ (.Y(_05663_),
    .B(_00007_),
    .A_N(_05662_));
 sg13g2_and2_1 _14680_ (.A(_02945_),
    .B(_05549_),
    .X(_05664_));
 sg13g2_a22oi_1 _14681_ (.Y(_05665_),
    .B1(_05663_),
    .B2(_05664_),
    .A2(_03639_),
    .A1(net8));
 sg13g2_o21ai_1 _14682_ (.B1(net6188),
    .Y(_05666_),
    .A1(net5788),
    .A2(net4188));
 sg13g2_a21oi_1 _14683_ (.A1(net5788),
    .A2(_05665_),
    .Y(_00554_),
    .B1(_05666_));
 sg13g2_mux4_1 _14684_ (.S0(net6079),
    .A0(\mem.mem[0][7] ),
    .A1(\mem.mem[1][7] ),
    .A2(\mem.mem[2][7] ),
    .A3(\mem.mem[3][7] ),
    .S1(net5936),
    .X(_05667_));
 sg13g2_nor2_2 _14685_ (.A(net5862),
    .B(_05667_),
    .Y(_05668_));
 sg13g2_mux2_1 _14686_ (.A0(\mem.mem[4][7] ),
    .A1(\mem.mem[5][7] ),
    .S(net6077),
    .X(_05669_));
 sg13g2_nor2_1 _14687_ (.A(net5391),
    .B(\mem.mem[7][7] ),
    .Y(_05670_));
 sg13g2_o21ai_1 _14688_ (.B1(net5934),
    .Y(_05671_),
    .A1(net6075),
    .A2(\mem.mem[6][7] ));
 sg13g2_o21ai_1 _14689_ (.B1(net5863),
    .Y(_05672_),
    .A1(_05670_),
    .A2(_05671_));
 sg13g2_a21oi_1 _14690_ (.A1(net5356),
    .A2(_05669_),
    .Y(_05673_),
    .B1(_05672_));
 sg13g2_nor3_1 _14691_ (.A(net5835),
    .B(_05668_),
    .C(_05673_),
    .Y(_05674_));
 sg13g2_mux4_1 _14692_ (.S0(net6083),
    .A0(\mem.mem[8][7] ),
    .A1(\mem.mem[9][7] ),
    .A2(\mem.mem[10][7] ),
    .A3(\mem.mem[11][7] ),
    .S1(net5939),
    .X(_05675_));
 sg13g2_nor2_1 _14693_ (.A(net5862),
    .B(_05675_),
    .Y(_05676_));
 sg13g2_mux2_1 _14694_ (.A0(\mem.mem[12][7] ),
    .A1(\mem.mem[13][7] ),
    .S(net6082),
    .X(_05677_));
 sg13g2_nor2_1 _14695_ (.A(net5403),
    .B(\mem.mem[15][7] ),
    .Y(_05678_));
 sg13g2_o21ai_1 _14696_ (.B1(net5958),
    .Y(_05679_),
    .A1(net6110),
    .A2(\mem.mem[14][7] ));
 sg13g2_o21ai_1 _14697_ (.B1(net5870),
    .Y(_05680_),
    .A1(_05678_),
    .A2(_05679_));
 sg13g2_a21oi_1 _14698_ (.A1(net5356),
    .A2(_05677_),
    .Y(_05681_),
    .B1(_05680_));
 sg13g2_nor3_2 _14699_ (.A(net5283),
    .B(_05676_),
    .C(_05681_),
    .Y(_05682_));
 sg13g2_nor2_1 _14700_ (.A(_05674_),
    .B(_05682_),
    .Y(_05683_));
 sg13g2_a21oi_1 _14701_ (.A1(net5407),
    .A2(_02876_),
    .Y(_05684_),
    .B1(net5362));
 sg13g2_o21ai_1 _14702_ (.B1(_05684_),
    .Y(_05685_),
    .A1(net5406),
    .A2(\mem.mem[23][7] ));
 sg13g2_mux2_1 _14703_ (.A0(\mem.mem[20][7] ),
    .A1(\mem.mem[21][7] ),
    .S(net6127),
    .X(_05686_));
 sg13g2_a21oi_1 _14704_ (.A1(net5363),
    .A2(_05686_),
    .Y(_05687_),
    .B1(net5331));
 sg13g2_mux2_1 _14705_ (.A0(\mem.mem[18][7] ),
    .A1(\mem.mem[19][7] ),
    .S(net6122),
    .X(_05688_));
 sg13g2_nand2_1 _14706_ (.Y(_05689_),
    .A(net5966),
    .B(_05688_));
 sg13g2_mux2_1 _14707_ (.A0(\mem.mem[16][7] ),
    .A1(\mem.mem[17][7] ),
    .S(net6123),
    .X(_05690_));
 sg13g2_a21oi_1 _14708_ (.A1(net5363),
    .A2(_05690_),
    .Y(_05691_),
    .B1(net5871));
 sg13g2_a221oi_1 _14709_ (.B2(_05691_),
    .C1(net5840),
    .B1(_05689_),
    .A1(_05685_),
    .Y(_05692_),
    .A2(_05687_));
 sg13g2_mux4_1 _14710_ (.S0(net6120),
    .A0(\mem.mem[24][7] ),
    .A1(\mem.mem[25][7] ),
    .A2(\mem.mem[26][7] ),
    .A3(\mem.mem[27][7] ),
    .S1(net5964),
    .X(_05693_));
 sg13g2_nor2_1 _14711_ (.A(net5872),
    .B(_05693_),
    .Y(_05694_));
 sg13g2_nor2_1 _14712_ (.A(net5415),
    .B(\mem.mem[29][7] ),
    .Y(_05695_));
 sg13g2_nor2_1 _14713_ (.A(net6151),
    .B(\mem.mem[28][7] ),
    .Y(_05696_));
 sg13g2_nor3_1 _14714_ (.A(net5988),
    .B(_05695_),
    .C(_05696_),
    .Y(_05697_));
 sg13g2_nor2_1 _14715_ (.A(net5415),
    .B(\mem.mem[31][7] ),
    .Y(_05698_));
 sg13g2_o21ai_1 _14716_ (.B1(net5988),
    .Y(_05699_),
    .A1(net6150),
    .A2(\mem.mem[30][7] ));
 sg13g2_o21ai_1 _14717_ (.B1(net5880),
    .Y(_05700_),
    .A1(_05698_),
    .A2(_05699_));
 sg13g2_o21ai_1 _14718_ (.B1(net5846),
    .Y(_05701_),
    .A1(_05697_),
    .A2(_05700_));
 sg13g2_o21ai_1 _14719_ (.B1(net5822),
    .Y(_05702_),
    .A1(_05694_),
    .A2(_05701_));
 sg13g2_o21ai_1 _14720_ (.B1(net5266),
    .Y(_05703_),
    .A1(_05692_),
    .A2(_05702_));
 sg13g2_a21oi_1 _14721_ (.A1(net5268),
    .A2(_05683_),
    .Y(_05704_),
    .B1(_05703_));
 sg13g2_nor2b_1 _14722_ (.A(net6166),
    .B_N(\mem.mem[38][7] ),
    .Y(_05705_));
 sg13g2_a21oi_1 _14723_ (.A1(net6166),
    .A2(\mem.mem[39][7] ),
    .Y(_05706_),
    .B1(_05705_));
 sg13g2_nand2_1 _14724_ (.Y(_05707_),
    .A(net5417),
    .B(\mem.mem[36][7] ));
 sg13g2_a21oi_1 _14725_ (.A1(net6158),
    .A2(\mem.mem[37][7] ),
    .Y(_05708_),
    .B1(net5992));
 sg13g2_a221oi_1 _14726_ (.B2(_05708_),
    .C1(net5342),
    .B1(_05707_),
    .A1(net5993),
    .Y(_05709_),
    .A2(_05706_));
 sg13g2_nand2_1 _14727_ (.Y(_05710_),
    .A(net5420),
    .B(\mem.mem[32][7] ));
 sg13g2_a21oi_1 _14728_ (.A1(net6167),
    .A2(\mem.mem[33][7] ),
    .Y(_05711_),
    .B1(net5993));
 sg13g2_nor2b_1 _14729_ (.A(net6160),
    .B_N(\mem.mem[34][7] ),
    .Y(_05712_));
 sg13g2_a21oi_1 _14730_ (.A1(net6167),
    .A2(\mem.mem[35][7] ),
    .Y(_05713_),
    .B1(_05712_));
 sg13g2_a221oi_1 _14731_ (.B2(net5993),
    .C1(net5881),
    .B1(_05713_),
    .A1(_05710_),
    .Y(_05714_),
    .A2(_05711_));
 sg13g2_nor3_1 _14732_ (.A(net5848),
    .B(_05709_),
    .C(_05714_),
    .Y(_05715_));
 sg13g2_mux4_1 _14733_ (.S0(net6170),
    .A0(\mem.mem[40][7] ),
    .A1(\mem.mem[41][7] ),
    .A2(\mem.mem[42][7] ),
    .A3(\mem.mem[43][7] ),
    .S1(net6001),
    .X(_05716_));
 sg13g2_mux2_1 _14734_ (.A0(\mem.mem[44][7] ),
    .A1(\mem.mem[45][7] ),
    .S(net6171),
    .X(_05717_));
 sg13g2_a21o_1 _14735_ (.A2(\mem.mem[46][7] ),
    .A1(net5421),
    .B1(net5367),
    .X(_05718_));
 sg13g2_a21oi_1 _14736_ (.A1(net6170),
    .A2(\mem.mem[47][7] ),
    .Y(_05719_),
    .B1(_05718_));
 sg13g2_o21ai_1 _14737_ (.B1(net5881),
    .Y(_05720_),
    .A1(net6001),
    .A2(_05717_));
 sg13g2_o21ai_1 _14738_ (.B1(net5847),
    .Y(_05721_),
    .A1(_05719_),
    .A2(_05720_));
 sg13g2_a21oi_1 _14739_ (.A1(net5345),
    .A2(_05716_),
    .Y(_05722_),
    .B1(_05721_));
 sg13g2_o21ai_1 _14740_ (.B1(net5274),
    .Y(_05723_),
    .A1(_05715_),
    .A2(_05722_));
 sg13g2_nand2_1 _14741_ (.Y(_05724_),
    .A(net5379),
    .B(\mem.mem[52][7] ));
 sg13g2_a21oi_1 _14742_ (.A1(net6026),
    .A2(\mem.mem[53][7] ),
    .Y(_05725_),
    .B1(net5902));
 sg13g2_and2_1 _14743_ (.A(net6026),
    .B(\mem.mem[55][7] ),
    .X(_05726_));
 sg13g2_a21oi_1 _14744_ (.A1(net5379),
    .A2(\mem.mem[54][7] ),
    .Y(_05727_),
    .B1(_05726_));
 sg13g2_a221oi_1 _14745_ (.B2(net5902),
    .C1(net5305),
    .B1(_05727_),
    .A1(_05724_),
    .Y(_05728_),
    .A2(_05725_));
 sg13g2_nand2_1 _14746_ (.Y(_05729_),
    .A(net5370),
    .B(\mem.mem[48][7] ));
 sg13g2_a21oi_1 _14747_ (.A1(net6010),
    .A2(\mem.mem[49][7] ),
    .Y(_05730_),
    .B1(net5889));
 sg13g2_nor2b_1 _14748_ (.A(net6010),
    .B_N(\mem.mem[50][7] ),
    .Y(_05731_));
 sg13g2_a21oi_1 _14749_ (.A1(net6010),
    .A2(\mem.mem[51][7] ),
    .Y(_05732_),
    .B1(_05731_));
 sg13g2_a221oi_1 _14750_ (.B2(net5889),
    .C1(net5850),
    .B1(_05732_),
    .A1(_05729_),
    .Y(_05733_),
    .A2(_05730_));
 sg13g2_nor3_1 _14751_ (.A(net5829),
    .B(_05728_),
    .C(_05733_),
    .Y(_05734_));
 sg13g2_mux4_1 _14752_ (.S0(net6032),
    .A0(\mem.mem[56][7] ),
    .A1(\mem.mem[57][7] ),
    .A2(\mem.mem[58][7] ),
    .A3(\mem.mem[59][7] ),
    .S1(net5905),
    .X(_05735_));
 sg13g2_a21oi_1 _14753_ (.A1(net6033),
    .A2(\mem.mem[63][7] ),
    .Y(_05736_),
    .B1(net5350));
 sg13g2_o21ai_1 _14754_ (.B1(_05736_),
    .Y(_05737_),
    .A1(net6033),
    .A2(_02877_));
 sg13g2_nand2_1 _14755_ (.Y(_05738_),
    .A(net6039),
    .B(\mem.mem[61][7] ));
 sg13g2_a21oi_1 _14756_ (.A1(net5378),
    .A2(\mem.mem[60][7] ),
    .Y(_05739_),
    .B1(net5906));
 sg13g2_a21oi_1 _14757_ (.A1(_05738_),
    .A2(_05739_),
    .Y(_05740_),
    .B1(net5305));
 sg13g2_a221oi_1 _14758_ (.B2(_05740_),
    .C1(net5279),
    .B1(_05737_),
    .A1(net5304),
    .Y(_05741_),
    .A2(_05735_));
 sg13g2_o21ai_1 _14759_ (.B1(net5817),
    .Y(_05742_),
    .A1(_05734_),
    .A2(_05741_));
 sg13g2_nand3_1 _14760_ (.B(_05723_),
    .C(_05742_),
    .A(net5809),
    .Y(_05743_));
 sg13g2_nor2_2 _14761_ (.A(net5808),
    .B(_05704_),
    .Y(_05744_));
 sg13g2_mux2_1 _14762_ (.A0(\mem.mem[76][7] ),
    .A1(\mem.mem[77][7] ),
    .S(net6022),
    .X(_05745_));
 sg13g2_nand2_1 _14763_ (.Y(_05746_),
    .A(net5349),
    .B(_05745_));
 sg13g2_mux2_1 _14764_ (.A0(\mem.mem[78][7] ),
    .A1(\mem.mem[79][7] ),
    .S(net6012),
    .X(_05747_));
 sg13g2_a21oi_1 _14765_ (.A1(net5890),
    .A2(_05747_),
    .Y(_05748_),
    .B1(net5300));
 sg13g2_mux4_1 _14766_ (.S0(net6022),
    .A0(\mem.mem[72][7] ),
    .A1(\mem.mem[73][7] ),
    .A2(\mem.mem[74][7] ),
    .A3(\mem.mem[75][7] ),
    .S1(net5897),
    .X(_05749_));
 sg13g2_o21ai_1 _14767_ (.B1(net5828),
    .Y(_05750_),
    .A1(net5853),
    .A2(_05749_));
 sg13g2_a21oi_1 _14768_ (.A1(_05746_),
    .A2(_05748_),
    .Y(_05751_),
    .B1(_05750_));
 sg13g2_mux4_1 _14769_ (.S0(net6006),
    .A0(\mem.mem[64][7] ),
    .A1(\mem.mem[65][7] ),
    .A2(\mem.mem[66][7] ),
    .A3(\mem.mem[67][7] ),
    .S1(net5886),
    .X(_05752_));
 sg13g2_nor2_1 _14770_ (.A(net5850),
    .B(_05752_),
    .Y(_05753_));
 sg13g2_mux2_1 _14771_ (.A0(\mem.mem[70][7] ),
    .A1(\mem.mem[71][7] ),
    .S(net6015),
    .X(_05754_));
 sg13g2_nand2b_1 _14772_ (.Y(_05755_),
    .B(net6015),
    .A_N(\mem.mem[69][7] ));
 sg13g2_o21ai_1 _14773_ (.B1(_05755_),
    .Y(_05756_),
    .A1(net6015),
    .A2(\mem.mem[68][7] ));
 sg13g2_o21ai_1 _14774_ (.B1(net5850),
    .Y(_05757_),
    .A1(net5892),
    .A2(_05756_));
 sg13g2_a21oi_1 _14775_ (.A1(net5892),
    .A2(_05754_),
    .Y(_05758_),
    .B1(_05757_));
 sg13g2_nor3_2 _14776_ (.A(net5827),
    .B(_05753_),
    .C(_05758_),
    .Y(_05759_));
 sg13g2_nor3_2 _14777_ (.A(net5816),
    .B(_05751_),
    .C(_05759_),
    .Y(_05760_));
 sg13g2_mux4_1 _14778_ (.S0(net6005),
    .A0(\mem.mem[80][7] ),
    .A1(\mem.mem[81][7] ),
    .A2(\mem.mem[82][7] ),
    .A3(\mem.mem[83][7] ),
    .S1(net5885),
    .X(_05761_));
 sg13g2_nor2_2 _14779_ (.A(net5850),
    .B(_05761_),
    .Y(_05762_));
 sg13g2_mux2_1 _14780_ (.A0(\mem.mem[86][7] ),
    .A1(\mem.mem[87][7] ),
    .S(net6009),
    .X(_05763_));
 sg13g2_nand2b_1 _14781_ (.Y(_05764_),
    .B(net6012),
    .A_N(\mem.mem[85][7] ));
 sg13g2_o21ai_1 _14782_ (.B1(_05764_),
    .Y(_05765_),
    .A1(net6012),
    .A2(\mem.mem[84][7] ));
 sg13g2_o21ai_1 _14783_ (.B1(net5851),
    .Y(_05766_),
    .A1(net5888),
    .A2(_05765_));
 sg13g2_a21oi_1 _14784_ (.A1(net5888),
    .A2(_05763_),
    .Y(_05767_),
    .B1(_05766_));
 sg13g2_nor3_2 _14785_ (.A(net5828),
    .B(_05762_),
    .C(_05767_),
    .Y(_05768_));
 sg13g2_mux4_1 _14786_ (.S0(net6046),
    .A0(\mem.mem[88][7] ),
    .A1(\mem.mem[89][7] ),
    .A2(\mem.mem[90][7] ),
    .A3(\mem.mem[91][7] ),
    .S1(net5916),
    .X(_05769_));
 sg13g2_nor2_1 _14787_ (.A(net5852),
    .B(_05769_),
    .Y(_05770_));
 sg13g2_nor2_1 _14788_ (.A(net5386),
    .B(\mem.mem[93][7] ),
    .Y(_05771_));
 sg13g2_nor2_1 _14789_ (.A(net6051),
    .B(\mem.mem[92][7] ),
    .Y(_05772_));
 sg13g2_nor3_1 _14790_ (.A(net5917),
    .B(_05771_),
    .C(_05772_),
    .Y(_05773_));
 sg13g2_nor2_1 _14791_ (.A(net5385),
    .B(\mem.mem[95][7] ),
    .Y(_05774_));
 sg13g2_o21ai_1 _14792_ (.B1(net5917),
    .Y(_05775_),
    .A1(net6051),
    .A2(\mem.mem[94][7] ));
 sg13g2_o21ai_1 _14793_ (.B1(net5860),
    .Y(_05776_),
    .A1(_05774_),
    .A2(_05775_));
 sg13g2_o21ai_1 _14794_ (.B1(net5831),
    .Y(_05777_),
    .A1(_05773_),
    .A2(_05776_));
 sg13g2_o21ai_1 _14795_ (.B1(net5816),
    .Y(_05778_),
    .A1(_05770_),
    .A2(_05777_));
 sg13g2_o21ai_1 _14796_ (.B1(net5264),
    .Y(_05779_),
    .A1(_05768_),
    .A2(_05778_));
 sg13g2_nor2_1 _14797_ (.A(_05760_),
    .B(_05779_),
    .Y(_05780_));
 sg13g2_nor2b_1 _14798_ (.A(net6070),
    .B_N(\mem.mem[102][7] ),
    .Y(_05781_));
 sg13g2_a21oi_1 _14799_ (.A1(net6068),
    .A2(\mem.mem[103][7] ),
    .Y(_05782_),
    .B1(_05781_));
 sg13g2_nand2_1 _14800_ (.Y(_05783_),
    .A(net5389),
    .B(\mem.mem[100][7] ));
 sg13g2_a21oi_1 _14801_ (.A1(net6068),
    .A2(\mem.mem[101][7] ),
    .Y(_05784_),
    .B1(net5929));
 sg13g2_a221oi_1 _14802_ (.B2(_05784_),
    .C1(net5316),
    .B1(_05783_),
    .A1(net5928),
    .Y(_05785_),
    .A2(_05782_));
 sg13g2_nand2_1 _14803_ (.Y(_05786_),
    .A(net5389),
    .B(\mem.mem[96][7] ));
 sg13g2_a21oi_1 _14804_ (.A1(net6070),
    .A2(\mem.mem[97][7] ),
    .Y(_05787_),
    .B1(net5929));
 sg13g2_nor2b_1 _14805_ (.A(net6069),
    .B_N(\mem.mem[98][7] ),
    .Y(_05788_));
 sg13g2_a21oi_1 _14806_ (.A1(net6069),
    .A2(\mem.mem[99][7] ),
    .Y(_05789_),
    .B1(_05788_));
 sg13g2_a221oi_1 _14807_ (.B2(net5929),
    .C1(net5864),
    .B1(_05789_),
    .A1(_05786_),
    .Y(_05790_),
    .A2(_05787_));
 sg13g2_nor3_1 _14808_ (.A(net5833),
    .B(_05785_),
    .C(_05790_),
    .Y(_05791_));
 sg13g2_mux4_1 _14809_ (.S0(net6063),
    .A0(\mem.mem[104][7] ),
    .A1(\mem.mem[105][7] ),
    .A2(\mem.mem[106][7] ),
    .A3(\mem.mem[107][7] ),
    .S1(net5927),
    .X(_05792_));
 sg13g2_mux2_1 _14810_ (.A0(\mem.mem[108][7] ),
    .A1(\mem.mem[109][7] ),
    .S(net6067),
    .X(_05793_));
 sg13g2_a21o_1 _14811_ (.A2(\mem.mem[110][7] ),
    .A1(net5388),
    .B1(net5355),
    .X(_05794_));
 sg13g2_a21oi_1 _14812_ (.A1(net6065),
    .A2(\mem.mem[111][7] ),
    .Y(_05795_),
    .B1(_05794_));
 sg13g2_o21ai_1 _14813_ (.B1(net5861),
    .Y(_05796_),
    .A1(net5926),
    .A2(_05793_));
 sg13g2_o21ai_1 _14814_ (.B1(net5833),
    .Y(_05797_),
    .A1(_05795_),
    .A2(_05796_));
 sg13g2_a21oi_1 _14815_ (.A1(net5315),
    .A2(_05792_),
    .Y(_05798_),
    .B1(_05797_));
 sg13g2_o21ai_1 _14816_ (.B1(net5268),
    .Y(_05799_),
    .A1(_05791_),
    .A2(_05798_));
 sg13g2_nand2_1 _14817_ (.Y(_05800_),
    .A(net5380),
    .B(\mem.mem[116][7] ));
 sg13g2_a21oi_1 _14818_ (.A1(net6035),
    .A2(\mem.mem[117][7] ),
    .Y(_05801_),
    .B1(net5909));
 sg13g2_and2_1 _14819_ (.A(net6036),
    .B(\mem.mem[119][7] ),
    .X(_05802_));
 sg13g2_a21oi_1 _14820_ (.A1(net5380),
    .A2(\mem.mem[118][7] ),
    .Y(_05803_),
    .B1(_05802_));
 sg13g2_a221oi_1 _14821_ (.B2(net5909),
    .C1(net5306),
    .B1(_05803_),
    .A1(_05800_),
    .Y(_05804_),
    .A2(_05801_));
 sg13g2_nand2_1 _14822_ (.Y(_05805_),
    .A(net5385),
    .B(\mem.mem[112][7] ));
 sg13g2_a21oi_1 _14823_ (.A1(net6050),
    .A2(\mem.mem[113][7] ),
    .Y(_05806_),
    .B1(net5919));
 sg13g2_nor2b_1 _14824_ (.A(net6050),
    .B_N(\mem.mem[114][7] ),
    .Y(_05807_));
 sg13g2_a21oi_1 _14825_ (.A1(net6050),
    .A2(\mem.mem[115][7] ),
    .Y(_05808_),
    .B1(_05807_));
 sg13g2_a221oi_1 _14826_ (.B2(net5919),
    .C1(net5857),
    .B1(_05808_),
    .A1(_05805_),
    .Y(_05809_),
    .A2(_05806_));
 sg13g2_nor3_1 _14827_ (.A(net5830),
    .B(_05804_),
    .C(_05809_),
    .Y(_05810_));
 sg13g2_mux4_1 _14828_ (.S0(net6041),
    .A0(\mem.mem[120][7] ),
    .A1(\mem.mem[121][7] ),
    .A2(\mem.mem[122][7] ),
    .A3(\mem.mem[123][7] ),
    .S1(net5911),
    .X(_05811_));
 sg13g2_a21oi_1 _14829_ (.A1(net6041),
    .A2(\mem.mem[127][7] ),
    .Y(_05812_),
    .B1(net5351));
 sg13g2_o21ai_1 _14830_ (.B1(_05812_),
    .Y(_05813_),
    .A1(net6041),
    .A2(_02878_));
 sg13g2_nand2_1 _14831_ (.Y(_05814_),
    .A(net6041),
    .B(\mem.mem[125][7] ));
 sg13g2_a21oi_1 _14832_ (.A1(net5381),
    .A2(\mem.mem[124][7] ),
    .Y(_05815_),
    .B1(net5912));
 sg13g2_a21oi_1 _14833_ (.A1(_05814_),
    .A2(_05815_),
    .Y(_05816_),
    .B1(net5307));
 sg13g2_a221oi_1 _14834_ (.B2(_05816_),
    .C1(net5280),
    .B1(_05813_),
    .A1(net5307),
    .Y(_05817_),
    .A2(_05811_));
 sg13g2_o21ai_1 _14835_ (.B1(net5818),
    .Y(_05818_),
    .A1(_05810_),
    .A2(_05817_));
 sg13g2_nand3_1 _14836_ (.B(_05799_),
    .C(_05818_),
    .A(net5809),
    .Y(_05819_));
 sg13g2_nor2_2 _14837_ (.A(net5262),
    .B(_05780_),
    .Y(_05820_));
 sg13g2_a22oi_1 _14838_ (.Y(_05821_),
    .B1(_05819_),
    .B2(_05820_),
    .A2(_05744_),
    .A1(_05743_));
 sg13g2_or2_1 _14839_ (.X(_05822_),
    .B(_05821_),
    .A(_00007_));
 sg13g2_mux4_1 _14840_ (.S0(net6132),
    .A0(\mem.mem[176][7] ),
    .A1(\mem.mem[177][7] ),
    .A2(\mem.mem[178][7] ),
    .A3(\mem.mem[179][7] ),
    .S1(net5973),
    .X(_05823_));
 sg13g2_mux2_1 _14841_ (.A0(\mem.mem[180][7] ),
    .A1(\mem.mem[181][7] ),
    .S(net6130),
    .X(_05824_));
 sg13g2_nor2_1 _14842_ (.A(net5411),
    .B(\mem.mem[183][7] ),
    .Y(_05825_));
 sg13g2_o21ai_1 _14843_ (.B1(net5975),
    .Y(_05826_),
    .A1(net6134),
    .A2(\mem.mem[182][7] ));
 sg13g2_o21ai_1 _14844_ (.B1(net5875),
    .Y(_05827_),
    .A1(_05825_),
    .A2(_05826_));
 sg13g2_a21oi_1 _14845_ (.A1(net5366),
    .A2(_05824_),
    .Y(_05828_),
    .B1(_05827_));
 sg13g2_nor2_1 _14846_ (.A(net5845),
    .B(_05828_),
    .Y(_05829_));
 sg13g2_o21ai_1 _14847_ (.B1(_05829_),
    .Y(_05830_),
    .A1(net5875),
    .A2(_05823_));
 sg13g2_mux4_1 _14848_ (.S0(net6096),
    .A0(\mem.mem[184][7] ),
    .A1(\mem.mem[185][7] ),
    .A2(\mem.mem[186][7] ),
    .A3(\mem.mem[187][7] ),
    .S1(net5950),
    .X(_05831_));
 sg13g2_mux2_1 _14849_ (.A0(\mem.mem[188][7] ),
    .A1(\mem.mem[189][7] ),
    .S(net6103),
    .X(_05832_));
 sg13g2_nor2_1 _14850_ (.A(net5400),
    .B(\mem.mem[191][7] ),
    .Y(_05833_));
 sg13g2_o21ai_1 _14851_ (.B1(net5952),
    .Y(_05834_),
    .A1(net6101),
    .A2(\mem.mem[190][7] ));
 sg13g2_o21ai_1 _14852_ (.B1(net5868),
    .Y(_05835_),
    .A1(_05833_),
    .A2(_05834_));
 sg13g2_a21oi_1 _14853_ (.A1(net5358),
    .A2(_05832_),
    .Y(_05836_),
    .B1(_05835_));
 sg13g2_nor2_1 _14854_ (.A(net5289),
    .B(_05836_),
    .Y(_05837_));
 sg13g2_o21ai_1 _14855_ (.B1(_05837_),
    .Y(_05838_),
    .A1(net5867),
    .A2(_05831_));
 sg13g2_nand3_1 _14856_ (.B(_05830_),
    .C(_05838_),
    .A(net5823),
    .Y(_05839_));
 sg13g2_mux4_1 _14857_ (.S0(net6086),
    .A0(\mem.mem[168][7] ),
    .A1(\mem.mem[169][7] ),
    .A2(\mem.mem[170][7] ),
    .A3(\mem.mem[171][7] ),
    .S1(net5945),
    .X(_05840_));
 sg13g2_nor2_1 _14858_ (.A(net5865),
    .B(_05840_),
    .Y(_05841_));
 sg13g2_nor2_1 _14859_ (.A(net5397),
    .B(\mem.mem[173][7] ),
    .Y(_05842_));
 sg13g2_nor2_1 _14860_ (.A(net6091),
    .B(\mem.mem[172][7] ),
    .Y(_05843_));
 sg13g2_nor3_1 _14861_ (.A(net5946),
    .B(_05842_),
    .C(_05843_),
    .Y(_05844_));
 sg13g2_nor2_1 _14862_ (.A(net5397),
    .B(\mem.mem[175][7] ),
    .Y(_05845_));
 sg13g2_o21ai_1 _14863_ (.B1(net5949),
    .Y(_05846_),
    .A1(net6091),
    .A2(\mem.mem[174][7] ));
 sg13g2_o21ai_1 _14864_ (.B1(net5866),
    .Y(_05847_),
    .A1(_05845_),
    .A2(_05846_));
 sg13g2_o21ai_1 _14865_ (.B1(net5838),
    .Y(_05848_),
    .A1(_05844_),
    .A2(_05847_));
 sg13g2_a21oi_1 _14866_ (.A1(net5387),
    .A2(_02879_),
    .Y(_05849_),
    .B1(net5353));
 sg13g2_o21ai_1 _14867_ (.B1(_05849_),
    .Y(_05850_),
    .A1(net5387),
    .A2(\mem.mem[167][7] ));
 sg13g2_mux2_1 _14868_ (.A0(\mem.mem[164][7] ),
    .A1(\mem.mem[165][7] ),
    .S(net6055),
    .X(_05851_));
 sg13g2_a21oi_1 _14869_ (.A1(net5353),
    .A2(_05851_),
    .Y(_05852_),
    .B1(net5312));
 sg13g2_mux2_1 _14870_ (.A0(\mem.mem[162][7] ),
    .A1(\mem.mem[163][7] ),
    .S(net6056),
    .X(_05853_));
 sg13g2_nand2_1 _14871_ (.Y(_05854_),
    .A(net5924),
    .B(_05853_));
 sg13g2_mux2_1 _14872_ (.A0(\mem.mem[160][7] ),
    .A1(\mem.mem[161][7] ),
    .S(net6055),
    .X(_05855_));
 sg13g2_a21oi_1 _14873_ (.A1(net5353),
    .A2(_05855_),
    .Y(_05856_),
    .B1(net5859));
 sg13g2_a221oi_1 _14874_ (.B2(_05856_),
    .C1(net5832),
    .B1(_05854_),
    .A1(_05850_),
    .Y(_05857_),
    .A2(_05852_));
 sg13g2_nor2_2 _14875_ (.A(net5820),
    .B(_05857_),
    .Y(_05858_));
 sg13g2_o21ai_1 _14876_ (.B1(_05858_),
    .Y(_05859_),
    .A1(_05841_),
    .A2(_05848_));
 sg13g2_nand3_1 _14877_ (.B(_05839_),
    .C(_05859_),
    .A(net5812),
    .Y(_05860_));
 sg13g2_mux4_1 _14878_ (.S0(net6114),
    .A0(\mem.mem[136][7] ),
    .A1(\mem.mem[137][7] ),
    .A2(\mem.mem[138][7] ),
    .A3(\mem.mem[139][7] ),
    .S1(net5959),
    .X(_05861_));
 sg13g2_nor2_1 _14879_ (.A(net5869),
    .B(_05861_),
    .Y(_05862_));
 sg13g2_nor2_1 _14880_ (.A(net5404),
    .B(\mem.mem[141][7] ),
    .Y(_05863_));
 sg13g2_nor2_1 _14881_ (.A(net6114),
    .B(\mem.mem[140][7] ),
    .Y(_05864_));
 sg13g2_nor3_1 _14882_ (.A(net5959),
    .B(_05863_),
    .C(_05864_),
    .Y(_05865_));
 sg13g2_nor2_1 _14883_ (.A(net5404),
    .B(\mem.mem[143][7] ),
    .Y(_05866_));
 sg13g2_o21ai_1 _14884_ (.B1(net5959),
    .Y(_05867_),
    .A1(net6114),
    .A2(\mem.mem[142][7] ));
 sg13g2_o21ai_1 _14885_ (.B1(net5870),
    .Y(_05868_),
    .A1(_05866_),
    .A2(_05867_));
 sg13g2_o21ai_1 _14886_ (.B1(net5841),
    .Y(_05869_),
    .A1(_05865_),
    .A2(_05868_));
 sg13g2_mux4_1 _14887_ (.S0(net6117),
    .A0(\mem.mem[128][7] ),
    .A1(\mem.mem[129][7] ),
    .A2(\mem.mem[130][7] ),
    .A3(\mem.mem[131][7] ),
    .S1(net5963),
    .X(_05870_));
 sg13g2_mux2_1 _14888_ (.A0(\mem.mem[132][7] ),
    .A1(\mem.mem[133][7] ),
    .S(net6119),
    .X(_05871_));
 sg13g2_nand2_1 _14889_ (.Y(_05872_),
    .A(net5362),
    .B(_05871_));
 sg13g2_mux2_1 _14890_ (.A0(\mem.mem[134][7] ),
    .A1(\mem.mem[135][7] ),
    .S(net6118),
    .X(_05873_));
 sg13g2_a21oi_1 _14891_ (.A1(net5964),
    .A2(_05873_),
    .Y(_05874_),
    .B1(net5332));
 sg13g2_a21oi_1 _14892_ (.A1(_05872_),
    .A2(_05874_),
    .Y(_05875_),
    .B1(net5840));
 sg13g2_o21ai_1 _14893_ (.B1(_05875_),
    .Y(_05876_),
    .A1(net5872),
    .A2(_05870_));
 sg13g2_o21ai_1 _14894_ (.B1(_05876_),
    .Y(_05877_),
    .A1(_05862_),
    .A2(_05869_));
 sg13g2_mux4_1 _14895_ (.S0(net6077),
    .A0(\mem.mem[144][7] ),
    .A1(\mem.mem[145][7] ),
    .A2(\mem.mem[146][7] ),
    .A3(\mem.mem[147][7] ),
    .S1(net5933),
    .X(_05878_));
 sg13g2_nor2_1 _14896_ (.A(net5869),
    .B(_05878_),
    .Y(_05879_));
 sg13g2_mux2_1 _14897_ (.A0(\mem.mem[148][7] ),
    .A1(\mem.mem[149][7] ),
    .S(net6106),
    .X(_05880_));
 sg13g2_nor2_1 _14898_ (.A(net5402),
    .B(\mem.mem[151][7] ),
    .Y(_05881_));
 sg13g2_o21ai_1 _14899_ (.B1(net5955),
    .Y(_05882_),
    .A1(net6105),
    .A2(\mem.mem[150][7] ));
 sg13g2_o21ai_1 _14900_ (.B1(net5869),
    .Y(_05883_),
    .A1(_05881_),
    .A2(_05882_));
 sg13g2_a21oi_1 _14901_ (.A1(net5361),
    .A2(_05880_),
    .Y(_05884_),
    .B1(_05883_));
 sg13g2_nor3_1 _14902_ (.A(net5841),
    .B(_05879_),
    .C(_05884_),
    .Y(_05885_));
 sg13g2_mux2_1 _14903_ (.A0(\mem.mem[156][7] ),
    .A1(\mem.mem[157][7] ),
    .S(net6107),
    .X(_05886_));
 sg13g2_mux2_1 _14904_ (.A0(\mem.mem[158][7] ),
    .A1(\mem.mem[159][7] ),
    .S(net6092),
    .X(_05887_));
 sg13g2_nand2_1 _14905_ (.Y(_05888_),
    .A(net5948),
    .B(_05887_));
 sg13g2_a21oi_2 _14906_ (.B1(net5329),
    .Y(_05889_),
    .A2(_05886_),
    .A1(net5361));
 sg13g2_mux2_1 _14907_ (.A0(\mem.mem[154][7] ),
    .A1(\mem.mem[155][7] ),
    .S(net6100),
    .X(_05890_));
 sg13g2_nand2_1 _14908_ (.Y(_05891_),
    .A(net5947),
    .B(_05890_));
 sg13g2_mux2_1 _14909_ (.A0(\mem.mem[152][7] ),
    .A1(\mem.mem[153][7] ),
    .S(net6092),
    .X(_05892_));
 sg13g2_a21oi_1 _14910_ (.A1(net5360),
    .A2(_05892_),
    .Y(_05893_),
    .B1(net5866));
 sg13g2_a221oi_1 _14911_ (.B2(_05893_),
    .C1(net5287),
    .B1(_05891_),
    .A1(_05888_),
    .Y(_05894_),
    .A2(_05889_));
 sg13g2_nor3_1 _14912_ (.A(net5271),
    .B(_05885_),
    .C(_05894_),
    .Y(_05895_));
 sg13g2_nor2_1 _14913_ (.A(net5814),
    .B(_05895_),
    .Y(_05896_));
 sg13g2_o21ai_1 _14914_ (.B1(_05896_),
    .Y(_05897_),
    .A1(net5822),
    .A2(_05877_));
 sg13g2_nand3_1 _14915_ (.B(_05860_),
    .C(_05897_),
    .A(net5262),
    .Y(_05898_));
 sg13g2_mux4_1 _14916_ (.S0(net6095),
    .A0(\mem.mem[192][7] ),
    .A1(\mem.mem[193][7] ),
    .A2(\mem.mem[194][7] ),
    .A3(\mem.mem[195][7] ),
    .S1(net5951),
    .X(_05899_));
 sg13g2_nand2_1 _14917_ (.Y(_05900_),
    .A(net5401),
    .B(\mem.mem[198][7] ));
 sg13g2_a21oi_1 _14918_ (.A1(net6096),
    .A2(\mem.mem[199][7] ),
    .Y(_05901_),
    .B1(net5359));
 sg13g2_nand2b_1 _14919_ (.Y(_05902_),
    .B(net6096),
    .A_N(\mem.mem[197][7] ));
 sg13g2_o21ai_1 _14920_ (.B1(_05902_),
    .Y(_05903_),
    .A1(net6096),
    .A2(\mem.mem[196][7] ));
 sg13g2_a221oi_1 _14921_ (.B2(net5359),
    .C1(net5326),
    .B1(_05903_),
    .A1(_05900_),
    .Y(_05904_),
    .A2(_05901_));
 sg13g2_a21oi_1 _14922_ (.A1(net5326),
    .A2(_05899_),
    .Y(_05905_),
    .B1(_05904_));
 sg13g2_mux4_1 _14923_ (.S0(net6087),
    .A0(\mem.mem[200][7] ),
    .A1(\mem.mem[201][7] ),
    .A2(\mem.mem[202][7] ),
    .A3(\mem.mem[203][7] ),
    .S1(net5944),
    .X(_05906_));
 sg13g2_nand2_1 _14924_ (.Y(_05907_),
    .A(net5324),
    .B(_05906_));
 sg13g2_mux4_1 _14925_ (.S0(net6095),
    .A0(\mem.mem[204][7] ),
    .A1(\mem.mem[205][7] ),
    .A2(\mem.mem[206][7] ),
    .A3(\mem.mem[207][7] ),
    .S1(net5951),
    .X(_05908_));
 sg13g2_a21oi_1 _14926_ (.A1(net5867),
    .A2(_05908_),
    .Y(_05909_),
    .B1(net5288));
 sg13g2_a22oi_1 _14927_ (.Y(_05910_),
    .B1(_05907_),
    .B2(_05909_),
    .A2(_05905_),
    .A1(net5288));
 sg13g2_mux4_1 _14928_ (.S0(net6136),
    .A0(\mem.mem[216][7] ),
    .A1(\mem.mem[217][7] ),
    .A2(\mem.mem[218][7] ),
    .A3(\mem.mem[219][7] ),
    .S1(net5976),
    .X(_05911_));
 sg13g2_nand2_1 _14929_ (.Y(_05912_),
    .A(net5335),
    .B(_05911_));
 sg13g2_mux4_1 _14930_ (.S0(net6161),
    .A0(\mem.mem[220][7] ),
    .A1(\mem.mem[221][7] ),
    .A2(\mem.mem[222][7] ),
    .A3(\mem.mem[223][7] ),
    .S1(net5995),
    .X(_05913_));
 sg13g2_a21oi_1 _14931_ (.A1(net5879),
    .A2(_05913_),
    .Y(_05914_),
    .B1(net5294));
 sg13g2_mux4_1 _14932_ (.S0(net6161),
    .A0(\mem.mem[208][7] ),
    .A1(\mem.mem[209][7] ),
    .A2(\mem.mem[210][7] ),
    .A3(\mem.mem[211][7] ),
    .S1(net5995),
    .X(_05915_));
 sg13g2_nand2_1 _14933_ (.Y(_05916_),
    .A(net5338),
    .B(_05915_));
 sg13g2_mux4_1 _14934_ (.S0(net6147),
    .A0(\mem.mem[212][7] ),
    .A1(\mem.mem[213][7] ),
    .A2(\mem.mem[214][7] ),
    .A3(\mem.mem[215][7] ),
    .S1(net5984),
    .X(_05917_));
 sg13g2_a21oi_1 _14935_ (.A1(net5879),
    .A2(_05917_),
    .Y(_05918_),
    .B1(net5844));
 sg13g2_a22oi_1 _14936_ (.Y(_05919_),
    .B1(_05916_),
    .B2(_05918_),
    .A2(_05914_),
    .A1(_05912_));
 sg13g2_mux4_1 _14937_ (.S0(net6138),
    .A0(\mem.mem[224][7] ),
    .A1(\mem.mem[225][7] ),
    .A2(\mem.mem[226][7] ),
    .A3(\mem.mem[227][7] ),
    .S1(net5978),
    .X(_05920_));
 sg13g2_mux4_1 _14938_ (.S0(net6138),
    .A0(\mem.mem[228][7] ),
    .A1(\mem.mem[229][7] ),
    .A2(\mem.mem[230][7] ),
    .A3(\mem.mem[231][7] ),
    .S1(net5978),
    .X(_05921_));
 sg13g2_nand2_1 _14939_ (.Y(_05922_),
    .A(net5878),
    .B(_05921_));
 sg13g2_a21oi_1 _14940_ (.A1(net5339),
    .A2(_05920_),
    .Y(_05923_),
    .B1(net5843));
 sg13g2_nor2b_1 _14941_ (.A(net6141),
    .B_N(\mem.mem[234][7] ),
    .Y(_05924_));
 sg13g2_a21oi_1 _14942_ (.A1(net6141),
    .A2(\mem.mem[235][7] ),
    .Y(_05925_),
    .B1(_05924_));
 sg13g2_nand2_1 _14943_ (.Y(_05926_),
    .A(net6141),
    .B(\mem.mem[233][7] ));
 sg13g2_nand2_1 _14944_ (.Y(_05927_),
    .A(net5414),
    .B(\mem.mem[232][7] ));
 sg13g2_nand3_1 _14945_ (.B(_05926_),
    .C(_05927_),
    .A(net5365),
    .Y(_05928_));
 sg13g2_a21oi_1 _14946_ (.A1(net5979),
    .A2(_05925_),
    .Y(_05929_),
    .B1(net5878));
 sg13g2_mux2_1 _14947_ (.A0(\mem.mem[236][7] ),
    .A1(\mem.mem[237][7] ),
    .S(net6145),
    .X(_05930_));
 sg13g2_and2_1 _14948_ (.A(net6145),
    .B(\mem.mem[239][7] ),
    .X(_05931_));
 sg13g2_a21oi_1 _14949_ (.A1(net5412),
    .A2(\mem.mem[238][7] ),
    .Y(_05932_),
    .B1(_05931_));
 sg13g2_a21oi_1 _14950_ (.A1(net5983),
    .A2(_05932_),
    .Y(_05933_),
    .B1(net5337));
 sg13g2_o21ai_1 _14951_ (.B1(_05933_),
    .Y(_05934_),
    .A1(net5983),
    .A2(_05930_));
 sg13g2_a21oi_1 _14952_ (.A1(_05928_),
    .A2(_05929_),
    .Y(_05935_),
    .B1(net5293));
 sg13g2_a22oi_1 _14953_ (.Y(_05936_),
    .B1(_05934_),
    .B2(_05935_),
    .A2(_05923_),
    .A1(_05922_));
 sg13g2_mux4_1 _14954_ (.S0(net6048),
    .A0(\mem.mem[240][7] ),
    .A1(\mem.mem[241][7] ),
    .A2(\mem.mem[242][7] ),
    .A3(\mem.mem[243][7] ),
    .S1(net5915),
    .X(_05937_));
 sg13g2_mux4_1 _14955_ (.S0(net6053),
    .A0(\mem.mem[244][7] ),
    .A1(\mem.mem[245][7] ),
    .A2(\mem.mem[246][7] ),
    .A3(\mem.mem[247][7] ),
    .S1(net5918),
    .X(_05938_));
 sg13g2_mux4_1 _14956_ (.S0(net6048),
    .A0(\mem.mem[248][7] ),
    .A1(\mem.mem[249][7] ),
    .A2(\mem.mem[250][7] ),
    .A3(\mem.mem[251][7] ),
    .S1(net5915),
    .X(_05939_));
 sg13g2_mux4_1 _14957_ (.S0(net5281),
    .A0(\mem.mem[252][7] ),
    .A1(_05938_),
    .A2(_05939_),
    .A3(_05937_),
    .S1(net5310),
    .X(_05940_));
 sg13g2_mux4_1 _14958_ (.S0(net5822),
    .A0(_05910_),
    .A1(_05919_),
    .A2(_05936_),
    .A3(_05940_),
    .S1(net5813),
    .X(_05941_));
 sg13g2_o21ai_1 _14959_ (.B1(_05898_),
    .Y(_05942_),
    .A1(net5262),
    .A2(_05941_));
 sg13g2_a21oi_2 _14960_ (.B1(_02944_),
    .Y(_05943_),
    .A2(_05942_),
    .A1(_00007_));
 sg13g2_a22oi_1 _14961_ (.Y(_05944_),
    .B1(_05822_),
    .B2(_05943_),
    .A2(_03639_),
    .A1(net9));
 sg13g2_o21ai_1 _14962_ (.B1(net6190),
    .Y(_05945_),
    .A1(net4200),
    .A2(net5789));
 sg13g2_a21oi_1 _14963_ (.A1(net5788),
    .A2(_05944_),
    .Y(_00555_),
    .B1(net4201));
 sg13g2_o21ai_1 _14964_ (.B1(net6185),
    .Y(_05946_),
    .A1(net5794),
    .A2(net4193));
 sg13g2_a21oi_1 _14965_ (.A1(net5794),
    .A2(_03944_),
    .Y(_00556_),
    .B1(_05946_));
 sg13g2_o21ai_1 _14966_ (.B1(net6183),
    .Y(_05947_),
    .A1(net5794),
    .A2(net4206));
 sg13g2_a21oi_1 _14967_ (.A1(net5794),
    .A2(_04215_),
    .Y(_00557_),
    .B1(_05947_));
 sg13g2_o21ai_1 _14968_ (.B1(net6185),
    .Y(_05948_),
    .A1(net5796),
    .A2(net4202));
 sg13g2_a21oi_1 _14969_ (.A1(net5794),
    .A2(_04561_),
    .Y(_00558_),
    .B1(net4203));
 sg13g2_o21ai_1 _14970_ (.B1(net6186),
    .Y(_05949_),
    .A1(net5794),
    .A2(net4194));
 sg13g2_a21oi_1 _14971_ (.A1(net5794),
    .A2(_04863_),
    .Y(_00559_),
    .B1(_05949_));
 sg13g2_o21ai_1 _14972_ (.B1(net6187),
    .Y(_05950_),
    .A1(net5795),
    .A2(net4199));
 sg13g2_a21oi_1 _14973_ (.A1(net5795),
    .A2(_05141_),
    .Y(_00560_),
    .B1(_05950_));
 sg13g2_o21ai_1 _14974_ (.B1(net6187),
    .Y(_05951_),
    .A1(net5795),
    .A2(net4192));
 sg13g2_a21oi_1 _14975_ (.A1(net5795),
    .A2(_05412_),
    .Y(_00561_),
    .B1(_05951_));
 sg13g2_o21ai_1 _14976_ (.B1(net6187),
    .Y(_05952_),
    .A1(net5796),
    .A2(net4189));
 sg13g2_a21oi_1 _14977_ (.A1(net5796),
    .A2(_05665_),
    .Y(_00562_),
    .B1(net4190));
 sg13g2_o21ai_1 _14978_ (.B1(net6188),
    .Y(_05953_),
    .A1(net4204),
    .A2(net5795));
 sg13g2_a21oi_1 _14979_ (.A1(net5795),
    .A2(_05944_),
    .Y(_00563_),
    .B1(_05953_));
 sg13g2_o21ai_1 _14980_ (.B1(net6183),
    .Y(_05954_),
    .A1(net5786),
    .A2(net4185));
 sg13g2_a21oi_1 _14981_ (.A1(net5786),
    .A2(_03944_),
    .Y(_00564_),
    .B1(_05954_));
 sg13g2_o21ai_1 _14982_ (.B1(net6183),
    .Y(_05955_),
    .A1(net5786),
    .A2(net4171));
 sg13g2_a21oi_1 _14983_ (.A1(net5786),
    .A2(_04215_),
    .Y(_00565_),
    .B1(_05955_));
 sg13g2_o21ai_1 _14984_ (.B1(net6183),
    .Y(_05956_),
    .A1(net5786),
    .A2(net4169));
 sg13g2_a21oi_1 _14985_ (.A1(net5786),
    .A2(_04561_),
    .Y(_00566_),
    .B1(_05956_));
 sg13g2_o21ai_1 _14986_ (.B1(net6184),
    .Y(_05957_),
    .A1(net5785),
    .A2(net3902));
 sg13g2_a21oi_1 _14987_ (.A1(net5785),
    .A2(_04863_),
    .Y(_00567_),
    .B1(_05957_));
 sg13g2_o21ai_1 _14988_ (.B1(net6188),
    .Y(_05958_),
    .A1(net5785),
    .A2(net4174));
 sg13g2_a21oi_1 _14989_ (.A1(net5785),
    .A2(_05141_),
    .Y(_00568_),
    .B1(_05958_));
 sg13g2_o21ai_1 _14990_ (.B1(net6188),
    .Y(_05959_),
    .A1(net5785),
    .A2(net3919));
 sg13g2_a21oi_1 _14991_ (.A1(\state[6] ),
    .A2(_05412_),
    .Y(_00569_),
    .B1(_05959_));
 sg13g2_o21ai_1 _14992_ (.B1(net6188),
    .Y(_05960_),
    .A1(net5785),
    .A2(net4177));
 sg13g2_a21oi_1 _14993_ (.A1(net5785),
    .A2(_05665_),
    .Y(_00570_),
    .B1(_05960_));
 sg13g2_o21ai_1 _14994_ (.B1(net6188),
    .Y(_05961_),
    .A1(net4175),
    .A2(net5785));
 sg13g2_a21oi_1 _14995_ (.A1(\state[6] ),
    .A2(_05944_),
    .Y(_00571_),
    .B1(_05961_));
 sg13g2_nand2_1 _14996_ (.Y(_05962_),
    .A(_02880_),
    .B(net6179));
 sg13g2_o21ai_1 _14997_ (.B1(_05962_),
    .Y(_05963_),
    .A1(_00019_),
    .A2(net6179));
 sg13g2_nand2_1 _14998_ (.Y(_05964_),
    .A(_02881_),
    .B(_03293_));
 sg13g2_a22oi_1 _14999_ (.Y(_05965_),
    .B1(_03293_),
    .B2(_02881_),
    .A2(_02884_),
    .A1(_02882_));
 sg13g2_o21ai_1 _15000_ (.B1(_05964_),
    .Y(_05966_),
    .A1(net5792),
    .A2(halted));
 sg13g2_o21ai_1 _15001_ (.B1(net5233),
    .Y(_05967_),
    .A1(net5790),
    .A2(_05963_));
 sg13g2_a21oi_1 _15002_ (.A1(net5790),
    .A2(_02906_),
    .Y(_05968_),
    .B1(_05967_));
 sg13g2_o21ai_1 _15003_ (.B1(net6184),
    .Y(_05969_),
    .A1(net4223),
    .A2(net5233));
 sg13g2_nor2_1 _15004_ (.A(_05968_),
    .B(_05969_),
    .Y(_00572_));
 sg13g2_nand2_1 _15005_ (.Y(_05970_),
    .A(_02881_),
    .B(_02909_));
 sg13g2_a21oi_1 _15006_ (.A1(_02841_),
    .A2(net6179),
    .Y(_05971_),
    .B1(net5790));
 sg13g2_a221oi_1 _15007_ (.B2(_05971_),
    .C1(_05966_),
    .B1(_05970_),
    .A1(net5790),
    .Y(_05972_),
    .A2(_02911_));
 sg13g2_o21ai_1 _15008_ (.B1(net6184),
    .Y(_05973_),
    .A1(net4230),
    .A2(net5233));
 sg13g2_nor2_1 _15009_ (.A(_05972_),
    .B(_05973_),
    .Y(_00573_));
 sg13g2_nand3_1 _15010_ (.B(\PC[1] ),
    .C(\PC[0] ),
    .A(\PC[2] ),
    .Y(_05974_));
 sg13g2_xnor2_1 _15011_ (.Y(_05975_),
    .A(\PC[2] ),
    .B(_02908_));
 sg13g2_a21oi_1 _15012_ (.A1(_02843_),
    .A2(net6179),
    .Y(_05976_),
    .B1(net5790));
 sg13g2_o21ai_1 _15013_ (.B1(_05976_),
    .Y(_05977_),
    .A1(net6179),
    .A2(_05975_));
 sg13g2_and2_1 _15014_ (.A(net5233),
    .B(_05977_),
    .X(_05978_));
 sg13g2_o21ai_1 _15015_ (.B1(net6184),
    .Y(_05979_),
    .A1(net4240),
    .A2(net5233));
 sg13g2_a21oi_1 _15016_ (.A1(net4237),
    .A2(_05978_),
    .Y(_00574_),
    .B1(_05979_));
 sg13g2_nand4_1 _15017_ (.B(\PC[2] ),
    .C(\PC[1] ),
    .A(\PC[3] ),
    .Y(_05980_),
    .D(\PC[0] ));
 sg13g2_nand2b_1 _15018_ (.Y(_05981_),
    .B(_05974_),
    .A_N(\PC[3] ));
 sg13g2_a21oi_1 _15019_ (.A1(_05980_),
    .A2(_05981_),
    .Y(_05982_),
    .B1(net6179));
 sg13g2_nor2_1 _15020_ (.A(net5),
    .B(_02881_),
    .Y(_05983_));
 sg13g2_nor3_1 _15021_ (.A(net5790),
    .B(_05982_),
    .C(_05983_),
    .Y(_05984_));
 sg13g2_nor3_1 _15022_ (.A(_03311_),
    .B(_05966_),
    .C(_05984_),
    .Y(_05985_));
 sg13g2_o21ai_1 _15023_ (.B1(net6184),
    .Y(_05986_),
    .A1(net4231),
    .A2(net5233));
 sg13g2_nor2_1 _15024_ (.A(_05985_),
    .B(_05986_),
    .Y(_00575_));
 sg13g2_xnor2_1 _15025_ (.Y(_05987_),
    .A(\PC[4] ),
    .B(_05980_));
 sg13g2_a21oi_1 _15026_ (.A1(_02857_),
    .A2(net6179),
    .Y(_05988_),
    .B1(net5791));
 sg13g2_o21ai_1 _15027_ (.B1(_05988_),
    .Y(_05989_),
    .A1(net6179),
    .A2(_05987_));
 sg13g2_nand3_1 _15028_ (.B(net5233),
    .C(_05989_),
    .A(_03317_),
    .Y(_05990_));
 sg13g2_o21ai_1 _15029_ (.B1(_05990_),
    .Y(_05991_),
    .A1(net4232),
    .A2(net5233));
 sg13g2_nor2_1 _15030_ (.A(net6175),
    .B(net4233),
    .Y(_00576_));
 sg13g2_nor2_1 _15031_ (.A(_00018_),
    .B(_05980_),
    .Y(_05992_));
 sg13g2_xnor2_1 _15032_ (.Y(_05993_),
    .A(_02832_),
    .B(_05992_));
 sg13g2_a21oi_1 _15033_ (.A1(_02865_),
    .A2(net6180),
    .Y(_05994_),
    .B1(net5792));
 sg13g2_o21ai_1 _15034_ (.B1(_05994_),
    .Y(_05995_),
    .A1(net6180),
    .A2(_05993_));
 sg13g2_and2_1 _15035_ (.A(_05965_),
    .B(_05995_),
    .X(_05996_));
 sg13g2_a221oi_1 _15036_ (.B2(_03323_),
    .C1(net6176),
    .B1(_05996_),
    .A1(_02832_),
    .Y(_00577_),
    .A2(_05966_));
 sg13g2_nor2_1 _15037_ (.A(_02893_),
    .B(_05980_),
    .Y(_05997_));
 sg13g2_xnor2_1 _15038_ (.Y(_05998_),
    .A(\PC[6] ),
    .B(_05997_));
 sg13g2_nand2_1 _15039_ (.Y(_05999_),
    .A(_02881_),
    .B(_05998_));
 sg13g2_a21oi_1 _15040_ (.A1(_02868_),
    .A2(net6180),
    .Y(_06000_),
    .B1(net5792));
 sg13g2_a221oi_1 _15041_ (.B2(_06000_),
    .C1(_05966_),
    .B1(_05999_),
    .A1(net5792),
    .Y(_06001_),
    .A2(_02925_));
 sg13g2_o21ai_1 _15042_ (.B1(net6188),
    .Y(_06002_),
    .A1(net4221),
    .A2(_05965_));
 sg13g2_nor2_1 _15043_ (.A(_06001_),
    .B(_06002_),
    .Y(_00578_));
 sg13g2_nand2b_1 _15044_ (.Y(_06003_),
    .B(_05997_),
    .A_N(_00017_));
 sg13g2_a21oi_1 _15045_ (.A1(\PC[7] ),
    .A2(_06003_),
    .Y(_06004_),
    .B1(net6180));
 sg13g2_o21ai_1 _15046_ (.B1(_06004_),
    .Y(_06005_),
    .A1(net4234),
    .A2(_06003_));
 sg13g2_a21oi_1 _15047_ (.A1(_02875_),
    .A2(net6180),
    .Y(_06006_),
    .B1(net5792));
 sg13g2_a21oi_1 _15048_ (.A1(_06005_),
    .A2(_06006_),
    .Y(_06007_),
    .B1(_05966_));
 sg13g2_a221oi_1 _15049_ (.B2(_03339_),
    .C1(net6175),
    .B1(_06007_),
    .A1(_02831_),
    .Y(_00579_),
    .A2(_05966_));
 sg13g2_nor2_1 _15050_ (.A(_02964_),
    .B(net5138),
    .Y(_06008_));
 sg13g2_nor2_1 _15051_ (.A(net3939),
    .B(net4755),
    .Y(_06009_));
 sg13g2_a21oi_1 _15052_ (.A1(net5451),
    .A2(net4755),
    .Y(_00588_),
    .B1(_06009_));
 sg13g2_nor2_1 _15053_ (.A(net3417),
    .B(net4754),
    .Y(_06010_));
 sg13g2_a21oi_1 _15054_ (.A1(net5497),
    .A2(net4754),
    .Y(_00589_),
    .B1(_06010_));
 sg13g2_nor2_1 _15055_ (.A(net3732),
    .B(net4755),
    .Y(_06011_));
 sg13g2_a21oi_1 _15056_ (.A1(net5541),
    .A2(net4755),
    .Y(_00590_),
    .B1(_06011_));
 sg13g2_nor2_1 _15057_ (.A(net4031),
    .B(net4754),
    .Y(_06012_));
 sg13g2_a21oi_1 _15058_ (.A1(net5586),
    .A2(net4754),
    .Y(_00591_),
    .B1(_06012_));
 sg13g2_nor2_1 _15059_ (.A(net3775),
    .B(net4754),
    .Y(_06013_));
 sg13g2_a21oi_1 _15060_ (.A1(net5631),
    .A2(net4754),
    .Y(_00592_),
    .B1(_06013_));
 sg13g2_nor2_1 _15061_ (.A(net4026),
    .B(net4755),
    .Y(_06014_));
 sg13g2_a21oi_1 _15062_ (.A1(net5675),
    .A2(net4755),
    .Y(_00593_),
    .B1(_06014_));
 sg13g2_nor2_1 _15063_ (.A(net4134),
    .B(net4755),
    .Y(_06015_));
 sg13g2_a21oi_1 _15064_ (.A1(net5721),
    .A2(net4755),
    .Y(_00594_),
    .B1(_06015_));
 sg13g2_nor2_1 _15065_ (.A(net3869),
    .B(net4754),
    .Y(_06016_));
 sg13g2_a21oi_1 _15066_ (.A1(net5766),
    .A2(net4754),
    .Y(_00595_),
    .B1(_06016_));
 sg13g2_a21o_1 _15067_ (.A2(_02884_),
    .A1(net5261),
    .B1(_03293_),
    .X(_06017_));
 sg13g2_o21ai_1 _15068_ (.B1(_02828_),
    .Y(_06018_),
    .A1(_03640_),
    .A2(_03943_));
 sg13g2_a21oi_1 _15069_ (.A1(net4205),
    .A2(_03944_),
    .Y(_06019_),
    .B1(net5260));
 sg13g2_nand2_1 _15070_ (.Y(_06020_),
    .A(_06018_),
    .B(_06019_));
 sg13g2_a21oi_1 _15071_ (.A1(net5260),
    .A2(_02880_),
    .Y(_06021_),
    .B1(net5231));
 sg13g2_a22oi_1 _15072_ (.Y(_06022_),
    .B1(_06020_),
    .B2(_06021_),
    .A2(net5231),
    .A1(\mem.data_in[0] ));
 sg13g2_nor2_1 _15073_ (.A(net6175),
    .B(_06022_),
    .Y(_00596_));
 sg13g2_a21oi_1 _15074_ (.A1(_03946_),
    .A2(_04214_),
    .Y(_06023_),
    .B1(_00016_));
 sg13g2_nand3_1 _15075_ (.B(_03946_),
    .C(_04214_),
    .A(_00016_),
    .Y(_06024_));
 sg13g2_nor2b_1 _15076_ (.A(_06023_),
    .B_N(_06024_),
    .Y(_06025_));
 sg13g2_xnor2_1 _15077_ (.Y(_06026_),
    .A(_06018_),
    .B(_06025_));
 sg13g2_nand2_1 _15078_ (.Y(_06027_),
    .A(\state[5] ),
    .B(_06026_));
 sg13g2_a21oi_1 _15079_ (.A1(_02841_),
    .A2(net5260),
    .Y(_06028_),
    .B1(net5232));
 sg13g2_a22oi_1 _15080_ (.Y(_06029_),
    .B1(_06027_),
    .B2(_06028_),
    .A2(net5232),
    .A1(net4225));
 sg13g2_nor2_1 _15081_ (.A(net6175),
    .B(net4226),
    .Y(_00597_));
 sg13g2_nand2_1 _15082_ (.Y(_06030_),
    .A(net4218),
    .B(net5231));
 sg13g2_a21oi_2 _15083_ (.B1(_06023_),
    .Y(_06031_),
    .A2(_06024_),
    .A1(_06018_));
 sg13g2_nand2_1 _15084_ (.Y(_06032_),
    .A(\mem_A[2] ),
    .B(_04561_));
 sg13g2_xnor2_1 _15085_ (.Y(_06033_),
    .A(\mem_A[2] ),
    .B(_04561_));
 sg13g2_xor2_1 _15086_ (.B(_06033_),
    .A(_06031_),
    .X(_06034_));
 sg13g2_a21oi_1 _15087_ (.A1(net5260),
    .A2(_02843_),
    .Y(_06035_),
    .B1(net5231));
 sg13g2_o21ai_1 _15088_ (.B1(_06035_),
    .Y(_06036_),
    .A1(net5260),
    .A2(_06034_));
 sg13g2_a21oi_1 _15089_ (.A1(_06030_),
    .A2(_06036_),
    .Y(_00598_),
    .B1(net6175));
 sg13g2_nor2_1 _15090_ (.A(\mem_A[3] ),
    .B(_04863_),
    .Y(_06037_));
 sg13g2_nand2_1 _15091_ (.Y(_06038_),
    .A(\mem_A[3] ),
    .B(_04863_));
 sg13g2_xnor2_1 _15092_ (.Y(_06039_),
    .A(\mem_A[3] ),
    .B(_04863_));
 sg13g2_o21ai_1 _15093_ (.B1(_06032_),
    .Y(_06040_),
    .A1(_06031_),
    .A2(_06033_));
 sg13g2_a21oi_1 _15094_ (.A1(_06039_),
    .A2(_06040_),
    .Y(_06041_),
    .B1(net5260));
 sg13g2_o21ai_1 _15095_ (.B1(_06041_),
    .Y(_06042_),
    .A1(_06039_),
    .A2(_06040_));
 sg13g2_a21oi_1 _15096_ (.A1(net5260),
    .A2(_02852_),
    .Y(_06043_),
    .B1(net5231));
 sg13g2_a22oi_1 _15097_ (.Y(_06044_),
    .B1(_06042_),
    .B2(_06043_),
    .A2(net5231),
    .A1(net4238));
 sg13g2_nor2_1 _15098_ (.A(net6175),
    .B(_06044_),
    .Y(_00599_));
 sg13g2_nor3_1 _15099_ (.A(_06031_),
    .B(_06033_),
    .C(_06039_),
    .Y(_06045_));
 sg13g2_o21ai_1 _15100_ (.B1(_06038_),
    .Y(_06046_),
    .A1(_06032_),
    .A2(_06037_));
 sg13g2_or2_1 _15101_ (.X(_06047_),
    .B(_06046_),
    .A(_06045_));
 sg13g2_nand2_1 _15102_ (.Y(_06048_),
    .A(\mem_A[4] ),
    .B(_05141_));
 sg13g2_xnor2_1 _15103_ (.Y(_06049_),
    .A(\mem_A[4] ),
    .B(_05141_));
 sg13g2_nand2b_1 _15104_ (.Y(_06050_),
    .B(_06047_),
    .A_N(_06049_));
 sg13g2_xor2_1 _15105_ (.B(_06049_),
    .A(_06047_),
    .X(_06051_));
 sg13g2_nand2_1 _15106_ (.Y(_06052_),
    .A(\state[5] ),
    .B(_06051_));
 sg13g2_a21oi_1 _15107_ (.A1(net5260),
    .A2(_02857_),
    .Y(_06053_),
    .B1(net5231));
 sg13g2_a22oi_1 _15108_ (.Y(_06054_),
    .B1(_06052_),
    .B2(_06053_),
    .A2(net5231),
    .A1(net4228));
 sg13g2_nor2_1 _15109_ (.A(net6175),
    .B(net4229),
    .Y(_00600_));
 sg13g2_nor2_1 _15110_ (.A(\mem_A[5] ),
    .B(_05412_),
    .Y(_06055_));
 sg13g2_xnor2_1 _15111_ (.Y(_06056_),
    .A(\mem_A[5] ),
    .B(_05412_));
 sg13g2_nand2_1 _15112_ (.Y(_06057_),
    .A(_06048_),
    .B(_06050_));
 sg13g2_xnor2_1 _15113_ (.Y(_06058_),
    .A(_06056_),
    .B(_06057_));
 sg13g2_a21oi_1 _15114_ (.A1(net5261),
    .A2(_02865_),
    .Y(_06059_),
    .B1(net5232));
 sg13g2_o21ai_1 _15115_ (.B1(_06059_),
    .Y(_06060_),
    .A1(net5261),
    .A2(_06058_));
 sg13g2_nand2_1 _15116_ (.Y(_06061_),
    .A(net4165),
    .B(net5232));
 sg13g2_a21oi_1 _15117_ (.A1(_06060_),
    .A2(_06061_),
    .Y(_00601_),
    .B1(net6175));
 sg13g2_nor2_1 _15118_ (.A(_06049_),
    .B(_06056_),
    .Y(_06062_));
 sg13g2_nor2_1 _15119_ (.A(_06048_),
    .B(_06055_),
    .Y(_06063_));
 sg13g2_a221oi_1 _15120_ (.B2(_06062_),
    .C1(_06063_),
    .B1(_06047_),
    .A1(\mem_A[5] ),
    .Y(_06064_),
    .A2(_05412_));
 sg13g2_nand2_1 _15121_ (.Y(_06065_),
    .A(\mem_A[6] ),
    .B(_05665_));
 sg13g2_xnor2_1 _15122_ (.Y(_06066_),
    .A(\mem_A[6] ),
    .B(_05665_));
 sg13g2_xnor2_1 _15123_ (.Y(_06067_),
    .A(_06064_),
    .B(_06066_));
 sg13g2_nand2_1 _15124_ (.Y(_06068_),
    .A(\state[5] ),
    .B(_06067_));
 sg13g2_a21oi_1 _15125_ (.A1(net5261),
    .A2(_02868_),
    .Y(_06069_),
    .B1(net5232));
 sg13g2_a22oi_1 _15126_ (.Y(_06070_),
    .B1(_06068_),
    .B2(_06069_),
    .A2(net5232),
    .A1(net4211));
 sg13g2_nor2_1 _15127_ (.A(net6176),
    .B(net4212),
    .Y(_00602_));
 sg13g2_o21ai_1 _15128_ (.B1(_06065_),
    .Y(_06071_),
    .A1(_06064_),
    .A2(_06066_));
 sg13g2_xor2_1 _15129_ (.B(_05944_),
    .A(\mem_A[7] ),
    .X(_06072_));
 sg13g2_xnor2_1 _15130_ (.Y(_06073_),
    .A(_06071_),
    .B(_06072_));
 sg13g2_a21o_1 _15131_ (.A2(_02875_),
    .A1(net5261),
    .B1(_06017_),
    .X(_06074_));
 sg13g2_a21o_1 _15132_ (.A2(_06073_),
    .A1(net4239),
    .B1(_06074_),
    .X(_06075_));
 sg13g2_nand2_1 _15133_ (.Y(_06076_),
    .A(net4251),
    .B(net5232));
 sg13g2_a21oi_1 _15134_ (.A1(_06075_),
    .A2(_06076_),
    .Y(_00603_),
    .B1(net6176));
 sg13g2_o21ai_1 _15135_ (.B1(net6183),
    .Y(_06077_),
    .A1(net5798),
    .A2(net4205));
 sg13g2_a21oi_1 _15136_ (.A1(net5798),
    .A2(_03944_),
    .Y(_00604_),
    .B1(_06077_));
 sg13g2_o21ai_1 _15137_ (.B1(net6183),
    .Y(_06078_),
    .A1(net5798),
    .A2(net4152));
 sg13g2_a21oi_1 _15138_ (.A1(net5798),
    .A2(_04215_),
    .Y(_00605_),
    .B1(_06078_));
 sg13g2_o21ai_1 _15139_ (.B1(net6182),
    .Y(_06079_),
    .A1(net5798),
    .A2(net4207));
 sg13g2_a21oi_1 _15140_ (.A1(net5798),
    .A2(_04561_),
    .Y(_00606_),
    .B1(_06079_));
 sg13g2_o21ai_1 _15141_ (.B1(net6182),
    .Y(_06080_),
    .A1(net5798),
    .A2(net4215));
 sg13g2_a21oi_1 _15142_ (.A1(net5798),
    .A2(_04863_),
    .Y(_00607_),
    .B1(_06080_));
 sg13g2_o21ai_1 _15143_ (.B1(net6182),
    .Y(_06081_),
    .A1(net5797),
    .A2(net4208));
 sg13g2_a21oi_1 _15144_ (.A1(net5797),
    .A2(_05141_),
    .Y(_00608_),
    .B1(_06081_));
 sg13g2_o21ai_1 _15145_ (.B1(net6189),
    .Y(_06082_),
    .A1(net5800),
    .A2(net4213));
 sg13g2_a21oi_1 _15146_ (.A1(net5797),
    .A2(_05412_),
    .Y(_00609_),
    .B1(net4214));
 sg13g2_o21ai_1 _15147_ (.B1(net6182),
    .Y(_06083_),
    .A1(net5797),
    .A2(net4210));
 sg13g2_a21oi_1 _15148_ (.A1(net5797),
    .A2(_05665_),
    .Y(_00610_),
    .B1(_06083_));
 sg13g2_o21ai_1 _15149_ (.B1(net6182),
    .Y(_06084_),
    .A1(net4209),
    .A2(net5797));
 sg13g2_a21oi_1 _15150_ (.A1(net5797),
    .A2(_05944_),
    .Y(_00611_),
    .B1(_06084_));
 sg13g2_nor2_1 _15151_ (.A(net5155),
    .B(_03467_),
    .Y(_06085_));
 sg13g2_nor2_1 _15152_ (.A(net3081),
    .B(net4753),
    .Y(_06086_));
 sg13g2_a21oi_1 _15153_ (.A1(net5424),
    .A2(net4753),
    .Y(_00612_),
    .B1(_06086_));
 sg13g2_nor2_1 _15154_ (.A(net4045),
    .B(net4752),
    .Y(_06087_));
 sg13g2_a21oi_1 _15155_ (.A1(net5468),
    .A2(net4752),
    .Y(_00613_),
    .B1(_06087_));
 sg13g2_nor2_1 _15156_ (.A(net3434),
    .B(net4753),
    .Y(_06088_));
 sg13g2_a21oi_1 _15157_ (.A1(net5515),
    .A2(net4753),
    .Y(_00614_),
    .B1(_06088_));
 sg13g2_nor2_1 _15158_ (.A(net4016),
    .B(net4753),
    .Y(_06089_));
 sg13g2_a21oi_1 _15159_ (.A1(net5558),
    .A2(net4753),
    .Y(_00615_),
    .B1(_06089_));
 sg13g2_nor2_1 _15160_ (.A(net4010),
    .B(net4752),
    .Y(_06090_));
 sg13g2_a21oi_1 _15161_ (.A1(net5605),
    .A2(net4752),
    .Y(_00616_),
    .B1(_06090_));
 sg13g2_nor2_1 _15162_ (.A(net3411),
    .B(net4752),
    .Y(_06091_));
 sg13g2_a21oi_1 _15163_ (.A1(net5650),
    .A2(net4752),
    .Y(_00617_),
    .B1(_06091_));
 sg13g2_nor2_1 _15164_ (.A(net3848),
    .B(net4752),
    .Y(_06092_));
 sg13g2_a21oi_1 _15165_ (.A1(net5696),
    .A2(net4752),
    .Y(_00618_),
    .B1(_06092_));
 sg13g2_nor2_1 _15166_ (.A(net3309),
    .B(net4753),
    .Y(_06093_));
 sg13g2_a21oi_1 _15167_ (.A1(net5745),
    .A2(net4753),
    .Y(_00619_),
    .B1(_06093_));
 sg13g2_nor2_1 _15168_ (.A(_02964_),
    .B(net5154),
    .Y(_06094_));
 sg13g2_nor2_1 _15169_ (.A(net3456),
    .B(net4750),
    .Y(_06095_));
 sg13g2_a21oi_1 _15170_ (.A1(net5428),
    .A2(net4750),
    .Y(_00620_),
    .B1(_06095_));
 sg13g2_nor2_1 _15171_ (.A(net3746),
    .B(net4751),
    .Y(_06096_));
 sg13g2_a21oi_1 _15172_ (.A1(net5475),
    .A2(net4751),
    .Y(_00621_),
    .B1(_06096_));
 sg13g2_nor2_1 _15173_ (.A(net4136),
    .B(net4751),
    .Y(_06097_));
 sg13g2_a21oi_1 _15174_ (.A1(net5518),
    .A2(net4751),
    .Y(_00622_),
    .B1(_06097_));
 sg13g2_nor2_1 _15175_ (.A(net3673),
    .B(net4751),
    .Y(_06098_));
 sg13g2_a21oi_1 _15176_ (.A1(net5565),
    .A2(net4751),
    .Y(_00623_),
    .B1(_06098_));
 sg13g2_nor2_1 _15177_ (.A(net3843),
    .B(net4751),
    .Y(_06099_));
 sg13g2_a21oi_1 _15178_ (.A1(net5610),
    .A2(net4751),
    .Y(_00624_),
    .B1(_06099_));
 sg13g2_nor2_1 _15179_ (.A(net3976),
    .B(net4750),
    .Y(_06100_));
 sg13g2_a21oi_1 _15180_ (.A1(net5655),
    .A2(net4750),
    .Y(_00625_),
    .B1(_06100_));
 sg13g2_nor2_1 _15181_ (.A(net4112),
    .B(net4750),
    .Y(_06101_));
 sg13g2_a21oi_1 _15182_ (.A1(net5700),
    .A2(net4750),
    .Y(_00626_),
    .B1(_06101_));
 sg13g2_nor2_1 _15183_ (.A(net3718),
    .B(net4750),
    .Y(_06102_));
 sg13g2_a21oi_1 _15184_ (.A1(net5745),
    .A2(net4750),
    .Y(_00627_),
    .B1(_06102_));
 sg13g2_nor2_1 _15185_ (.A(_03364_),
    .B(_03467_),
    .Y(_06103_));
 sg13g2_nor2_1 _15186_ (.A(net3533),
    .B(net5061),
    .Y(_06104_));
 sg13g2_a21oi_1 _15187_ (.A1(net5459),
    .A2(net5061),
    .Y(_00628_),
    .B1(_06104_));
 sg13g2_nor2_1 _15188_ (.A(net3726),
    .B(net5062),
    .Y(_06105_));
 sg13g2_a21oi_1 _15189_ (.A1(net5510),
    .A2(net5062),
    .Y(_00629_),
    .B1(_06105_));
 sg13g2_nor2_1 _15190_ (.A(net3741),
    .B(_06103_),
    .Y(_06106_));
 sg13g2_a21oi_1 _15191_ (.A1(net5551),
    .A2(net5062),
    .Y(_00630_),
    .B1(_06106_));
 sg13g2_nor2_1 _15192_ (.A(net4083),
    .B(net5062),
    .Y(_06107_));
 sg13g2_a21oi_1 _15193_ (.A1(net5595),
    .A2(net5062),
    .Y(_00631_),
    .B1(_06107_));
 sg13g2_nor2_1 _15194_ (.A(net3497),
    .B(net5062),
    .Y(_06108_));
 sg13g2_a21oi_1 _15195_ (.A1(net5641),
    .A2(net5062),
    .Y(_00632_),
    .B1(_06108_));
 sg13g2_nor2_1 _15196_ (.A(net3933),
    .B(net5061),
    .Y(_06109_));
 sg13g2_a21oi_1 _15197_ (.A1(net5686),
    .A2(net5061),
    .Y(_00633_),
    .B1(_06109_));
 sg13g2_nor2_1 _15198_ (.A(net3107),
    .B(net5061),
    .Y(_06110_));
 sg13g2_a21oi_1 _15199_ (.A1(net5730),
    .A2(net5061),
    .Y(_00634_),
    .B1(_06110_));
 sg13g2_nor2_1 _15200_ (.A(net3403),
    .B(net5061),
    .Y(_06111_));
 sg13g2_a21oi_1 _15201_ (.A1(net5778),
    .A2(net5061),
    .Y(_00635_),
    .B1(_06111_));
 sg13g2_nand2_1 _15202_ (.Y(_06112_),
    .A(_02963_),
    .B(_03363_));
 sg13g2_nand2_1 _15203_ (.Y(_06113_),
    .A(net3000),
    .B(net5059));
 sg13g2_o21ai_1 _15204_ (.B1(_06113_),
    .Y(_00636_),
    .A1(net5449),
    .A2(net5059));
 sg13g2_nand2_1 _15205_ (.Y(_06114_),
    .A(net2946),
    .B(net5059));
 sg13g2_o21ai_1 _15206_ (.B1(_06114_),
    .Y(_00637_),
    .A1(net5496),
    .A2(net5059));
 sg13g2_nand2_1 _15207_ (.Y(_06115_),
    .A(net2845),
    .B(net5059));
 sg13g2_o21ai_1 _15208_ (.B1(_06115_),
    .Y(_00638_),
    .A1(net5552),
    .A2(net5059));
 sg13g2_nand2_1 _15209_ (.Y(_06116_),
    .A(net2806),
    .B(net5060));
 sg13g2_o21ai_1 _15210_ (.B1(_06116_),
    .Y(_00639_),
    .A1(net5595),
    .A2(net5060));
 sg13g2_nand2_1 _15211_ (.Y(_06117_),
    .A(net2494),
    .B(net5060));
 sg13g2_o21ai_1 _15212_ (.B1(_06117_),
    .Y(_00640_),
    .A1(net5640),
    .A2(net5060));
 sg13g2_nand2_1 _15213_ (.Y(_06118_),
    .A(net3207),
    .B(net5060));
 sg13g2_o21ai_1 _15214_ (.B1(_06118_),
    .Y(_00641_),
    .A1(net5687),
    .A2(net5060));
 sg13g2_nand2_1 _15215_ (.Y(_06119_),
    .A(net2858),
    .B(net5060));
 sg13g2_o21ai_1 _15216_ (.B1(_06119_),
    .Y(_00642_),
    .A1(net5730),
    .A2(net5060));
 sg13g2_nand2_1 _15217_ (.Y(_06120_),
    .A(net3236),
    .B(net5059));
 sg13g2_o21ai_1 _15218_ (.B1(_06120_),
    .Y(_00643_),
    .A1(net5765),
    .A2(net5059));
 sg13g2_nor2_1 _15219_ (.A(_02981_),
    .B(net5210),
    .Y(_06121_));
 sg13g2_nor2_1 _15220_ (.A(net3897),
    .B(net5057),
    .Y(_06122_));
 sg13g2_a21oi_1 _15221_ (.A1(net5449),
    .A2(net5057),
    .Y(_00644_),
    .B1(_06122_));
 sg13g2_nor2_1 _15222_ (.A(net4110),
    .B(net5057),
    .Y(_06123_));
 sg13g2_a21oi_1 _15223_ (.A1(net5495),
    .A2(net5057),
    .Y(_00645_),
    .B1(_06123_));
 sg13g2_nor2_1 _15224_ (.A(net3913),
    .B(net5057),
    .Y(_06124_));
 sg13g2_a21oi_1 _15225_ (.A1(net5553),
    .A2(net5057),
    .Y(_00646_),
    .B1(_06124_));
 sg13g2_nor2_1 _15226_ (.A(net3387),
    .B(net5058),
    .Y(_06125_));
 sg13g2_a21oi_1 _15227_ (.A1(net5595),
    .A2(net5058),
    .Y(_00647_),
    .B1(_06125_));
 sg13g2_nor2_1 _15228_ (.A(net3223),
    .B(net5058),
    .Y(_06126_));
 sg13g2_a21oi_1 _15229_ (.A1(net5640),
    .A2(net5058),
    .Y(_00648_),
    .B1(_06126_));
 sg13g2_nor2_1 _15230_ (.A(net3783),
    .B(net5058),
    .Y(_06127_));
 sg13g2_a21oi_1 _15231_ (.A1(net5687),
    .A2(net5058),
    .Y(_00649_),
    .B1(_06127_));
 sg13g2_nor2_1 _15232_ (.A(net3833),
    .B(net5058),
    .Y(_06128_));
 sg13g2_a21oi_1 _15233_ (.A1(net5731),
    .A2(net5058),
    .Y(_00650_),
    .B1(_06128_));
 sg13g2_nor2_1 _15234_ (.A(net3683),
    .B(net5057),
    .Y(_06129_));
 sg13g2_a21oi_1 _15235_ (.A1(net5765),
    .A2(net5057),
    .Y(_00651_),
    .B1(_06129_));
 sg13g2_nor2_1 _15236_ (.A(_03017_),
    .B(net5210),
    .Y(_06130_));
 sg13g2_nor2_1 _15237_ (.A(net3839),
    .B(net5055),
    .Y(_06131_));
 sg13g2_a21oi_1 _15238_ (.A1(net5452),
    .A2(net5055),
    .Y(_00652_),
    .B1(_06131_));
 sg13g2_nor2_1 _15239_ (.A(net3489),
    .B(net5055),
    .Y(_06132_));
 sg13g2_a21oi_1 _15240_ (.A1(net5495),
    .A2(net5055),
    .Y(_00653_),
    .B1(_06132_));
 sg13g2_nor2_1 _15241_ (.A(net3955),
    .B(net5055),
    .Y(_06133_));
 sg13g2_a21oi_1 _15242_ (.A1(net5552),
    .A2(net5055),
    .Y(_00654_),
    .B1(_06133_));
 sg13g2_nor2_1 _15243_ (.A(net3666),
    .B(net5056),
    .Y(_06134_));
 sg13g2_a21oi_1 _15244_ (.A1(net5595),
    .A2(net5056),
    .Y(_00655_),
    .B1(_06134_));
 sg13g2_nor2_1 _15245_ (.A(net3842),
    .B(net5056),
    .Y(_06135_));
 sg13g2_a21oi_1 _15246_ (.A1(net5642),
    .A2(net5056),
    .Y(_00656_),
    .B1(_06135_));
 sg13g2_nor2_1 _15247_ (.A(net4120),
    .B(net5056),
    .Y(_06136_));
 sg13g2_a21oi_1 _15248_ (.A1(net5686),
    .A2(net5056),
    .Y(_00657_),
    .B1(_06136_));
 sg13g2_nor2_1 _15249_ (.A(net3896),
    .B(net5056),
    .Y(_06137_));
 sg13g2_a21oi_1 _15250_ (.A1(net5731),
    .A2(net5056),
    .Y(_00658_),
    .B1(_06137_));
 sg13g2_nor2_1 _15251_ (.A(net3799),
    .B(net5055),
    .Y(_06138_));
 sg13g2_a21oi_1 _15252_ (.A1(net5765),
    .A2(net5055),
    .Y(_00659_),
    .B1(_06138_));
 sg13g2_nor2_2 _15253_ (.A(_02941_),
    .B(_02947_),
    .Y(_06139_));
 sg13g2_nand2b_2 _15254_ (.Y(_06140_),
    .B(_02946_),
    .A_N(_02941_));
 sg13g2_nor2_1 _15255_ (.A(_03467_),
    .B(_06140_),
    .Y(_06141_));
 sg13g2_nor2_1 _15256_ (.A(net3675),
    .B(net5204),
    .Y(_06142_));
 sg13g2_a21oi_1 _15257_ (.A1(net5432),
    .A2(net5204),
    .Y(_00660_),
    .B1(_06142_));
 sg13g2_nor2_1 _15258_ (.A(net3988),
    .B(net5205),
    .Y(_06143_));
 sg13g2_a21oi_1 _15259_ (.A1(net5477),
    .A2(net5205),
    .Y(_00661_),
    .B1(_06143_));
 sg13g2_nor2_1 _15260_ (.A(net3806),
    .B(net5205),
    .Y(_06144_));
 sg13g2_a21oi_1 _15261_ (.A1(net5522),
    .A2(net5205),
    .Y(_00662_),
    .B1(_06144_));
 sg13g2_nor2_1 _15262_ (.A(net3432),
    .B(net5204),
    .Y(_06145_));
 sg13g2_a21oi_1 _15263_ (.A1(net5567),
    .A2(net5204),
    .Y(_00663_),
    .B1(_06145_));
 sg13g2_nor2_1 _15264_ (.A(net3545),
    .B(net5205),
    .Y(_06146_));
 sg13g2_a21oi_1 _15265_ (.A1(net5611),
    .A2(net5205),
    .Y(_00664_),
    .B1(_06146_));
 sg13g2_nor2_1 _15266_ (.A(net3699),
    .B(net5204),
    .Y(_06147_));
 sg13g2_a21oi_1 _15267_ (.A1(net5660),
    .A2(net5204),
    .Y(_00665_),
    .B1(_06147_));
 sg13g2_nor2_1 _15268_ (.A(net3408),
    .B(net5205),
    .Y(_06148_));
 sg13g2_a21oi_1 _15269_ (.A1(net5710),
    .A2(net5205),
    .Y(_00666_),
    .B1(_06148_));
 sg13g2_nor2_1 _15270_ (.A(net4048),
    .B(net5204),
    .Y(_06149_));
 sg13g2_a21oi_1 _15271_ (.A1(net5748),
    .A2(net5204),
    .Y(_00667_),
    .B1(_06149_));
 sg13g2_nand2_1 _15272_ (.Y(_06150_),
    .A(net5239),
    .B(_06139_));
 sg13g2_nand2_1 _15273_ (.Y(_06151_),
    .A(net2758),
    .B(net5054));
 sg13g2_o21ai_1 _15274_ (.B1(_06151_),
    .Y(_00668_),
    .A1(net5431),
    .A2(net5054));
 sg13g2_nand2_1 _15275_ (.Y(_06152_),
    .A(net2417),
    .B(net5054));
 sg13g2_o21ai_1 _15276_ (.B1(_06152_),
    .Y(_00669_),
    .A1(net5479),
    .A2(net5054));
 sg13g2_nand2_1 _15277_ (.Y(_06153_),
    .A(net2613),
    .B(net5054));
 sg13g2_o21ai_1 _15278_ (.B1(_06153_),
    .Y(_00670_),
    .A1(net5521),
    .A2(net5054));
 sg13g2_nand2_1 _15279_ (.Y(_06154_),
    .A(net3338),
    .B(net5053));
 sg13g2_o21ai_1 _15280_ (.B1(_06154_),
    .Y(_00671_),
    .A1(net5566),
    .A2(net5053));
 sg13g2_nand2_1 _15281_ (.Y(_06155_),
    .A(net2618),
    .B(net5053));
 sg13g2_o21ai_1 _15282_ (.B1(_06155_),
    .Y(_00672_),
    .A1(net5611),
    .A2(net5053));
 sg13g2_nand2_1 _15283_ (.Y(_06156_),
    .A(net3158),
    .B(net5053));
 sg13g2_o21ai_1 _15284_ (.B1(_06156_),
    .Y(_00673_),
    .A1(net5656),
    .A2(net5053));
 sg13g2_nand2_1 _15285_ (.Y(_06157_),
    .A(net2442),
    .B(net5054));
 sg13g2_o21ai_1 _15286_ (.B1(_06157_),
    .Y(_00674_),
    .A1(net5703),
    .A2(net5054));
 sg13g2_nand2_1 _15287_ (.Y(_06158_),
    .A(net3371),
    .B(net5053));
 sg13g2_o21ai_1 _15288_ (.B1(_06158_),
    .Y(_00675_),
    .A1(net5749),
    .A2(net5053));
 sg13g2_nor2_1 _15289_ (.A(_02940_),
    .B(net5228),
    .Y(_06159_));
 sg13g2_nor3_2 _15290_ (.A(_02940_),
    .B(net5228),
    .C(net5240),
    .Y(_06160_));
 sg13g2_nor2_1 _15291_ (.A(net3327),
    .B(net5201),
    .Y(_06161_));
 sg13g2_a21oi_1 _15292_ (.A1(net5458),
    .A2(net5201),
    .Y(_00676_),
    .B1(_06161_));
 sg13g2_nor2_1 _15293_ (.A(net4065),
    .B(net5201),
    .Y(_06162_));
 sg13g2_a21oi_1 _15294_ (.A1(net5505),
    .A2(net5201),
    .Y(_00677_),
    .B1(_06162_));
 sg13g2_nor2_1 _15295_ (.A(net3448),
    .B(net5201),
    .Y(_06163_));
 sg13g2_a21oi_1 _15296_ (.A1(net5549),
    .A2(net5201),
    .Y(_00678_),
    .B1(_06163_));
 sg13g2_nor2_1 _15297_ (.A(net4098),
    .B(net5200),
    .Y(_06164_));
 sg13g2_a21oi_1 _15298_ (.A1(net5592),
    .A2(net5200),
    .Y(_00679_),
    .B1(_06164_));
 sg13g2_nor2_1 _15299_ (.A(net4093),
    .B(net5200),
    .Y(_06165_));
 sg13g2_a21oi_1 _15300_ (.A1(net5638),
    .A2(net5200),
    .Y(_00680_),
    .B1(_06165_));
 sg13g2_nor2_1 _15301_ (.A(net3925),
    .B(net5200),
    .Y(_06166_));
 sg13g2_a21oi_1 _15302_ (.A1(net5683),
    .A2(net5200),
    .Y(_00681_),
    .B1(_06166_));
 sg13g2_nor2_1 _15303_ (.A(net3345),
    .B(net5200),
    .Y(_06167_));
 sg13g2_a21oi_1 _15304_ (.A1(net5728),
    .A2(net5200),
    .Y(_00682_),
    .B1(_06167_));
 sg13g2_nor2_1 _15305_ (.A(net3324),
    .B(net5201),
    .Y(_06168_));
 sg13g2_a21oi_1 _15306_ (.A1(net5776),
    .A2(net5201),
    .Y(_00683_),
    .B1(_06168_));
 sg13g2_nand2_1 _15307_ (.Y(_06169_),
    .A(_03200_),
    .B(net5203));
 sg13g2_nand2_1 _15308_ (.Y(_06170_),
    .A(net2305),
    .B(net5052));
 sg13g2_o21ai_1 _15309_ (.B1(_06170_),
    .Y(_00684_),
    .A1(net5457),
    .A2(net5052));
 sg13g2_nand2_1 _15310_ (.Y(_06171_),
    .A(net3097),
    .B(net5052));
 sg13g2_o21ai_1 _15311_ (.B1(_06171_),
    .Y(_00685_),
    .A1(net5504),
    .A2(net5052));
 sg13g2_nand2_1 _15312_ (.Y(_06172_),
    .A(net2574),
    .B(net5052));
 sg13g2_o21ai_1 _15313_ (.B1(_06172_),
    .Y(_00686_),
    .A1(net5548),
    .A2(net5052));
 sg13g2_nand2_1 _15314_ (.Y(_06173_),
    .A(net3246),
    .B(net5052));
 sg13g2_o21ai_1 _15315_ (.B1(_06173_),
    .Y(_00687_),
    .A1(net5593),
    .A2(net5052));
 sg13g2_nand2_1 _15316_ (.Y(_06174_),
    .A(net2308),
    .B(net5051));
 sg13g2_o21ai_1 _15317_ (.B1(_06174_),
    .Y(_00688_),
    .A1(net5636),
    .A2(net5051));
 sg13g2_nand2_1 _15318_ (.Y(_06175_),
    .A(net2405),
    .B(net5051));
 sg13g2_o21ai_1 _15319_ (.B1(_06175_),
    .Y(_00689_),
    .A1(net5682),
    .A2(net5051));
 sg13g2_nand2_1 _15320_ (.Y(_06176_),
    .A(net3139),
    .B(net5051));
 sg13g2_o21ai_1 _15321_ (.B1(_06176_),
    .Y(_00690_),
    .A1(net5726),
    .A2(net5051));
 sg13g2_nand2_1 _15322_ (.Y(_06177_),
    .A(net2294),
    .B(net5051));
 sg13g2_o21ai_1 _15323_ (.B1(_06177_),
    .Y(_00691_),
    .A1(net5773),
    .A2(net5051));
 sg13g2_nor2_1 _15324_ (.A(_02940_),
    .B(net5230),
    .Y(_06178_));
 sg13g2_nand2_1 _15325_ (.Y(_06179_),
    .A(_02963_),
    .B(net5199));
 sg13g2_nand2_1 _15326_ (.Y(_06180_),
    .A(net3028),
    .B(net5050));
 sg13g2_o21ai_1 _15327_ (.B1(_06180_),
    .Y(_00692_),
    .A1(net5459),
    .A2(net5050));
 sg13g2_nand2_1 _15328_ (.Y(_06181_),
    .A(net3074),
    .B(net5049));
 sg13g2_o21ai_1 _15329_ (.B1(_06181_),
    .Y(_00693_),
    .A1(net5503),
    .A2(net5049));
 sg13g2_nand2_1 _15330_ (.Y(_06182_),
    .A(net2549),
    .B(net5050));
 sg13g2_o21ai_1 _15331_ (.B1(_06182_),
    .Y(_00694_),
    .A1(net5545),
    .A2(net5050));
 sg13g2_nand2_1 _15332_ (.Y(_06183_),
    .A(net2795),
    .B(net5049));
 sg13g2_o21ai_1 _15333_ (.B1(_06183_),
    .Y(_00695_),
    .A1(net5589),
    .A2(net5049));
 sg13g2_nand2_1 _15334_ (.Y(_06184_),
    .A(net2400),
    .B(net5050));
 sg13g2_o21ai_1 _15335_ (.B1(_06184_),
    .Y(_00696_),
    .A1(net5643),
    .A2(net5050));
 sg13g2_nand2_1 _15336_ (.Y(_06185_),
    .A(net3372),
    .B(net5049));
 sg13g2_o21ai_1 _15337_ (.B1(_06185_),
    .Y(_00697_),
    .A1(net5684),
    .A2(net5049));
 sg13g2_nand2_1 _15338_ (.Y(_06186_),
    .A(net3279),
    .B(_06179_));
 sg13g2_o21ai_1 _15339_ (.B1(_06186_),
    .Y(_00698_),
    .A1(net5733),
    .A2(net5050));
 sg13g2_nand2_1 _15340_ (.Y(_06187_),
    .A(net3161),
    .B(net5049));
 sg13g2_o21ai_1 _15341_ (.B1(_06187_),
    .Y(_00699_),
    .A1(net5775),
    .A2(net5049));
 sg13g2_nand2_1 _15342_ (.Y(_06188_),
    .A(_03139_),
    .B(net5198));
 sg13g2_nand2_1 _15343_ (.Y(_06189_),
    .A(net2464),
    .B(net5047));
 sg13g2_o21ai_1 _15344_ (.B1(_06189_),
    .Y(_00700_),
    .A1(net5460),
    .A2(net5047));
 sg13g2_nand2_1 _15345_ (.Y(_06190_),
    .A(net2576),
    .B(net5048));
 sg13g2_o21ai_1 _15346_ (.B1(_06190_),
    .Y(_00701_),
    .A1(net5509),
    .A2(net5048));
 sg13g2_nand2_1 _15347_ (.Y(_06191_),
    .A(net2763),
    .B(net5048));
 sg13g2_o21ai_1 _15348_ (.B1(_06191_),
    .Y(_00702_),
    .A1(net5554),
    .A2(net5048));
 sg13g2_nand2_1 _15349_ (.Y(_06192_),
    .A(net2798),
    .B(net5048));
 sg13g2_o21ai_1 _15350_ (.B1(_06192_),
    .Y(_00703_),
    .A1(net5601),
    .A2(net5048));
 sg13g2_nand2_1 _15351_ (.Y(_06193_),
    .A(net3012),
    .B(net5048));
 sg13g2_o21ai_1 _15352_ (.B1(_06193_),
    .Y(_00704_),
    .A1(net5645),
    .A2(net5048));
 sg13g2_nand2_1 _15353_ (.Y(_06194_),
    .A(net2930),
    .B(net5047));
 sg13g2_o21ai_1 _15354_ (.B1(_06194_),
    .Y(_00705_),
    .A1(net5683),
    .A2(net5047));
 sg13g2_nand2_1 _15355_ (.Y(_06195_),
    .A(net2627),
    .B(net5047));
 sg13g2_o21ai_1 _15356_ (.B1(_06195_),
    .Y(_00706_),
    .A1(net5734),
    .A2(net5047));
 sg13g2_nand2_1 _15357_ (.Y(_06196_),
    .A(net2438),
    .B(net5047));
 sg13g2_o21ai_1 _15358_ (.B1(_06196_),
    .Y(_00707_),
    .A1(net5779),
    .A2(net5047));
 sg13g2_nand2b_2 _15359_ (.Y(_06197_),
    .B(net5220),
    .A_N(_02940_));
 sg13g2_nand4_1 _15360_ (.B(net5803),
    .C(net5220),
    .A(net5801),
    .Y(_06198_),
    .D(net5238));
 sg13g2_nand2_1 _15361_ (.Y(_06199_),
    .A(net3152),
    .B(net5044));
 sg13g2_o21ai_1 _15362_ (.B1(_06199_),
    .Y(_00708_),
    .A1(net5444),
    .A2(net5044));
 sg13g2_nand2_1 _15363_ (.Y(_06200_),
    .A(net2722),
    .B(net5044));
 sg13g2_o21ai_1 _15364_ (.B1(_06200_),
    .Y(_00709_),
    .A1(net5491),
    .A2(net5044));
 sg13g2_nand2_1 _15365_ (.Y(_06201_),
    .A(net2784),
    .B(net5044));
 sg13g2_o21ai_1 _15366_ (.B1(_06201_),
    .Y(_00710_),
    .A1(net5536),
    .A2(_06198_));
 sg13g2_nand2_1 _15367_ (.Y(_06202_),
    .A(net3147),
    .B(net5043));
 sg13g2_o21ai_1 _15368_ (.B1(_06202_),
    .Y(_00711_),
    .A1(net5579),
    .A2(net5043));
 sg13g2_nand2_1 _15369_ (.Y(_06203_),
    .A(net3267),
    .B(net5044));
 sg13g2_o21ai_1 _15370_ (.B1(_06203_),
    .Y(_00712_),
    .A1(net5633),
    .A2(net5043));
 sg13g2_nand2_1 _15371_ (.Y(_06204_),
    .A(net2922),
    .B(net5043));
 sg13g2_o21ai_1 _15372_ (.B1(_06204_),
    .Y(_00713_),
    .A1(net5678),
    .A2(net5043));
 sg13g2_nand2_1 _15373_ (.Y(_06205_),
    .A(net2559),
    .B(net5043));
 sg13g2_o21ai_1 _15374_ (.B1(_06205_),
    .Y(_00714_),
    .A1(net5723),
    .A2(net5044));
 sg13g2_nand2_1 _15375_ (.Y(_06206_),
    .A(net2371),
    .B(net5043));
 sg13g2_o21ai_1 _15376_ (.B1(_06206_),
    .Y(_00715_),
    .A1(net5770),
    .A2(net5043));
 sg13g2_nor2_2 _15377_ (.A(_03160_),
    .B(_03180_),
    .Y(_06207_));
 sg13g2_nand2_1 _15378_ (.Y(_06208_),
    .A(_03211_),
    .B(net5197));
 sg13g2_nand2_1 _15379_ (.Y(_06209_),
    .A(net3281),
    .B(net5042));
 sg13g2_o21ai_1 _15380_ (.B1(_06209_),
    .Y(_00716_),
    .A1(net5455),
    .A2(net5042));
 sg13g2_nand2_1 _15381_ (.Y(_06210_),
    .A(net3797),
    .B(net5042));
 sg13g2_o21ai_1 _15382_ (.B1(_06210_),
    .Y(_00717_),
    .A1(net5502),
    .A2(net5042));
 sg13g2_nand2_1 _15383_ (.Y(_06211_),
    .A(net3005),
    .B(net5041));
 sg13g2_o21ai_1 _15384_ (.B1(_06211_),
    .Y(_00718_),
    .A1(net5546),
    .A2(net5041));
 sg13g2_nand2_1 _15385_ (.Y(_06212_),
    .A(net3014),
    .B(net5042));
 sg13g2_o21ai_1 _15386_ (.B1(_06212_),
    .Y(_00719_),
    .A1(net5589),
    .A2(net5042));
 sg13g2_nand2_1 _15387_ (.Y(_06213_),
    .A(net2248),
    .B(net5042));
 sg13g2_o21ai_1 _15388_ (.B1(_06213_),
    .Y(_00720_),
    .A1(net5634),
    .A2(net5042));
 sg13g2_nand2_1 _15389_ (.Y(_06214_),
    .A(net2976),
    .B(net5041));
 sg13g2_o21ai_1 _15390_ (.B1(_06214_),
    .Y(_00721_),
    .A1(net5685),
    .A2(net5041));
 sg13g2_nand2_1 _15391_ (.Y(_06215_),
    .A(net3259),
    .B(net5041));
 sg13g2_o21ai_1 _15392_ (.B1(_06215_),
    .Y(_00722_),
    .A1(net5725),
    .A2(net5041));
 sg13g2_nand2_1 _15393_ (.Y(_06216_),
    .A(net2756),
    .B(net5041));
 sg13g2_o21ai_1 _15394_ (.B1(_06216_),
    .Y(_00723_),
    .A1(net5777),
    .A2(net5041));
 sg13g2_nand2_1 _15395_ (.Y(_06217_),
    .A(_03139_),
    .B(net5217));
 sg13g2_nand2_1 _15396_ (.Y(_06218_),
    .A(net2953),
    .B(net5039));
 sg13g2_o21ai_1 _15397_ (.B1(_06218_),
    .Y(_00724_),
    .A1(net5425),
    .A2(net5039));
 sg13g2_nand2_1 _15398_ (.Y(_06219_),
    .A(net2449),
    .B(net5039));
 sg13g2_o21ai_1 _15399_ (.B1(_06219_),
    .Y(_00725_),
    .A1(net5470),
    .A2(net5039));
 sg13g2_nand2_1 _15400_ (.Y(_06220_),
    .A(net3009),
    .B(net5040));
 sg13g2_o21ai_1 _15401_ (.B1(_06220_),
    .Y(_00726_),
    .A1(net5513),
    .A2(_06217_));
 sg13g2_nand2_1 _15402_ (.Y(_06221_),
    .A(net3098),
    .B(net5040));
 sg13g2_o21ai_1 _15403_ (.B1(_06221_),
    .Y(_00727_),
    .A1(net5558),
    .A2(net5040));
 sg13g2_nand2_1 _15404_ (.Y(_06222_),
    .A(net2997),
    .B(net5040));
 sg13g2_o21ai_1 _15405_ (.B1(_06222_),
    .Y(_00728_),
    .A1(net5606),
    .A2(net5040));
 sg13g2_nand2_1 _15406_ (.Y(_06223_),
    .A(net3530),
    .B(net5040));
 sg13g2_o21ai_1 _15407_ (.B1(_06223_),
    .Y(_00729_),
    .A1(net5649),
    .A2(net5040));
 sg13g2_nand2_1 _15408_ (.Y(_06224_),
    .A(net2590),
    .B(net5039));
 sg13g2_o21ai_1 _15409_ (.B1(_06224_),
    .Y(_00730_),
    .A1(net5697),
    .A2(net5039));
 sg13g2_nand2_1 _15410_ (.Y(_06225_),
    .A(net2566),
    .B(net5039));
 sg13g2_o21ai_1 _15411_ (.B1(_06225_),
    .Y(_00731_),
    .A1(net5741),
    .A2(net5039));
 sg13g2_nand2_1 _15412_ (.Y(_06226_),
    .A(_02967_),
    .B(net5238));
 sg13g2_nand2_1 _15413_ (.Y(_06227_),
    .A(net3109),
    .B(net5037));
 sg13g2_o21ai_1 _15414_ (.B1(_06227_),
    .Y(_00732_),
    .A1(net5460),
    .A2(net5037));
 sg13g2_nand2_1 _15415_ (.Y(_06228_),
    .A(net2491),
    .B(net5037));
 sg13g2_o21ai_1 _15416_ (.B1(_06228_),
    .Y(_00733_),
    .A1(net5508),
    .A2(net5037));
 sg13g2_nand2_1 _15417_ (.Y(_06229_),
    .A(net2212),
    .B(net5037));
 sg13g2_o21ai_1 _15418_ (.B1(_06229_),
    .Y(_00734_),
    .A1(net5553),
    .A2(net5037));
 sg13g2_nand2_1 _15419_ (.Y(_06230_),
    .A(net3095),
    .B(net5037));
 sg13g2_o21ai_1 _15420_ (.B1(_06230_),
    .Y(_00735_),
    .A1(net5597),
    .A2(net5037));
 sg13g2_nand2_1 _15421_ (.Y(_06231_),
    .A(net2970),
    .B(net5038));
 sg13g2_o21ai_1 _15422_ (.B1(_06231_),
    .Y(_00736_),
    .A1(net5646),
    .A2(net5038));
 sg13g2_nand2_1 _15423_ (.Y(_06232_),
    .A(net2415),
    .B(net5038));
 sg13g2_o21ai_1 _15424_ (.B1(_06232_),
    .Y(_00737_),
    .A1(net5690),
    .A2(net5038));
 sg13g2_nand2_1 _15425_ (.Y(_06233_),
    .A(net3033),
    .B(net5038));
 sg13g2_o21ai_1 _15426_ (.B1(_06233_),
    .Y(_00738_),
    .A1(net5735),
    .A2(net5038));
 sg13g2_nand2_1 _15427_ (.Y(_06234_),
    .A(net2460),
    .B(net5038));
 sg13g2_o21ai_1 _15428_ (.B1(_06234_),
    .Y(_00739_),
    .A1(net5780),
    .A2(net5038));
 sg13g2_nand2_1 _15429_ (.Y(_06235_),
    .A(net5253),
    .B(net5196));
 sg13g2_nand2_1 _15430_ (.Y(_06236_),
    .A(net2661),
    .B(net5036));
 sg13g2_o21ai_1 _15431_ (.B1(_06236_),
    .Y(_00740_),
    .A1(net5454),
    .A2(net5036));
 sg13g2_nand2_1 _15432_ (.Y(_06237_),
    .A(net2645),
    .B(net5035));
 sg13g2_o21ai_1 _15433_ (.B1(_06237_),
    .Y(_00741_),
    .A1(net5501),
    .A2(net5035));
 sg13g2_nand2_1 _15434_ (.Y(_06238_),
    .A(net3146),
    .B(net5036));
 sg13g2_o21ai_1 _15435_ (.B1(_06238_),
    .Y(_00742_),
    .A1(net5547),
    .A2(net5036));
 sg13g2_nand2_1 _15436_ (.Y(_06239_),
    .A(net2878),
    .B(net5035));
 sg13g2_o21ai_1 _15437_ (.B1(_06239_),
    .Y(_00743_),
    .A1(net5590),
    .A2(net5035));
 sg13g2_nand2_1 _15438_ (.Y(_06240_),
    .A(net2918),
    .B(net5036));
 sg13g2_o21ai_1 _15439_ (.B1(_06240_),
    .Y(_00744_),
    .A1(net5633),
    .A2(net5036));
 sg13g2_nand2_1 _15440_ (.Y(_06241_),
    .A(net2521),
    .B(net5036));
 sg13g2_o21ai_1 _15441_ (.B1(_06241_),
    .Y(_00745_),
    .A1(net5679),
    .A2(net5036));
 sg13g2_nand2_1 _15442_ (.Y(_06242_),
    .A(net2928),
    .B(net5035));
 sg13g2_o21ai_1 _15443_ (.B1(_06242_),
    .Y(_00746_),
    .A1(net5723),
    .A2(net5035));
 sg13g2_nand2_1 _15444_ (.Y(_06243_),
    .A(net2198),
    .B(net5035));
 sg13g2_o21ai_1 _15445_ (.B1(_06243_),
    .Y(_00747_),
    .A1(net5771),
    .A2(net5035));
 sg13g2_nand2_1 _15446_ (.Y(_06244_),
    .A(_03211_),
    .B(_03363_));
 sg13g2_nand2_1 _15447_ (.Y(_06245_),
    .A(net3180),
    .B(net5033));
 sg13g2_o21ai_1 _15448_ (.B1(_06245_),
    .Y(_00748_),
    .A1(net5459),
    .A2(net5033));
 sg13g2_nand2_1 _15449_ (.Y(_06246_),
    .A(net2474),
    .B(net5034));
 sg13g2_o21ai_1 _15450_ (.B1(_06246_),
    .Y(_00749_),
    .A1(net5510),
    .A2(net5034));
 sg13g2_nand2_1 _15451_ (.Y(_06247_),
    .A(net2545),
    .B(net5034));
 sg13g2_o21ai_1 _15452_ (.B1(_06247_),
    .Y(_00750_),
    .A1(net5551),
    .A2(net5034));
 sg13g2_nand2_1 _15453_ (.Y(_06248_),
    .A(net2612),
    .B(net5034));
 sg13g2_o21ai_1 _15454_ (.B1(_06248_),
    .Y(_00751_),
    .A1(net5595),
    .A2(_06244_));
 sg13g2_nand2_1 _15455_ (.Y(_06249_),
    .A(net2942),
    .B(net5034));
 sg13g2_o21ai_1 _15456_ (.B1(_06249_),
    .Y(_00752_),
    .A1(net5640),
    .A2(net5034));
 sg13g2_nand2_1 _15457_ (.Y(_06250_),
    .A(net3197),
    .B(net5033));
 sg13g2_o21ai_1 _15458_ (.B1(_06250_),
    .Y(_00753_),
    .A1(net5686),
    .A2(net5033));
 sg13g2_nand2_1 _15459_ (.Y(_06251_),
    .A(net3343),
    .B(net5033));
 sg13g2_o21ai_1 _15460_ (.B1(_06251_),
    .Y(_00754_),
    .A1(net5730),
    .A2(net5033));
 sg13g2_nand2_1 _15461_ (.Y(_06252_),
    .A(net2264),
    .B(net5033));
 sg13g2_o21ai_1 _15462_ (.B1(_06252_),
    .Y(_00755_),
    .A1(net5778),
    .A2(net5033));
 sg13g2_nor2_1 _15463_ (.A(net5227),
    .B(net5258),
    .Y(_06253_));
 sg13g2_nand2_1 _15464_ (.Y(_06254_),
    .A(net5239),
    .B(net5194));
 sg13g2_nand2_1 _15465_ (.Y(_06255_),
    .A(net3132),
    .B(net5031));
 sg13g2_o21ai_1 _15466_ (.B1(_06255_),
    .Y(_00756_),
    .A1(net5440),
    .A2(net5032));
 sg13g2_nand2_1 _15467_ (.Y(_06256_),
    .A(net2739),
    .B(net5031));
 sg13g2_o21ai_1 _15468_ (.B1(_06256_),
    .Y(_00757_),
    .A1(net5485),
    .A2(net5031));
 sg13g2_nand2_1 _15469_ (.Y(_06257_),
    .A(net2445),
    .B(net5032));
 sg13g2_o21ai_1 _15470_ (.B1(_06257_),
    .Y(_00758_),
    .A1(net5532),
    .A2(net5032));
 sg13g2_nand2_1 _15471_ (.Y(_06258_),
    .A(net2457),
    .B(_06254_));
 sg13g2_o21ai_1 _15472_ (.B1(_06258_),
    .Y(_00759_),
    .A1(net5576),
    .A2(net5032));
 sg13g2_nand2_1 _15473_ (.Y(_06259_),
    .A(net3023),
    .B(net5032));
 sg13g2_o21ai_1 _15474_ (.B1(_06259_),
    .Y(_00760_),
    .A1(net5621),
    .A2(net5032));
 sg13g2_nand2_1 _15475_ (.Y(_06260_),
    .A(net2834),
    .B(net5031));
 sg13g2_o21ai_1 _15476_ (.B1(_06260_),
    .Y(_00761_),
    .A1(net5665),
    .A2(net5031));
 sg13g2_nand2_1 _15477_ (.Y(_06261_),
    .A(net2697),
    .B(net5031));
 sg13g2_o21ai_1 _15478_ (.B1(_06261_),
    .Y(_00762_),
    .A1(net5710),
    .A2(net5031));
 sg13g2_nand2_1 _15479_ (.Y(_06262_),
    .A(net2775),
    .B(net5032));
 sg13g2_o21ai_1 _15480_ (.B1(_06262_),
    .Y(_00763_),
    .A1(net5758),
    .A2(net5031));
 sg13g2_nor3_1 _15481_ (.A(net5229),
    .B(net5240),
    .C(_03160_),
    .Y(_06263_));
 sg13g2_nor2_1 _15482_ (.A(net3936),
    .B(net5192),
    .Y(_06264_));
 sg13g2_a21oi_1 _15483_ (.A1(net5446),
    .A2(net5192),
    .Y(_00764_),
    .B1(_06264_));
 sg13g2_nor2_1 _15484_ (.A(net3686),
    .B(net5193),
    .Y(_06265_));
 sg13g2_a21oi_1 _15485_ (.A1(net5490),
    .A2(net5193),
    .Y(_00765_),
    .B1(_06265_));
 sg13g2_nor2_1 _15486_ (.A(net3738),
    .B(net5192),
    .Y(_06266_));
 sg13g2_a21oi_1 _15487_ (.A1(net5540),
    .A2(net5192),
    .Y(_00766_),
    .B1(_06266_));
 sg13g2_nor2_1 _15488_ (.A(net3658),
    .B(net5193),
    .Y(_06267_));
 sg13g2_a21oi_1 _15489_ (.A1(net5584),
    .A2(net5193),
    .Y(_00767_),
    .B1(_06267_));
 sg13g2_nor2_1 _15490_ (.A(net4100),
    .B(net5192),
    .Y(_06268_));
 sg13g2_a21oi_1 _15491_ (.A1(net5626),
    .A2(net5192),
    .Y(_00768_),
    .B1(_06268_));
 sg13g2_nor2_1 _15492_ (.A(net3708),
    .B(net5192),
    .Y(_06269_));
 sg13g2_a21oi_1 _15493_ (.A1(net5674),
    .A2(net5192),
    .Y(_00769_),
    .B1(_06269_));
 sg13g2_nor2_1 _15494_ (.A(net4043),
    .B(net5193),
    .Y(_06270_));
 sg13g2_a21oi_1 _15495_ (.A1(net5719),
    .A2(net5193),
    .Y(_00770_),
    .B1(_06270_));
 sg13g2_nor2_1 _15496_ (.A(net3805),
    .B(net5193),
    .Y(_06271_));
 sg13g2_a21oi_1 _15497_ (.A1(net5761),
    .A2(net5193),
    .Y(_00771_),
    .B1(_06271_));
 sg13g2_nand2_1 _15498_ (.Y(_06272_),
    .A(net5224),
    .B(net5243));
 sg13g2_nand2_1 _15499_ (.Y(_06273_),
    .A(net2376),
    .B(net5029));
 sg13g2_o21ai_1 _15500_ (.B1(_06273_),
    .Y(_00772_),
    .A1(net5430),
    .A2(net5029));
 sg13g2_nand2_1 _15501_ (.Y(_06274_),
    .A(net2380),
    .B(net5030));
 sg13g2_o21ai_1 _15502_ (.B1(_06274_),
    .Y(_00773_),
    .A1(net5474),
    .A2(net5030));
 sg13g2_nand2_1 _15503_ (.Y(_06275_),
    .A(net2992),
    .B(net5029));
 sg13g2_o21ai_1 _15504_ (.B1(_06275_),
    .Y(_00774_),
    .A1(net5520),
    .A2(net5029));
 sg13g2_nand2_1 _15505_ (.Y(_06276_),
    .A(net2454),
    .B(net5030));
 sg13g2_o21ai_1 _15506_ (.B1(_06276_),
    .Y(_00775_),
    .A1(net5563),
    .A2(net5030));
 sg13g2_nand2_1 _15507_ (.Y(_06277_),
    .A(net2764),
    .B(net5029));
 sg13g2_o21ai_1 _15508_ (.B1(_06277_),
    .Y(_00776_),
    .A1(net5610),
    .A2(net5029));
 sg13g2_nand2_1 _15509_ (.Y(_06278_),
    .A(net2307),
    .B(net5030));
 sg13g2_o21ai_1 _15510_ (.B1(_06278_),
    .Y(_00777_),
    .A1(net5656),
    .A2(net5030));
 sg13g2_nand2_1 _15511_ (.Y(_06279_),
    .A(net2674),
    .B(net5029));
 sg13g2_o21ai_1 _15512_ (.B1(_06279_),
    .Y(_00778_),
    .A1(net5701),
    .A2(net5029));
 sg13g2_nand2_1 _15513_ (.Y(_06280_),
    .A(net2859),
    .B(net5030));
 sg13g2_o21ai_1 _15514_ (.B1(_06280_),
    .Y(_00779_),
    .A1(net5746),
    .A2(net5030));
 sg13g2_nand2_1 _15515_ (.Y(_06281_),
    .A(net5224),
    .B(net5242));
 sg13g2_nand2_1 _15516_ (.Y(_06282_),
    .A(net2547),
    .B(net5028));
 sg13g2_o21ai_1 _15517_ (.B1(_06282_),
    .Y(_00780_),
    .A1(net5430),
    .A2(net5028));
 sg13g2_nand2_1 _15518_ (.Y(_06283_),
    .A(net2424),
    .B(net5027));
 sg13g2_o21ai_1 _15519_ (.B1(_06283_),
    .Y(_00781_),
    .A1(net5474),
    .A2(net5027));
 sg13g2_nand2_1 _15520_ (.Y(_06284_),
    .A(net2204),
    .B(_06281_));
 sg13g2_o21ai_1 _15521_ (.B1(_06284_),
    .Y(_00782_),
    .A1(net5520),
    .A2(net5028));
 sg13g2_nand2_1 _15522_ (.Y(_06285_),
    .A(net3183),
    .B(net5027));
 sg13g2_o21ai_1 _15523_ (.B1(_06285_),
    .Y(_00783_),
    .A1(net5563),
    .A2(net5027));
 sg13g2_nand2_1 _15524_ (.Y(_06286_),
    .A(net2283),
    .B(net5028));
 sg13g2_o21ai_1 _15525_ (.B1(_06286_),
    .Y(_00784_),
    .A1(net5610),
    .A2(net5028));
 sg13g2_nand2_1 _15526_ (.Y(_06287_),
    .A(net2328),
    .B(net5027));
 sg13g2_o21ai_1 _15527_ (.B1(_06287_),
    .Y(_00785_),
    .A1(net5656),
    .A2(net5027));
 sg13g2_nand2_1 _15528_ (.Y(_06288_),
    .A(net2642),
    .B(net5028));
 sg13g2_o21ai_1 _15529_ (.B1(_06288_),
    .Y(_00786_),
    .A1(net5701),
    .A2(net5028));
 sg13g2_nand2_1 _15530_ (.Y(_06289_),
    .A(net2496),
    .B(net5027));
 sg13g2_o21ai_1 _15531_ (.B1(_06289_),
    .Y(_00787_),
    .A1(net5746),
    .A2(net5027));
 sg13g2_nor2_1 _15532_ (.A(_02939_),
    .B(net5142),
    .Y(_06290_));
 sg13g2_nor2_1 _15533_ (.A(net4099),
    .B(net4749),
    .Y(_06291_));
 sg13g2_a21oi_1 _15534_ (.A1(net5453),
    .A2(net4749),
    .Y(_00788_),
    .B1(_06291_));
 sg13g2_nor2_1 _15535_ (.A(net3498),
    .B(net4748),
    .Y(_06292_));
 sg13g2_a21oi_1 _15536_ (.A1(net5492),
    .A2(net4748),
    .Y(_00789_),
    .B1(_06292_));
 sg13g2_nor2_1 _15537_ (.A(net3443),
    .B(net4749),
    .Y(_06293_));
 sg13g2_a21oi_1 _15538_ (.A1(net5543),
    .A2(net4749),
    .Y(_00790_),
    .B1(_06293_));
 sg13g2_nor2_1 _15539_ (.A(net4097),
    .B(net4748),
    .Y(_06294_));
 sg13g2_a21oi_1 _15540_ (.A1(net5581),
    .A2(net4748),
    .Y(_00791_),
    .B1(_06294_));
 sg13g2_nor2_1 _15541_ (.A(net3325),
    .B(net4749),
    .Y(_06295_));
 sg13g2_a21oi_1 _15542_ (.A1(net5628),
    .A2(net4749),
    .Y(_00792_),
    .B1(_06295_));
 sg13g2_nor2_1 _15543_ (.A(net3968),
    .B(net4748),
    .Y(_06296_));
 sg13g2_a21oi_1 _15544_ (.A1(net5672),
    .A2(net4748),
    .Y(_00793_),
    .B1(_06296_));
 sg13g2_nor2_1 _15545_ (.A(net4157),
    .B(net4748),
    .Y(_06297_));
 sg13g2_a21oi_1 _15546_ (.A1(net5722),
    .A2(net4748),
    .Y(_00794_),
    .B1(_06297_));
 sg13g2_nor2_1 _15547_ (.A(net4014),
    .B(net4749),
    .Y(_06298_));
 sg13g2_a21oi_1 _15548_ (.A1(net5764),
    .A2(net4749),
    .Y(_00795_),
    .B1(_06298_));
 sg13g2_nor2_2 _15549_ (.A(net5222),
    .B(_03467_),
    .Y(_06299_));
 sg13g2_nor2_1 _15550_ (.A(net3587),
    .B(net5026),
    .Y(_06300_));
 sg13g2_a21oi_1 _15551_ (.A1(net5460),
    .A2(net5026),
    .Y(_00796_),
    .B1(_06300_));
 sg13g2_nor2_1 _15552_ (.A(net3648),
    .B(net5026),
    .Y(_06301_));
 sg13g2_a21oi_1 _15553_ (.A1(net5507),
    .A2(net5026),
    .Y(_00797_),
    .B1(_06301_));
 sg13g2_nor2_1 _15554_ (.A(net3735),
    .B(net5025),
    .Y(_06302_));
 sg13g2_a21oi_1 _15555_ (.A1(net5554),
    .A2(net5025),
    .Y(_00798_),
    .B1(_06302_));
 sg13g2_nor2_1 _15556_ (.A(net3603),
    .B(net5025),
    .Y(_06303_));
 sg13g2_a21oi_1 _15557_ (.A1(net5601),
    .A2(net5025),
    .Y(_00799_),
    .B1(_06303_));
 sg13g2_nor2_1 _15558_ (.A(net3482),
    .B(net5025),
    .Y(_06304_));
 sg13g2_a21oi_1 _15559_ (.A1(net5644),
    .A2(net5025),
    .Y(_00800_),
    .B1(_06304_));
 sg13g2_nor2_1 _15560_ (.A(net3593),
    .B(net5026),
    .Y(_06305_));
 sg13g2_a21oi_1 _15561_ (.A1(net5688),
    .A2(net5026),
    .Y(_00801_),
    .B1(_06305_));
 sg13g2_nor2_1 _15562_ (.A(net2712),
    .B(net5025),
    .Y(_06306_));
 sg13g2_a21oi_1 _15563_ (.A1(net5734),
    .A2(net5025),
    .Y(_00802_),
    .B1(_06306_));
 sg13g2_nor2_1 _15564_ (.A(net2867),
    .B(net5026),
    .Y(_06307_));
 sg13g2_a21oi_1 _15565_ (.A1(net5781),
    .A2(_06299_),
    .Y(_00803_),
    .B1(_06307_));
 sg13g2_nand2b_2 _15566_ (.Y(_06308_),
    .B(net5246),
    .A_N(_02941_));
 sg13g2_o21ai_1 _15567_ (.B1(net1),
    .Y(_06309_),
    .A1(\mem.out_strobe ),
    .A2(net2138));
 sg13g2_a21oi_1 _15568_ (.A1(net2138),
    .A2(_06308_),
    .Y(_00804_),
    .B1(_06309_));
 sg13g2_nor2_1 _15569_ (.A(_00015_),
    .B(_06308_),
    .Y(_06310_));
 sg13g2_o21ai_1 _15570_ (.B1(net6181),
    .Y(_06311_),
    .A1(net4248),
    .A2(net5226));
 sg13g2_a21oi_1 _15571_ (.A1(net5427),
    .A2(_06310_),
    .Y(_00805_),
    .B1(_06311_));
 sg13g2_o21ai_1 _15572_ (.B1(net6181),
    .Y(_06312_),
    .A1(net4246),
    .A2(net5226));
 sg13g2_a21oi_1 _15573_ (.A1(net5472),
    .A2(net5226),
    .Y(_00806_),
    .B1(_06312_));
 sg13g2_o21ai_1 _15574_ (.B1(net6181),
    .Y(_06313_),
    .A1(net4242),
    .A2(net5226));
 sg13g2_a21oi_1 _15575_ (.A1(net5516),
    .A2(net5226),
    .Y(_00807_),
    .B1(_06313_));
 sg13g2_o21ai_1 _15576_ (.B1(net6181),
    .Y(_06314_),
    .A1(net4245),
    .A2(net5226));
 sg13g2_a21oi_1 _15577_ (.A1(net5560),
    .A2(net5225),
    .Y(_00808_),
    .B1(_06314_));
 sg13g2_o21ai_1 _15578_ (.B1(net6181),
    .Y(_06315_),
    .A1(net4243),
    .A2(net5225));
 sg13g2_a21oi_1 _15579_ (.A1(net5608),
    .A2(net5226),
    .Y(_00809_),
    .B1(_06315_));
 sg13g2_o21ai_1 _15580_ (.B1(net6181),
    .Y(_06316_),
    .A1(net4241),
    .A2(net5225));
 sg13g2_a21oi_1 _15581_ (.A1(net5652),
    .A2(net5225),
    .Y(_00810_),
    .B1(_06316_));
 sg13g2_o21ai_1 _15582_ (.B1(net6181),
    .Y(_06317_),
    .A1(net4247),
    .A2(net5225));
 sg13g2_a21oi_1 _15583_ (.A1(net5699),
    .A2(net5225),
    .Y(_00811_),
    .B1(_06317_));
 sg13g2_o21ai_1 _15584_ (.B1(net6181),
    .Y(_06318_),
    .A1(net4250),
    .A2(net5225));
 sg13g2_a21oi_1 _15585_ (.A1(net5744),
    .A2(net5225),
    .Y(_00812_),
    .B1(_06318_));
 sg13g2_nor2_1 _15586_ (.A(_03120_),
    .B(_03364_),
    .Y(_06319_));
 sg13g2_nor2_1 _15587_ (.A(net4133),
    .B(net5023),
    .Y(_06320_));
 sg13g2_a21oi_1 _15588_ (.A1(net5452),
    .A2(net5023),
    .Y(_00813_),
    .B1(_06320_));
 sg13g2_nor2_1 _15589_ (.A(net3971),
    .B(net5023),
    .Y(_06321_));
 sg13g2_a21oi_1 _15590_ (.A1(net5497),
    .A2(net5023),
    .Y(_00814_),
    .B1(_06321_));
 sg13g2_nor2_1 _15591_ (.A(net4030),
    .B(net5023),
    .Y(_06322_));
 sg13g2_a21oi_1 _15592_ (.A1(net5541),
    .A2(net5023),
    .Y(_00815_),
    .B1(_06322_));
 sg13g2_nor2_1 _15593_ (.A(net3954),
    .B(net5024),
    .Y(_06323_));
 sg13g2_a21oi_1 _15594_ (.A1(net5598),
    .A2(net5024),
    .Y(_00816_),
    .B1(_06323_));
 sg13g2_nor2_1 _15595_ (.A(net3500),
    .B(net5024),
    .Y(_06324_));
 sg13g2_a21oi_1 _15596_ (.A1(net5642),
    .A2(net5024),
    .Y(_00817_),
    .B1(_06324_));
 sg13g2_nor2_1 _15597_ (.A(net3871),
    .B(net5024),
    .Y(_06325_));
 sg13g2_a21oi_1 _15598_ (.A1(net5692),
    .A2(net5024),
    .Y(_00818_),
    .B1(_06325_));
 sg13g2_nor2_1 _15599_ (.A(net4129),
    .B(net5024),
    .Y(_06326_));
 sg13g2_a21oi_1 _15600_ (.A1(net5737),
    .A2(net5024),
    .Y(_00819_),
    .B1(_06326_));
 sg13g2_nor2_1 _15601_ (.A(net4090),
    .B(net5023),
    .Y(_06327_));
 sg13g2_a21oi_1 _15602_ (.A1(net5767),
    .A2(net5023),
    .Y(_00820_),
    .B1(_06327_));
 sg13g2_nand2_1 _15603_ (.Y(_06328_),
    .A(net5224),
    .B(net5239));
 sg13g2_nand2_1 _15604_ (.Y(_06329_),
    .A(net2973),
    .B(net5021));
 sg13g2_o21ai_1 _15605_ (.B1(_06329_),
    .Y(_00821_),
    .A1(net5430),
    .A2(net5021));
 sg13g2_nand2_1 _15606_ (.Y(_06330_),
    .A(net3379),
    .B(net5022));
 sg13g2_o21ai_1 _15607_ (.B1(_06330_),
    .Y(_00822_),
    .A1(net5479),
    .A2(net5022));
 sg13g2_nand2_1 _15608_ (.Y(_06331_),
    .A(net3045),
    .B(net5022));
 sg13g2_o21ai_1 _15609_ (.B1(_06331_),
    .Y(_00823_),
    .A1(net5520),
    .A2(net5021));
 sg13g2_nand2_1 _15610_ (.Y(_06332_),
    .A(net2573),
    .B(net5022));
 sg13g2_o21ai_1 _15611_ (.B1(_06332_),
    .Y(_00824_),
    .A1(net5563),
    .A2(_06328_));
 sg13g2_nand2_1 _15612_ (.Y(_06333_),
    .A(net2651),
    .B(net5021));
 sg13g2_o21ai_1 _15613_ (.B1(_06333_),
    .Y(_00825_),
    .A1(net5609),
    .A2(net5021));
 sg13g2_nand2_1 _15614_ (.Y(_06334_),
    .A(net3421),
    .B(net5022));
 sg13g2_o21ai_1 _15615_ (.B1(_06334_),
    .Y(_00826_),
    .A1(net5656),
    .A2(net5022));
 sg13g2_nand2_1 _15616_ (.Y(_06335_),
    .A(net2224),
    .B(net5021));
 sg13g2_o21ai_1 _15617_ (.B1(_06335_),
    .Y(_00827_),
    .A1(net5701),
    .A2(net5021));
 sg13g2_nand2_1 _15618_ (.Y(_06336_),
    .A(net2287),
    .B(net5021));
 sg13g2_o21ai_1 _15619_ (.B1(_06336_),
    .Y(_00828_),
    .A1(net5746),
    .A2(net5022));
 sg13g2_nor2_1 _15620_ (.A(net5155),
    .B(net5241),
    .Y(_06337_));
 sg13g2_nor2_1 _15621_ (.A(net4058),
    .B(net4746),
    .Y(_06338_));
 sg13g2_a21oi_1 _15622_ (.A1(net5424),
    .A2(net4746),
    .Y(_00829_),
    .B1(_06338_));
 sg13g2_nor2_1 _15623_ (.A(net3610),
    .B(net4747),
    .Y(_06339_));
 sg13g2_a21oi_1 _15624_ (.A1(net5468),
    .A2(net4747),
    .Y(_00830_),
    .B1(_06339_));
 sg13g2_nor2_1 _15625_ (.A(net3938),
    .B(net4747),
    .Y(_06340_));
 sg13g2_a21oi_1 _15626_ (.A1(net5513),
    .A2(net4747),
    .Y(_00831_),
    .B1(_06340_));
 sg13g2_nor2_1 _15627_ (.A(net3979),
    .B(net4747),
    .Y(_06341_));
 sg13g2_a21oi_1 _15628_ (.A1(net5558),
    .A2(net4747),
    .Y(_00832_),
    .B1(_06341_));
 sg13g2_nor2_1 _15629_ (.A(net3771),
    .B(net4747),
    .Y(_06342_));
 sg13g2_a21oi_1 _15630_ (.A1(net5604),
    .A2(net4747),
    .Y(_00833_),
    .B1(_06342_));
 sg13g2_nor2_1 _15631_ (.A(net3684),
    .B(net4746),
    .Y(_06343_));
 sg13g2_a21oi_1 _15632_ (.A1(net5650),
    .A2(net4746),
    .Y(_00834_),
    .B1(_06343_));
 sg13g2_nor2_1 _15633_ (.A(net3422),
    .B(net4746),
    .Y(_06344_));
 sg13g2_a21oi_1 _15634_ (.A1(net5696),
    .A2(net4746),
    .Y(_00835_),
    .B1(_06344_));
 sg13g2_nor2_1 _15635_ (.A(net3731),
    .B(net4746),
    .Y(_06345_));
 sg13g2_a21oi_1 _15636_ (.A1(net5741),
    .A2(net4746),
    .Y(_00836_),
    .B1(_06345_));
 sg13g2_nand2_1 _15637_ (.Y(_06346_),
    .A(net5224),
    .B(net5245));
 sg13g2_nand2_1 _15638_ (.Y(_06347_),
    .A(net2174),
    .B(net5019));
 sg13g2_o21ai_1 _15639_ (.B1(_06347_),
    .Y(_00837_),
    .A1(net5430),
    .A2(net5019));
 sg13g2_nand2_1 _15640_ (.Y(_06348_),
    .A(net2546),
    .B(net5020));
 sg13g2_o21ai_1 _15641_ (.B1(_06348_),
    .Y(_00838_),
    .A1(net5478),
    .A2(net5020));
 sg13g2_nand2_1 _15642_ (.Y(_06349_),
    .A(net2965),
    .B(net5019));
 sg13g2_o21ai_1 _15643_ (.B1(_06349_),
    .Y(_00839_),
    .A1(net5519),
    .A2(net5019));
 sg13g2_nand2_1 _15644_ (.Y(_06350_),
    .A(net3002),
    .B(net5020));
 sg13g2_o21ai_1 _15645_ (.B1(_06350_),
    .Y(_00840_),
    .A1(net5566),
    .A2(net5020));
 sg13g2_nand2_1 _15646_ (.Y(_06351_),
    .A(net2887),
    .B(net5019));
 sg13g2_o21ai_1 _15647_ (.B1(_06351_),
    .Y(_00841_),
    .A1(net5609),
    .A2(net5019));
 sg13g2_nand2_1 _15648_ (.Y(_06352_),
    .A(net2648),
    .B(net5020));
 sg13g2_o21ai_1 _15649_ (.B1(_06352_),
    .Y(_00842_),
    .A1(net5657),
    .A2(net5020));
 sg13g2_nand2_1 _15650_ (.Y(_06353_),
    .A(net2312),
    .B(net5019));
 sg13g2_o21ai_1 _15651_ (.B1(_06353_),
    .Y(_00843_),
    .A1(net5701),
    .A2(net5019));
 sg13g2_nand2_1 _15652_ (.Y(_06354_),
    .A(net2326),
    .B(net5020));
 sg13g2_o21ai_1 _15653_ (.B1(_06354_),
    .Y(_00844_),
    .A1(net5747),
    .A2(net5020));
 sg13g2_nand2_1 _15654_ (.Y(_06355_),
    .A(net5223),
    .B(net5251));
 sg13g2_nand2_1 _15655_ (.Y(_06356_),
    .A(net2961),
    .B(net5017));
 sg13g2_o21ai_1 _15656_ (.B1(_06356_),
    .Y(_00845_),
    .A1(net5428),
    .A2(net5017));
 sg13g2_nand2_1 _15657_ (.Y(_06357_),
    .A(net2996),
    .B(net5018));
 sg13g2_o21ai_1 _15658_ (.B1(_06357_),
    .Y(_00846_),
    .A1(net5474),
    .A2(net5018));
 sg13g2_nand2_1 _15659_ (.Y(_06358_),
    .A(net3318),
    .B(net5017));
 sg13g2_o21ai_1 _15660_ (.B1(_06358_),
    .Y(_00847_),
    .A1(net5519),
    .A2(net5017));
 sg13g2_nand2_1 _15661_ (.Y(_06359_),
    .A(net2222),
    .B(net5018));
 sg13g2_o21ai_1 _15662_ (.B1(_06359_),
    .Y(_00848_),
    .A1(net5563),
    .A2(net5018));
 sg13g2_nand2_1 _15663_ (.Y(_06360_),
    .A(net3113),
    .B(net5017));
 sg13g2_o21ai_1 _15664_ (.B1(_06360_),
    .Y(_00849_),
    .A1(net5609),
    .A2(net5017));
 sg13g2_nand2_1 _15665_ (.Y(_06361_),
    .A(net2632),
    .B(net5018));
 sg13g2_o21ai_1 _15666_ (.B1(_06361_),
    .Y(_00850_),
    .A1(net5657),
    .A2(net5018));
 sg13g2_nand2_1 _15667_ (.Y(_06362_),
    .A(net2746),
    .B(net5017));
 sg13g2_o21ai_1 _15668_ (.B1(_06362_),
    .Y(_00851_),
    .A1(net5701),
    .A2(net5017));
 sg13g2_nand2_1 _15669_ (.Y(_06363_),
    .A(net3096),
    .B(net5018));
 sg13g2_o21ai_1 _15670_ (.B1(_06363_),
    .Y(_00852_),
    .A1(net5746),
    .A2(net5018));
 sg13g2_nand2_1 _15671_ (.Y(_06364_),
    .A(net5223),
    .B(net5246));
 sg13g2_nand2_1 _15672_ (.Y(_06365_),
    .A(net2810),
    .B(net5015));
 sg13g2_o21ai_1 _15673_ (.B1(_06365_),
    .Y(_00853_),
    .A1(net5433),
    .A2(net5015));
 sg13g2_nand2_1 _15674_ (.Y(_06366_),
    .A(net2303),
    .B(net5016));
 sg13g2_o21ai_1 _15675_ (.B1(_06366_),
    .Y(_00854_),
    .A1(net5475),
    .A2(net5016));
 sg13g2_nand2_1 _15676_ (.Y(_06367_),
    .A(net3164),
    .B(net5015));
 sg13g2_o21ai_1 _15677_ (.B1(_06367_),
    .Y(_00855_),
    .A1(net5519),
    .A2(net5015));
 sg13g2_nand2_1 _15678_ (.Y(_06368_),
    .A(net2293),
    .B(net5016));
 sg13g2_o21ai_1 _15679_ (.B1(_06368_),
    .Y(_00856_),
    .A1(net5564),
    .A2(net5016));
 sg13g2_nand2_1 _15680_ (.Y(_06369_),
    .A(net2325),
    .B(net5015));
 sg13g2_o21ai_1 _15681_ (.B1(_06369_),
    .Y(_00857_),
    .A1(net5613),
    .A2(net5015));
 sg13g2_nand2_1 _15682_ (.Y(_06370_),
    .A(net3024),
    .B(net5016));
 sg13g2_o21ai_1 _15683_ (.B1(_06370_),
    .Y(_00858_),
    .A1(net5657),
    .A2(net5016));
 sg13g2_nand2_1 _15684_ (.Y(_06371_),
    .A(net3135),
    .B(net5015));
 sg13g2_o21ai_1 _15685_ (.B1(_06371_),
    .Y(_00859_),
    .A1(net5702),
    .A2(net5015));
 sg13g2_nand2_1 _15686_ (.Y(_06372_),
    .A(net2599),
    .B(net5016));
 sg13g2_o21ai_1 _15687_ (.B1(_06372_),
    .Y(_00860_),
    .A1(net5747),
    .A2(net5016));
 sg13g2_nor3_1 _15688_ (.A(net5229),
    .B(net5259),
    .C(net5241),
    .Y(_06373_));
 sg13g2_nor2_1 _15689_ (.A(net4040),
    .B(net5190),
    .Y(_06374_));
 sg13g2_a21oi_1 _15690_ (.A1(net5433),
    .A2(net5190),
    .Y(_00861_),
    .B1(_06374_));
 sg13g2_nor2_1 _15691_ (.A(net3650),
    .B(net5191),
    .Y(_06375_));
 sg13g2_a21oi_1 _15692_ (.A1(net5475),
    .A2(net5191),
    .Y(_00862_),
    .B1(_06375_));
 sg13g2_nor2_1 _15693_ (.A(net3949),
    .B(net5190),
    .Y(_06376_));
 sg13g2_a21oi_1 _15694_ (.A1(net5519),
    .A2(net5190),
    .Y(_00863_),
    .B1(_06376_));
 sg13g2_nor2_1 _15695_ (.A(net3572),
    .B(net5191),
    .Y(_06377_));
 sg13g2_a21oi_1 _15696_ (.A1(net5564),
    .A2(net5191),
    .Y(_00864_),
    .B1(_06377_));
 sg13g2_nor2_1 _15697_ (.A(net3959),
    .B(net5190),
    .Y(_06378_));
 sg13g2_a21oi_1 _15698_ (.A1(net5613),
    .A2(net5190),
    .Y(_00865_),
    .B1(_06378_));
 sg13g2_nor2_1 _15699_ (.A(net3886),
    .B(net5191),
    .Y(_06379_));
 sg13g2_a21oi_1 _15700_ (.A1(net5657),
    .A2(net5191),
    .Y(_00866_),
    .B1(_06379_));
 sg13g2_nor2_1 _15701_ (.A(net3698),
    .B(net5190),
    .Y(_06380_));
 sg13g2_a21oi_1 _15702_ (.A1(net5702),
    .A2(net5190),
    .Y(_00867_),
    .B1(_06380_));
 sg13g2_nor2_1 _15703_ (.A(net3926),
    .B(net5191),
    .Y(_06381_));
 sg13g2_a21oi_1 _15704_ (.A1(net5747),
    .A2(net5191),
    .Y(_00868_),
    .B1(_06381_));
 sg13g2_nand2_1 _15705_ (.Y(_06382_),
    .A(net5216),
    .B(net5248));
 sg13g2_nand2_1 _15706_ (.Y(_06383_),
    .A(net2148),
    .B(net5014));
 sg13g2_o21ai_1 _15707_ (.B1(_06383_),
    .Y(_00869_),
    .A1(net5437),
    .A2(net5014));
 sg13g2_nand2_1 _15708_ (.Y(_06384_),
    .A(net2606),
    .B(net5014));
 sg13g2_o21ai_1 _15709_ (.B1(_06384_),
    .Y(_00870_),
    .A1(net5482),
    .A2(net5014));
 sg13g2_nand2_1 _15710_ (.Y(_06385_),
    .A(net2978),
    .B(net5014));
 sg13g2_o21ai_1 _15711_ (.B1(_06385_),
    .Y(_00871_),
    .A1(net5528),
    .A2(net5014));
 sg13g2_nand2_1 _15712_ (.Y(_06386_),
    .A(net2619),
    .B(net5013));
 sg13g2_o21ai_1 _15713_ (.B1(_06386_),
    .Y(_00872_),
    .A1(net5569),
    .A2(net5013));
 sg13g2_nand2_1 _15714_ (.Y(_06387_),
    .A(net2710),
    .B(net5014));
 sg13g2_o21ai_1 _15715_ (.B1(_06387_),
    .Y(_00873_),
    .A1(net5617),
    .A2(net5014));
 sg13g2_nand2_1 _15716_ (.Y(_06388_),
    .A(net3212),
    .B(net5013));
 sg13g2_o21ai_1 _15717_ (.B1(_06388_),
    .Y(_00874_),
    .A1(net5662),
    .A2(net5013));
 sg13g2_nand2_1 _15718_ (.Y(_06389_),
    .A(net2270),
    .B(net5013));
 sg13g2_o21ai_1 _15719_ (.B1(_06389_),
    .Y(_00875_),
    .A1(net5706),
    .A2(net5013));
 sg13g2_nand2_1 _15720_ (.Y(_06390_),
    .A(net2886),
    .B(net5013));
 sg13g2_o21ai_1 _15721_ (.B1(_06390_),
    .Y(_00876_),
    .A1(net5752),
    .A2(net5013));
 sg13g2_nor3_1 _15722_ (.A(net5259),
    .B(net5227),
    .C(net5252),
    .Y(_06391_));
 sg13g2_nor2_1 _15723_ (.A(net4108),
    .B(net5189),
    .Y(_06392_));
 sg13g2_a21oi_1 _15724_ (.A1(net5437),
    .A2(net5189),
    .Y(_00877_),
    .B1(_06392_));
 sg13g2_nor2_1 _15725_ (.A(net3656),
    .B(net5189),
    .Y(_06393_));
 sg13g2_a21oi_1 _15726_ (.A1(net5482),
    .A2(net5189),
    .Y(_00878_),
    .B1(_06393_));
 sg13g2_nor2_1 _15727_ (.A(net3589),
    .B(net5189),
    .Y(_06394_));
 sg13g2_a21oi_1 _15728_ (.A1(net5528),
    .A2(net5189),
    .Y(_00879_),
    .B1(_06394_));
 sg13g2_nor2_1 _15729_ (.A(net3529),
    .B(net5188),
    .Y(_06395_));
 sg13g2_a21oi_1 _15730_ (.A1(net5571),
    .A2(net5188),
    .Y(_00880_),
    .B1(_06395_));
 sg13g2_nor2_1 _15731_ (.A(net4029),
    .B(net5189),
    .Y(_06396_));
 sg13g2_a21oi_1 _15732_ (.A1(net5616),
    .A2(net5189),
    .Y(_00881_),
    .B1(_06396_));
 sg13g2_nor2_1 _15733_ (.A(net3370),
    .B(net5188),
    .Y(_06397_));
 sg13g2_a21oi_1 _15734_ (.A1(net5662),
    .A2(net5188),
    .Y(_00882_),
    .B1(_06397_));
 sg13g2_nor2_1 _15735_ (.A(net3542),
    .B(net5188),
    .Y(_06398_));
 sg13g2_a21oi_1 _15736_ (.A1(net5706),
    .A2(net5188),
    .Y(_00883_),
    .B1(_06398_));
 sg13g2_nor2_1 _15737_ (.A(net3986),
    .B(net5188),
    .Y(_06399_));
 sg13g2_a21oi_1 _15738_ (.A1(net5752),
    .A2(net5188),
    .Y(_00884_),
    .B1(_06399_));
 sg13g2_nor3_1 _15739_ (.A(net5259),
    .B(net5227),
    .C(net5254),
    .Y(_06400_));
 sg13g2_nor2_1 _15740_ (.A(net2777),
    .B(net5187),
    .Y(_06401_));
 sg13g2_a21oi_1 _15741_ (.A1(net5437),
    .A2(net5187),
    .Y(_00885_),
    .B1(_06401_));
 sg13g2_nor2_1 _15742_ (.A(net3636),
    .B(net5187),
    .Y(_06402_));
 sg13g2_a21oi_1 _15743_ (.A1(net5482),
    .A2(net5187),
    .Y(_00886_),
    .B1(_06402_));
 sg13g2_nor2_1 _15744_ (.A(net4111),
    .B(net5187),
    .Y(_06403_));
 sg13g2_a21oi_1 _15745_ (.A1(net5528),
    .A2(net5187),
    .Y(_00887_),
    .B1(_06403_));
 sg13g2_nor2_1 _15746_ (.A(net3635),
    .B(net5186),
    .Y(_06404_));
 sg13g2_a21oi_1 _15747_ (.A1(net5569),
    .A2(net5186),
    .Y(_00888_),
    .B1(_06404_));
 sg13g2_nor2_1 _15748_ (.A(net3546),
    .B(net5187),
    .Y(_06405_));
 sg13g2_a21oi_1 _15749_ (.A1(net5616),
    .A2(net5187),
    .Y(_00889_),
    .B1(_06405_));
 sg13g2_nor2_1 _15750_ (.A(net3711),
    .B(net5186),
    .Y(_06406_));
 sg13g2_a21oi_1 _15751_ (.A1(net5662),
    .A2(net5186),
    .Y(_00890_),
    .B1(_06406_));
 sg13g2_nor2_1 _15752_ (.A(net3763),
    .B(net5186),
    .Y(_06407_));
 sg13g2_a21oi_1 _15753_ (.A1(net5706),
    .A2(net5186),
    .Y(_00891_),
    .B1(_06407_));
 sg13g2_nor2_1 _15754_ (.A(net3614),
    .B(net5186),
    .Y(_06408_));
 sg13g2_a21oi_1 _15755_ (.A1(net5752),
    .A2(net5186),
    .Y(_00892_),
    .B1(_06408_));
 sg13g2_nand3_1 _15756_ (.B(net5220),
    .C(net5248),
    .A(_02966_),
    .Y(_06409_));
 sg13g2_nand2_1 _15757_ (.Y(_06410_),
    .A(net2681),
    .B(net5012));
 sg13g2_o21ai_1 _15758_ (.B1(_06410_),
    .Y(_00893_),
    .A1(net5438),
    .A2(net5012));
 sg13g2_nand2_1 _15759_ (.Y(_06411_),
    .A(net3064),
    .B(net5012));
 sg13g2_o21ai_1 _15760_ (.B1(_06411_),
    .Y(_00894_),
    .A1(net5482),
    .A2(net5012));
 sg13g2_nand2_1 _15761_ (.Y(_06412_),
    .A(net2972),
    .B(net5012));
 sg13g2_o21ai_1 _15762_ (.B1(_06412_),
    .Y(_00895_),
    .A1(net5529),
    .A2(net5012));
 sg13g2_nand2_1 _15763_ (.Y(_06413_),
    .A(net2755),
    .B(net5011));
 sg13g2_o21ai_1 _15764_ (.B1(_06413_),
    .Y(_00896_),
    .A1(net5573),
    .A2(net5011));
 sg13g2_nand2_1 _15765_ (.Y(_06414_),
    .A(net3543),
    .B(_06409_));
 sg13g2_o21ai_1 _15766_ (.B1(_06414_),
    .Y(_00897_),
    .A1(net5618),
    .A2(net5012));
 sg13g2_nand2_1 _15767_ (.Y(_06415_),
    .A(net2273),
    .B(net5011));
 sg13g2_o21ai_1 _15768_ (.B1(_06415_),
    .Y(_00898_),
    .A1(net5671),
    .A2(net5011));
 sg13g2_nand2_1 _15769_ (.Y(_06416_),
    .A(net2993),
    .B(net5011));
 sg13g2_o21ai_1 _15770_ (.B1(_06416_),
    .Y(_00899_),
    .A1(net5707),
    .A2(net5011));
 sg13g2_nand2_1 _15771_ (.Y(_06417_),
    .A(net3254),
    .B(net5011));
 sg13g2_o21ai_1 _15772_ (.B1(_06417_),
    .Y(_00900_),
    .A1(net5753),
    .A2(net5011));
 sg13g2_nand2_1 _15773_ (.Y(_06418_),
    .A(net5235),
    .B(net5215));
 sg13g2_nand2_1 _15774_ (.Y(_06419_),
    .A(net2133),
    .B(net5009));
 sg13g2_o21ai_1 _15775_ (.B1(_06419_),
    .Y(_00901_),
    .A1(net5437),
    .A2(net5009));
 sg13g2_nand2_1 _15776_ (.Y(_06420_),
    .A(net2365),
    .B(net5010));
 sg13g2_o21ai_1 _15777_ (.B1(_06420_),
    .Y(_00902_),
    .A1(net5483),
    .A2(net5010));
 sg13g2_nand2_1 _15778_ (.Y(_06421_),
    .A(net2354),
    .B(net5009));
 sg13g2_o21ai_1 _15779_ (.B1(_06421_),
    .Y(_00903_),
    .A1(net5528),
    .A2(net5009));
 sg13g2_nand2_1 _15780_ (.Y(_06422_),
    .A(net3354),
    .B(net5008));
 sg13g2_o21ai_1 _15781_ (.B1(_06422_),
    .Y(_00904_),
    .A1(net5572),
    .A2(net5009));
 sg13g2_nand2_1 _15782_ (.Y(_06423_),
    .A(net2860),
    .B(net5008));
 sg13g2_o21ai_1 _15783_ (.B1(_06423_),
    .Y(_00905_),
    .A1(net5618),
    .A2(net5009));
 sg13g2_nand2_1 _15784_ (.Y(_06424_),
    .A(net2368),
    .B(net5008));
 sg13g2_o21ai_1 _15785_ (.B1(_06424_),
    .Y(_00906_),
    .A1(net5663),
    .A2(net5008));
 sg13g2_nand2_1 _15786_ (.Y(_06425_),
    .A(net2323),
    .B(net5008));
 sg13g2_o21ai_1 _15787_ (.B1(_06425_),
    .Y(_00907_),
    .A1(net5706),
    .A2(net5008));
 sg13g2_nand2_1 _15788_ (.Y(_06426_),
    .A(net2692),
    .B(net5008));
 sg13g2_o21ai_1 _15789_ (.B1(_06426_),
    .Y(_00908_),
    .A1(net5752),
    .A2(net5008));
 sg13g2_nand2_1 _15790_ (.Y(_06427_),
    .A(net5234),
    .B(net5215));
 sg13g2_nand2_1 _15791_ (.Y(_06428_),
    .A(net3355),
    .B(net5007));
 sg13g2_o21ai_1 _15792_ (.B1(_06428_),
    .Y(_00909_),
    .A1(net5437),
    .A2(net5007));
 sg13g2_nand2_1 _15793_ (.Y(_06429_),
    .A(net3048),
    .B(net5007));
 sg13g2_o21ai_1 _15794_ (.B1(_06429_),
    .Y(_00910_),
    .A1(net5483),
    .A2(net5007));
 sg13g2_nand2_1 _15795_ (.Y(_06430_),
    .A(net3290),
    .B(net5006));
 sg13g2_o21ai_1 _15796_ (.B1(_06430_),
    .Y(_00911_),
    .A1(net5528),
    .A2(net5006));
 sg13g2_nand2_1 _15797_ (.Y(_06431_),
    .A(net2945),
    .B(net5005));
 sg13g2_o21ai_1 _15798_ (.B1(_06431_),
    .Y(_00912_),
    .A1(net5572),
    .A2(net5005));
 sg13g2_nand2_1 _15799_ (.Y(_06432_),
    .A(net2885),
    .B(net5006));
 sg13g2_o21ai_1 _15800_ (.B1(_06432_),
    .Y(_00913_),
    .A1(net5618),
    .A2(net5006));
 sg13g2_nand2_1 _15801_ (.Y(_06433_),
    .A(net2450),
    .B(net5005));
 sg13g2_o21ai_1 _15802_ (.B1(_06433_),
    .Y(_00914_),
    .A1(net5662),
    .A2(net5005));
 sg13g2_nand2_1 _15803_ (.Y(_06434_),
    .A(net3186),
    .B(net5005));
 sg13g2_o21ai_1 _15804_ (.B1(_06434_),
    .Y(_00915_),
    .A1(net5706),
    .A2(net5005));
 sg13g2_nand2_1 _15805_ (.Y(_06435_),
    .A(net2819),
    .B(net5005));
 sg13g2_o21ai_1 _15806_ (.B1(_06435_),
    .Y(_00916_),
    .A1(net5752),
    .A2(net5005));
 sg13g2_nand2_1 _15807_ (.Y(_06436_),
    .A(net5236),
    .B(net5216));
 sg13g2_nor2_1 _15808_ (.A(\mem.data_in[0] ),
    .B(net5004),
    .Y(_06437_));
 sg13g2_a21oi_1 _15809_ (.A1(_02886_),
    .A2(net5004),
    .Y(_00917_),
    .B1(_06437_));
 sg13g2_nand2_1 _15810_ (.Y(_06438_),
    .A(net3288),
    .B(net5004));
 sg13g2_o21ai_1 _15811_ (.B1(_06438_),
    .Y(_00918_),
    .A1(net5483),
    .A2(net5004));
 sg13g2_nand2_1 _15812_ (.Y(_06439_),
    .A(net2825),
    .B(net5003));
 sg13g2_o21ai_1 _15813_ (.B1(_06439_),
    .Y(_00919_),
    .A1(net5528),
    .A2(net5002));
 sg13g2_nand2_1 _15814_ (.Y(_06440_),
    .A(net3077),
    .B(net5003));
 sg13g2_o21ai_1 _15815_ (.B1(_06440_),
    .Y(_00920_),
    .A1(net5572),
    .A2(net5002));
 sg13g2_nand2_1 _15816_ (.Y(_06441_),
    .A(net2761),
    .B(net5003));
 sg13g2_o21ai_1 _15817_ (.B1(_06441_),
    .Y(_00921_),
    .A1(net5618),
    .A2(net5003));
 sg13g2_nand2_1 _15818_ (.Y(_06442_),
    .A(net2607),
    .B(net5002));
 sg13g2_o21ai_1 _15819_ (.B1(_06442_),
    .Y(_00922_),
    .A1(net5663),
    .A2(net5002));
 sg13g2_nand2_1 _15820_ (.Y(_06443_),
    .A(net2319),
    .B(net5002));
 sg13g2_o21ai_1 _15821_ (.B1(_06443_),
    .Y(_00923_),
    .A1(net5706),
    .A2(net5002));
 sg13g2_nand2_1 _15822_ (.Y(_06444_),
    .A(net2876),
    .B(net5002));
 sg13g2_o21ai_1 _15823_ (.B1(_06444_),
    .Y(_00924_),
    .A1(net5752),
    .A2(net5002));
 sg13g2_nand2_1 _15824_ (.Y(_06445_),
    .A(net5237),
    .B(net5216));
 sg13g2_nand2_1 _15825_ (.Y(_06446_),
    .A(net2302),
    .B(net5001));
 sg13g2_o21ai_1 _15826_ (.B1(_06446_),
    .Y(_00925_),
    .A1(net5437),
    .A2(net5001));
 sg13g2_nand2_1 _15827_ (.Y(_06447_),
    .A(net2471),
    .B(net5001));
 sg13g2_o21ai_1 _15828_ (.B1(_06447_),
    .Y(_00926_),
    .A1(net5482),
    .A2(net5001));
 sg13g2_nand2_1 _15829_ (.Y(_06448_),
    .A(net2750),
    .B(net4999));
 sg13g2_o21ai_1 _15830_ (.B1(_06448_),
    .Y(_00927_),
    .A1(net5528),
    .A2(net5000));
 sg13g2_nand2_1 _15831_ (.Y(_06449_),
    .A(net2384),
    .B(net5000));
 sg13g2_o21ai_1 _15832_ (.B1(_06449_),
    .Y(_00928_),
    .A1(net5572),
    .A2(net4999));
 sg13g2_nand2_1 _15833_ (.Y(_06450_),
    .A(net2733),
    .B(net5000));
 sg13g2_o21ai_1 _15834_ (.B1(_06450_),
    .Y(_00929_),
    .A1(net5618),
    .A2(net5000));
 sg13g2_nand2_1 _15835_ (.Y(_06451_),
    .A(net2458),
    .B(net4999));
 sg13g2_o21ai_1 _15836_ (.B1(_06451_),
    .Y(_00930_),
    .A1(net5663),
    .A2(net4999));
 sg13g2_nand2_1 _15837_ (.Y(_06452_),
    .A(net2317),
    .B(net4999));
 sg13g2_o21ai_1 _15838_ (.B1(_06452_),
    .Y(_00931_),
    .A1(net5706),
    .A2(net4999));
 sg13g2_nand2_1 _15839_ (.Y(_06453_),
    .A(net2888),
    .B(net4999));
 sg13g2_o21ai_1 _15840_ (.B1(_06453_),
    .Y(_00932_),
    .A1(net5752),
    .A2(net4999));
 sg13g2_nand2_1 _15841_ (.Y(_06454_),
    .A(net5244),
    .B(net5215));
 sg13g2_nand2_1 _15842_ (.Y(_06455_),
    .A(net2332),
    .B(net4997));
 sg13g2_o21ai_1 _15843_ (.B1(_06455_),
    .Y(_00933_),
    .A1(net5436),
    .A2(net4997));
 sg13g2_nand2_1 _15844_ (.Y(_06456_),
    .A(net2240),
    .B(net4997));
 sg13g2_o21ai_1 _15845_ (.B1(_06456_),
    .Y(_00934_),
    .A1(net5478),
    .A2(net4997));
 sg13g2_nand2_1 _15846_ (.Y(_06457_),
    .A(net3004),
    .B(net4998));
 sg13g2_o21ai_1 _15847_ (.B1(_06457_),
    .Y(_00935_),
    .A1(net5526),
    .A2(net4998));
 sg13g2_nand2_1 _15848_ (.Y(_06458_),
    .A(net2343),
    .B(net4997));
 sg13g2_o21ai_1 _15849_ (.B1(_06458_),
    .Y(_00936_),
    .A1(net5571),
    .A2(net4997));
 sg13g2_nand2_1 _15850_ (.Y(_06459_),
    .A(net2540),
    .B(net4998));
 sg13g2_o21ai_1 _15851_ (.B1(_06459_),
    .Y(_00937_),
    .A1(net5616),
    .A2(net4998));
 sg13g2_nand2_1 _15852_ (.Y(_06460_),
    .A(net3137),
    .B(net4997));
 sg13g2_o21ai_1 _15853_ (.B1(_06460_),
    .Y(_00938_),
    .A1(net5658),
    .A2(net4997));
 sg13g2_nand2_1 _15854_ (.Y(_06461_),
    .A(net2909),
    .B(net4998));
 sg13g2_o21ai_1 _15855_ (.B1(_06461_),
    .Y(_00939_),
    .A1(net5708),
    .A2(net4998));
 sg13g2_nand2_1 _15856_ (.Y(_06462_),
    .A(net3653),
    .B(net4998));
 sg13g2_o21ai_1 _15857_ (.B1(_06462_),
    .Y(_00940_),
    .A1(net5754),
    .A2(net4998));
 sg13g2_nand2_1 _15858_ (.Y(_06463_),
    .A(net5239),
    .B(net5215));
 sg13g2_nand2_1 _15859_ (.Y(_06464_),
    .A(net2790),
    .B(net4995));
 sg13g2_o21ai_1 _15860_ (.B1(_06464_),
    .Y(_00941_),
    .A1(net5436),
    .A2(net4995));
 sg13g2_nand2_1 _15861_ (.Y(_06465_),
    .A(net2543),
    .B(net4995));
 sg13g2_o21ai_1 _15862_ (.B1(_06465_),
    .Y(_00942_),
    .A1(net5478),
    .A2(net4995));
 sg13g2_nand2_1 _15863_ (.Y(_06466_),
    .A(net2964),
    .B(net4996));
 sg13g2_o21ai_1 _15864_ (.B1(_06466_),
    .Y(_00943_),
    .A1(net5526),
    .A2(net4996));
 sg13g2_nand2_1 _15865_ (.Y(_06467_),
    .A(net2659),
    .B(net4995));
 sg13g2_o21ai_1 _15866_ (.B1(_06467_),
    .Y(_00944_),
    .A1(net5571),
    .A2(net4995));
 sg13g2_nand2_1 _15867_ (.Y(_06468_),
    .A(net2800),
    .B(net4996));
 sg13g2_o21ai_1 _15868_ (.B1(_06468_),
    .Y(_00945_),
    .A1(net5616),
    .A2(net4996));
 sg13g2_nand2_1 _15869_ (.Y(_06469_),
    .A(net3178),
    .B(net4995));
 sg13g2_o21ai_1 _15870_ (.B1(_06469_),
    .Y(_00946_),
    .A1(net5657),
    .A2(net4995));
 sg13g2_nand2_1 _15871_ (.Y(_06470_),
    .A(net2616),
    .B(net4996));
 sg13g2_o21ai_1 _15872_ (.B1(_06470_),
    .Y(_00947_),
    .A1(net5708),
    .A2(net4996));
 sg13g2_nand2_1 _15873_ (.Y(_06471_),
    .A(net2562),
    .B(net4996));
 sg13g2_o21ai_1 _15874_ (.B1(_06471_),
    .Y(_00948_),
    .A1(net5754),
    .A2(net4996));
 sg13g2_nand2_1 _15875_ (.Y(_06472_),
    .A(net5242),
    .B(net5215));
 sg13g2_nand2_1 _15876_ (.Y(_06473_),
    .A(net3119),
    .B(net4993));
 sg13g2_o21ai_1 _15877_ (.B1(_06473_),
    .Y(_00949_),
    .A1(net5436),
    .A2(net4993));
 sg13g2_nand2_1 _15878_ (.Y(_06474_),
    .A(net2621),
    .B(net4994));
 sg13g2_o21ai_1 _15879_ (.B1(_06474_),
    .Y(_00950_),
    .A1(net5478),
    .A2(net4994));
 sg13g2_nand2_1 _15880_ (.Y(_06475_),
    .A(net2958),
    .B(net4993));
 sg13g2_o21ai_1 _15881_ (.B1(_06475_),
    .Y(_00951_),
    .A1(net5526),
    .A2(net4994));
 sg13g2_nand2_1 _15882_ (.Y(_06476_),
    .A(net2537),
    .B(net4994));
 sg13g2_o21ai_1 _15883_ (.B1(_06476_),
    .Y(_00952_),
    .A1(net5567),
    .A2(net4994));
 sg13g2_nand2_1 _15884_ (.Y(_06477_),
    .A(net3204),
    .B(net4993));
 sg13g2_o21ai_1 _15885_ (.B1(_06477_),
    .Y(_00953_),
    .A1(net5616),
    .A2(net4993));
 sg13g2_nand2_1 _15886_ (.Y(_06478_),
    .A(net2740),
    .B(net4994));
 sg13g2_o21ai_1 _15887_ (.B1(_06478_),
    .Y(_00954_),
    .A1(net5657),
    .A2(net4994));
 sg13g2_nand2_1 _15888_ (.Y(_06479_),
    .A(net3340),
    .B(net4993));
 sg13g2_o21ai_1 _15889_ (.B1(_06479_),
    .Y(_00955_),
    .A1(net5708),
    .A2(net4993));
 sg13g2_nand2_1 _15890_ (.Y(_06480_),
    .A(net3182),
    .B(_06472_));
 sg13g2_o21ai_1 _15891_ (.B1(_06480_),
    .Y(_00956_),
    .A1(net5754),
    .A2(net4993));
 sg13g2_nand2_1 _15892_ (.Y(_06481_),
    .A(net5243),
    .B(net5215));
 sg13g2_nand2_1 _15893_ (.Y(_06482_),
    .A(net3739),
    .B(net4991));
 sg13g2_o21ai_1 _15894_ (.B1(_06482_),
    .Y(_00957_),
    .A1(net5432),
    .A2(net4991));
 sg13g2_nand2_1 _15895_ (.Y(_06483_),
    .A(net3060),
    .B(net4991));
 sg13g2_o21ai_1 _15896_ (.B1(_06483_),
    .Y(_00958_),
    .A1(net5478),
    .A2(net4991));
 sg13g2_nand2_1 _15897_ (.Y(_06484_),
    .A(net2759),
    .B(net4992));
 sg13g2_o21ai_1 _15898_ (.B1(_06484_),
    .Y(_00959_),
    .A1(net5526),
    .A2(net4992));
 sg13g2_nand2_1 _15899_ (.Y(_06485_),
    .A(net2425),
    .B(net4991));
 sg13g2_o21ai_1 _15900_ (.B1(_06485_),
    .Y(_00960_),
    .A1(net5567),
    .A2(net4991));
 sg13g2_nand2_1 _15901_ (.Y(_06486_),
    .A(net3599),
    .B(net4992));
 sg13g2_o21ai_1 _15902_ (.B1(_06486_),
    .Y(_00961_),
    .A1(net5616),
    .A2(net4992));
 sg13g2_nand2_1 _15903_ (.Y(_06487_),
    .A(net2653),
    .B(net4991));
 sg13g2_o21ai_1 _15904_ (.B1(_06487_),
    .Y(_00962_),
    .A1(net5657),
    .A2(net4991));
 sg13g2_nand2_1 _15905_ (.Y(_06488_),
    .A(net3203),
    .B(net4992));
 sg13g2_o21ai_1 _15906_ (.B1(_06488_),
    .Y(_00963_),
    .A1(net5708),
    .A2(net4992));
 sg13g2_nand2_1 _15907_ (.Y(_06489_),
    .A(net3256),
    .B(net4992));
 sg13g2_o21ai_1 _15908_ (.B1(_06489_),
    .Y(_00964_),
    .A1(net5754),
    .A2(net4992));
 sg13g2_nand2_1 _15909_ (.Y(_06490_),
    .A(net5216),
    .B(net5245));
 sg13g2_nand2_1 _15910_ (.Y(_06491_),
    .A(net2261),
    .B(net4990));
 sg13g2_o21ai_1 _15911_ (.B1(_06491_),
    .Y(_00965_),
    .A1(net5436),
    .A2(net4990));
 sg13g2_nand2_1 _15912_ (.Y(_06492_),
    .A(net2231),
    .B(net4989));
 sg13g2_o21ai_1 _15913_ (.B1(_06492_),
    .Y(_00966_),
    .A1(net5477),
    .A2(net4989));
 sg13g2_nand2_1 _15914_ (.Y(_06493_),
    .A(net2440),
    .B(net4990));
 sg13g2_o21ai_1 _15915_ (.B1(_06493_),
    .Y(_00967_),
    .A1(net5526),
    .A2(net4990));
 sg13g2_nand2_1 _15916_ (.Y(_06494_),
    .A(net3263),
    .B(net4989));
 sg13g2_o21ai_1 _15917_ (.B1(_06494_),
    .Y(_00968_),
    .A1(net5571),
    .A2(net4989));
 sg13g2_nand2_1 _15918_ (.Y(_06495_),
    .A(net2522),
    .B(net4989));
 sg13g2_o21ai_1 _15919_ (.B1(_06495_),
    .Y(_00969_),
    .A1(net5618),
    .A2(net4989));
 sg13g2_nand2_1 _15920_ (.Y(_06496_),
    .A(net3061),
    .B(net4989));
 sg13g2_o21ai_1 _15921_ (.B1(_06496_),
    .Y(_00970_),
    .A1(net5659),
    .A2(net4989));
 sg13g2_nand2_1 _15922_ (.Y(_06497_),
    .A(net2209),
    .B(net4990));
 sg13g2_o21ai_1 _15923_ (.B1(_06497_),
    .Y(_00971_),
    .A1(net5708),
    .A2(net4990));
 sg13g2_nand2_1 _15924_ (.Y(_06498_),
    .A(net2227),
    .B(net4990));
 sg13g2_o21ai_1 _15925_ (.B1(_06498_),
    .Y(_00972_),
    .A1(net5754),
    .A2(net4990));
 sg13g2_nor2_1 _15926_ (.A(_02981_),
    .B(net5142),
    .Y(_06499_));
 sg13g2_nor2_1 _15927_ (.A(net4070),
    .B(net4745),
    .Y(_06500_));
 sg13g2_a21oi_1 _15928_ (.A1(net5453),
    .A2(net4745),
    .Y(_00973_),
    .B1(_06500_));
 sg13g2_nor2_1 _15929_ (.A(net3766),
    .B(net4744),
    .Y(_06501_));
 sg13g2_a21oi_1 _15930_ (.A1(net5492),
    .A2(net4744),
    .Y(_00974_),
    .B1(_06501_));
 sg13g2_nor2_1 _15931_ (.A(net3750),
    .B(net4745),
    .Y(_06502_));
 sg13g2_a21oi_1 _15932_ (.A1(net5543),
    .A2(net4745),
    .Y(_00975_),
    .B1(_06502_));
 sg13g2_nor2_1 _15933_ (.A(net3915),
    .B(net4744),
    .Y(_06503_));
 sg13g2_a21oi_1 _15934_ (.A1(net5581),
    .A2(net4744),
    .Y(_00976_),
    .B1(_06503_));
 sg13g2_nor2_1 _15935_ (.A(net3825),
    .B(net4745),
    .Y(_06504_));
 sg13g2_a21oi_1 _15936_ (.A1(net5628),
    .A2(net4745),
    .Y(_00977_),
    .B1(_06504_));
 sg13g2_nor2_1 _15937_ (.A(net4107),
    .B(net4744),
    .Y(_06505_));
 sg13g2_a21oi_1 _15938_ (.A1(net5671),
    .A2(net4744),
    .Y(_00978_),
    .B1(_06505_));
 sg13g2_nor2_1 _15939_ (.A(net3602),
    .B(net4744),
    .Y(_06506_));
 sg13g2_a21oi_1 _15940_ (.A1(net5718),
    .A2(net4744),
    .Y(_00979_),
    .B1(_06506_));
 sg13g2_nor2_1 _15941_ (.A(net4081),
    .B(net4745),
    .Y(_06507_));
 sg13g2_a21oi_1 _15942_ (.A1(net5764),
    .A2(net4745),
    .Y(_00980_),
    .B1(_06507_));
 sg13g2_nand2_1 _15943_ (.Y(_06508_),
    .A(net5215),
    .B(net5246));
 sg13g2_nand2_1 _15944_ (.Y(_06509_),
    .A(net2141),
    .B(_06508_));
 sg13g2_o21ai_1 _15945_ (.B1(_06509_),
    .Y(_00981_),
    .A1(net5438),
    .A2(net4988));
 sg13g2_nand2_1 _15946_ (.Y(_06510_),
    .A(net2822),
    .B(net4987));
 sg13g2_o21ai_1 _15947_ (.B1(_06510_),
    .Y(_00982_),
    .A1(net5479),
    .A2(net4987));
 sg13g2_nand2_1 _15948_ (.Y(_06511_),
    .A(net3011),
    .B(net4988));
 sg13g2_o21ai_1 _15949_ (.B1(_06511_),
    .Y(_00983_),
    .A1(net5526),
    .A2(net4988));
 sg13g2_nand2_1 _15950_ (.Y(_06512_),
    .A(net2178),
    .B(net4987));
 sg13g2_o21ai_1 _15951_ (.B1(_06512_),
    .Y(_00984_),
    .A1(net5572),
    .A2(net4987));
 sg13g2_nand2_1 _15952_ (.Y(_06513_),
    .A(net3276),
    .B(net4987));
 sg13g2_o21ai_1 _15953_ (.B1(_06513_),
    .Y(_00985_),
    .A1(net5617),
    .A2(net4987));
 sg13g2_nand2_1 _15954_ (.Y(_06514_),
    .A(net2735),
    .B(net4988));
 sg13g2_o21ai_1 _15955_ (.B1(_06514_),
    .Y(_00986_),
    .A1(net5659),
    .A2(net4988));
 sg13g2_nand2_1 _15956_ (.Y(_06515_),
    .A(net2727),
    .B(net4987));
 sg13g2_o21ai_1 _15957_ (.B1(_06515_),
    .Y(_00987_),
    .A1(net5708),
    .A2(net4987));
 sg13g2_nand2_1 _15958_ (.Y(_06516_),
    .A(net3126),
    .B(net4988));
 sg13g2_o21ai_1 _15959_ (.B1(_06516_),
    .Y(_00988_),
    .A1(net5754),
    .A2(net4988));
 sg13g2_nor3_1 _15960_ (.A(net5259),
    .B(net5227),
    .C(net5241),
    .Y(_06517_));
 sg13g2_nor2_1 _15961_ (.A(net4142),
    .B(net5185),
    .Y(_06518_));
 sg13g2_a21oi_1 _15962_ (.A1(net5438),
    .A2(_06517_),
    .Y(_00989_),
    .B1(_06518_));
 sg13g2_nor2_1 _15963_ (.A(net3473),
    .B(net5184),
    .Y(_06519_));
 sg13g2_a21oi_1 _15964_ (.A1(net5477),
    .A2(net5184),
    .Y(_00990_),
    .B1(_06519_));
 sg13g2_nor2_1 _15965_ (.A(net3840),
    .B(net5185),
    .Y(_06520_));
 sg13g2_a21oi_1 _15966_ (.A1(net5526),
    .A2(net5185),
    .Y(_00991_),
    .B1(_06520_));
 sg13g2_nor2_1 _15967_ (.A(net3462),
    .B(net5184),
    .Y(_06521_));
 sg13g2_a21oi_1 _15968_ (.A1(net5572),
    .A2(net5184),
    .Y(_00992_),
    .B1(_06521_));
 sg13g2_nor2_1 _15969_ (.A(net4086),
    .B(net5184),
    .Y(_06522_));
 sg13g2_a21oi_1 _15970_ (.A1(net5617),
    .A2(net5184),
    .Y(_00993_),
    .B1(_06522_));
 sg13g2_nor2_1 _15971_ (.A(net3721),
    .B(net5185),
    .Y(_06523_));
 sg13g2_a21oi_1 _15972_ (.A1(net5659),
    .A2(net5185),
    .Y(_00994_),
    .B1(_06523_));
 sg13g2_nor2_1 _15973_ (.A(net3633),
    .B(net5184),
    .Y(_06524_));
 sg13g2_a21oi_1 _15974_ (.A1(net5708),
    .A2(net5184),
    .Y(_00995_),
    .B1(_06524_));
 sg13g2_nor2_1 _15975_ (.A(net3478),
    .B(net5185),
    .Y(_06525_));
 sg13g2_a21oi_1 _15976_ (.A1(net5754),
    .A2(net5185),
    .Y(_00996_),
    .B1(_06525_));
 sg13g2_nand2_1 _15977_ (.Y(_06526_),
    .A(net5213),
    .B(net5248));
 sg13g2_nand2_1 _15978_ (.Y(_06527_),
    .A(net2473),
    .B(net4986));
 sg13g2_o21ai_1 _15979_ (.B1(_06527_),
    .Y(_00997_),
    .A1(net5434),
    .A2(net4986));
 sg13g2_nand2_1 _15980_ (.Y(_06528_),
    .A(net2383),
    .B(net4985));
 sg13g2_o21ai_1 _15981_ (.B1(_06528_),
    .Y(_00998_),
    .A1(net5476),
    .A2(net4985));
 sg13g2_nand2_1 _15982_ (.Y(_06529_),
    .A(net3397),
    .B(net4986));
 sg13g2_o21ai_1 _15983_ (.B1(_06529_),
    .Y(_00999_),
    .A1(net5531),
    .A2(net4986));
 sg13g2_nand2_1 _15984_ (.Y(_06530_),
    .A(net2406),
    .B(net4985));
 sg13g2_o21ai_1 _15985_ (.B1(_06530_),
    .Y(_01000_),
    .A1(net5564),
    .A2(net4985));
 sg13g2_nand2_1 _15986_ (.Y(_06531_),
    .A(net2532),
    .B(_06526_));
 sg13g2_o21ai_1 _15987_ (.B1(_06531_),
    .Y(_01001_),
    .A1(net5614),
    .A2(net4986));
 sg13g2_nand2_1 _15988_ (.Y(_06532_),
    .A(net2708),
    .B(net4985));
 sg13g2_o21ai_1 _15989_ (.B1(_06532_),
    .Y(_01002_),
    .A1(net5658),
    .A2(net4985));
 sg13g2_nand2_1 _15990_ (.Y(_06533_),
    .A(net3480),
    .B(net4986));
 sg13g2_o21ai_1 _15991_ (.B1(_06533_),
    .Y(_01003_),
    .A1(net5704),
    .A2(net4986));
 sg13g2_nand2_1 _15992_ (.Y(_06534_),
    .A(net2257),
    .B(net4985));
 sg13g2_o21ai_1 _15993_ (.B1(_06534_),
    .Y(_01004_),
    .A1(net5745),
    .A2(net4985));
 sg13g2_nand2_1 _15994_ (.Y(_06535_),
    .A(_03139_),
    .B(net5213));
 sg13g2_nand2_1 _15995_ (.Y(_06536_),
    .A(net3157),
    .B(net4984));
 sg13g2_o21ai_1 _15996_ (.B1(_06536_),
    .Y(_01005_),
    .A1(net5434),
    .A2(net4984));
 sg13g2_nand2_1 _15997_ (.Y(_06537_),
    .A(net2828),
    .B(net4983));
 sg13g2_o21ai_1 _15998_ (.B1(_06537_),
    .Y(_01006_),
    .A1(net5476),
    .A2(net4983));
 sg13g2_nand2_1 _15999_ (.Y(_06538_),
    .A(net2907),
    .B(net4984));
 sg13g2_o21ai_1 _16000_ (.B1(_06538_),
    .Y(_01007_),
    .A1(net5531),
    .A2(net4984));
 sg13g2_nand2_1 _16001_ (.Y(_06539_),
    .A(net2414),
    .B(net4983));
 sg13g2_o21ai_1 _16002_ (.B1(_06539_),
    .Y(_01008_),
    .A1(net5564),
    .A2(net4983));
 sg13g2_nand2_1 _16003_ (.Y(_06540_),
    .A(net3177),
    .B(_06535_));
 sg13g2_o21ai_1 _16004_ (.B1(_06540_),
    .Y(_01009_),
    .A1(net5614),
    .A2(net4984));
 sg13g2_nand2_1 _16005_ (.Y(_06541_),
    .A(net2431),
    .B(net4983));
 sg13g2_o21ai_1 _16006_ (.B1(_06541_),
    .Y(_01010_),
    .A1(net5658),
    .A2(net4983));
 sg13g2_nand2_1 _16007_ (.Y(_06542_),
    .A(net3336),
    .B(net4984));
 sg13g2_o21ai_1 _16008_ (.B1(_06542_),
    .Y(_01011_),
    .A1(net5704),
    .A2(net4984));
 sg13g2_nand2_1 _16009_ (.Y(_06543_),
    .A(net2602),
    .B(net4983));
 sg13g2_o21ai_1 _16010_ (.B1(_06543_),
    .Y(_01012_),
    .A1(net5745),
    .A2(net4983));
 sg13g2_nand2_1 _16011_ (.Y(_06544_),
    .A(_03079_),
    .B(net5213));
 sg13g2_nand2_1 _16012_ (.Y(_06545_),
    .A(net2176),
    .B(net4982));
 sg13g2_o21ai_1 _16013_ (.B1(_06545_),
    .Y(_01013_),
    .A1(net5434),
    .A2(net4982));
 sg13g2_nand2_1 _16014_ (.Y(_06546_),
    .A(net3019),
    .B(net4981));
 sg13g2_o21ai_1 _16015_ (.B1(_06546_),
    .Y(_01014_),
    .A1(net5475),
    .A2(net4981));
 sg13g2_nand2_1 _16016_ (.Y(_06547_),
    .A(net2348),
    .B(net4982));
 sg13g2_o21ai_1 _16017_ (.B1(_06547_),
    .Y(_01015_),
    .A1(net5519),
    .A2(net4982));
 sg13g2_nand2_1 _16018_ (.Y(_06548_),
    .A(net2210),
    .B(net4981));
 sg13g2_o21ai_1 _16019_ (.B1(_06548_),
    .Y(_01016_),
    .A1(net5564),
    .A2(net4981));
 sg13g2_nand2_1 _16020_ (.Y(_06549_),
    .A(net2447),
    .B(net4982));
 sg13g2_o21ai_1 _16021_ (.B1(_06549_),
    .Y(_01017_),
    .A1(net5614),
    .A2(net4982));
 sg13g2_nand2_1 _16022_ (.Y(_06550_),
    .A(net2620),
    .B(net4981));
 sg13g2_o21ai_1 _16023_ (.B1(_06550_),
    .Y(_01018_),
    .A1(net5658),
    .A2(net4981));
 sg13g2_nand2_1 _16024_ (.Y(_06551_),
    .A(net2495),
    .B(net4982));
 sg13g2_o21ai_1 _16025_ (.B1(_06551_),
    .Y(_01019_),
    .A1(net5704),
    .A2(net4982));
 sg13g2_nand2_1 _16026_ (.Y(_06552_),
    .A(net2773),
    .B(net4981));
 sg13g2_o21ai_1 _16027_ (.B1(_06552_),
    .Y(_01020_),
    .A1(net5749),
    .A2(net4981));
 sg13g2_nand2_2 _16028_ (.Y(_06553_),
    .A(net5253),
    .B(net5213));
 sg13g2_nand2_1 _16029_ (.Y(_06554_),
    .A(net2533),
    .B(net4980));
 sg13g2_o21ai_1 _16030_ (.B1(_06554_),
    .Y(_01021_),
    .A1(net5434),
    .A2(net4980));
 sg13g2_nand2_1 _16031_ (.Y(_06555_),
    .A(net2584),
    .B(net4979));
 sg13g2_o21ai_1 _16032_ (.B1(_06555_),
    .Y(_01022_),
    .A1(net5475),
    .A2(net4979));
 sg13g2_nand2_1 _16033_ (.Y(_06556_),
    .A(net2723),
    .B(net4980));
 sg13g2_o21ai_1 _16034_ (.B1(_06556_),
    .Y(_01023_),
    .A1(net5519),
    .A2(net4980));
 sg13g2_nand2_1 _16035_ (.Y(_06557_),
    .A(net3111),
    .B(net4979));
 sg13g2_o21ai_1 _16036_ (.B1(_06557_),
    .Y(_01024_),
    .A1(net5564),
    .A2(net4979));
 sg13g2_nand2_1 _16037_ (.Y(_06558_),
    .A(net2695),
    .B(net4980));
 sg13g2_o21ai_1 _16038_ (.B1(_06558_),
    .Y(_01025_),
    .A1(net5616),
    .A2(net4980));
 sg13g2_nand2_1 _16039_ (.Y(_06559_),
    .A(net2863),
    .B(net4979));
 sg13g2_o21ai_1 _16040_ (.B1(_06559_),
    .Y(_01026_),
    .A1(net5658),
    .A2(net4979));
 sg13g2_nand2_1 _16041_ (.Y(_06560_),
    .A(net3044),
    .B(net4980));
 sg13g2_o21ai_1 _16042_ (.B1(_06560_),
    .Y(_01027_),
    .A1(net5704),
    .A2(net4980));
 sg13g2_nand2_1 _16043_ (.Y(_06561_),
    .A(net2760),
    .B(net4979));
 sg13g2_o21ai_1 _16044_ (.B1(_06561_),
    .Y(_01028_),
    .A1(net5749),
    .A2(net4979));
 sg13g2_nand2_1 _16045_ (.Y(_06562_),
    .A(net5235),
    .B(net5213));
 sg13g2_nand2_1 _16046_ (.Y(_06563_),
    .A(net2200),
    .B(net4978));
 sg13g2_o21ai_1 _16047_ (.B1(_06563_),
    .Y(_01029_),
    .A1(net5434),
    .A2(net4977));
 sg13g2_nand2_1 _16048_ (.Y(_06564_),
    .A(net3523),
    .B(net4977));
 sg13g2_o21ai_1 _16049_ (.B1(_06564_),
    .Y(_01030_),
    .A1(net5481),
    .A2(net4977));
 sg13g2_nand2_1 _16050_ (.Y(_06565_),
    .A(net2497),
    .B(net4978));
 sg13g2_o21ai_1 _16051_ (.B1(_06565_),
    .Y(_01031_),
    .A1(net5518),
    .A2(net4978));
 sg13g2_nand2_1 _16052_ (.Y(_06566_),
    .A(net2411),
    .B(net4978));
 sg13g2_o21ai_1 _16053_ (.B1(_06566_),
    .Y(_01032_),
    .A1(net5565),
    .A2(net4978));
 sg13g2_nand2_1 _16054_ (.Y(_06567_),
    .A(net2950),
    .B(net4977));
 sg13g2_o21ai_1 _16055_ (.B1(_06567_),
    .Y(_01033_),
    .A1(net5614),
    .A2(net4978));
 sg13g2_nand2_1 _16056_ (.Y(_06568_),
    .A(net2904),
    .B(net4978));
 sg13g2_o21ai_1 _16057_ (.B1(_06568_),
    .Y(_01034_),
    .A1(net5654),
    .A2(net4978));
 sg13g2_nand2_1 _16058_ (.Y(_06569_),
    .A(net2796),
    .B(net4977));
 sg13g2_o21ai_1 _16059_ (.B1(_06569_),
    .Y(_01035_),
    .A1(net5704),
    .A2(net4977));
 sg13g2_nand2_1 _16060_ (.Y(_06570_),
    .A(net3315),
    .B(net4977));
 sg13g2_o21ai_1 _16061_ (.B1(_06570_),
    .Y(_01036_),
    .A1(net5751),
    .A2(net4977));
 sg13g2_nand2_1 _16062_ (.Y(_06571_),
    .A(net5234),
    .B(net5213));
 sg13g2_nand2_1 _16063_ (.Y(_06572_),
    .A(net3406),
    .B(_06571_));
 sg13g2_o21ai_1 _16064_ (.B1(_06572_),
    .Y(_01037_),
    .A1(net5434),
    .A2(net4976));
 sg13g2_nand2_1 _16065_ (.Y(_06573_),
    .A(net2911),
    .B(net4975));
 sg13g2_o21ai_1 _16066_ (.B1(_06573_),
    .Y(_01038_),
    .A1(net5480),
    .A2(net4975));
 sg13g2_nand2_1 _16067_ (.Y(_06574_),
    .A(net2957),
    .B(net4976));
 sg13g2_o21ai_1 _16068_ (.B1(_06574_),
    .Y(_01039_),
    .A1(net5518),
    .A2(net4976));
 sg13g2_nand2_1 _16069_ (.Y(_06575_),
    .A(net3073),
    .B(net4976));
 sg13g2_o21ai_1 _16070_ (.B1(_06575_),
    .Y(_01040_),
    .A1(net5564),
    .A2(net4976));
 sg13g2_nand2_1 _16071_ (.Y(_06576_),
    .A(net2635),
    .B(net4975));
 sg13g2_o21ai_1 _16072_ (.B1(_06576_),
    .Y(_01041_),
    .A1(net5614),
    .A2(net4975));
 sg13g2_nand2_1 _16073_ (.Y(_06577_),
    .A(net3187),
    .B(net4976));
 sg13g2_o21ai_1 _16074_ (.B1(_06577_),
    .Y(_01042_),
    .A1(net5654),
    .A2(net4976));
 sg13g2_nand2_1 _16075_ (.Y(_06578_),
    .A(net2443),
    .B(net4975));
 sg13g2_o21ai_1 _16076_ (.B1(_06578_),
    .Y(_01043_),
    .A1(net5704),
    .A2(net4975));
 sg13g2_nand2_1 _16077_ (.Y(_06579_),
    .A(net2690),
    .B(net4975));
 sg13g2_o21ai_1 _16078_ (.B1(_06579_),
    .Y(_01044_),
    .A1(net5751),
    .A2(net4975));
 sg13g2_nand2_1 _16079_ (.Y(_06580_),
    .A(net5236),
    .B(net5213));
 sg13g2_nor2_1 _16080_ (.A(\mem.data_in[0] ),
    .B(net4973),
    .Y(_06581_));
 sg13g2_a21oi_1 _16081_ (.A1(_02887_),
    .A2(net4973),
    .Y(_01045_),
    .B1(_06581_));
 sg13g2_nand2_1 _16082_ (.Y(_06582_),
    .A(net3145),
    .B(net4973));
 sg13g2_o21ai_1 _16083_ (.B1(_06582_),
    .Y(_01046_),
    .A1(net5480),
    .A2(net4973));
 sg13g2_nand2_1 _16084_ (.Y(_06583_),
    .A(net2300),
    .B(net4974));
 sg13g2_o21ai_1 _16085_ (.B1(_06583_),
    .Y(_01047_),
    .A1(net5518),
    .A2(net4974));
 sg13g2_nand2_1 _16086_ (.Y(_06584_),
    .A(net2482),
    .B(net4974));
 sg13g2_o21ai_1 _16087_ (.B1(_06584_),
    .Y(_01048_),
    .A1(net5564),
    .A2(net4974));
 sg13g2_nand2_1 _16088_ (.Y(_06585_),
    .A(net2594),
    .B(net4973));
 sg13g2_o21ai_1 _16089_ (.B1(_06585_),
    .Y(_01049_),
    .A1(net5614),
    .A2(net4973));
 sg13g2_nand2_1 _16090_ (.Y(_06586_),
    .A(net2994),
    .B(net4974));
 sg13g2_o21ai_1 _16091_ (.B1(_06586_),
    .Y(_01050_),
    .A1(net5654),
    .A2(net4974));
 sg13g2_nand2_1 _16092_ (.Y(_06587_),
    .A(net2682),
    .B(net4973));
 sg13g2_o21ai_1 _16093_ (.B1(_06587_),
    .Y(_01051_),
    .A1(net5704),
    .A2(net4973));
 sg13g2_nand2_1 _16094_ (.Y(_06588_),
    .A(net2940),
    .B(_06580_));
 sg13g2_o21ai_1 _16095_ (.B1(_06588_),
    .Y(_01052_),
    .A1(net5751),
    .A2(net4974));
 sg13g2_nor2_1 _16096_ (.A(_02964_),
    .B(net5143),
    .Y(_06589_));
 sg13g2_nor2_1 _16097_ (.A(net3632),
    .B(net4742),
    .Y(_06590_));
 sg13g2_a21oi_1 _16098_ (.A1(net5448),
    .A2(net4742),
    .Y(_01053_),
    .B1(_06590_));
 sg13g2_nor2_1 _16099_ (.A(net3634),
    .B(net4743),
    .Y(_06591_));
 sg13g2_a21oi_1 _16100_ (.A1(net5492),
    .A2(net4743),
    .Y(_01054_),
    .B1(_06591_));
 sg13g2_nor2_1 _16101_ (.A(net4180),
    .B(net4743),
    .Y(_06592_));
 sg13g2_a21oi_1 _16102_ (.A1(net5543),
    .A2(_06589_),
    .Y(_01055_),
    .B1(_06592_));
 sg13g2_nor2_1 _16103_ (.A(net3559),
    .B(net4742),
    .Y(_06593_));
 sg13g2_a21oi_1 _16104_ (.A1(net5581),
    .A2(net4742),
    .Y(_01056_),
    .B1(_06593_));
 sg13g2_nor2_1 _16105_ (.A(net3720),
    .B(net4742),
    .Y(_06594_));
 sg13g2_a21oi_1 _16106_ (.A1(net5628),
    .A2(net4742),
    .Y(_01057_),
    .B1(_06594_));
 sg13g2_nor2_1 _16107_ (.A(net3793),
    .B(net4743),
    .Y(_06595_));
 sg13g2_a21oi_1 _16108_ (.A1(net5671),
    .A2(net4743),
    .Y(_01058_),
    .B1(_06595_));
 sg13g2_nor2_1 _16109_ (.A(net4144),
    .B(net4743),
    .Y(_06596_));
 sg13g2_a21oi_1 _16110_ (.A1(net5717),
    .A2(net4743),
    .Y(_01059_),
    .B1(_06596_));
 sg13g2_nor2_1 _16111_ (.A(net3671),
    .B(net4742),
    .Y(_06597_));
 sg13g2_a21oi_1 _16112_ (.A1(net5764),
    .A2(net4742),
    .Y(_01060_),
    .B1(_06597_));
 sg13g2_nand2_1 _16113_ (.Y(_06598_),
    .A(net5244),
    .B(net5214));
 sg13g2_nand2_1 _16114_ (.Y(_06599_),
    .A(net2391),
    .B(net4971));
 sg13g2_o21ai_1 _16115_ (.B1(_06599_),
    .Y(_01061_),
    .A1(net5435),
    .A2(net4971));
 sg13g2_nand2_1 _16116_ (.Y(_06600_),
    .A(net3100),
    .B(net4971));
 sg13g2_o21ai_1 _16117_ (.B1(_06600_),
    .Y(_01062_),
    .A1(net5481),
    .A2(net4972));
 sg13g2_nand2_1 _16118_ (.Y(_06601_),
    .A(net3231),
    .B(net4972));
 sg13g2_o21ai_1 _16119_ (.B1(_06601_),
    .Y(_01063_),
    .A1(net5525),
    .A2(net4972));
 sg13g2_nand2_1 _16120_ (.Y(_06602_),
    .A(net3245),
    .B(net4971));
 sg13g2_o21ai_1 _16121_ (.B1(_06602_),
    .Y(_01064_),
    .A1(net5570),
    .A2(net4971));
 sg13g2_nand2_1 _16122_ (.Y(_06603_),
    .A(net2902),
    .B(net4972));
 sg13g2_o21ai_1 _16123_ (.B1(_06603_),
    .Y(_01065_),
    .A1(net5615),
    .A2(_06598_));
 sg13g2_nand2_1 _16124_ (.Y(_06604_),
    .A(net2804),
    .B(net4971));
 sg13g2_o21ai_1 _16125_ (.B1(_06604_),
    .Y(_01066_),
    .A1(net5662),
    .A2(net4971));
 sg13g2_nand2_1 _16126_ (.Y(_06605_),
    .A(net2274),
    .B(net4971));
 sg13g2_o21ai_1 _16127_ (.B1(_06605_),
    .Y(_01067_),
    .A1(net5705),
    .A2(net4972));
 sg13g2_nand2_1 _16128_ (.Y(_06606_),
    .A(net2730),
    .B(net4972));
 sg13g2_o21ai_1 _16129_ (.B1(_06606_),
    .Y(_01068_),
    .A1(net5750),
    .A2(net4972));
 sg13g2_nand2_1 _16130_ (.Y(_06607_),
    .A(net5239),
    .B(net5214));
 sg13g2_nand2_1 _16131_ (.Y(_06608_),
    .A(net2636),
    .B(net4969));
 sg13g2_o21ai_1 _16132_ (.B1(_06608_),
    .Y(_01069_),
    .A1(net5434),
    .A2(net4969));
 sg13g2_nand2_1 _16133_ (.Y(_06609_),
    .A(net3020),
    .B(net4970));
 sg13g2_o21ai_1 _16134_ (.B1(_06609_),
    .Y(_01070_),
    .A1(net5481),
    .A2(net4970));
 sg13g2_nand2_1 _16135_ (.Y(_06610_),
    .A(net2678),
    .B(net4970));
 sg13g2_o21ai_1 _16136_ (.B1(_06610_),
    .Y(_01071_),
    .A1(net5525),
    .A2(net4970));
 sg13g2_nand2_1 _16137_ (.Y(_06611_),
    .A(net2295),
    .B(net4969));
 sg13g2_o21ai_1 _16138_ (.B1(_06611_),
    .Y(_01072_),
    .A1(net5570),
    .A2(net4969));
 sg13g2_nand2_1 _16139_ (.Y(_06612_),
    .A(net2948),
    .B(_06607_));
 sg13g2_o21ai_1 _16140_ (.B1(_06612_),
    .Y(_01073_),
    .A1(net5615),
    .A2(net4970));
 sg13g2_nand2_1 _16141_ (.Y(_06613_),
    .A(net3123),
    .B(net4969));
 sg13g2_o21ai_1 _16142_ (.B1(_06613_),
    .Y(_01074_),
    .A1(net5662),
    .A2(net4969));
 sg13g2_nand2_1 _16143_ (.Y(_06614_),
    .A(net3243),
    .B(net4969));
 sg13g2_o21ai_1 _16144_ (.B1(_06614_),
    .Y(_01075_),
    .A1(net5707),
    .A2(net4969));
 sg13g2_nand2_1 _16145_ (.Y(_06615_),
    .A(net2638),
    .B(net4970));
 sg13g2_o21ai_1 _16146_ (.B1(_06615_),
    .Y(_01076_),
    .A1(net5751),
    .A2(net4970));
 sg13g2_nand2_1 _16147_ (.Y(_06616_),
    .A(net5242),
    .B(net5214));
 sg13g2_nand2_1 _16148_ (.Y(_06617_),
    .A(net3099),
    .B(net4967));
 sg13g2_o21ai_1 _16149_ (.B1(_06617_),
    .Y(_01077_),
    .A1(net5435),
    .A2(net4967));
 sg13g2_nand2_1 _16150_ (.Y(_06618_),
    .A(net3377),
    .B(net4968));
 sg13g2_o21ai_1 _16151_ (.B1(_06618_),
    .Y(_01078_),
    .A1(net5481),
    .A2(net4968));
 sg13g2_nand2_1 _16152_ (.Y(_06619_),
    .A(net2717),
    .B(net4968));
 sg13g2_o21ai_1 _16153_ (.B1(_06619_),
    .Y(_01079_),
    .A1(net5524),
    .A2(net4968));
 sg13g2_nand2_1 _16154_ (.Y(_06620_),
    .A(net2919),
    .B(net4967));
 sg13g2_o21ai_1 _16155_ (.B1(_06620_),
    .Y(_01080_),
    .A1(net5570),
    .A2(net4967));
 sg13g2_nand2_1 _16156_ (.Y(_06621_),
    .A(net2217),
    .B(net4968));
 sg13g2_o21ai_1 _16157_ (.B1(_06621_),
    .Y(_01081_),
    .A1(net5615),
    .A2(_06616_));
 sg13g2_nand2_1 _16158_ (.Y(_06622_),
    .A(net2239),
    .B(net4967));
 sg13g2_o21ai_1 _16159_ (.B1(_06622_),
    .Y(_01082_),
    .A1(net5661),
    .A2(net4967));
 sg13g2_nand2_1 _16160_ (.Y(_06623_),
    .A(net2939),
    .B(net4967));
 sg13g2_o21ai_1 _16161_ (.B1(_06623_),
    .Y(_01083_),
    .A1(net5705),
    .A2(net4967));
 sg13g2_nand2_1 _16162_ (.Y(_06624_),
    .A(net2203),
    .B(net4968));
 sg13g2_o21ai_1 _16163_ (.B1(_06624_),
    .Y(_01084_),
    .A1(net5751),
    .A2(net4968));
 sg13g2_nand2_1 _16164_ (.Y(_06625_),
    .A(net5243),
    .B(net5214));
 sg13g2_nand2_1 _16165_ (.Y(_06626_),
    .A(net2499),
    .B(net4965));
 sg13g2_o21ai_1 _16166_ (.B1(_06626_),
    .Y(_01085_),
    .A1(net5435),
    .A2(net4965));
 sg13g2_nand2_1 _16167_ (.Y(_06627_),
    .A(net2536),
    .B(net4966));
 sg13g2_o21ai_1 _16168_ (.B1(_06627_),
    .Y(_01086_),
    .A1(net5480),
    .A2(net4966));
 sg13g2_nand2_1 _16169_ (.Y(_06628_),
    .A(net3175),
    .B(net4965));
 sg13g2_o21ai_1 _16170_ (.B1(_06628_),
    .Y(_01087_),
    .A1(net5525),
    .A2(net4965));
 sg13g2_nand2_1 _16171_ (.Y(_06629_),
    .A(net2279),
    .B(net4966));
 sg13g2_o21ai_1 _16172_ (.B1(_06629_),
    .Y(_01088_),
    .A1(net5570),
    .A2(net4966));
 sg13g2_nand2_1 _16173_ (.Y(_06630_),
    .A(net2943),
    .B(_06625_));
 sg13g2_o21ai_1 _16174_ (.B1(_06630_),
    .Y(_01089_),
    .A1(net5615),
    .A2(net4966));
 sg13g2_nand2_1 _16175_ (.Y(_06631_),
    .A(net2631),
    .B(net4966));
 sg13g2_o21ai_1 _16176_ (.B1(_06631_),
    .Y(_01090_),
    .A1(net5662),
    .A2(net4966));
 sg13g2_nand2_1 _16177_ (.Y(_06632_),
    .A(net2560),
    .B(net4965));
 sg13g2_o21ai_1 _16178_ (.B1(_06632_),
    .Y(_01091_),
    .A1(net5705),
    .A2(net4965));
 sg13g2_nand2_1 _16179_ (.Y(_06633_),
    .A(net3055),
    .B(net4965));
 sg13g2_o21ai_1 _16180_ (.B1(_06633_),
    .Y(_01092_),
    .A1(net5750),
    .A2(net4965));
 sg13g2_nand2_1 _16181_ (.Y(_06634_),
    .A(net5214),
    .B(net5245));
 sg13g2_nand2_1 _16182_ (.Y(_06635_),
    .A(net2962),
    .B(net4963));
 sg13g2_o21ai_1 _16183_ (.B1(_06635_),
    .Y(_01093_),
    .A1(net5435),
    .A2(net4963));
 sg13g2_nand2_1 _16184_ (.Y(_06636_),
    .A(net2747),
    .B(net4964));
 sg13g2_o21ai_1 _16185_ (.B1(_06636_),
    .Y(_01094_),
    .A1(net5480),
    .A2(net4964));
 sg13g2_nand2_1 _16186_ (.Y(_06637_),
    .A(net2539),
    .B(net4962));
 sg13g2_o21ai_1 _16187_ (.B1(_06637_),
    .Y(_01095_),
    .A1(net5524),
    .A2(net4962));
 sg13g2_nand2_1 _16188_ (.Y(_06638_),
    .A(net2246),
    .B(net4964));
 sg13g2_o21ai_1 _16189_ (.B1(_06638_),
    .Y(_01096_),
    .A1(net5569),
    .A2(net4964));
 sg13g2_nand2_1 _16190_ (.Y(_06639_),
    .A(net3031),
    .B(net4963));
 sg13g2_o21ai_1 _16191_ (.B1(_06639_),
    .Y(_01097_),
    .A1(net5615),
    .A2(net4962));
 sg13g2_nand2_1 _16192_ (.Y(_06640_),
    .A(net2504),
    .B(net4962));
 sg13g2_o21ai_1 _16193_ (.B1(_06640_),
    .Y(_01098_),
    .A1(net5661),
    .A2(net4962));
 sg13g2_nand2_1 _16194_ (.Y(_06641_),
    .A(net2237),
    .B(net4962));
 sg13g2_o21ai_1 _16195_ (.B1(_06641_),
    .Y(_01099_),
    .A1(net5705),
    .A2(net4962));
 sg13g2_nand2_1 _16196_ (.Y(_06642_),
    .A(net2637),
    .B(net4963));
 sg13g2_o21ai_1 _16197_ (.B1(_06642_),
    .Y(_01100_),
    .A1(net5750),
    .A2(net4962));
 sg13g2_nand2_1 _16198_ (.Y(_06643_),
    .A(net5251),
    .B(net5214));
 sg13g2_nand2_1 _16199_ (.Y(_06644_),
    .A(net2868),
    .B(net4959));
 sg13g2_o21ai_1 _16200_ (.B1(_06644_),
    .Y(_01101_),
    .A1(net5435),
    .A2(net4959));
 sg13g2_nand2_1 _16201_ (.Y(_06645_),
    .A(net2291),
    .B(net4961));
 sg13g2_o21ai_1 _16202_ (.B1(_06645_),
    .Y(_01102_),
    .A1(net5480),
    .A2(net4961));
 sg13g2_nand2_1 _16203_ (.Y(_06646_),
    .A(net2979),
    .B(net4959));
 sg13g2_o21ai_1 _16204_ (.B1(_06646_),
    .Y(_01103_),
    .A1(net5524),
    .A2(net4959));
 sg13g2_nand2_1 _16205_ (.Y(_06647_),
    .A(net3144),
    .B(net4961));
 sg13g2_o21ai_1 _16206_ (.B1(_06647_),
    .Y(_01104_),
    .A1(net5569),
    .A2(net4961));
 sg13g2_nand2_1 _16207_ (.Y(_06648_),
    .A(net2390),
    .B(net4960));
 sg13g2_o21ai_1 _16208_ (.B1(_06648_),
    .Y(_01105_),
    .A1(net5615),
    .A2(net4959));
 sg13g2_nand2_1 _16209_ (.Y(_06649_),
    .A(net3191),
    .B(net4960));
 sg13g2_o21ai_1 _16210_ (.B1(_06649_),
    .Y(_01106_),
    .A1(net5661),
    .A2(net4959));
 sg13g2_nand2_1 _16211_ (.Y(_06650_),
    .A(net2275),
    .B(net4960));
 sg13g2_o21ai_1 _16212_ (.B1(_06650_),
    .Y(_01107_),
    .A1(net5705),
    .A2(net4960));
 sg13g2_nand2_1 _16213_ (.Y(_06651_),
    .A(net2359),
    .B(net4959));
 sg13g2_o21ai_1 _16214_ (.B1(_06651_),
    .Y(_01108_),
    .A1(net5750),
    .A2(net4959));
 sg13g2_nand2_1 _16215_ (.Y(_06652_),
    .A(net5214),
    .B(net5246));
 sg13g2_nand2_1 _16216_ (.Y(_06653_),
    .A(net3086),
    .B(net4956));
 sg13g2_o21ai_1 _16217_ (.B1(_06653_),
    .Y(_01109_),
    .A1(net5435),
    .A2(net4956));
 sg13g2_nand2_1 _16218_ (.Y(_06654_),
    .A(net2165),
    .B(net4958));
 sg13g2_o21ai_1 _16219_ (.B1(_06654_),
    .Y(_01110_),
    .A1(net5480),
    .A2(net4958));
 sg13g2_nand2_1 _16220_ (.Y(_06655_),
    .A(net2789),
    .B(net4956));
 sg13g2_o21ai_1 _16221_ (.B1(_06655_),
    .Y(_01111_),
    .A1(net5524),
    .A2(net4956));
 sg13g2_nand2_1 _16222_ (.Y(_06656_),
    .A(net3322),
    .B(net4958));
 sg13g2_o21ai_1 _16223_ (.B1(_06656_),
    .Y(_01112_),
    .A1(net5569),
    .A2(net4958));
 sg13g2_nand2_1 _16224_ (.Y(_06657_),
    .A(net3868),
    .B(net4957));
 sg13g2_o21ai_1 _16225_ (.B1(_06657_),
    .Y(_01113_),
    .A1(net5614),
    .A2(net4956));
 sg13g2_nand2_1 _16226_ (.Y(_06658_),
    .A(net3196),
    .B(net4957));
 sg13g2_o21ai_1 _16227_ (.B1(_06658_),
    .Y(_01114_),
    .A1(net5664),
    .A2(net4957));
 sg13g2_nand2_1 _16228_ (.Y(_06659_),
    .A(net2190),
    .B(net4957));
 sg13g2_o21ai_1 _16229_ (.B1(_06659_),
    .Y(_01115_),
    .A1(net5705),
    .A2(net4956));
 sg13g2_nand2_1 _16230_ (.Y(_06660_),
    .A(net2335),
    .B(net4956));
 sg13g2_o21ai_1 _16231_ (.B1(_06660_),
    .Y(_01116_),
    .A1(net5750),
    .A2(net4956));
 sg13g2_nor2_2 _16232_ (.A(_02947_),
    .B(_03331_),
    .Y(_06661_));
 sg13g2_nor2_1 _16233_ (.A(net3485),
    .B(net4739),
    .Y(_06662_));
 sg13g2_a21oi_1 _16234_ (.A1(net5435),
    .A2(net4739),
    .Y(_01117_),
    .B1(_06662_));
 sg13g2_nor2_1 _16235_ (.A(net3942),
    .B(net4741),
    .Y(_06663_));
 sg13g2_a21oi_1 _16236_ (.A1(net5480),
    .A2(net4741),
    .Y(_01118_),
    .B1(_06663_));
 sg13g2_nor2_1 _16237_ (.A(net3761),
    .B(net4739),
    .Y(_06664_));
 sg13g2_a21oi_1 _16238_ (.A1(net5524),
    .A2(net4739),
    .Y(_01119_),
    .B1(_06664_));
 sg13g2_nor2_1 _16239_ (.A(net3932),
    .B(net4741),
    .Y(_06665_));
 sg13g2_a21oi_1 _16240_ (.A1(net5569),
    .A2(net4741),
    .Y(_01120_),
    .B1(_06665_));
 sg13g2_nor2_1 _16241_ (.A(net3787),
    .B(net4740),
    .Y(_06666_));
 sg13g2_a21oi_1 _16242_ (.A1(net5615),
    .A2(net4740),
    .Y(_01121_),
    .B1(_06666_));
 sg13g2_nor2_1 _16243_ (.A(net4036),
    .B(net4740),
    .Y(_06667_));
 sg13g2_a21oi_1 _16244_ (.A1(net5661),
    .A2(net4740),
    .Y(_01122_),
    .B1(_06667_));
 sg13g2_nor2_1 _16245_ (.A(net3690),
    .B(net4739),
    .Y(_06668_));
 sg13g2_a21oi_1 _16246_ (.A1(net5705),
    .A2(net4739),
    .Y(_01123_),
    .B1(_06668_));
 sg13g2_nor2_1 _16247_ (.A(net3410),
    .B(net4739),
    .Y(_06669_));
 sg13g2_a21oi_1 _16248_ (.A1(net5750),
    .A2(net4739),
    .Y(_01124_),
    .B1(_06669_));
 sg13g2_nand3_1 _16249_ (.B(_03159_),
    .C(net5249),
    .A(net5220),
    .Y(_06670_));
 sg13g2_nand2_1 _16250_ (.Y(_06671_),
    .A(net2233),
    .B(net4955));
 sg13g2_o21ai_1 _16251_ (.B1(_06671_),
    .Y(_01125_),
    .A1(net5450),
    .A2(net4955));
 sg13g2_nand2_1 _16252_ (.Y(_06672_),
    .A(net3049),
    .B(net4954));
 sg13g2_o21ai_1 _16253_ (.B1(_06672_),
    .Y(_01126_),
    .A1(net5495),
    .A2(net4954));
 sg13g2_nand2_1 _16254_ (.Y(_06673_),
    .A(net3269),
    .B(net4954));
 sg13g2_o21ai_1 _16255_ (.B1(_06673_),
    .Y(_01127_),
    .A1(net5543),
    .A2(net4954));
 sg13g2_nand2_1 _16256_ (.Y(_06674_),
    .A(net2676),
    .B(net4955));
 sg13g2_o21ai_1 _16257_ (.B1(_06674_),
    .Y(_01128_),
    .A1(net5584),
    .A2(net4955));
 sg13g2_nand2_1 _16258_ (.Y(_06675_),
    .A(net3265),
    .B(net4954));
 sg13g2_o21ai_1 _16259_ (.B1(_06675_),
    .Y(_01129_),
    .A1(net5630),
    .A2(net4954));
 sg13g2_nand2_1 _16260_ (.Y(_06676_),
    .A(net2719),
    .B(net4954));
 sg13g2_o21ai_1 _16261_ (.B1(_06676_),
    .Y(_01130_),
    .A1(net5675),
    .A2(net4954));
 sg13g2_nand2_1 _16262_ (.Y(_06677_),
    .A(net2147),
    .B(net4955));
 sg13g2_o21ai_1 _16263_ (.B1(_06677_),
    .Y(_01131_),
    .A1(net5720),
    .A2(net4955));
 sg13g2_nand2_1 _16264_ (.Y(_06678_),
    .A(net2511),
    .B(net4955));
 sg13g2_o21ai_1 _16265_ (.B1(_06678_),
    .Y(_01132_),
    .A1(net5765),
    .A2(net4955));
 sg13g2_nor2_1 _16266_ (.A(net5143),
    .B(_03467_),
    .Y(_06679_));
 sg13g2_nor2_1 _16267_ (.A(net3331),
    .B(net4737),
    .Y(_06680_));
 sg13g2_a21oi_1 _16268_ (.A1(net5448),
    .A2(net4737),
    .Y(_01133_),
    .B1(_06680_));
 sg13g2_nor2_1 _16269_ (.A(net3570),
    .B(net4737),
    .Y(_06681_));
 sg13g2_a21oi_1 _16270_ (.A1(net5492),
    .A2(net4737),
    .Y(_01134_),
    .B1(_06681_));
 sg13g2_nor2_1 _16271_ (.A(net3449),
    .B(net4738),
    .Y(_06682_));
 sg13g2_a21oi_1 _16272_ (.A1(net5539),
    .A2(net4738),
    .Y(_01135_),
    .B1(_06682_));
 sg13g2_nor2_1 _16273_ (.A(net3337),
    .B(net4738),
    .Y(_06683_));
 sg13g2_a21oi_1 _16274_ (.A1(net5582),
    .A2(net4738),
    .Y(_01136_),
    .B1(_06683_));
 sg13g2_nor2_1 _16275_ (.A(net3989),
    .B(net4738),
    .Y(_06684_));
 sg13g2_a21oi_1 _16276_ (.A1(net5629),
    .A2(net4738),
    .Y(_01137_),
    .B1(_06684_));
 sg13g2_nor2_1 _16277_ (.A(net3962),
    .B(net4737),
    .Y(_06685_));
 sg13g2_a21oi_1 _16278_ (.A1(net5672),
    .A2(net4737),
    .Y(_01138_),
    .B1(_06685_));
 sg13g2_nor2_1 _16279_ (.A(net3821),
    .B(net4737),
    .Y(_06686_));
 sg13g2_a21oi_1 _16280_ (.A1(net5718),
    .A2(net4737),
    .Y(_01139_),
    .B1(_06686_));
 sg13g2_nor2_1 _16281_ (.A(net3670),
    .B(net4738),
    .Y(_06687_));
 sg13g2_a21oi_1 _16282_ (.A1(net5763),
    .A2(net4738),
    .Y(_01140_),
    .B1(_06687_));
 sg13g2_nor2_1 _16283_ (.A(net5254),
    .B(net5139),
    .Y(_06688_));
 sg13g2_nor2_1 _16284_ (.A(net3538),
    .B(net4736),
    .Y(_06689_));
 sg13g2_a21oi_1 _16285_ (.A1(net5450),
    .A2(net4736),
    .Y(_01141_),
    .B1(_06689_));
 sg13g2_nor2_1 _16286_ (.A(net3659),
    .B(net4735),
    .Y(_06690_));
 sg13g2_a21oi_1 _16287_ (.A1(net5490),
    .A2(net4735),
    .Y(_01142_),
    .B1(_06690_));
 sg13g2_nor2_1 _16288_ (.A(net3964),
    .B(net4735),
    .Y(_06691_));
 sg13g2_a21oi_1 _16289_ (.A1(net5540),
    .A2(net4735),
    .Y(_01143_),
    .B1(_06691_));
 sg13g2_nor2_1 _16290_ (.A(net3882),
    .B(net4736),
    .Y(_06692_));
 sg13g2_a21oi_1 _16291_ (.A1(net5585),
    .A2(net4736),
    .Y(_01144_),
    .B1(_06692_));
 sg13g2_nor2_1 _16292_ (.A(net3597),
    .B(net4735),
    .Y(_06693_));
 sg13g2_a21oi_1 _16293_ (.A1(net5626),
    .A2(net4735),
    .Y(_01145_),
    .B1(_06693_));
 sg13g2_nor2_1 _16294_ (.A(net3774),
    .B(net4735),
    .Y(_06694_));
 sg13g2_a21oi_1 _16295_ (.A1(net5675),
    .A2(net4735),
    .Y(_01146_),
    .B1(_06694_));
 sg13g2_nor2_1 _16296_ (.A(net3935),
    .B(net4736),
    .Y(_06695_));
 sg13g2_a21oi_1 _16297_ (.A1(net5720),
    .A2(net4736),
    .Y(_01147_),
    .B1(_06695_));
 sg13g2_nor2_1 _16298_ (.A(net3794),
    .B(net4736),
    .Y(_06696_));
 sg13g2_a21oi_1 _16299_ (.A1(net5768),
    .A2(net4736),
    .Y(_01148_),
    .B1(_06696_));
 sg13g2_nor2_1 _16300_ (.A(_03120_),
    .B(net5139),
    .Y(_06697_));
 sg13g2_nor2_1 _16301_ (.A(net3704),
    .B(net4734),
    .Y(_06698_));
 sg13g2_a21oi_1 _16302_ (.A1(net5449),
    .A2(net4734),
    .Y(_01149_),
    .B1(_06698_));
 sg13g2_nor2_1 _16303_ (.A(net3314),
    .B(net4733),
    .Y(_06699_));
 sg13g2_a21oi_1 _16304_ (.A1(net5490),
    .A2(net4733),
    .Y(_01150_),
    .B1(_06699_));
 sg13g2_nor2_1 _16305_ (.A(net4019),
    .B(net4733),
    .Y(_06700_));
 sg13g2_a21oi_1 _16306_ (.A1(net5540),
    .A2(net4733),
    .Y(_01151_),
    .B1(_06700_));
 sg13g2_nor2_1 _16307_ (.A(net3561),
    .B(net4734),
    .Y(_06701_));
 sg13g2_a21oi_1 _16308_ (.A1(net5585),
    .A2(net4734),
    .Y(_01152_),
    .B1(_06701_));
 sg13g2_nor2_1 _16309_ (.A(net4041),
    .B(net4733),
    .Y(_06702_));
 sg13g2_a21oi_1 _16310_ (.A1(net5626),
    .A2(net4733),
    .Y(_01153_),
    .B1(_06702_));
 sg13g2_nor2_1 _16311_ (.A(net3874),
    .B(net4733),
    .Y(_06703_));
 sg13g2_a21oi_1 _16312_ (.A1(net5674),
    .A2(net4733),
    .Y(_01154_),
    .B1(_06703_));
 sg13g2_nor2_1 _16313_ (.A(net3472),
    .B(net4734),
    .Y(_06704_));
 sg13g2_a21oi_1 _16314_ (.A1(net5720),
    .A2(net4734),
    .Y(_01155_),
    .B1(_06704_));
 sg13g2_nor2_1 _16315_ (.A(net3754),
    .B(net4734),
    .Y(_06705_));
 sg13g2_a21oi_1 _16316_ (.A1(net5768),
    .A2(net4734),
    .Y(_01156_),
    .B1(_06705_));
 sg13g2_nor2_1 _16317_ (.A(_03109_),
    .B(net5139),
    .Y(_06706_));
 sg13g2_nor2_1 _16318_ (.A(net3729),
    .B(net4731),
    .Y(_06707_));
 sg13g2_a21oi_1 _16319_ (.A1(net5449),
    .A2(net4731),
    .Y(_01157_),
    .B1(_06707_));
 sg13g2_nor2_1 _16320_ (.A(net3459),
    .B(net4731),
    .Y(_06708_));
 sg13g2_a21oi_1 _16321_ (.A1(net5495),
    .A2(net4731),
    .Y(_01158_),
    .B1(_06708_));
 sg13g2_nor2_1 _16322_ (.A(net4080),
    .B(net4731),
    .Y(_06709_));
 sg13g2_a21oi_1 _16323_ (.A1(net5540),
    .A2(net4731),
    .Y(_01159_),
    .B1(_06709_));
 sg13g2_nor2_1 _16324_ (.A(net3198),
    .B(net4731),
    .Y(_06710_));
 sg13g2_a21oi_1 _16325_ (.A1(net5585),
    .A2(net4731),
    .Y(_01160_),
    .B1(_06710_));
 sg13g2_nor2_1 _16326_ (.A(net4131),
    .B(net4732),
    .Y(_06711_));
 sg13g2_a21oi_1 _16327_ (.A1(net5640),
    .A2(net4732),
    .Y(_01161_),
    .B1(_06711_));
 sg13g2_nor2_1 _16328_ (.A(net3931),
    .B(net4732),
    .Y(_06712_));
 sg13g2_a21oi_1 _16329_ (.A1(net5686),
    .A2(net4732),
    .Y(_01162_),
    .B1(_06712_));
 sg13g2_nor2_1 _16330_ (.A(net3567),
    .B(net4732),
    .Y(_06713_));
 sg13g2_a21oi_1 _16331_ (.A1(net5731),
    .A2(net4732),
    .Y(_01163_),
    .B1(_06713_));
 sg13g2_nor2_1 _16332_ (.A(net3518),
    .B(net4732),
    .Y(_06714_));
 sg13g2_a21oi_1 _16333_ (.A1(net5778),
    .A2(net4732),
    .Y(_01164_),
    .B1(_06714_));
 sg13g2_nor2_1 _16334_ (.A(net5139),
    .B(_03201_),
    .Y(_06715_));
 sg13g2_nor2_1 _16335_ (.A(net3999),
    .B(net4729),
    .Y(_06716_));
 sg13g2_a21oi_1 _16336_ (.A1(net5449),
    .A2(net4729),
    .Y(_01165_),
    .B1(_06716_));
 sg13g2_nor2_1 _16337_ (.A(net3435),
    .B(net4729),
    .Y(_06717_));
 sg13g2_a21oi_1 _16338_ (.A1(net5495),
    .A2(net4729),
    .Y(_01166_),
    .B1(_06717_));
 sg13g2_nor2_1 _16339_ (.A(net3649),
    .B(net4729),
    .Y(_06718_));
 sg13g2_a21oi_1 _16340_ (.A1(net5540),
    .A2(net4729),
    .Y(_01167_),
    .B1(_06718_));
 sg13g2_nor2_1 _16341_ (.A(net4114),
    .B(net4730),
    .Y(_06719_));
 sg13g2_a21oi_1 _16342_ (.A1(net5585),
    .A2(net4730),
    .Y(_01168_),
    .B1(_06719_));
 sg13g2_nor2_1 _16343_ (.A(net3427),
    .B(net4729),
    .Y(_06720_));
 sg13g2_a21oi_1 _16344_ (.A1(net5634),
    .A2(net4729),
    .Y(_01169_),
    .B1(_06720_));
 sg13g2_nor2_1 _16345_ (.A(net4050),
    .B(_06715_),
    .Y(_06721_));
 sg13g2_a21oi_1 _16346_ (.A1(net5686),
    .A2(net4730),
    .Y(_01170_),
    .B1(_06721_));
 sg13g2_nor2_1 _16347_ (.A(net4150),
    .B(net4730),
    .Y(_06722_));
 sg13g2_a21oi_1 _16348_ (.A1(net5730),
    .A2(net4730),
    .Y(_01171_),
    .B1(_06722_));
 sg13g2_nor2_1 _16349_ (.A(net4089),
    .B(net4730),
    .Y(_06723_));
 sg13g2_a21oi_1 _16350_ (.A1(net5778),
    .A2(net4730),
    .Y(_01172_),
    .B1(_06723_));
 sg13g2_nor2_1 _16351_ (.A(_03067_),
    .B(net5139),
    .Y(_06724_));
 sg13g2_nor2_1 _16352_ (.A(net3924),
    .B(net4728),
    .Y(_06725_));
 sg13g2_a21oi_1 _16353_ (.A1(net5449),
    .A2(net4728),
    .Y(_01173_),
    .B1(_06725_));
 sg13g2_nor2_1 _16354_ (.A(net3321),
    .B(net4727),
    .Y(_06726_));
 sg13g2_a21oi_1 _16355_ (.A1(net5490),
    .A2(net4727),
    .Y(_01174_),
    .B1(_06726_));
 sg13g2_nor2_1 _16356_ (.A(net3798),
    .B(net4727),
    .Y(_06727_));
 sg13g2_a21oi_1 _16357_ (.A1(net5540),
    .A2(net4727),
    .Y(_01175_),
    .B1(_06727_));
 sg13g2_nor2_1 _16358_ (.A(net3075),
    .B(net4728),
    .Y(_06728_));
 sg13g2_a21oi_1 _16359_ (.A1(net5584),
    .A2(net4728),
    .Y(_01176_),
    .B1(_06728_));
 sg13g2_nor2_1 _16360_ (.A(net4004),
    .B(net4727),
    .Y(_06729_));
 sg13g2_a21oi_1 _16361_ (.A1(net5634),
    .A2(net4727),
    .Y(_01177_),
    .B1(_06729_));
 sg13g2_nor2_1 _16362_ (.A(net3333),
    .B(net4727),
    .Y(_06730_));
 sg13g2_a21oi_1 _16363_ (.A1(net5686),
    .A2(net4727),
    .Y(_01178_),
    .B1(_06730_));
 sg13g2_nor2_1 _16364_ (.A(net4068),
    .B(net4728),
    .Y(_06731_));
 sg13g2_a21oi_1 _16365_ (.A1(net5731),
    .A2(net4728),
    .Y(_01179_),
    .B1(_06731_));
 sg13g2_nor2_1 _16366_ (.A(net3466),
    .B(net4728),
    .Y(_06732_));
 sg13g2_a21oi_1 _16367_ (.A1(net5778),
    .A2(net4728),
    .Y(_01180_),
    .B1(_06732_));
 sg13g2_nand3_1 _16368_ (.B(net5238),
    .C(_03159_),
    .A(net5220),
    .Y(_06733_));
 sg13g2_nand2_1 _16369_ (.Y(_06734_),
    .A(net2954),
    .B(net4953));
 sg13g2_o21ai_1 _16370_ (.B1(_06734_),
    .Y(_01181_),
    .A1(net5449),
    .A2(net4953));
 sg13g2_nand2_1 _16371_ (.Y(_06735_),
    .A(net2988),
    .B(net4953));
 sg13g2_o21ai_1 _16372_ (.B1(_06735_),
    .Y(_01182_),
    .A1(net5495),
    .A2(net4953));
 sg13g2_nand2_1 _16373_ (.Y(_06736_),
    .A(net3115),
    .B(net4952));
 sg13g2_o21ai_1 _16374_ (.B1(_06736_),
    .Y(_01183_),
    .A1(net5553),
    .A2(net4952));
 sg13g2_nand2_1 _16375_ (.Y(_06737_),
    .A(net3206),
    .B(net4953));
 sg13g2_o21ai_1 _16376_ (.B1(_06737_),
    .Y(_01184_),
    .A1(net5584),
    .A2(net4953));
 sg13g2_nand2_1 _16377_ (.Y(_06738_),
    .A(net3251),
    .B(net4952));
 sg13g2_o21ai_1 _16378_ (.B1(_06738_),
    .Y(_01185_),
    .A1(net5634),
    .A2(net4952));
 sg13g2_nand2_1 _16379_ (.Y(_06739_),
    .A(net2654),
    .B(net4952));
 sg13g2_o21ai_1 _16380_ (.B1(_06739_),
    .Y(_01186_),
    .A1(net5686),
    .A2(net4952));
 sg13g2_nand2_1 _16381_ (.Y(_06740_),
    .A(net3037),
    .B(net4953));
 sg13g2_o21ai_1 _16382_ (.B1(_06740_),
    .Y(_01187_),
    .A1(net5731),
    .A2(_06733_));
 sg13g2_nand2_1 _16383_ (.Y(_06741_),
    .A(net3195),
    .B(net4952));
 sg13g2_o21ai_1 _16384_ (.B1(_06741_),
    .Y(_01188_),
    .A1(net5778),
    .A2(net4952));
 sg13g2_nor2_1 _16385_ (.A(_02939_),
    .B(net5138),
    .Y(_06742_));
 sg13g2_nor2_1 _16386_ (.A(net3424),
    .B(net4726),
    .Y(_06743_));
 sg13g2_a21oi_1 _16387_ (.A1(net5451),
    .A2(net4726),
    .Y(_01189_),
    .B1(_06743_));
 sg13g2_nor2_1 _16388_ (.A(net4077),
    .B(net4725),
    .Y(_06744_));
 sg13g2_a21oi_1 _16389_ (.A1(net5492),
    .A2(net4725),
    .Y(_01190_),
    .B1(_06744_));
 sg13g2_nor2_1 _16390_ (.A(net3651),
    .B(net4726),
    .Y(_06745_));
 sg13g2_a21oi_1 _16391_ (.A1(net5542),
    .A2(net4726),
    .Y(_01191_),
    .B1(_06745_));
 sg13g2_nor2_1 _16392_ (.A(net3588),
    .B(net4725),
    .Y(_06746_));
 sg13g2_a21oi_1 _16393_ (.A1(net5586),
    .A2(net4725),
    .Y(_01192_),
    .B1(_06746_));
 sg13g2_nor2_1 _16394_ (.A(net3722),
    .B(net4725),
    .Y(_06747_));
 sg13g2_a21oi_1 _16395_ (.A1(net5631),
    .A2(net4725),
    .Y(_01193_),
    .B1(_06747_));
 sg13g2_nor2_1 _16396_ (.A(net4011),
    .B(net4726),
    .Y(_06748_));
 sg13g2_a21oi_1 _16397_ (.A1(net5675),
    .A2(net4726),
    .Y(_01194_),
    .B1(_06748_));
 sg13g2_nor2_1 _16398_ (.A(net3596),
    .B(net4726),
    .Y(_06749_));
 sg13g2_a21oi_1 _16399_ (.A1(net5722),
    .A2(net4726),
    .Y(_01195_),
    .B1(_06749_));
 sg13g2_nor2_1 _16400_ (.A(net3737),
    .B(net4725),
    .Y(_06750_));
 sg13g2_a21oi_1 _16401_ (.A1(net5766),
    .A2(net4725),
    .Y(_01196_),
    .B1(_06750_));
 sg13g2_nor2_1 _16402_ (.A(_03017_),
    .B(net5139),
    .Y(_06751_));
 sg13g2_nor2_1 _16403_ (.A(net3420),
    .B(net4724),
    .Y(_06752_));
 sg13g2_a21oi_1 _16404_ (.A1(net5451),
    .A2(net4724),
    .Y(_01197_),
    .B1(_06752_));
 sg13g2_nor2_1 _16405_ (.A(net4028),
    .B(net4723),
    .Y(_06753_));
 sg13g2_a21oi_1 _16406_ (.A1(net5497),
    .A2(net4723),
    .Y(_01198_),
    .B1(_06753_));
 sg13g2_nor2_1 _16407_ (.A(net3824),
    .B(net4724),
    .Y(_06754_));
 sg13g2_a21oi_1 _16408_ (.A1(net5542),
    .A2(net4724),
    .Y(_01199_),
    .B1(_06754_));
 sg13g2_nor2_1 _16409_ (.A(net3767),
    .B(net4723),
    .Y(_06755_));
 sg13g2_a21oi_1 _16410_ (.A1(net5586),
    .A2(net4723),
    .Y(_01200_),
    .B1(_06755_));
 sg13g2_nor2_1 _16411_ (.A(net3464),
    .B(net4723),
    .Y(_06756_));
 sg13g2_a21oi_1 _16412_ (.A1(net5631),
    .A2(net4723),
    .Y(_01201_),
    .B1(_06756_));
 sg13g2_nor2_1 _16413_ (.A(net3326),
    .B(net4724),
    .Y(_06757_));
 sg13g2_a21oi_1 _16414_ (.A1(net5675),
    .A2(net4724),
    .Y(_01202_),
    .B1(_06757_));
 sg13g2_nor2_1 _16415_ (.A(net4074),
    .B(net4724),
    .Y(_06758_));
 sg13g2_a21oi_1 _16416_ (.A1(net5722),
    .A2(net4724),
    .Y(_01203_),
    .B1(_06758_));
 sg13g2_nor2_1 _16417_ (.A(net3551),
    .B(net4723),
    .Y(_06759_));
 sg13g2_a21oi_1 _16418_ (.A1(net5766),
    .A2(net4723),
    .Y(_01204_),
    .B1(_06759_));
 sg13g2_nor2_1 _16419_ (.A(_02981_),
    .B(net5138),
    .Y(_06760_));
 sg13g2_nor2_1 _16420_ (.A(net3845),
    .B(net4722),
    .Y(_06761_));
 sg13g2_a21oi_1 _16421_ (.A1(net5451),
    .A2(net4722),
    .Y(_01205_),
    .B1(_06761_));
 sg13g2_nor2_1 _16422_ (.A(net3696),
    .B(net4721),
    .Y(_06762_));
 sg13g2_a21oi_1 _16423_ (.A1(net5497),
    .A2(net4721),
    .Y(_01206_),
    .B1(_06762_));
 sg13g2_nor2_1 _16424_ (.A(net3373),
    .B(net4722),
    .Y(_06763_));
 sg13g2_a21oi_1 _16425_ (.A1(net5541),
    .A2(net4722),
    .Y(_01207_),
    .B1(_06763_));
 sg13g2_nor2_1 _16426_ (.A(net3956),
    .B(net4721),
    .Y(_06764_));
 sg13g2_a21oi_1 _16427_ (.A1(net5586),
    .A2(net4721),
    .Y(_01208_),
    .B1(_06764_));
 sg13g2_nor2_1 _16428_ (.A(net3350),
    .B(net4721),
    .Y(_06765_));
 sg13g2_a21oi_1 _16429_ (.A1(net5631),
    .A2(net4721),
    .Y(_01209_),
    .B1(_06765_));
 sg13g2_nor2_1 _16430_ (.A(net3757),
    .B(net4722),
    .Y(_06766_));
 sg13g2_a21oi_1 _16431_ (.A1(net5675),
    .A2(net4722),
    .Y(_01210_),
    .B1(_06766_));
 sg13g2_nor2_1 _16432_ (.A(net3927),
    .B(net4722),
    .Y(_06767_));
 sg13g2_a21oi_1 _16433_ (.A1(net5721),
    .A2(net4722),
    .Y(_01211_),
    .B1(_06767_));
 sg13g2_nor2_1 _16434_ (.A(net3604),
    .B(net4721),
    .Y(_06768_));
 sg13g2_a21oi_1 _16435_ (.A1(net5766),
    .A2(net4721),
    .Y(_01212_),
    .B1(_06768_));
 sg13g2_nor2_1 _16436_ (.A(net5143),
    .B(_03212_),
    .Y(_06769_));
 sg13g2_nor2_1 _16437_ (.A(net4123),
    .B(net4720),
    .Y(_06770_));
 sg13g2_a21oi_1 _16438_ (.A1(net5448),
    .A2(net4720),
    .Y(_01213_),
    .B1(_06770_));
 sg13g2_nor2_1 _16439_ (.A(net3847),
    .B(net4720),
    .Y(_06771_));
 sg13g2_a21oi_1 _16440_ (.A1(net5493),
    .A2(net4720),
    .Y(_01214_),
    .B1(_06771_));
 sg13g2_nor2_1 _16441_ (.A(net3364),
    .B(net4719),
    .Y(_06772_));
 sg13g2_a21oi_1 _16442_ (.A1(net5539),
    .A2(net4720),
    .Y(_01215_),
    .B1(_06772_));
 sg13g2_nor2_1 _16443_ (.A(net3952),
    .B(net4719),
    .Y(_06773_));
 sg13g2_a21oi_1 _16444_ (.A1(net5582),
    .A2(net4719),
    .Y(_01216_),
    .B1(_06773_));
 sg13g2_nor2_1 _16445_ (.A(net3645),
    .B(net4719),
    .Y(_06774_));
 sg13g2_a21oi_1 _16446_ (.A1(net5629),
    .A2(_06769_),
    .Y(_01217_),
    .B1(_06774_));
 sg13g2_nor2_1 _16447_ (.A(net4017),
    .B(net4719),
    .Y(_06775_));
 sg13g2_a21oi_1 _16448_ (.A1(net5672),
    .A2(net4719),
    .Y(_01218_),
    .B1(_06775_));
 sg13g2_nor2_1 _16449_ (.A(net3873),
    .B(net4720),
    .Y(_06776_));
 sg13g2_a21oi_1 _16450_ (.A1(net5717),
    .A2(net4720),
    .Y(_01219_),
    .B1(_06776_));
 sg13g2_nor2_1 _16451_ (.A(net3592),
    .B(net4719),
    .Y(_06777_));
 sg13g2_a21oi_1 _16452_ (.A1(net5763),
    .A2(net4719),
    .Y(_01220_),
    .B1(_06777_));
 sg13g2_nor2_1 _16453_ (.A(net5138),
    .B(_03467_),
    .Y(_06778_));
 sg13g2_nor2_1 _16454_ (.A(net4164),
    .B(net4717),
    .Y(_06779_));
 sg13g2_a21oi_1 _16455_ (.A1(net5451),
    .A2(net4717),
    .Y(_01221_),
    .B1(_06779_));
 sg13g2_nor2_1 _16456_ (.A(net4055),
    .B(net4718),
    .Y(_06780_));
 sg13g2_a21oi_1 _16457_ (.A1(net5493),
    .A2(net4718),
    .Y(_01222_),
    .B1(_06780_));
 sg13g2_nor2_1 _16458_ (.A(net3870),
    .B(net4717),
    .Y(_06781_));
 sg13g2_a21oi_1 _16459_ (.A1(net5542),
    .A2(net4717),
    .Y(_01223_),
    .B1(_06781_));
 sg13g2_nor2_1 _16460_ (.A(net2743),
    .B(net4718),
    .Y(_06782_));
 sg13g2_a21oi_1 _16461_ (.A1(net5581),
    .A2(net4718),
    .Y(_01224_),
    .B1(_06782_));
 sg13g2_nor2_1 _16462_ (.A(net3492),
    .B(net4718),
    .Y(_06783_));
 sg13g2_a21oi_1 _16463_ (.A1(net5630),
    .A2(net4718),
    .Y(_01225_),
    .B1(_06783_));
 sg13g2_nor2_1 _16464_ (.A(net3359),
    .B(net4717),
    .Y(_06784_));
 sg13g2_a21oi_1 _16465_ (.A1(net5676),
    .A2(net4717),
    .Y(_01226_),
    .B1(_06784_));
 sg13g2_nor2_1 _16466_ (.A(net4125),
    .B(net4717),
    .Y(_06785_));
 sg13g2_a21oi_1 _16467_ (.A1(net5721),
    .A2(net4717),
    .Y(_01227_),
    .B1(_06785_));
 sg13g2_nor2_1 _16468_ (.A(net3743),
    .B(_06778_),
    .Y(_06786_));
 sg13g2_a21oi_1 _16469_ (.A1(net5766),
    .A2(net4718),
    .Y(_01228_),
    .B1(_06786_));
 sg13g2_nor2_1 _16470_ (.A(net5138),
    .B(_03212_),
    .Y(_06787_));
 sg13g2_nor2_1 _16471_ (.A(net3744),
    .B(net4716),
    .Y(_06788_));
 sg13g2_a21oi_1 _16472_ (.A1(net5451),
    .A2(net4716),
    .Y(_01229_),
    .B1(_06788_));
 sg13g2_nor2_1 _16473_ (.A(net3661),
    .B(net4715),
    .Y(_06789_));
 sg13g2_a21oi_1 _16474_ (.A1(net5493),
    .A2(net4715),
    .Y(_01230_),
    .B1(_06789_));
 sg13g2_nor2_1 _16475_ (.A(net3672),
    .B(net4716),
    .Y(_06790_));
 sg13g2_a21oi_1 _16476_ (.A1(net5542),
    .A2(net4716),
    .Y(_01231_),
    .B1(_06790_));
 sg13g2_nor2_1 _16477_ (.A(net4148),
    .B(net4715),
    .Y(_06791_));
 sg13g2_a21oi_1 _16478_ (.A1(net5581),
    .A2(net4715),
    .Y(_01232_),
    .B1(_06791_));
 sg13g2_nor2_1 _16479_ (.A(net3445),
    .B(net4715),
    .Y(_06792_));
 sg13g2_a21oi_1 _16480_ (.A1(net5631),
    .A2(net4715),
    .Y(_01233_),
    .B1(_06792_));
 sg13g2_nor2_1 _16481_ (.A(net4084),
    .B(net4716),
    .Y(_06793_));
 sg13g2_a21oi_1 _16482_ (.A1(net5676),
    .A2(net4716),
    .Y(_01234_),
    .B1(_06793_));
 sg13g2_nor2_1 _16483_ (.A(net3414),
    .B(net4716),
    .Y(_06794_));
 sg13g2_a21oi_1 _16484_ (.A1(net5721),
    .A2(net4716),
    .Y(_01235_),
    .B1(_06794_));
 sg13g2_nor2_1 _16485_ (.A(net4022),
    .B(net4715),
    .Y(_06795_));
 sg13g2_a21oi_1 _16486_ (.A1(net5766),
    .A2(net4715),
    .Y(_01236_),
    .B1(_06795_));
 sg13g2_nor2_1 _16487_ (.A(net5138),
    .B(_03375_),
    .Y(_06796_));
 sg13g2_nor2_1 _16488_ (.A(net3413),
    .B(net4713),
    .Y(_06797_));
 sg13g2_a21oi_1 _16489_ (.A1(net5451),
    .A2(net4713),
    .Y(_01237_),
    .B1(_06797_));
 sg13g2_nor2_1 _16490_ (.A(net3486),
    .B(net4714),
    .Y(_06798_));
 sg13g2_a21oi_1 _16491_ (.A1(net5492),
    .A2(net4714),
    .Y(_01238_),
    .B1(_06798_));
 sg13g2_nor2_1 _16492_ (.A(net3552),
    .B(_06796_),
    .Y(_06799_));
 sg13g2_a21oi_1 _16493_ (.A1(net5542),
    .A2(net4713),
    .Y(_01239_),
    .B1(_06799_));
 sg13g2_nor2_1 _16494_ (.A(net3361),
    .B(net4714),
    .Y(_06800_));
 sg13g2_a21oi_1 _16495_ (.A1(net5581),
    .A2(net4714),
    .Y(_01240_),
    .B1(_06800_));
 sg13g2_nor2_1 _16496_ (.A(net3601),
    .B(net4714),
    .Y(_06801_));
 sg13g2_a21oi_1 _16497_ (.A1(net5630),
    .A2(net4714),
    .Y(_01241_),
    .B1(_06801_));
 sg13g2_nor2_1 _16498_ (.A(net3577),
    .B(net4713),
    .Y(_06802_));
 sg13g2_a21oi_1 _16499_ (.A1(net5676),
    .A2(net4713),
    .Y(_01242_),
    .B1(_06802_));
 sg13g2_nor2_1 _16500_ (.A(net3409),
    .B(net4713),
    .Y(_06803_));
 sg13g2_a21oi_1 _16501_ (.A1(net5721),
    .A2(net4713),
    .Y(_01243_),
    .B1(_06803_));
 sg13g2_nor2_1 _16502_ (.A(net4012),
    .B(net4713),
    .Y(_06804_));
 sg13g2_a21oi_1 _16503_ (.A1(net5766),
    .A2(net4714),
    .Y(_01244_),
    .B1(_06804_));
 sg13g2_nor2_1 _16504_ (.A(net5240),
    .B(net5138),
    .Y(_06805_));
 sg13g2_nor2_1 _16505_ (.A(net3558),
    .B(net4712),
    .Y(_06806_));
 sg13g2_a21oi_1 _16506_ (.A1(net5451),
    .A2(net4712),
    .Y(_01245_),
    .B1(_06806_));
 sg13g2_nor2_1 _16507_ (.A(net3640),
    .B(net4711),
    .Y(_06807_));
 sg13g2_a21oi_1 _16508_ (.A1(net5492),
    .A2(net4711),
    .Y(_01246_),
    .B1(_06807_));
 sg13g2_nor2_1 _16509_ (.A(net4154),
    .B(net4712),
    .Y(_06808_));
 sg13g2_a21oi_1 _16510_ (.A1(net5542),
    .A2(net4712),
    .Y(_01247_),
    .B1(_06808_));
 sg13g2_nor2_1 _16511_ (.A(net3674),
    .B(net4711),
    .Y(_06809_));
 sg13g2_a21oi_1 _16512_ (.A1(net5581),
    .A2(net4711),
    .Y(_01248_),
    .B1(_06809_));
 sg13g2_nor2_1 _16513_ (.A(net3921),
    .B(net4711),
    .Y(_06810_));
 sg13g2_a21oi_1 _16514_ (.A1(net5630),
    .A2(net4711),
    .Y(_01249_),
    .B1(_06810_));
 sg13g2_nor2_1 _16515_ (.A(net3681),
    .B(net4712),
    .Y(_06811_));
 sg13g2_a21oi_1 _16516_ (.A1(net5676),
    .A2(net4712),
    .Y(_01250_),
    .B1(_06811_));
 sg13g2_nor2_1 _16517_ (.A(net3525),
    .B(net4712),
    .Y(_06812_));
 sg13g2_a21oi_1 _16518_ (.A1(net5721),
    .A2(net4712),
    .Y(_01251_),
    .B1(_06812_));
 sg13g2_nor2_1 _16519_ (.A(net3590),
    .B(net4711),
    .Y(_06813_));
 sg13g2_a21oi_1 _16520_ (.A1(net5766),
    .A2(net4711),
    .Y(_01252_),
    .B1(_06813_));
 sg13g2_nand2_1 _16521_ (.Y(_06814_),
    .A(net5212),
    .B(net5249));
 sg13g2_nand2_1 _16522_ (.Y(_06815_),
    .A(net2999),
    .B(net4951));
 sg13g2_o21ai_1 _16523_ (.B1(_06815_),
    .Y(_01253_),
    .A1(net5446),
    .A2(net4951));
 sg13g2_nand2_1 _16524_ (.Y(_06816_),
    .A(net2565),
    .B(net4951));
 sg13g2_o21ai_1 _16525_ (.B1(_06816_),
    .Y(_01254_),
    .A1(net5494),
    .A2(net4951));
 sg13g2_nand2_1 _16526_ (.Y(_06817_),
    .A(net2652),
    .B(net4950));
 sg13g2_o21ai_1 _16527_ (.B1(_06817_),
    .Y(_01255_),
    .A1(net5538),
    .A2(net4950));
 sg13g2_nor2_1 _16528_ (.A(\mem.data_in[3] ),
    .B(net4951),
    .Y(_06818_));
 sg13g2_a21oi_1 _16529_ (.A1(_02856_),
    .A2(net4951),
    .Y(_01256_),
    .B1(_06818_));
 sg13g2_nand2_1 _16530_ (.Y(_06819_),
    .A(net2604),
    .B(net4950));
 sg13g2_o21ai_1 _16531_ (.B1(_06819_),
    .Y(_01257_),
    .A1(net5620),
    .A2(net4950));
 sg13g2_nand2_1 _16532_ (.Y(_06820_),
    .A(net3084),
    .B(net4950));
 sg13g2_o21ai_1 _16533_ (.B1(_06820_),
    .Y(_01258_),
    .A1(net5670),
    .A2(net4950));
 sg13g2_nand2_1 _16534_ (.Y(_06821_),
    .A(net3426),
    .B(net4951));
 sg13g2_o21ai_1 _16535_ (.B1(_06821_),
    .Y(_01259_),
    .A1(net5718),
    .A2(_06814_));
 sg13g2_nand2_1 _16536_ (.Y(_06822_),
    .A(net2851),
    .B(net4950));
 sg13g2_o21ai_1 _16537_ (.B1(_06822_),
    .Y(_01260_),
    .A1(net5762),
    .A2(net4950));
 sg13g2_nor3_1 _16538_ (.A(net5229),
    .B(net5252),
    .C(net5258),
    .Y(_06823_));
 sg13g2_nor2_1 _16539_ (.A(net3626),
    .B(net5183),
    .Y(_06824_));
 sg13g2_a21oi_1 _16540_ (.A1(net5446),
    .A2(net5183),
    .Y(_01261_),
    .B1(_06824_));
 sg13g2_nor2_1 _16541_ (.A(net4061),
    .B(net5182),
    .Y(_06825_));
 sg13g2_a21oi_1 _16542_ (.A1(net5494),
    .A2(net5182),
    .Y(_01262_),
    .B1(_06825_));
 sg13g2_nor2_1 _16543_ (.A(net3471),
    .B(net5183),
    .Y(_06826_));
 sg13g2_a21oi_1 _16544_ (.A1(net5538),
    .A2(net5182),
    .Y(_01263_),
    .B1(_06826_));
 sg13g2_nor2_1 _16545_ (.A(net3966),
    .B(net5182),
    .Y(_06827_));
 sg13g2_a21oi_1 _16546_ (.A1(net5583),
    .A2(net5182),
    .Y(_01264_),
    .B1(_06827_));
 sg13g2_nor2_1 _16547_ (.A(net3917),
    .B(net5182),
    .Y(_06828_));
 sg13g2_a21oi_1 _16548_ (.A1(net5620),
    .A2(net5182),
    .Y(_01265_),
    .B1(_06828_));
 sg13g2_nor2_1 _16549_ (.A(net3740),
    .B(net5182),
    .Y(_06829_));
 sg13g2_a21oi_1 _16550_ (.A1(net5670),
    .A2(net5183),
    .Y(_01266_),
    .B1(_06829_));
 sg13g2_nor2_1 _16551_ (.A(net4071),
    .B(_06823_),
    .Y(_06830_));
 sg13g2_a21oi_1 _16552_ (.A1(net5718),
    .A2(net5183),
    .Y(_01267_),
    .B1(_06830_));
 sg13g2_nor2_1 _16553_ (.A(net3514),
    .B(net5183),
    .Y(_06831_));
 sg13g2_a21oi_1 _16554_ (.A1(net5762),
    .A2(net5183),
    .Y(_01268_),
    .B1(_06831_));
 sg13g2_nor3_1 _16555_ (.A(net5229),
    .B(net5254),
    .C(net5258),
    .Y(_06832_));
 sg13g2_nor2_1 _16556_ (.A(net3727),
    .B(net5181),
    .Y(_06833_));
 sg13g2_a21oi_1 _16557_ (.A1(net5446),
    .A2(net5181),
    .Y(_01269_),
    .B1(_06833_));
 sg13g2_nor2_1 _16558_ (.A(net4059),
    .B(net5180),
    .Y(_06834_));
 sg13g2_a21oi_1 _16559_ (.A1(net5487),
    .A2(net5180),
    .Y(_01270_),
    .B1(_06834_));
 sg13g2_nor2_1 _16560_ (.A(net4118),
    .B(net5180),
    .Y(_06835_));
 sg13g2_a21oi_1 _16561_ (.A1(net5534),
    .A2(net5180),
    .Y(_01271_),
    .B1(_06835_));
 sg13g2_nor2_1 _16562_ (.A(net3447),
    .B(net5180),
    .Y(_06836_));
 sg13g2_a21oi_1 _16563_ (.A1(net5583),
    .A2(net5180),
    .Y(_01272_),
    .B1(_06836_));
 sg13g2_nor2_1 _16564_ (.A(net3685),
    .B(_06832_),
    .Y(_06837_));
 sg13g2_a21oi_1 _16565_ (.A1(net5620),
    .A2(net5181),
    .Y(_01273_),
    .B1(_06837_));
 sg13g2_nor2_1 _16566_ (.A(net3341),
    .B(net5181),
    .Y(_06838_));
 sg13g2_a21oi_1 _16567_ (.A1(net5670),
    .A2(net5181),
    .Y(_01274_),
    .B1(_06838_));
 sg13g2_nor2_1 _16568_ (.A(net3453),
    .B(net5181),
    .Y(_06839_));
 sg13g2_a21oi_1 _16569_ (.A1(net5717),
    .A2(net5181),
    .Y(_01275_),
    .B1(_06839_));
 sg13g2_nor2_1 _16570_ (.A(net3834),
    .B(net5180),
    .Y(_06840_));
 sg13g2_a21oi_1 _16571_ (.A1(net5762),
    .A2(net5180),
    .Y(_01276_),
    .B1(_06840_));
 sg13g2_nand2_1 _16572_ (.Y(_06841_),
    .A(net5253),
    .B(net5212));
 sg13g2_nand2_1 _16573_ (.Y(_06842_),
    .A(net3247),
    .B(net4949));
 sg13g2_o21ai_1 _16574_ (.B1(_06842_),
    .Y(_01277_),
    .A1(net5446),
    .A2(net4948));
 sg13g2_nand2_1 _16575_ (.Y(_06843_),
    .A(net3301),
    .B(net4948));
 sg13g2_o21ai_1 _16576_ (.B1(_06843_),
    .Y(_01278_),
    .A1(net5494),
    .A2(net4948));
 sg13g2_nand2_1 _16577_ (.Y(_06844_),
    .A(net2266),
    .B(_06841_));
 sg13g2_o21ai_1 _16578_ (.B1(_06844_),
    .Y(_01279_),
    .A1(net5538),
    .A2(net4948));
 sg13g2_nand2_1 _16579_ (.Y(_06845_),
    .A(net3362),
    .B(net4948));
 sg13g2_o21ai_1 _16580_ (.B1(_06845_),
    .Y(_01280_),
    .A1(net5583),
    .A2(net4948));
 sg13g2_nand2_1 _16581_ (.Y(_06846_),
    .A(net3487),
    .B(net4949));
 sg13g2_o21ai_1 _16582_ (.B1(_06846_),
    .Y(_01281_),
    .A1(net5620),
    .A2(net4949));
 sg13g2_nand2_1 _16583_ (.Y(_06847_),
    .A(net3291),
    .B(net4949));
 sg13g2_o21ai_1 _16584_ (.B1(_06847_),
    .Y(_01282_),
    .A1(net5670),
    .A2(net4949));
 sg13g2_nand2_1 _16585_ (.Y(_06848_),
    .A(net2582),
    .B(net4949));
 sg13g2_o21ai_1 _16586_ (.B1(_06848_),
    .Y(_01283_),
    .A1(net5717),
    .A2(net4949));
 sg13g2_nand2_1 _16587_ (.Y(_06849_),
    .A(net2605),
    .B(net4948));
 sg13g2_o21ai_1 _16588_ (.B1(_06849_),
    .Y(_01284_),
    .A1(net5762),
    .A2(net4948));
 sg13g2_nand2_1 _16589_ (.Y(_06850_),
    .A(_03108_),
    .B(net5212));
 sg13g2_nand2_1 _16590_ (.Y(_06851_),
    .A(net3105),
    .B(net4947));
 sg13g2_o21ai_1 _16591_ (.B1(_06851_),
    .Y(_01285_),
    .A1(net5446),
    .A2(net4947));
 sg13g2_nand2_1 _16592_ (.Y(_06852_),
    .A(net2701),
    .B(net4947));
 sg13g2_o21ai_1 _16593_ (.B1(_06852_),
    .Y(_01286_),
    .A1(net5494),
    .A2(net4947));
 sg13g2_nand2_1 _16594_ (.Y(_06853_),
    .A(net2463),
    .B(net4947));
 sg13g2_o21ai_1 _16595_ (.B1(_06853_),
    .Y(_01287_),
    .A1(net5539),
    .A2(net4947));
 sg13g2_nand2_1 _16596_ (.Y(_06854_),
    .A(net2146),
    .B(net4946));
 sg13g2_o21ai_1 _16597_ (.B1(_06854_),
    .Y(_01288_),
    .A1(net5583),
    .A2(net4947));
 sg13g2_nand2_1 _16598_ (.Y(_06855_),
    .A(net2144),
    .B(net4946));
 sg13g2_o21ai_1 _16599_ (.B1(_06855_),
    .Y(_01289_),
    .A1(net5630),
    .A2(_06850_));
 sg13g2_nand2_1 _16600_ (.Y(_06856_),
    .A(net3181),
    .B(net4946));
 sg13g2_o21ai_1 _16601_ (.B1(_06856_),
    .Y(_01290_),
    .A1(net5674),
    .A2(net4946));
 sg13g2_nand2_1 _16602_ (.Y(_06857_),
    .A(net3303),
    .B(net4946));
 sg13g2_o21ai_1 _16603_ (.B1(_06857_),
    .Y(_01291_),
    .A1(net5719),
    .A2(net4946));
 sg13g2_nand2_1 _16604_ (.Y(_06858_),
    .A(net2149),
    .B(net4946));
 sg13g2_o21ai_1 _16605_ (.B1(_06858_),
    .Y(_01292_),
    .A1(net5765),
    .A2(net4946));
 sg13g2_nor2_1 _16606_ (.A(net5143),
    .B(_03375_),
    .Y(_06859_));
 sg13g2_nor2_1 _16607_ (.A(net3584),
    .B(net4709),
    .Y(_06860_));
 sg13g2_a21oi_1 _16608_ (.A1(net5448),
    .A2(net4709),
    .Y(_01293_),
    .B1(_06860_));
 sg13g2_nor2_1 _16609_ (.A(net3598),
    .B(net4709),
    .Y(_06861_));
 sg13g2_a21oi_1 _16610_ (.A1(net5493),
    .A2(net4709),
    .Y(_01294_),
    .B1(_06861_));
 sg13g2_nor2_1 _16611_ (.A(net3510),
    .B(net4710),
    .Y(_06862_));
 sg13g2_a21oi_1 _16612_ (.A1(net5539),
    .A2(net4710),
    .Y(_01295_),
    .B1(_06862_));
 sg13g2_nor2_1 _16613_ (.A(net3531),
    .B(net4710),
    .Y(_06863_));
 sg13g2_a21oi_1 _16614_ (.A1(net5582),
    .A2(net4710),
    .Y(_01296_),
    .B1(_06863_));
 sg13g2_nor2_1 _16615_ (.A(net3522),
    .B(net4710),
    .Y(_06864_));
 sg13g2_a21oi_1 _16616_ (.A1(net5628),
    .A2(net4710),
    .Y(_01297_),
    .B1(_06864_));
 sg13g2_nor2_1 _16617_ (.A(net3641),
    .B(net4709),
    .Y(_06865_));
 sg13g2_a21oi_1 _16618_ (.A1(net5671),
    .A2(net4709),
    .Y(_01298_),
    .B1(_06865_));
 sg13g2_nor2_1 _16619_ (.A(net3516),
    .B(net4709),
    .Y(_06866_));
 sg13g2_a21oi_1 _16620_ (.A1(net5718),
    .A2(net4709),
    .Y(_01299_),
    .B1(_06866_));
 sg13g2_nor2_1 _16621_ (.A(net3412),
    .B(net4710),
    .Y(_06867_));
 sg13g2_a21oi_1 _16622_ (.A1(net5763),
    .A2(net4710),
    .Y(_01300_),
    .B1(_06867_));
 sg13g2_nand2_1 _16623_ (.Y(_06868_),
    .A(_03066_),
    .B(net5212));
 sg13g2_nand2_1 _16624_ (.Y(_06869_),
    .A(net2855),
    .B(net4944));
 sg13g2_o21ai_1 _16625_ (.B1(_06869_),
    .Y(_01301_),
    .A1(net5447),
    .A2(net4944));
 sg13g2_nand2_1 _16626_ (.Y(_06870_),
    .A(net2208),
    .B(net4945));
 sg13g2_o21ai_1 _16627_ (.B1(_06870_),
    .Y(_01302_),
    .A1(net5494),
    .A2(net4944));
 sg13g2_nand2_1 _16628_ (.Y(_06871_),
    .A(net2803),
    .B(net4944));
 sg13g2_o21ai_1 _16629_ (.B1(_06871_),
    .Y(_01303_),
    .A1(net5538),
    .A2(net4944));
 sg13g2_nand2_1 _16630_ (.Y(_06872_),
    .A(net3112),
    .B(net4944));
 sg13g2_o21ai_1 _16631_ (.B1(_06872_),
    .Y(_01304_),
    .A1(net5583),
    .A2(net4944));
 sg13g2_nand2_1 _16632_ (.Y(_06873_),
    .A(net3059),
    .B(net4945));
 sg13g2_o21ai_1 _16633_ (.B1(_06873_),
    .Y(_01305_),
    .A1(net5630),
    .A2(net4945));
 sg13g2_nand2_1 _16634_ (.Y(_06874_),
    .A(net2466),
    .B(net4945));
 sg13g2_o21ai_1 _16635_ (.B1(_06874_),
    .Y(_01306_),
    .A1(net5674),
    .A2(net4945));
 sg13g2_nand2_1 _16636_ (.Y(_06875_),
    .A(net3311),
    .B(net4945));
 sg13g2_o21ai_1 _16637_ (.B1(_06875_),
    .Y(_01307_),
    .A1(net5719),
    .A2(_06868_));
 sg13g2_nand2_1 _16638_ (.Y(_06876_),
    .A(net3027),
    .B(net4945));
 sg13g2_o21ai_1 _16639_ (.B1(_06876_),
    .Y(_01308_),
    .A1(net5763),
    .A2(net4944));
 sg13g2_nand2_1 _16640_ (.Y(_06877_),
    .A(net5238),
    .B(net5212));
 sg13g2_nand2_1 _16641_ (.Y(_06878_),
    .A(net2512),
    .B(net4942));
 sg13g2_o21ai_1 _16642_ (.B1(_06878_),
    .Y(_01309_),
    .A1(net5446),
    .A2(net4942));
 sg13g2_nand2_1 _16643_ (.Y(_06879_),
    .A(net3008),
    .B(net4942));
 sg13g2_o21ai_1 _16644_ (.B1(_06879_),
    .Y(_01310_),
    .A1(net5494),
    .A2(net4942));
 sg13g2_nand2_1 _16645_ (.Y(_06880_),
    .A(net2514),
    .B(net4942));
 sg13g2_o21ai_1 _16646_ (.B1(_06880_),
    .Y(_01311_),
    .A1(net5538),
    .A2(net4942));
 sg13g2_nand2_1 _16647_ (.Y(_06881_),
    .A(net2873),
    .B(net4943));
 sg13g2_o21ai_1 _16648_ (.B1(_06881_),
    .Y(_01312_),
    .A1(net5583),
    .A2(net4942));
 sg13g2_nand2_1 _16649_ (.Y(_06882_),
    .A(net2567),
    .B(net4943));
 sg13g2_o21ai_1 _16650_ (.B1(_06882_),
    .Y(_01313_),
    .A1(net5630),
    .A2(_06877_));
 sg13g2_nand2_1 _16651_ (.Y(_06883_),
    .A(net3310),
    .B(net4943));
 sg13g2_o21ai_1 _16652_ (.B1(_06883_),
    .Y(_01314_),
    .A1(net5674),
    .A2(net4943));
 sg13g2_nand2_1 _16653_ (.Y(_06884_),
    .A(net3784),
    .B(net4943));
 sg13g2_o21ai_1 _16654_ (.B1(_06884_),
    .Y(_01315_),
    .A1(net5719),
    .A2(net4943));
 sg13g2_nand2_1 _16655_ (.Y(_06885_),
    .A(net3038),
    .B(net4942));
 sg13g2_o21ai_1 _16656_ (.B1(_06885_),
    .Y(_01316_),
    .A1(net5763),
    .A2(net4943));
 sg13g2_nand2_1 _16657_ (.Y(_06886_),
    .A(_02938_),
    .B(net5211));
 sg13g2_nand2_1 _16658_ (.Y(_06887_),
    .A(net2493),
    .B(net4940));
 sg13g2_o21ai_1 _16659_ (.B1(_06887_),
    .Y(_01317_),
    .A1(net5441),
    .A2(net4940));
 sg13g2_nand2_1 _16660_ (.Y(_06888_),
    .A(net3184),
    .B(net4941));
 sg13g2_o21ai_1 _16661_ (.B1(_06888_),
    .Y(_01318_),
    .A1(net5489),
    .A2(net4941));
 sg13g2_nand2_1 _16662_ (.Y(_06889_),
    .A(net3418),
    .B(net4940));
 sg13g2_o21ai_1 _16663_ (.B1(_06889_),
    .Y(_01319_),
    .A1(net5535),
    .A2(net4940));
 sg13g2_nand2_1 _16664_ (.Y(_06890_),
    .A(net3400),
    .B(net4941));
 sg13g2_o21ai_1 _16665_ (.B1(_06890_),
    .Y(_01320_),
    .A1(net5580),
    .A2(net4941));
 sg13g2_nand2_1 _16666_ (.Y(_06891_),
    .A(net3094),
    .B(net4940));
 sg13g2_o21ai_1 _16667_ (.B1(_06891_),
    .Y(_01321_),
    .A1(net5626),
    .A2(net4940));
 sg13g2_nand2_1 _16668_ (.Y(_06892_),
    .A(net2901),
    .B(net4940));
 sg13g2_o21ai_1 _16669_ (.B1(_06892_),
    .Y(_01322_),
    .A1(net5668),
    .A2(net4940));
 sg13g2_nand2_1 _16670_ (.Y(_06893_),
    .A(net2890),
    .B(net4941));
 sg13g2_o21ai_1 _16671_ (.B1(_06893_),
    .Y(_01323_),
    .A1(net5716),
    .A2(net4941));
 sg13g2_nand2_1 _16672_ (.Y(_06894_),
    .A(net2256),
    .B(net4941));
 sg13g2_o21ai_1 _16673_ (.B1(_06894_),
    .Y(_01324_),
    .A1(net5761),
    .A2(net4941));
 sg13g2_nand2_1 _16674_ (.Y(_06895_),
    .A(_03016_),
    .B(net5211));
 sg13g2_nand2_1 _16675_ (.Y(_06896_),
    .A(net3035),
    .B(net4939));
 sg13g2_o21ai_1 _16676_ (.B1(_06896_),
    .Y(_01325_),
    .A1(net5441),
    .A2(net4939));
 sg13g2_nand2_1 _16677_ (.Y(_06897_),
    .A(net2436),
    .B(net4938));
 sg13g2_o21ai_1 _16678_ (.B1(_06897_),
    .Y(_01326_),
    .A1(net5489),
    .A2(net4938));
 sg13g2_nand2_1 _16679_ (.Y(_06898_),
    .A(net3457),
    .B(_06895_));
 sg13g2_o21ai_1 _16680_ (.B1(_06898_),
    .Y(_01327_),
    .A1(net5540),
    .A2(net4939));
 sg13g2_nand2_1 _16681_ (.Y(_06899_),
    .A(net2709),
    .B(net4939));
 sg13g2_o21ai_1 _16682_ (.B1(_06899_),
    .Y(_01328_),
    .A1(net5580),
    .A2(net4939));
 sg13g2_nand2_1 _16683_ (.Y(_06900_),
    .A(net2626),
    .B(net4938));
 sg13g2_o21ai_1 _16684_ (.B1(_06900_),
    .Y(_01329_),
    .A1(net5626),
    .A2(net4938));
 sg13g2_nand2_1 _16685_ (.Y(_06901_),
    .A(net3193),
    .B(net4938));
 sg13g2_o21ai_1 _16686_ (.B1(_06901_),
    .Y(_01330_),
    .A1(net5668),
    .A2(net4938));
 sg13g2_nand2_1 _16687_ (.Y(_06902_),
    .A(net3219),
    .B(net4938));
 sg13g2_o21ai_1 _16688_ (.B1(_06902_),
    .Y(_01331_),
    .A1(net5716),
    .A2(net4938));
 sg13g2_nand2_1 _16689_ (.Y(_06903_),
    .A(net3101),
    .B(net4939));
 sg13g2_o21ai_1 _16690_ (.B1(_06903_),
    .Y(_01332_),
    .A1(net5761),
    .A2(net4939));
 sg13g2_nand2_1 _16691_ (.Y(_06904_),
    .A(_02980_),
    .B(net5211));
 sg13g2_nand2_1 _16692_ (.Y(_06905_),
    .A(net2226),
    .B(net4936));
 sg13g2_o21ai_1 _16693_ (.B1(_06905_),
    .Y(_01333_),
    .A1(net5441),
    .A2(net4936));
 sg13g2_nand2_1 _16694_ (.Y(_06906_),
    .A(net2941),
    .B(net4937));
 sg13g2_o21ai_1 _16695_ (.B1(_06906_),
    .Y(_01334_),
    .A1(net5489),
    .A2(net4937));
 sg13g2_nand2_1 _16696_ (.Y(_06907_),
    .A(net2529),
    .B(net4936));
 sg13g2_o21ai_1 _16697_ (.B1(_06907_),
    .Y(_01335_),
    .A1(net5535),
    .A2(net4936));
 sg13g2_nand2_1 _16698_ (.Y(_06908_),
    .A(net3953),
    .B(net4937));
 sg13g2_o21ai_1 _16699_ (.B1(_06908_),
    .Y(_01336_),
    .A1(net5580),
    .A2(net4937));
 sg13g2_nand2_1 _16700_ (.Y(_06909_),
    .A(net2588),
    .B(net4936));
 sg13g2_o21ai_1 _16701_ (.B1(_06909_),
    .Y(_01337_),
    .A1(net5626),
    .A2(net4936));
 sg13g2_nand2_1 _16702_ (.Y(_06910_),
    .A(net2908),
    .B(net4936));
 sg13g2_o21ai_1 _16703_ (.B1(_06910_),
    .Y(_01338_),
    .A1(net5668),
    .A2(net4936));
 sg13g2_nand2_1 _16704_ (.Y(_06911_),
    .A(net2725),
    .B(net4937));
 sg13g2_o21ai_1 _16705_ (.B1(_06911_),
    .Y(_01339_),
    .A1(net5716),
    .A2(net4937));
 sg13g2_nand2_1 _16706_ (.Y(_06912_),
    .A(net2136),
    .B(net4937));
 sg13g2_o21ai_1 _16707_ (.B1(_06912_),
    .Y(_01340_),
    .A1(net5761),
    .A2(net4937));
 sg13g2_nand2_1 _16708_ (.Y(_06913_),
    .A(net5243),
    .B(net5211));
 sg13g2_nand2_1 _16709_ (.Y(_06914_),
    .A(net2985),
    .B(net4934));
 sg13g2_o21ai_1 _16710_ (.B1(_06914_),
    .Y(_01341_),
    .A1(net5441),
    .A2(net4934));
 sg13g2_nand2_1 _16711_ (.Y(_06915_),
    .A(net2783),
    .B(net4935));
 sg13g2_o21ai_1 _16712_ (.B1(_06915_),
    .Y(_01342_),
    .A1(net5489),
    .A2(net4935));
 sg13g2_nand2_1 _16713_ (.Y(_06916_),
    .A(net2622),
    .B(net4934));
 sg13g2_o21ai_1 _16714_ (.B1(_06916_),
    .Y(_01343_),
    .A1(net5535),
    .A2(net4934));
 sg13g2_nand2_1 _16715_ (.Y(_06917_),
    .A(net2923),
    .B(net4935));
 sg13g2_o21ai_1 _16716_ (.B1(_06917_),
    .Y(_01344_),
    .A1(net5580),
    .A2(net4935));
 sg13g2_nand2_1 _16717_ (.Y(_06918_),
    .A(net3232),
    .B(net4934));
 sg13g2_o21ai_1 _16718_ (.B1(_06918_),
    .Y(_01345_),
    .A1(net5626),
    .A2(net4934));
 sg13g2_nand2_1 _16719_ (.Y(_06919_),
    .A(net2628),
    .B(net4934));
 sg13g2_o21ai_1 _16720_ (.B1(_06919_),
    .Y(_01346_),
    .A1(net5668),
    .A2(net4934));
 sg13g2_nand2_1 _16721_ (.Y(_06920_),
    .A(net3041),
    .B(net4935));
 sg13g2_o21ai_1 _16722_ (.B1(_06920_),
    .Y(_01347_),
    .A1(net5716),
    .A2(net4935));
 sg13g2_nand2_1 _16723_ (.Y(_06921_),
    .A(net2779),
    .B(net4935));
 sg13g2_o21ai_1 _16724_ (.B1(_06921_),
    .Y(_01348_),
    .A1(net5761),
    .A2(net4935));
 sg13g2_nand2_1 _16725_ (.Y(_06922_),
    .A(net5211),
    .B(_03466_));
 sg13g2_nand2_1 _16726_ (.Y(_06923_),
    .A(net2265),
    .B(net4933));
 sg13g2_o21ai_1 _16727_ (.B1(_06923_),
    .Y(_01349_),
    .A1(net5447),
    .A2(net4933));
 sg13g2_nand2_1 _16728_ (.Y(_06924_),
    .A(net3582),
    .B(net4932));
 sg13g2_o21ai_1 _16729_ (.B1(_06924_),
    .Y(_01350_),
    .A1(net5496),
    .A2(net4932));
 sg13g2_nand2_1 _16730_ (.Y(_06925_),
    .A(net3200),
    .B(net4932));
 sg13g2_o21ai_1 _16731_ (.B1(_06925_),
    .Y(_01351_),
    .A1(net5538),
    .A2(net4933));
 sg13g2_nand2_1 _16732_ (.Y(_06926_),
    .A(net3072),
    .B(_06922_));
 sg13g2_o21ai_1 _16733_ (.B1(_06926_),
    .Y(_01352_),
    .A1(net5584),
    .A2(net4932));
 sg13g2_nand2_1 _16734_ (.Y(_06927_),
    .A(net2311),
    .B(net4933));
 sg13g2_o21ai_1 _16735_ (.B1(_06927_),
    .Y(_01353_),
    .A1(net5620),
    .A2(net4933));
 sg13g2_nand2_1 _16736_ (.Y(_06928_),
    .A(net3168),
    .B(net4933));
 sg13g2_o21ai_1 _16737_ (.B1(_06928_),
    .Y(_01354_),
    .A1(net5670),
    .A2(net4933));
 sg13g2_nand2_1 _16738_ (.Y(_06929_),
    .A(net2991),
    .B(net4932));
 sg13g2_o21ai_1 _16739_ (.B1(_06929_),
    .Y(_01355_),
    .A1(net5719),
    .A2(net4932));
 sg13g2_nand2_1 _16740_ (.Y(_06930_),
    .A(net2159),
    .B(net4932));
 sg13g2_o21ai_1 _16741_ (.B1(_06930_),
    .Y(_01356_),
    .A1(net5765),
    .A2(net4932));
 sg13g2_nand2_1 _16742_ (.Y(_06931_),
    .A(net5251),
    .B(net5211));
 sg13g2_nand2_1 _16743_ (.Y(_06932_),
    .A(net2333),
    .B(net4930));
 sg13g2_o21ai_1 _16744_ (.B1(_06932_),
    .Y(_01357_),
    .A1(net5447),
    .A2(net4930));
 sg13g2_nand2_1 _16745_ (.Y(_06933_),
    .A(net2765),
    .B(net4931));
 sg13g2_o21ai_1 _16746_ (.B1(_06933_),
    .Y(_01358_),
    .A1(net5496),
    .A2(net4931));
 sg13g2_nand2_1 _16747_ (.Y(_06934_),
    .A(net2408),
    .B(net4930));
 sg13g2_o21ai_1 _16748_ (.B1(_06934_),
    .Y(_01359_),
    .A1(net5538),
    .A2(net4930));
 sg13g2_nand2_1 _16749_ (.Y(_06935_),
    .A(net3394),
    .B(net4931));
 sg13g2_o21ai_1 _16750_ (.B1(_06935_),
    .Y(_01360_),
    .A1(net5584),
    .A2(net4931));
 sg13g2_nand2_1 _16751_ (.Y(_06936_),
    .A(net2778),
    .B(net4930));
 sg13g2_o21ai_1 _16752_ (.B1(_06936_),
    .Y(_01361_),
    .A1(net5620),
    .A2(net4930));
 sg13g2_nand2_1 _16753_ (.Y(_06937_),
    .A(net3334),
    .B(net4930));
 sg13g2_o21ai_1 _16754_ (.B1(_06937_),
    .Y(_01362_),
    .A1(net5674),
    .A2(net4930));
 sg13g2_nand2_1 _16755_ (.Y(_06938_),
    .A(net2524),
    .B(net4931));
 sg13g2_o21ai_1 _16756_ (.B1(_06938_),
    .Y(_01363_),
    .A1(net5719),
    .A2(net4931));
 sg13g2_nand2_1 _16757_ (.Y(_06939_),
    .A(net3348),
    .B(net4931));
 sg13g2_o21ai_1 _16758_ (.B1(_06939_),
    .Y(_01364_),
    .A1(net5765),
    .A2(net4931));
 sg13g2_nand2_1 _16759_ (.Y(_06940_),
    .A(net5211),
    .B(net5247));
 sg13g2_nand2_1 _16760_ (.Y(_06941_),
    .A(net2470),
    .B(net4928));
 sg13g2_o21ai_1 _16761_ (.B1(_06941_),
    .Y(_01365_),
    .A1(net5446),
    .A2(net4928));
 sg13g2_nand2_1 _16762_ (.Y(_06942_),
    .A(net2158),
    .B(net4929));
 sg13g2_o21ai_1 _16763_ (.B1(_06942_),
    .Y(_01366_),
    .A1(net5489),
    .A2(net4929));
 sg13g2_nand2_1 _16764_ (.Y(_06943_),
    .A(net2772),
    .B(net4928));
 sg13g2_o21ai_1 _16765_ (.B1(_06943_),
    .Y(_01367_),
    .A1(net5538),
    .A2(net4928));
 sg13g2_nand2_1 _16766_ (.Y(_06944_),
    .A(net2900),
    .B(net4929));
 sg13g2_o21ai_1 _16767_ (.B1(_06944_),
    .Y(_01368_),
    .A1(net5584),
    .A2(net4929));
 sg13g2_nand2_1 _16768_ (.Y(_06945_),
    .A(net3255),
    .B(net4928));
 sg13g2_o21ai_1 _16769_ (.B1(_06945_),
    .Y(_01369_),
    .A1(net5620),
    .A2(net4928));
 sg13g2_nand2_1 _16770_ (.Y(_06946_),
    .A(net2608),
    .B(net4928));
 sg13g2_o21ai_1 _16771_ (.B1(_06946_),
    .Y(_01370_),
    .A1(net5674),
    .A2(net4928));
 sg13g2_nand2_1 _16772_ (.Y(_06947_),
    .A(net2289),
    .B(net4929));
 sg13g2_o21ai_1 _16773_ (.B1(_06947_),
    .Y(_01371_),
    .A1(net5719),
    .A2(net4929));
 sg13g2_nand2_1 _16774_ (.Y(_06948_),
    .A(net2216),
    .B(net4929));
 sg13g2_o21ai_1 _16775_ (.B1(_06948_),
    .Y(_01372_),
    .A1(net5761),
    .A2(net4929));
 sg13g2_nor2_1 _16776_ (.A(net5240),
    .B(net5143),
    .Y(_06949_));
 sg13g2_nor2_1 _16777_ (.A(net4109),
    .B(net4707),
    .Y(_06950_));
 sg13g2_a21oi_1 _16778_ (.A1(net5448),
    .A2(net4707),
    .Y(_01373_),
    .B1(_06950_));
 sg13g2_nor2_1 _16779_ (.A(net3892),
    .B(net4707),
    .Y(_06951_));
 sg13g2_a21oi_1 _16780_ (.A1(net5493),
    .A2(net4707),
    .Y(_01374_),
    .B1(_06951_));
 sg13g2_nor2_1 _16781_ (.A(net3693),
    .B(net4708),
    .Y(_06952_));
 sg13g2_a21oi_1 _16782_ (.A1(net5539),
    .A2(net4708),
    .Y(_01375_),
    .B1(_06952_));
 sg13g2_nor2_1 _16783_ (.A(net3458),
    .B(net4708),
    .Y(_06953_));
 sg13g2_a21oi_1 _16784_ (.A1(net5582),
    .A2(net4708),
    .Y(_01376_),
    .B1(_06953_));
 sg13g2_nor2_1 _16785_ (.A(net4079),
    .B(net4708),
    .Y(_06954_));
 sg13g2_a21oi_1 _16786_ (.A1(net5628),
    .A2(net4708),
    .Y(_01377_),
    .B1(_06954_));
 sg13g2_nor2_1 _16787_ (.A(net3829),
    .B(net4707),
    .Y(_06955_));
 sg13g2_a21oi_1 _16788_ (.A1(net5671),
    .A2(net4707),
    .Y(_01378_),
    .B1(_06955_));
 sg13g2_nor2_1 _16789_ (.A(net3764),
    .B(net4707),
    .Y(_06956_));
 sg13g2_a21oi_1 _16790_ (.A1(net5718),
    .A2(net4707),
    .Y(_01379_),
    .B1(_06956_));
 sg13g2_nor2_1 _16791_ (.A(net3975),
    .B(net4708),
    .Y(_06957_));
 sg13g2_a21oi_1 _16792_ (.A1(net5763),
    .A2(net4708),
    .Y(_01380_),
    .B1(_06957_));
 sg13g2_nand2_2 _16793_ (.Y(_06958_),
    .A(net5248),
    .B(net5194));
 sg13g2_nand2_1 _16794_ (.Y(_06959_),
    .A(net3759),
    .B(net4926));
 sg13g2_o21ai_1 _16795_ (.B1(_06959_),
    .Y(_01381_),
    .A1(net5431),
    .A2(net4926));
 sg13g2_nand2_1 _16796_ (.Y(_06960_),
    .A(net3150),
    .B(net4927));
 sg13g2_o21ai_1 _16797_ (.B1(_06960_),
    .Y(_01382_),
    .A1(net5485),
    .A2(net4927));
 sg13g2_nand2_1 _16798_ (.Y(_06961_),
    .A(net2655),
    .B(net4926));
 sg13g2_o21ai_1 _16799_ (.B1(_06961_),
    .Y(_01383_),
    .A1(net5532),
    .A2(net4926));
 sg13g2_nand2_1 _16800_ (.Y(_06962_),
    .A(net2603),
    .B(net4927));
 sg13g2_o21ai_1 _16801_ (.B1(_06962_),
    .Y(_01384_),
    .A1(net5575),
    .A2(_06958_));
 sg13g2_nand2_1 _16802_ (.Y(_06963_),
    .A(net2700),
    .B(net4926));
 sg13g2_o21ai_1 _16803_ (.B1(_06963_),
    .Y(_01385_),
    .A1(net5623),
    .A2(net4926));
 sg13g2_nand2_1 _16804_ (.Y(_06964_),
    .A(net2551),
    .B(net4927));
 sg13g2_o21ai_1 _16805_ (.B1(_06964_),
    .Y(_01386_),
    .A1(net5666),
    .A2(net4927));
 sg13g2_nand2_1 _16806_ (.Y(_06965_),
    .A(net3142),
    .B(net4927));
 sg13g2_o21ai_1 _16807_ (.B1(_06965_),
    .Y(_01387_),
    .A1(net5710),
    .A2(net4927));
 sg13g2_nand2_1 _16808_ (.Y(_06966_),
    .A(net2180),
    .B(net4926));
 sg13g2_o21ai_1 _16809_ (.B1(_06966_),
    .Y(_01388_),
    .A1(net5757),
    .A2(net4926));
 sg13g2_nor3_2 _16810_ (.A(net5227),
    .B(_03140_),
    .C(net5258),
    .Y(_06967_));
 sg13g2_nor2_1 _16811_ (.A(net3396),
    .B(net5178),
    .Y(_06968_));
 sg13g2_a21oi_1 _16812_ (.A1(net5440),
    .A2(net5178),
    .Y(_01389_),
    .B1(_06968_));
 sg13g2_nor2_1 _16813_ (.A(net4033),
    .B(net5179),
    .Y(_06969_));
 sg13g2_a21oi_1 _16814_ (.A1(net5485),
    .A2(net5179),
    .Y(_01390_),
    .B1(_06969_));
 sg13g2_nor2_1 _16815_ (.A(net3937),
    .B(net5178),
    .Y(_06970_));
 sg13g2_a21oi_1 _16816_ (.A1(net5532),
    .A2(net5178),
    .Y(_01391_),
    .B1(_06970_));
 sg13g2_nor2_1 _16817_ (.A(net4047),
    .B(net5179),
    .Y(_06971_));
 sg13g2_a21oi_1 _16818_ (.A1(net5575),
    .A2(net5179),
    .Y(_01392_),
    .B1(_06971_));
 sg13g2_nor2_1 _16819_ (.A(net3519),
    .B(net5178),
    .Y(_06972_));
 sg13g2_a21oi_1 _16820_ (.A1(net5623),
    .A2(net5178),
    .Y(_01393_),
    .B1(_06972_));
 sg13g2_nor2_1 _16821_ (.A(net3854),
    .B(net5179),
    .Y(_06973_));
 sg13g2_a21oi_1 _16822_ (.A1(net5666),
    .A2(net5179),
    .Y(_01394_),
    .B1(_06973_));
 sg13g2_nor2_1 _16823_ (.A(net3736),
    .B(net5179),
    .Y(_06974_));
 sg13g2_a21oi_1 _16824_ (.A1(net5711),
    .A2(net5179),
    .Y(_01395_),
    .B1(_06974_));
 sg13g2_nor2_1 _16825_ (.A(net3852),
    .B(net5178),
    .Y(_06975_));
 sg13g2_a21oi_1 _16826_ (.A1(net5757),
    .A2(net5178),
    .Y(_01396_),
    .B1(_06975_));
 sg13g2_nor3_2 _16827_ (.A(net5227),
    .B(_03080_),
    .C(net5258),
    .Y(_06976_));
 sg13g2_nor2_1 _16828_ (.A(net3652),
    .B(net5176),
    .Y(_06977_));
 sg13g2_a21oi_1 _16829_ (.A1(net5440),
    .A2(net5176),
    .Y(_01397_),
    .B1(_06977_));
 sg13g2_nor2_1 _16830_ (.A(net3476),
    .B(net5176),
    .Y(_06978_));
 sg13g2_a21oi_1 _16831_ (.A1(net5485),
    .A2(net5176),
    .Y(_01398_),
    .B1(_06978_));
 sg13g2_nor2_1 _16832_ (.A(net3475),
    .B(net5176),
    .Y(_06979_));
 sg13g2_a21oi_1 _16833_ (.A1(net5532),
    .A2(net5176),
    .Y(_01399_),
    .B1(_06979_));
 sg13g2_nor2_1 _16834_ (.A(net3367),
    .B(net5177),
    .Y(_06980_));
 sg13g2_a21oi_1 _16835_ (.A1(net5575),
    .A2(_06976_),
    .Y(_01400_),
    .B1(_06980_));
 sg13g2_nor2_1 _16836_ (.A(net3851),
    .B(net5176),
    .Y(_06981_));
 sg13g2_a21oi_1 _16837_ (.A1(net5623),
    .A2(net5177),
    .Y(_01401_),
    .B1(_06981_));
 sg13g2_nor2_1 _16838_ (.A(net4095),
    .B(net5177),
    .Y(_06982_));
 sg13g2_a21oi_1 _16839_ (.A1(net5666),
    .A2(net5177),
    .Y(_01402_),
    .B1(_06982_));
 sg13g2_nor2_1 _16840_ (.A(net3987),
    .B(net5177),
    .Y(_06983_));
 sg13g2_a21oi_1 _16841_ (.A1(net5711),
    .A2(net5177),
    .Y(_01403_),
    .B1(_06983_));
 sg13g2_nor2_1 _16842_ (.A(net3165),
    .B(net5177),
    .Y(_06984_));
 sg13g2_a21oi_1 _16843_ (.A1(net5757),
    .A2(net5176),
    .Y(_01404_),
    .B1(_06984_));
 sg13g2_nand2_2 _16844_ (.Y(_06985_),
    .A(_03119_),
    .B(net5194));
 sg13g2_nand2_1 _16845_ (.Y(_06986_),
    .A(net3266),
    .B(net4924));
 sg13g2_o21ai_1 _16846_ (.B1(_06986_),
    .Y(_01405_),
    .A1(net5440),
    .A2(net4924));
 sg13g2_nand2_1 _16847_ (.Y(_06987_),
    .A(net2367),
    .B(net4924));
 sg13g2_o21ai_1 _16848_ (.B1(_06987_),
    .Y(_01406_),
    .A1(net5485),
    .A2(net4924));
 sg13g2_nand2_1 _16849_ (.Y(_06988_),
    .A(net3018),
    .B(net4924));
 sg13g2_o21ai_1 _16850_ (.B1(_06988_),
    .Y(_01407_),
    .A1(net5532),
    .A2(net4924));
 sg13g2_nand2_1 _16851_ (.Y(_06989_),
    .A(net2375),
    .B(_06985_));
 sg13g2_o21ai_1 _16852_ (.B1(_06989_),
    .Y(_01408_),
    .A1(net5575),
    .A2(net4925));
 sg13g2_nand2_1 _16853_ (.Y(_06990_),
    .A(net2614),
    .B(net4925));
 sg13g2_o21ai_1 _16854_ (.B1(_06990_),
    .Y(_01409_),
    .A1(net5623),
    .A2(net4925));
 sg13g2_nand2_1 _16855_ (.Y(_06991_),
    .A(net2921),
    .B(net4925));
 sg13g2_o21ai_1 _16856_ (.B1(_06991_),
    .Y(_01410_),
    .A1(net5666),
    .A2(net4925));
 sg13g2_nand2_1 _16857_ (.Y(_06992_),
    .A(net2548),
    .B(net4925));
 sg13g2_o21ai_1 _16858_ (.B1(_06992_),
    .Y(_01411_),
    .A1(net5711),
    .A2(net4925));
 sg13g2_nand2_1 _16859_ (.Y(_06993_),
    .A(net3117),
    .B(net4924));
 sg13g2_o21ai_1 _16860_ (.B1(_06993_),
    .Y(_01412_),
    .A1(net5757),
    .A2(net4924));
 sg13g2_nand2_1 _16861_ (.Y(_06994_),
    .A(net5235),
    .B(net5195));
 sg13g2_nand2_1 _16862_ (.Y(_06995_),
    .A(net2579),
    .B(net4922));
 sg13g2_o21ai_1 _16863_ (.B1(_06995_),
    .Y(_01413_),
    .A1(net5440),
    .A2(net4922));
 sg13g2_nand2_1 _16864_ (.Y(_06996_),
    .A(net2726),
    .B(_06994_));
 sg13g2_o21ai_1 _16865_ (.B1(_06996_),
    .Y(_01414_),
    .A1(net5488),
    .A2(net4923));
 sg13g2_nand2_1 _16866_ (.Y(_06997_),
    .A(net2963),
    .B(net4922));
 sg13g2_o21ai_1 _16867_ (.B1(_06997_),
    .Y(_01415_),
    .A1(net5532),
    .A2(net4922));
 sg13g2_nand2_1 _16868_ (.Y(_06998_),
    .A(net2163),
    .B(net4922));
 sg13g2_o21ai_1 _16869_ (.B1(_06998_),
    .Y(_01416_),
    .A1(net5577),
    .A2(net4922));
 sg13g2_nand2_1 _16870_ (.Y(_06999_),
    .A(net2762),
    .B(net4923));
 sg13g2_o21ai_1 _16871_ (.B1(_06999_),
    .Y(_01417_),
    .A1(net5622),
    .A2(net4923));
 sg13g2_nand2_1 _16872_ (.Y(_07000_),
    .A(net2877),
    .B(net4923));
 sg13g2_o21ai_1 _16873_ (.B1(_07000_),
    .Y(_01418_),
    .A1(net5665),
    .A2(net4923));
 sg13g2_nand2_1 _16874_ (.Y(_07001_),
    .A(net3162),
    .B(net4923));
 sg13g2_o21ai_1 _16875_ (.B1(_07001_),
    .Y(_01419_),
    .A1(net5712),
    .A2(net4923));
 sg13g2_nand2_1 _16876_ (.Y(_07002_),
    .A(net2166),
    .B(net4922));
 sg13g2_o21ai_1 _16877_ (.B1(_07002_),
    .Y(_01420_),
    .A1(net5757),
    .A2(net4922));
 sg13g2_nand2_1 _16878_ (.Y(_07003_),
    .A(net5234),
    .B(net5195));
 sg13g2_nand2_1 _16879_ (.Y(_07004_),
    .A(net2684),
    .B(net4920));
 sg13g2_o21ai_1 _16880_ (.B1(_07004_),
    .Y(_01421_),
    .A1(net5440),
    .A2(net4920));
 sg13g2_nand2_1 _16881_ (.Y(_07005_),
    .A(net2751),
    .B(_07003_));
 sg13g2_o21ai_1 _16882_ (.B1(_07005_),
    .Y(_01422_),
    .A1(net5487),
    .A2(net4921));
 sg13g2_nand2_1 _16883_ (.Y(_07006_),
    .A(net2716),
    .B(net4920));
 sg13g2_o21ai_1 _16884_ (.B1(_07006_),
    .Y(_01423_),
    .A1(net5532),
    .A2(net4920));
 sg13g2_nand2_1 _16885_ (.Y(_07007_),
    .A(net2429),
    .B(net4920));
 sg13g2_o21ai_1 _16886_ (.B1(_07007_),
    .Y(_01424_),
    .A1(net5577),
    .A2(net4920));
 sg13g2_nand2_1 _16887_ (.Y(_07008_),
    .A(net2388),
    .B(net4921));
 sg13g2_o21ai_1 _16888_ (.B1(_07008_),
    .Y(_01425_),
    .A1(net5622),
    .A2(net4921));
 sg13g2_nand2_1 _16889_ (.Y(_07009_),
    .A(net2797),
    .B(net4921));
 sg13g2_o21ai_1 _16890_ (.B1(_07009_),
    .Y(_01426_),
    .A1(net5665),
    .A2(net4921));
 sg13g2_nand2_1 _16891_ (.Y(_07010_),
    .A(net3202),
    .B(net4921));
 sg13g2_o21ai_1 _16892_ (.B1(_07010_),
    .Y(_01427_),
    .A1(net5712),
    .A2(net4921));
 sg13g2_nand2_1 _16893_ (.Y(_07011_),
    .A(net3239),
    .B(net4920));
 sg13g2_o21ai_1 _16894_ (.B1(_07011_),
    .Y(_01428_),
    .A1(net5757),
    .A2(net4920));
 sg13g2_nand2_1 _16895_ (.Y(_07012_),
    .A(net5236),
    .B(net5195));
 sg13g2_nand2_1 _16896_ (.Y(_07013_),
    .A(net2313),
    .B(net4918));
 sg13g2_o21ai_1 _16897_ (.B1(_07013_),
    .Y(_01429_),
    .A1(net5441),
    .A2(net4918));
 sg13g2_nand2_1 _16898_ (.Y(_07014_),
    .A(net2301),
    .B(net4919));
 sg13g2_o21ai_1 _16899_ (.B1(_07014_),
    .Y(_01430_),
    .A1(net5487),
    .A2(net4919));
 sg13g2_nand2_1 _16900_ (.Y(_07015_),
    .A(net2874),
    .B(net4918));
 sg13g2_o21ai_1 _16901_ (.B1(_07015_),
    .Y(_01431_),
    .A1(net5521),
    .A2(net4918));
 sg13g2_nand2_1 _16902_ (.Y(_07016_),
    .A(net2170),
    .B(net4918));
 sg13g2_o21ai_1 _16903_ (.B1(_07016_),
    .Y(_01432_),
    .A1(net5587),
    .A2(net4918));
 sg13g2_nand2_1 _16904_ (.Y(_07017_),
    .A(net2805),
    .B(net4919));
 sg13g2_o21ai_1 _16905_ (.B1(_07017_),
    .Y(_01433_),
    .A1(net5622),
    .A2(net4919));
 sg13g2_nand2_1 _16906_ (.Y(_07018_),
    .A(net2485),
    .B(net4919));
 sg13g2_o21ai_1 _16907_ (.B1(_07018_),
    .Y(_01434_),
    .A1(net5665),
    .A2(net4919));
 sg13g2_nand2_1 _16908_ (.Y(_07019_),
    .A(net3258),
    .B(net4918));
 sg13g2_o21ai_1 _16909_ (.B1(_07019_),
    .Y(_01435_),
    .A1(net5712),
    .A2(net4918));
 sg13g2_nor2_1 _16910_ (.A(\mem.data_in[7] ),
    .B(net4919),
    .Y(_07020_));
 sg13g2_a21oi_1 _16911_ (.A1(_02879_),
    .A2(net4919),
    .Y(_01436_),
    .B1(_07020_));
 sg13g2_nand2_1 _16912_ (.Y(_07021_),
    .A(net5237),
    .B(net5194));
 sg13g2_nand2_1 _16913_ (.Y(_07022_),
    .A(net3138),
    .B(net4916));
 sg13g2_o21ai_1 _16914_ (.B1(_07022_),
    .Y(_01437_),
    .A1(net5441),
    .A2(net4916));
 sg13g2_nand2_1 _16915_ (.Y(_07023_),
    .A(net3169),
    .B(net4917));
 sg13g2_o21ai_1 _16916_ (.B1(_07023_),
    .Y(_01438_),
    .A1(net5487),
    .A2(net4917));
 sg13g2_nand2_1 _16917_ (.Y(_07024_),
    .A(net2492),
    .B(net4916));
 sg13g2_o21ai_1 _16918_ (.B1(_07024_),
    .Y(_01439_),
    .A1(net5532),
    .A2(net4916));
 sg13g2_nand2_1 _16919_ (.Y(_07025_),
    .A(net3148),
    .B(net4916));
 sg13g2_o21ai_1 _16920_ (.B1(_07025_),
    .Y(_01440_),
    .A1(net5577),
    .A2(net4916));
 sg13g2_nand2_1 _16921_ (.Y(_07026_),
    .A(net3260),
    .B(net4917));
 sg13g2_o21ai_1 _16922_ (.B1(_07026_),
    .Y(_01441_),
    .A1(net5622),
    .A2(net4917));
 sg13g2_nand2_1 _16923_ (.Y(_07027_),
    .A(net2553),
    .B(net4917));
 sg13g2_o21ai_1 _16924_ (.B1(_07027_),
    .Y(_01442_),
    .A1(net5665),
    .A2(net4917));
 sg13g2_nand2_1 _16925_ (.Y(_07028_),
    .A(net3192),
    .B(net4916));
 sg13g2_o21ai_1 _16926_ (.B1(_07028_),
    .Y(_01443_),
    .A1(net5712),
    .A2(net4916));
 sg13g2_nand2_1 _16927_ (.Y(_07029_),
    .A(net3351),
    .B(net4917));
 sg13g2_o21ai_1 _16928_ (.B1(_07029_),
    .Y(_01444_),
    .A1(net5758),
    .A2(net4917));
 sg13g2_nand2_1 _16929_ (.Y(_07030_),
    .A(net5244),
    .B(net5194));
 sg13g2_nand2_1 _16930_ (.Y(_07031_),
    .A(net2488),
    .B(net4914));
 sg13g2_o21ai_1 _16931_ (.B1(_07031_),
    .Y(_01445_),
    .A1(net5440),
    .A2(net4914));
 sg13g2_nand2_1 _16932_ (.Y(_07032_),
    .A(net2816),
    .B(net4915));
 sg13g2_o21ai_1 _16933_ (.B1(_07032_),
    .Y(_01446_),
    .A1(net5485),
    .A2(net4915));
 sg13g2_nand2_1 _16934_ (.Y(_07033_),
    .A(net2412),
    .B(net4915));
 sg13g2_o21ai_1 _16935_ (.B1(_07033_),
    .Y(_01447_),
    .A1(net5533),
    .A2(net4915));
 sg13g2_nand2_1 _16936_ (.Y(_07034_),
    .A(net2153),
    .B(_07030_));
 sg13g2_o21ai_1 _16937_ (.B1(_07034_),
    .Y(_01448_),
    .A1(net5576),
    .A2(net4915));
 sg13g2_nand2_1 _16938_ (.Y(_07035_),
    .A(net2617),
    .B(net4915));
 sg13g2_o21ai_1 _16939_ (.B1(_07035_),
    .Y(_01449_),
    .A1(net5621),
    .A2(net4915));
 sg13g2_nand2_1 _16940_ (.Y(_07036_),
    .A(net3375),
    .B(net4914));
 sg13g2_o21ai_1 _16941_ (.B1(_07036_),
    .Y(_01450_),
    .A1(net5665),
    .A2(net4914));
 sg13g2_nand2_1 _16942_ (.Y(_07037_),
    .A(net3488),
    .B(net4914));
 sg13g2_o21ai_1 _16943_ (.B1(_07037_),
    .Y(_01451_),
    .A1(net5711),
    .A2(net4914));
 sg13g2_nand2_1 _16944_ (.Y(_07038_),
    .A(net3208),
    .B(net4914));
 sg13g2_o21ai_1 _16945_ (.B1(_07038_),
    .Y(_01452_),
    .A1(net5758),
    .A2(net4914));
 sg13g2_nand2_1 _16946_ (.Y(_07039_),
    .A(net5249),
    .B(_03363_));
 sg13g2_nor2_1 _16947_ (.A(\mem.data_in[0] ),
    .B(net4912),
    .Y(_07040_));
 sg13g2_a21oi_1 _16948_ (.A1(_02885_),
    .A2(net4912),
    .Y(_01453_),
    .B1(_07040_));
 sg13g2_nand2_1 _16949_ (.Y(_07041_),
    .A(net2854),
    .B(net4912));
 sg13g2_o21ai_1 _16950_ (.B1(_07041_),
    .Y(_01454_),
    .A1(net5498),
    .A2(net4912));
 sg13g2_nand2_1 _16951_ (.Y(_07042_),
    .A(net3174),
    .B(net4912));
 sg13g2_o21ai_1 _16952_ (.B1(_07042_),
    .Y(_01455_),
    .A1(net5541),
    .A2(net4912));
 sg13g2_nand2_1 _16953_ (.Y(_07043_),
    .A(net2929),
    .B(net4913));
 sg13g2_o21ai_1 _16954_ (.B1(_07043_),
    .Y(_01456_),
    .A1(net5596),
    .A2(net4913));
 sg13g2_nand2_1 _16955_ (.Y(_07044_),
    .A(net2296),
    .B(net4913));
 sg13g2_o21ai_1 _16956_ (.B1(_07044_),
    .Y(_01457_),
    .A1(net5641),
    .A2(net4913));
 sg13g2_nand2_1 _16957_ (.Y(_07045_),
    .A(net2278),
    .B(net4913));
 sg13g2_o21ai_1 _16958_ (.B1(_07045_),
    .Y(_01458_),
    .A1(net5692),
    .A2(net4913));
 sg13g2_nand2_1 _16959_ (.Y(_07046_),
    .A(net3106),
    .B(net4913));
 sg13g2_o21ai_1 _16960_ (.B1(_07046_),
    .Y(_01459_),
    .A1(net5732),
    .A2(net4913));
 sg13g2_nand2_1 _16961_ (.Y(_07047_),
    .A(net2331),
    .B(net4912));
 sg13g2_o21ai_1 _16962_ (.B1(_07047_),
    .Y(_01460_),
    .A1(net5767),
    .A2(net4912));
 sg13g2_nand2_1 _16963_ (.Y(_07048_),
    .A(net5242),
    .B(net5194));
 sg13g2_nand2_1 _16964_ (.Y(_07049_),
    .A(net2949),
    .B(net4910));
 sg13g2_o21ai_1 _16965_ (.B1(_07049_),
    .Y(_01461_),
    .A1(net5442),
    .A2(net4910));
 sg13g2_nand2_1 _16966_ (.Y(_07050_),
    .A(net2903),
    .B(net4911));
 sg13g2_o21ai_1 _16967_ (.B1(_07050_),
    .Y(_01462_),
    .A1(net5485),
    .A2(net4911));
 sg13g2_nand2_1 _16968_ (.Y(_07051_),
    .A(net3036),
    .B(_07048_));
 sg13g2_o21ai_1 _16969_ (.B1(_07051_),
    .Y(_01463_),
    .A1(net5533),
    .A2(net4911));
 sg13g2_nand2_1 _16970_ (.Y(_07052_),
    .A(net2143),
    .B(net4910));
 sg13g2_o21ai_1 _16971_ (.B1(_07052_),
    .Y(_01464_),
    .A1(net5575),
    .A2(net4910));
 sg13g2_nand2_1 _16972_ (.Y(_07053_),
    .A(net2745),
    .B(net4910));
 sg13g2_o21ai_1 _16973_ (.B1(_07053_),
    .Y(_01465_),
    .A1(net5623),
    .A2(net4910));
 sg13g2_nand2_1 _16974_ (.Y(_07054_),
    .A(net2720),
    .B(net4911));
 sg13g2_o21ai_1 _16975_ (.B1(_07054_),
    .Y(_01466_),
    .A1(net5666),
    .A2(net4911));
 sg13g2_nand2_1 _16976_ (.Y(_07055_),
    .A(net2526),
    .B(net4911));
 sg13g2_o21ai_1 _16977_ (.B1(_07055_),
    .Y(_01467_),
    .A1(net5710),
    .A2(net4911));
 sg13g2_nand2_1 _16978_ (.Y(_07056_),
    .A(net2925),
    .B(net4910));
 sg13g2_o21ai_1 _16979_ (.B1(_07056_),
    .Y(_01468_),
    .A1(net5757),
    .A2(net4910));
 sg13g2_nand2_1 _16980_ (.Y(_07057_),
    .A(net5243),
    .B(net5194));
 sg13g2_nand2_1 _16981_ (.Y(_07058_),
    .A(net2552),
    .B(net4909));
 sg13g2_o21ai_1 _16982_ (.B1(_07058_),
    .Y(_01469_),
    .A1(net5440),
    .A2(net4908));
 sg13g2_nand2_1 _16983_ (.Y(_07059_),
    .A(net2507),
    .B(net4908));
 sg13g2_o21ai_1 _16984_ (.B1(_07059_),
    .Y(_01470_),
    .A1(net5485),
    .A2(net4908));
 sg13g2_nand2_1 _16985_ (.Y(_07060_),
    .A(net3039),
    .B(net4909));
 sg13g2_o21ai_1 _16986_ (.B1(_07060_),
    .Y(_01471_),
    .A1(net5533),
    .A2(net4909));
 sg13g2_nand2_1 _16987_ (.Y(_07061_),
    .A(net2856),
    .B(net4909));
 sg13g2_o21ai_1 _16988_ (.B1(_07061_),
    .Y(_01472_),
    .A1(net5576),
    .A2(net4908));
 sg13g2_nand2_1 _16989_ (.Y(_07062_),
    .A(net3312),
    .B(net4909));
 sg13g2_o21ai_1 _16990_ (.B1(_07062_),
    .Y(_01473_),
    .A1(net5623),
    .A2(net4909));
 sg13g2_nand2_1 _16991_ (.Y(_07063_),
    .A(net2787),
    .B(net4908));
 sg13g2_o21ai_1 _16992_ (.B1(_07063_),
    .Y(_01474_),
    .A1(net5666),
    .A2(net4908));
 sg13g2_nand2_1 _16993_ (.Y(_07064_),
    .A(net2852),
    .B(net4908));
 sg13g2_o21ai_1 _16994_ (.B1(_07064_),
    .Y(_01475_),
    .A1(net5710),
    .A2(net4908));
 sg13g2_nand2_1 _16995_ (.Y(_07065_),
    .A(net2535),
    .B(net4909));
 sg13g2_o21ai_1 _16996_ (.B1(_07065_),
    .Y(_01476_),
    .A1(net5757),
    .A2(net4909));
 sg13g2_nand2_1 _16997_ (.Y(_07066_),
    .A(net5245),
    .B(net5195));
 sg13g2_nand2_1 _16998_ (.Y(_07067_),
    .A(net2671),
    .B(net4906));
 sg13g2_o21ai_1 _16999_ (.B1(_07067_),
    .Y(_01477_),
    .A1(net5441),
    .A2(net4906));
 sg13g2_nand2_1 _17000_ (.Y(_07068_),
    .A(net3381),
    .B(net4907));
 sg13g2_o21ai_1 _17001_ (.B1(_07068_),
    .Y(_01478_),
    .A1(net5487),
    .A2(net4907));
 sg13g2_nand2_1 _17002_ (.Y(_07069_),
    .A(net2344),
    .B(net4906));
 sg13g2_o21ai_1 _17003_ (.B1(_07069_),
    .Y(_01479_),
    .A1(net5534),
    .A2(net4906));
 sg13g2_nand2_1 _17004_ (.Y(_07070_),
    .A(net2135),
    .B(_07066_));
 sg13g2_o21ai_1 _17005_ (.B1(_07070_),
    .Y(_01480_),
    .A1(net5577),
    .A2(net4907));
 sg13g2_nand2_1 _17006_ (.Y(_07071_),
    .A(net3063),
    .B(net4906));
 sg13g2_o21ai_1 _17007_ (.B1(_07071_),
    .Y(_01481_),
    .A1(net5621),
    .A2(net4906));
 sg13g2_nand2_1 _17008_ (.Y(_07072_),
    .A(net3188),
    .B(net4907));
 sg13g2_o21ai_1 _17009_ (.B1(_07072_),
    .Y(_01482_),
    .A1(net5669),
    .A2(net4907));
 sg13g2_nand2_1 _17010_ (.Y(_07073_),
    .A(net3021),
    .B(net4907));
 sg13g2_o21ai_1 _17011_ (.B1(_07073_),
    .Y(_01483_),
    .A1(net5713),
    .A2(net4907));
 sg13g2_nand2_1 _17012_ (.Y(_07074_),
    .A(net2285),
    .B(net4906));
 sg13g2_o21ai_1 _17013_ (.B1(_07074_),
    .Y(_01484_),
    .A1(net5758),
    .A2(net4906));
 sg13g2_nand2_1 _17014_ (.Y(_07075_),
    .A(net5251),
    .B(net5195));
 sg13g2_nand2_1 _17015_ (.Y(_07076_),
    .A(net2938),
    .B(net4905));
 sg13g2_o21ai_1 _17016_ (.B1(_07076_),
    .Y(_01485_),
    .A1(net5442),
    .A2(net4905));
 sg13g2_nand2_1 _17017_ (.Y(_07077_),
    .A(net2694),
    .B(net4905));
 sg13g2_o21ai_1 _17018_ (.B1(_07077_),
    .Y(_01486_),
    .A1(net5487),
    .A2(net4905));
 sg13g2_nand2_1 _17019_ (.Y(_07078_),
    .A(net2410),
    .B(net4905));
 sg13g2_o21ai_1 _17020_ (.B1(_07078_),
    .Y(_01487_),
    .A1(net5534),
    .A2(net4905));
 sg13g2_nand2_1 _17021_ (.Y(_07079_),
    .A(net3438),
    .B(net4905));
 sg13g2_o21ai_1 _17022_ (.B1(_07079_),
    .Y(_01488_),
    .A1(net5577),
    .A2(_07075_));
 sg13g2_nand2_1 _17023_ (.Y(_07080_),
    .A(net2680),
    .B(net4904));
 sg13g2_o21ai_1 _17024_ (.B1(_07080_),
    .Y(_01489_),
    .A1(net5621),
    .A2(net4904));
 sg13g2_nand2_1 _17025_ (.Y(_07081_),
    .A(net3108),
    .B(net4904));
 sg13g2_o21ai_1 _17026_ (.B1(_07081_),
    .Y(_01490_),
    .A1(net5669),
    .A2(net4904));
 sg13g2_nand2_1 _17027_ (.Y(_07082_),
    .A(net3468),
    .B(net4904));
 sg13g2_o21ai_1 _17028_ (.B1(_07082_),
    .Y(_01491_),
    .A1(net5713),
    .A2(net4904));
 sg13g2_nand2_1 _17029_ (.Y(_07083_),
    .A(net3271),
    .B(net4904));
 sg13g2_o21ai_1 _17030_ (.B1(_07083_),
    .Y(_01492_),
    .A1(net5758),
    .A2(net4904));
 sg13g2_nand2_1 _17031_ (.Y(_07084_),
    .A(net5246),
    .B(net5194));
 sg13g2_nand2_1 _17032_ (.Y(_07085_),
    .A(net2363),
    .B(net4902));
 sg13g2_o21ai_1 _17033_ (.B1(_07085_),
    .Y(_01493_),
    .A1(net5442),
    .A2(net4902));
 sg13g2_nand2_1 _17034_ (.Y(_07086_),
    .A(net2624),
    .B(net4903));
 sg13g2_o21ai_1 _17035_ (.B1(_07086_),
    .Y(_01494_),
    .A1(net5487),
    .A2(net4903));
 sg13g2_nand2_1 _17036_ (.Y(_07087_),
    .A(net2936),
    .B(net4902));
 sg13g2_o21ai_1 _17037_ (.B1(_07087_),
    .Y(_01495_),
    .A1(net5534),
    .A2(net4902));
 sg13g2_nand2_1 _17038_ (.Y(_07088_),
    .A(net3298),
    .B(net4902));
 sg13g2_o21ai_1 _17039_ (.B1(_07088_),
    .Y(_01496_),
    .A1(net5577),
    .A2(net4902));
 sg13g2_nand2_1 _17040_ (.Y(_07089_),
    .A(net2752),
    .B(net4902));
 sg13g2_o21ai_1 _17041_ (.B1(_07089_),
    .Y(_01497_),
    .A1(net5621),
    .A2(net4903));
 sg13g2_nand2_1 _17042_ (.Y(_07090_),
    .A(net2827),
    .B(net4903));
 sg13g2_o21ai_1 _17043_ (.B1(_07090_),
    .Y(_01498_),
    .A1(net5665),
    .A2(net4903));
 sg13g2_nand2_1 _17044_ (.Y(_07091_),
    .A(net3176),
    .B(net4903));
 sg13g2_o21ai_1 _17045_ (.B1(_07091_),
    .Y(_01499_),
    .A1(net5712),
    .A2(net4903));
 sg13g2_nand2_1 _17046_ (.Y(_07092_),
    .A(net2809),
    .B(net4902));
 sg13g2_o21ai_1 _17047_ (.B1(_07092_),
    .Y(_01500_),
    .A1(net5758),
    .A2(_07084_));
 sg13g2_nor3_1 _17048_ (.A(net5227),
    .B(net5240),
    .C(net5258),
    .Y(_07093_));
 sg13g2_nor2_1 _17049_ (.A(net3495),
    .B(net5175),
    .Y(_07094_));
 sg13g2_a21oi_1 _17050_ (.A1(net5441),
    .A2(net5175),
    .Y(_01501_),
    .B1(_07094_));
 sg13g2_nor2_1 _17051_ (.A(net3691),
    .B(net5174),
    .Y(_07095_));
 sg13g2_a21oi_1 _17052_ (.A1(net5487),
    .A2(net5174),
    .Y(_01502_),
    .B1(_07095_));
 sg13g2_nor2_1 _17053_ (.A(net4153),
    .B(net5174),
    .Y(_07096_));
 sg13g2_a21oi_1 _17054_ (.A1(net5534),
    .A2(net5174),
    .Y(_01503_),
    .B1(_07096_));
 sg13g2_nor2_1 _17055_ (.A(net4149),
    .B(net5175),
    .Y(_07097_));
 sg13g2_a21oi_1 _17056_ (.A1(net5577),
    .A2(net5175),
    .Y(_01504_),
    .B1(_07097_));
 sg13g2_nor2_1 _17057_ (.A(net4091),
    .B(net5175),
    .Y(_07098_));
 sg13g2_a21oi_1 _17058_ (.A1(net5620),
    .A2(net5175),
    .Y(_01505_),
    .B1(_07098_));
 sg13g2_nor2_1 _17059_ (.A(net4168),
    .B(net5174),
    .Y(_07099_));
 sg13g2_a21oi_1 _17060_ (.A1(net5665),
    .A2(net5174),
    .Y(_01506_),
    .B1(_07099_));
 sg13g2_nor2_1 _17061_ (.A(net3849),
    .B(net5174),
    .Y(_07100_));
 sg13g2_a21oi_1 _17062_ (.A1(net5712),
    .A2(net5174),
    .Y(_01507_),
    .B1(_07100_));
 sg13g2_nor2_1 _17063_ (.A(net3857),
    .B(net5175),
    .Y(_07101_));
 sg13g2_a21oi_1 _17064_ (.A1(net5758),
    .A2(net5175),
    .Y(_01508_),
    .B1(_07101_));
 sg13g2_nand2_1 _17065_ (.Y(_02126_),
    .A(net5249),
    .B(net5196));
 sg13g2_nand2_1 _17066_ (.Y(_02127_),
    .A(net2731),
    .B(net4900));
 sg13g2_o21ai_1 _17067_ (.B1(_02127_),
    .Y(_01509_),
    .A1(net5454),
    .A2(net4900));
 sg13g2_nand2_1 _17068_ (.Y(_02128_),
    .A(net3006),
    .B(net4900));
 sg13g2_o21ai_1 _17069_ (.B1(_02128_),
    .Y(_01510_),
    .A1(net5500),
    .A2(_02126_));
 sg13g2_nand2_1 _17070_ (.Y(_02129_),
    .A(net2629),
    .B(net4901));
 sg13g2_o21ai_1 _17071_ (.B1(_02129_),
    .Y(_01511_),
    .A1(net5547),
    .A2(net4901));
 sg13g2_nand2_1 _17072_ (.Y(_02130_),
    .A(net2980),
    .B(net4901));
 sg13g2_o21ai_1 _17073_ (.B1(_02130_),
    .Y(_01512_),
    .A1(net5588),
    .A2(net4900));
 sg13g2_nand2_1 _17074_ (.Y(_02131_),
    .A(net2744),
    .B(net4901));
 sg13g2_o21ai_1 _17075_ (.B1(_02131_),
    .Y(_01513_),
    .A1(net5633),
    .A2(net4901));
 sg13g2_nand2_1 _17076_ (.Y(_02132_),
    .A(net2687),
    .B(net4901));
 sg13g2_o21ai_1 _17077_ (.B1(_02132_),
    .Y(_01514_),
    .A1(net5679),
    .A2(net4901));
 sg13g2_nand2_1 _17078_ (.Y(_02133_),
    .A(net2527),
    .B(net4900));
 sg13g2_o21ai_1 _17079_ (.B1(_02133_),
    .Y(_01515_),
    .A1(net5723),
    .A2(net4900));
 sg13g2_nand2_1 _17080_ (.Y(_02134_),
    .A(net2610),
    .B(net4900));
 sg13g2_o21ai_1 _17081_ (.B1(_02134_),
    .Y(_01516_),
    .A1(net5771),
    .A2(net4900));
 sg13g2_nand2_1 _17082_ (.Y(_02135_),
    .A(_03139_),
    .B(net5196));
 sg13g2_nand2_1 _17083_ (.Y(_02136_),
    .A(net2688),
    .B(net4898));
 sg13g2_o21ai_1 _17084_ (.B1(_02136_),
    .Y(_01517_),
    .A1(net5454),
    .A2(net4898));
 sg13g2_nand2_1 _17085_ (.Y(_02137_),
    .A(net2205),
    .B(net4898));
 sg13g2_o21ai_1 _17086_ (.B1(_02137_),
    .Y(_01518_),
    .A1(net5500),
    .A2(net4898));
 sg13g2_nand2_1 _17087_ (.Y(_02138_),
    .A(net2643),
    .B(_02135_));
 sg13g2_o21ai_1 _17088_ (.B1(_02138_),
    .Y(_01519_),
    .A1(net5547),
    .A2(net4899));
 sg13g2_nand2_1 _17089_ (.Y(_02139_),
    .A(net2484),
    .B(net4899));
 sg13g2_o21ai_1 _17090_ (.B1(_02139_),
    .Y(_01520_),
    .A1(net5588),
    .A2(net4899));
 sg13g2_nand2_1 _17091_ (.Y(_02140_),
    .A(net3067),
    .B(net4899));
 sg13g2_o21ai_1 _17092_ (.B1(_02140_),
    .Y(_01521_),
    .A1(net5633),
    .A2(net4899));
 sg13g2_nand2_1 _17093_ (.Y(_02141_),
    .A(net2615),
    .B(net4899));
 sg13g2_o21ai_1 _17094_ (.B1(_02141_),
    .Y(_01522_),
    .A1(net5678),
    .A2(net4899));
 sg13g2_nand2_1 _17095_ (.Y(_02142_),
    .A(net2821),
    .B(net4898));
 sg13g2_o21ai_1 _17096_ (.B1(_02142_),
    .Y(_01523_),
    .A1(net5723),
    .A2(net4898));
 sg13g2_nand2_1 _17097_ (.Y(_02143_),
    .A(net2875),
    .B(net4898));
 sg13g2_o21ai_1 _17098_ (.B1(_02143_),
    .Y(_01524_),
    .A1(net5771),
    .A2(net4898));
 sg13g2_nand2_1 _17099_ (.Y(_02144_),
    .A(_03079_),
    .B(net5196));
 sg13g2_nand2_1 _17100_ (.Y(_02145_),
    .A(net2683),
    .B(net4897));
 sg13g2_o21ai_1 _17101_ (.B1(_02145_),
    .Y(_01525_),
    .A1(net5454),
    .A2(net4897));
 sg13g2_nand2_1 _17102_ (.Y(_02146_),
    .A(net2381),
    .B(net4896));
 sg13g2_o21ai_1 _17103_ (.B1(_02146_),
    .Y(_01526_),
    .A1(net5500),
    .A2(net4896));
 sg13g2_nand2_1 _17104_ (.Y(_02147_),
    .A(net2386),
    .B(net4897));
 sg13g2_o21ai_1 _17105_ (.B1(_02147_),
    .Y(_01527_),
    .A1(net5544),
    .A2(net4897));
 sg13g2_nand2_1 _17106_ (.Y(_02148_),
    .A(net2581),
    .B(net4896));
 sg13g2_o21ai_1 _17107_ (.B1(_02148_),
    .Y(_01528_),
    .A1(net5590),
    .A2(net4896));
 sg13g2_nand2_1 _17108_ (.Y(_02149_),
    .A(net2776),
    .B(net4897));
 sg13g2_o21ai_1 _17109_ (.B1(_02149_),
    .Y(_01529_),
    .A1(net5633),
    .A2(net4897));
 sg13g2_nand2_1 _17110_ (.Y(_02150_),
    .A(net2934),
    .B(net4897));
 sg13g2_o21ai_1 _17111_ (.B1(_02150_),
    .Y(_01530_),
    .A1(net5679),
    .A2(net4897));
 sg13g2_nand2_1 _17112_ (.Y(_02151_),
    .A(net2670),
    .B(net4896));
 sg13g2_o21ai_1 _17113_ (.B1(_02151_),
    .Y(_01531_),
    .A1(net5723),
    .A2(net4896));
 sg13g2_nand2_1 _17114_ (.Y(_02152_),
    .A(net3043),
    .B(net4896));
 sg13g2_o21ai_1 _17115_ (.B1(_02152_),
    .Y(_01532_),
    .A1(net5771),
    .A2(net4896));
 sg13g2_nor2_1 _17116_ (.A(net5252),
    .B(net5210),
    .Y(_02153_));
 sg13g2_nor2_1 _17117_ (.A(net3657),
    .B(net4894),
    .Y(_02154_));
 sg13g2_a21oi_1 _17118_ (.A1(net5452),
    .A2(net4894),
    .Y(_01533_),
    .B1(_02154_));
 sg13g2_nor2_1 _17119_ (.A(net4075),
    .B(net4894),
    .Y(_02155_));
 sg13g2_a21oi_1 _17120_ (.A1(net5498),
    .A2(net4894),
    .Y(_01534_),
    .B1(_02155_));
 sg13g2_nor2_1 _17121_ (.A(net3574),
    .B(net4894),
    .Y(_02156_));
 sg13g2_a21oi_1 _17122_ (.A1(net5541),
    .A2(net4894),
    .Y(_01535_),
    .B1(_02156_));
 sg13g2_nor2_1 _17123_ (.A(net3391),
    .B(net4895),
    .Y(_02157_));
 sg13g2_a21oi_1 _17124_ (.A1(net5598),
    .A2(net4895),
    .Y(_01536_),
    .B1(_02157_));
 sg13g2_nor2_1 _17125_ (.A(net3643),
    .B(net4895),
    .Y(_02158_));
 sg13g2_a21oi_1 _17126_ (.A1(net5641),
    .A2(net4895),
    .Y(_01537_),
    .B1(_02158_));
 sg13g2_nor2_1 _17127_ (.A(net3701),
    .B(net4895),
    .Y(_02159_));
 sg13g2_a21oi_1 _17128_ (.A1(net5692),
    .A2(net4895),
    .Y(_01538_),
    .B1(_02159_));
 sg13g2_nor2_1 _17129_ (.A(net3353),
    .B(net4895),
    .Y(_02160_));
 sg13g2_a21oi_1 _17130_ (.A1(net5732),
    .A2(net4895),
    .Y(_01539_),
    .B1(_02160_));
 sg13g2_nor2_1 _17131_ (.A(net3585),
    .B(net4894),
    .Y(_02161_));
 sg13g2_a21oi_1 _17132_ (.A1(net5767),
    .A2(net4894),
    .Y(_01540_),
    .B1(_02161_));
 sg13g2_nand2_1 _17133_ (.Y(_02162_),
    .A(net5235),
    .B(net5197));
 sg13g2_nand2_1 _17134_ (.Y(_02163_),
    .A(net2575),
    .B(net4893));
 sg13g2_o21ai_1 _17135_ (.B1(_02163_),
    .Y(_01541_),
    .A1(net5455),
    .A2(net4893));
 sg13g2_nand2_1 _17136_ (.Y(_02164_),
    .A(net3242),
    .B(net4892));
 sg13g2_o21ai_1 _17137_ (.B1(_02164_),
    .Y(_01542_),
    .A1(net5500),
    .A2(net4892));
 sg13g2_nand2_1 _17138_ (.Y(_02165_),
    .A(net3225),
    .B(net4893));
 sg13g2_o21ai_1 _17139_ (.B1(_02165_),
    .Y(_01543_),
    .A1(net5545),
    .A2(net4893));
 sg13g2_nand2_1 _17140_ (.Y(_02166_),
    .A(net2134),
    .B(net4893));
 sg13g2_o21ai_1 _17141_ (.B1(_02166_),
    .Y(_01544_),
    .A1(net5588),
    .A2(net4893));
 sg13g2_nand2_1 _17142_ (.Y(_02167_),
    .A(net2385),
    .B(net4892));
 sg13g2_o21ai_1 _17143_ (.B1(_02167_),
    .Y(_01545_),
    .A1(net5634),
    .A2(net4892));
 sg13g2_nand2_1 _17144_ (.Y(_02168_),
    .A(net2595),
    .B(net4892));
 sg13g2_o21ai_1 _17145_ (.B1(_02168_),
    .Y(_01546_),
    .A1(net5680),
    .A2(net4892));
 sg13g2_nand2_1 _17146_ (.Y(_02169_),
    .A(net2472),
    .B(net4892));
 sg13g2_o21ai_1 _17147_ (.B1(_02169_),
    .Y(_01547_),
    .A1(net5725),
    .A2(net4892));
 sg13g2_nand2_1 _17148_ (.Y(_02170_),
    .A(net2151),
    .B(net4893));
 sg13g2_o21ai_1 _17149_ (.B1(_02170_),
    .Y(_01548_),
    .A1(net5770),
    .A2(net4893));
 sg13g2_nand2_1 _17150_ (.Y(_02171_),
    .A(net5234),
    .B(net5196));
 sg13g2_nand2_1 _17151_ (.Y(_02172_),
    .A(net2703),
    .B(net4891));
 sg13g2_o21ai_1 _17152_ (.B1(_02172_),
    .Y(_01549_),
    .A1(net5455),
    .A2(net4891));
 sg13g2_nand2_1 _17153_ (.Y(_02173_),
    .A(net2542),
    .B(net4890));
 sg13g2_o21ai_1 _17154_ (.B1(_02173_),
    .Y(_01550_),
    .A1(net5501),
    .A2(net4890));
 sg13g2_nand2_1 _17155_ (.Y(_02174_),
    .A(net2721),
    .B(net4891));
 sg13g2_o21ai_1 _17156_ (.B1(_02174_),
    .Y(_01551_),
    .A1(net5544),
    .A2(net4891));
 sg13g2_nand2_1 _17157_ (.Y(_02175_),
    .A(net2749),
    .B(net4891));
 sg13g2_o21ai_1 _17158_ (.B1(_02175_),
    .Y(_01552_),
    .A1(net5588),
    .A2(net4891));
 sg13g2_nand2_1 _17159_ (.Y(_02176_),
    .A(net3285),
    .B(net4890));
 sg13g2_o21ai_1 _17160_ (.B1(_02176_),
    .Y(_01553_),
    .A1(net5634),
    .A2(net4890));
 sg13g2_nand2_1 _17161_ (.Y(_02177_),
    .A(net3032),
    .B(net4890));
 sg13g2_o21ai_1 _17162_ (.B1(_02177_),
    .Y(_01554_),
    .A1(net5680),
    .A2(net4890));
 sg13g2_nand2_1 _17163_ (.Y(_02178_),
    .A(net3320),
    .B(net4890));
 sg13g2_o21ai_1 _17164_ (.B1(_02178_),
    .Y(_01555_),
    .A1(net5725),
    .A2(net4890));
 sg13g2_nand2_1 _17165_ (.Y(_02179_),
    .A(net2846),
    .B(net4891));
 sg13g2_o21ai_1 _17166_ (.B1(_02179_),
    .Y(_01556_),
    .A1(net5771),
    .A2(net4891));
 sg13g2_nand2_1 _17167_ (.Y(_02180_),
    .A(_03066_),
    .B(net5196));
 sg13g2_nand2_1 _17168_ (.Y(_02181_),
    .A(net2427),
    .B(net4889));
 sg13g2_o21ai_1 _17169_ (.B1(_02181_),
    .Y(_01557_),
    .A1(net5455),
    .A2(net4889));
 sg13g2_nand2_1 _17170_ (.Y(_02182_),
    .A(net2644),
    .B(net4888));
 sg13g2_o21ai_1 _17171_ (.B1(_02182_),
    .Y(_01558_),
    .A1(net5502),
    .A2(net4888));
 sg13g2_nand2_1 _17172_ (.Y(_02183_),
    .A(net2592),
    .B(net4889));
 sg13g2_o21ai_1 _17173_ (.B1(_02183_),
    .Y(_01559_),
    .A1(net5545),
    .A2(net4889));
 sg13g2_nand2_1 _17174_ (.Y(_02184_),
    .A(net2232),
    .B(net4889));
 sg13g2_o21ai_1 _17175_ (.B1(_02184_),
    .Y(_01560_),
    .A1(net5590),
    .A2(net4889));
 sg13g2_nand2_1 _17176_ (.Y(_02185_),
    .A(net2866),
    .B(net4888));
 sg13g2_o21ai_1 _17177_ (.B1(_02185_),
    .Y(_01561_),
    .A1(net5635),
    .A2(net4888));
 sg13g2_nand2_1 _17178_ (.Y(_02186_),
    .A(net2503),
    .B(net4888));
 sg13g2_o21ai_1 _17179_ (.B1(_02186_),
    .Y(_01562_),
    .A1(net5680),
    .A2(net4888));
 sg13g2_nand2_1 _17180_ (.Y(_02187_),
    .A(net2705),
    .B(net4888));
 sg13g2_o21ai_1 _17181_ (.B1(_02187_),
    .Y(_01563_),
    .A1(net5725),
    .A2(net4888));
 sg13g2_nand2_1 _17182_ (.Y(_02188_),
    .A(net3253),
    .B(net4889));
 sg13g2_o21ai_1 _17183_ (.B1(_02188_),
    .Y(_01564_),
    .A1(net5772),
    .A2(net4889));
 sg13g2_nand2_1 _17184_ (.Y(_02189_),
    .A(net5238),
    .B(net5196));
 sg13g2_nand2_1 _17185_ (.Y(_02190_),
    .A(net2554),
    .B(net4887));
 sg13g2_o21ai_1 _17186_ (.B1(_02190_),
    .Y(_01565_),
    .A1(net5455),
    .A2(_02189_));
 sg13g2_nand2_1 _17187_ (.Y(_02191_),
    .A(net3214),
    .B(net4886));
 sg13g2_o21ai_1 _17188_ (.B1(_02191_),
    .Y(_01566_),
    .A1(net5502),
    .A2(net4886));
 sg13g2_nand2_1 _17189_ (.Y(_02192_),
    .A(net3121),
    .B(net4887));
 sg13g2_o21ai_1 _17190_ (.B1(_02192_),
    .Y(_01567_),
    .A1(net5545),
    .A2(net4887));
 sg13g2_nand2_1 _17191_ (.Y(_02193_),
    .A(net3272),
    .B(net4887));
 sg13g2_o21ai_1 _17192_ (.B1(_02193_),
    .Y(_01568_),
    .A1(net5589),
    .A2(net4887));
 sg13g2_nand2_1 _17193_ (.Y(_02194_),
    .A(net2228),
    .B(net4887));
 sg13g2_o21ai_1 _17194_ (.B1(_02194_),
    .Y(_01569_),
    .A1(net5634),
    .A2(net4887));
 sg13g2_nand2_1 _17195_ (.Y(_02195_),
    .A(net2817),
    .B(net4886));
 sg13g2_o21ai_1 _17196_ (.B1(_02195_),
    .Y(_01570_),
    .A1(net5680),
    .A2(net4886));
 sg13g2_nand2_1 _17197_ (.Y(_02196_),
    .A(net2586),
    .B(net4886));
 sg13g2_o21ai_1 _17198_ (.B1(_02196_),
    .Y(_01571_),
    .A1(net5725),
    .A2(net4886));
 sg13g2_nand2_1 _17199_ (.Y(_02197_),
    .A(net2665),
    .B(net4886));
 sg13g2_o21ai_1 _17200_ (.B1(_02197_),
    .Y(_01572_),
    .A1(net5772),
    .A2(net4886));
 sg13g2_nand2_1 _17201_ (.Y(_02198_),
    .A(net5244),
    .B(net5197));
 sg13g2_nand2_1 _17202_ (.Y(_02199_),
    .A(net2715),
    .B(_02198_));
 sg13g2_o21ai_1 _17203_ (.B1(_02199_),
    .Y(_01573_),
    .A1(net5454),
    .A2(net4885));
 sg13g2_nand2_1 _17204_ (.Y(_02200_),
    .A(net2395),
    .B(net4884));
 sg13g2_o21ai_1 _17205_ (.B1(_02200_),
    .Y(_01574_),
    .A1(net5500),
    .A2(net4884));
 sg13g2_nand2_1 _17206_ (.Y(_02201_),
    .A(net2724),
    .B(net4885));
 sg13g2_o21ai_1 _17207_ (.B1(_02201_),
    .Y(_01575_),
    .A1(net5544),
    .A2(net4885));
 sg13g2_nand2_1 _17208_ (.Y(_02202_),
    .A(net2181),
    .B(net4885));
 sg13g2_o21ai_1 _17209_ (.B1(_02202_),
    .Y(_01576_),
    .A1(net5588),
    .A2(net4884));
 sg13g2_nand2_1 _17210_ (.Y(_02203_),
    .A(net2172),
    .B(net4885));
 sg13g2_o21ai_1 _17211_ (.B1(_02203_),
    .Y(_01577_),
    .A1(net5633),
    .A2(net4885));
 sg13g2_nand2_1 _17212_ (.Y(_02204_),
    .A(net3080),
    .B(net4885));
 sg13g2_o21ai_1 _17213_ (.B1(_02204_),
    .Y(_01578_),
    .A1(net5679),
    .A2(net4884));
 sg13g2_nand2_1 _17214_ (.Y(_02205_),
    .A(net2728),
    .B(net4884));
 sg13g2_o21ai_1 _17215_ (.B1(_02205_),
    .Y(_01579_),
    .A1(net5724),
    .A2(net4884));
 sg13g2_nand2_1 _17216_ (.Y(_02206_),
    .A(net2448),
    .B(net4884));
 sg13g2_o21ai_1 _17217_ (.B1(_02206_),
    .Y(_01580_),
    .A1(net5770),
    .A2(net4884));
 sg13g2_nand2_1 _17218_ (.Y(_02207_),
    .A(_03016_),
    .B(net5196));
 sg13g2_nand2_1 _17219_ (.Y(_02208_),
    .A(net2640),
    .B(net4883));
 sg13g2_o21ai_1 _17220_ (.B1(_02208_),
    .Y(_01581_),
    .A1(net5454),
    .A2(net4883));
 sg13g2_nand2_1 _17221_ (.Y(_02209_),
    .A(net2969),
    .B(net4882));
 sg13g2_o21ai_1 _17222_ (.B1(_02209_),
    .Y(_01582_),
    .A1(net5500),
    .A2(net4882));
 sg13g2_nand2_1 _17223_ (.Y(_02210_),
    .A(net2486),
    .B(net4883));
 sg13g2_o21ai_1 _17224_ (.B1(_02210_),
    .Y(_01583_),
    .A1(net5544),
    .A2(net4883));
 sg13g2_nand2_1 _17225_ (.Y(_02211_),
    .A(net2916),
    .B(net4882));
 sg13g2_o21ai_1 _17226_ (.B1(_02211_),
    .Y(_01584_),
    .A1(net5588),
    .A2(net4882));
 sg13g2_nand2_1 _17227_ (.Y(_02212_),
    .A(net2518),
    .B(net4883));
 sg13g2_o21ai_1 _17228_ (.B1(_02212_),
    .Y(_01585_),
    .A1(net5633),
    .A2(net4883));
 sg13g2_nand2_1 _17229_ (.Y(_02213_),
    .A(net3360),
    .B(net4883));
 sg13g2_o21ai_1 _17230_ (.B1(_02213_),
    .Y(_01586_),
    .A1(net5679),
    .A2(net4883));
 sg13g2_nand2_1 _17231_ (.Y(_02214_),
    .A(net2998),
    .B(net4882));
 sg13g2_o21ai_1 _17232_ (.B1(_02214_),
    .Y(_01587_),
    .A1(net5724),
    .A2(net4882));
 sg13g2_nand2_1 _17233_ (.Y(_02215_),
    .A(net3129),
    .B(net4882));
 sg13g2_o21ai_1 _17234_ (.B1(_02215_),
    .Y(_01588_),
    .A1(net5770),
    .A2(net4882));
 sg13g2_nand2_2 _17235_ (.Y(_02216_),
    .A(_02980_),
    .B(net5197));
 sg13g2_nand2_1 _17236_ (.Y(_02217_),
    .A(net2184),
    .B(net4881));
 sg13g2_o21ai_1 _17237_ (.B1(_02217_),
    .Y(_01589_),
    .A1(net5454),
    .A2(net4881));
 sg13g2_nand2_1 _17238_ (.Y(_02218_),
    .A(net2407),
    .B(net4880));
 sg13g2_o21ai_1 _17239_ (.B1(_02218_),
    .Y(_01590_),
    .A1(net5500),
    .A2(net4880));
 sg13g2_nand2_1 _17240_ (.Y(_02219_),
    .A(net2699),
    .B(net4881));
 sg13g2_o21ai_1 _17241_ (.B1(_02219_),
    .Y(_01591_),
    .A1(net5544),
    .A2(net4881));
 sg13g2_nand2_1 _17242_ (.Y(_02220_),
    .A(net2201),
    .B(net4880));
 sg13g2_o21ai_1 _17243_ (.B1(_02220_),
    .Y(_01592_),
    .A1(net5588),
    .A2(net4880));
 sg13g2_nand2_1 _17244_ (.Y(_02221_),
    .A(net2188),
    .B(net4881));
 sg13g2_o21ai_1 _17245_ (.B1(_02221_),
    .Y(_01593_),
    .A1(net5635),
    .A2(net4881));
 sg13g2_nand2_1 _17246_ (.Y(_02222_),
    .A(net2639),
    .B(net4881));
 sg13g2_o21ai_1 _17247_ (.B1(_02222_),
    .Y(_01594_),
    .A1(net5679),
    .A2(net4881));
 sg13g2_nand2_1 _17248_ (.Y(_02223_),
    .A(net2734),
    .B(net4880));
 sg13g2_o21ai_1 _17249_ (.B1(_02223_),
    .Y(_01595_),
    .A1(net5724),
    .A2(net4880));
 sg13g2_nand2_1 _17250_ (.Y(_02224_),
    .A(net2782),
    .B(net4880));
 sg13g2_o21ai_1 _17251_ (.B1(_02224_),
    .Y(_01596_),
    .A1(net5770),
    .A2(net4880));
 sg13g2_nand2_1 _17252_ (.Y(_02225_),
    .A(net5243),
    .B(net5197));
 sg13g2_nand2_1 _17253_ (.Y(_02226_),
    .A(net3040),
    .B(net4879));
 sg13g2_o21ai_1 _17254_ (.B1(_02226_),
    .Y(_01597_),
    .A1(net5454),
    .A2(net4879));
 sg13g2_nand2_1 _17255_ (.Y(_02227_),
    .A(net2792),
    .B(net4878));
 sg13g2_o21ai_1 _17256_ (.B1(_02227_),
    .Y(_01598_),
    .A1(net5500),
    .A2(net4878));
 sg13g2_nand2_1 _17257_ (.Y(_02228_),
    .A(net2585),
    .B(net4879));
 sg13g2_o21ai_1 _17258_ (.B1(_02228_),
    .Y(_01599_),
    .A1(net5544),
    .A2(net4879));
 sg13g2_nand2_1 _17259_ (.Y(_02229_),
    .A(net3302),
    .B(net4878));
 sg13g2_o21ai_1 _17260_ (.B1(_02229_),
    .Y(_01600_),
    .A1(net5588),
    .A2(net4878));
 sg13g2_nand2_1 _17261_ (.Y(_02230_),
    .A(net2364),
    .B(net4879));
 sg13g2_o21ai_1 _17262_ (.B1(_02230_),
    .Y(_01601_),
    .A1(net5635),
    .A2(net4879));
 sg13g2_nand2_1 _17263_ (.Y(_02231_),
    .A(net2669),
    .B(net4879));
 sg13g2_o21ai_1 _17264_ (.B1(_02231_),
    .Y(_01602_),
    .A1(net5679),
    .A2(net4879));
 sg13g2_nand2_1 _17265_ (.Y(_02232_),
    .A(net2418),
    .B(net4878));
 sg13g2_o21ai_1 _17266_ (.B1(_02232_),
    .Y(_01603_),
    .A1(net5724),
    .A2(net4878));
 sg13g2_nand2_1 _17267_ (.Y(_02233_),
    .A(net3297),
    .B(net4878));
 sg13g2_o21ai_1 _17268_ (.B1(_02233_),
    .Y(_01604_),
    .A1(net5770),
    .A2(net4878));
 sg13g2_nand2_1 _17269_ (.Y(_02234_),
    .A(net5245),
    .B(net5197));
 sg13g2_nand2_1 _17270_ (.Y(_02235_),
    .A(net3268),
    .B(net4877));
 sg13g2_o21ai_1 _17271_ (.B1(_02235_),
    .Y(_01605_),
    .A1(net5455),
    .A2(net4877));
 sg13g2_nand2_1 _17272_ (.Y(_02236_),
    .A(net2831),
    .B(net4877));
 sg13g2_o21ai_1 _17273_ (.B1(_02236_),
    .Y(_01606_),
    .A1(net5502),
    .A2(net4877));
 sg13g2_nand2_1 _17274_ (.Y(_02237_),
    .A(net2662),
    .B(net4876));
 sg13g2_o21ai_1 _17275_ (.B1(_02237_),
    .Y(_01607_),
    .A1(net5546),
    .A2(net4876));
 sg13g2_nand2_1 _17276_ (.Y(_02238_),
    .A(net2145),
    .B(net4877));
 sg13g2_o21ai_1 _17277_ (.B1(_02238_),
    .Y(_01608_),
    .A1(net5589),
    .A2(net4877));
 sg13g2_nand2_1 _17278_ (.Y(_02239_),
    .A(net2413),
    .B(net4877));
 sg13g2_o21ai_1 _17279_ (.B1(_02239_),
    .Y(_01609_),
    .A1(net5634),
    .A2(net4877));
 sg13g2_nand2_1 _17280_ (.Y(_02240_),
    .A(net2191),
    .B(net4876));
 sg13g2_o21ai_1 _17281_ (.B1(_02240_),
    .Y(_01610_),
    .A1(net5685),
    .A2(net4876));
 sg13g2_nand2_1 _17282_ (.Y(_02241_),
    .A(net2451),
    .B(net4876));
 sg13g2_o21ai_1 _17283_ (.B1(_02241_),
    .Y(_01611_),
    .A1(net5729),
    .A2(net4876));
 sg13g2_nand2_1 _17284_ (.Y(_02242_),
    .A(net2150),
    .B(net4876));
 sg13g2_o21ai_1 _17285_ (.B1(_02242_),
    .Y(_01612_),
    .A1(net5777),
    .A2(net4876));
 sg13g2_nor2_1 _17286_ (.A(net5254),
    .B(net5210),
    .Y(_02243_));
 sg13g2_nor2_1 _17287_ (.A(net3899),
    .B(net4874),
    .Y(_02244_));
 sg13g2_a21oi_1 _17288_ (.A1(net5452),
    .A2(net4874),
    .Y(_01613_),
    .B1(_02244_));
 sg13g2_nor2_1 _17289_ (.A(net4094),
    .B(net4874),
    .Y(_02245_));
 sg13g2_a21oi_1 _17290_ (.A1(net5497),
    .A2(net4874),
    .Y(_01614_),
    .B1(_02245_));
 sg13g2_nor2_1 _17291_ (.A(net3883),
    .B(net4874),
    .Y(_02246_));
 sg13g2_a21oi_1 _17292_ (.A1(net5541),
    .A2(net4874),
    .Y(_01615_),
    .B1(_02246_));
 sg13g2_nor2_1 _17293_ (.A(net3407),
    .B(net4875),
    .Y(_02247_));
 sg13g2_a21oi_1 _17294_ (.A1(net5598),
    .A2(net4875),
    .Y(_01616_),
    .B1(_02247_));
 sg13g2_nor2_1 _17295_ (.A(net3808),
    .B(net4875),
    .Y(_02248_));
 sg13g2_a21oi_1 _17296_ (.A1(net5641),
    .A2(net4875),
    .Y(_01617_),
    .B1(_02248_));
 sg13g2_nor2_1 _17297_ (.A(net3442),
    .B(net4875),
    .Y(_02249_));
 sg13g2_a21oi_1 _17298_ (.A1(net5687),
    .A2(net4875),
    .Y(_01618_),
    .B1(_02249_));
 sg13g2_nor2_1 _17299_ (.A(net3562),
    .B(net4875),
    .Y(_02250_));
 sg13g2_a21oi_1 _17300_ (.A1(net5732),
    .A2(net4875),
    .Y(_01619_),
    .B1(_02250_));
 sg13g2_nor2_1 _17301_ (.A(net3573),
    .B(net4874),
    .Y(_02251_));
 sg13g2_a21oi_1 _17302_ (.A1(net5767),
    .A2(net4874),
    .Y(_01620_),
    .B1(_02251_));
 sg13g2_nand2_1 _17303_ (.Y(_02252_),
    .A(net5247),
    .B(net5197));
 sg13g2_nand2_1 _17304_ (.Y(_02253_),
    .A(net3215),
    .B(net4872));
 sg13g2_o21ai_1 _17305_ (.B1(_02253_),
    .Y(_01621_),
    .A1(net5443),
    .A2(net4872));
 sg13g2_nand2_1 _17306_ (.Y(_02254_),
    .A(net2419),
    .B(net4873));
 sg13g2_o21ai_1 _17307_ (.B1(_02254_),
    .Y(_01622_),
    .A1(net5502),
    .A2(net4873));
 sg13g2_nand2_1 _17308_ (.Y(_02255_),
    .A(net2898),
    .B(net4872));
 sg13g2_o21ai_1 _17309_ (.B1(_02255_),
    .Y(_01623_),
    .A1(net5546),
    .A2(net4872));
 sg13g2_nand2_1 _17310_ (.Y(_02256_),
    .A(net2862),
    .B(net4872));
 sg13g2_o21ai_1 _17311_ (.B1(_02256_),
    .Y(_01624_),
    .A1(net5589),
    .A2(net4872));
 sg13g2_nand2_1 _17312_ (.Y(_02257_),
    .A(net2500),
    .B(net4873));
 sg13g2_o21ai_1 _17313_ (.B1(_02257_),
    .Y(_01625_),
    .A1(net5635),
    .A2(net4873));
 sg13g2_nand2_1 _17314_ (.Y(_02258_),
    .A(net2891),
    .B(net4873));
 sg13g2_o21ai_1 _17315_ (.B1(_02258_),
    .Y(_01626_),
    .A1(net5680),
    .A2(net4873));
 sg13g2_nand2_1 _17316_ (.Y(_02259_),
    .A(net2569),
    .B(net4873));
 sg13g2_o21ai_1 _17317_ (.B1(_02259_),
    .Y(_01627_),
    .A1(net5729),
    .A2(net4873));
 sg13g2_nand2_1 _17318_ (.Y(_02260_),
    .A(net3085),
    .B(net4872));
 sg13g2_o21ai_1 _17319_ (.B1(_02260_),
    .Y(_01628_),
    .A1(net5772),
    .A2(net4872));
 sg13g2_nor3_2 _17320_ (.A(net5241),
    .B(net5258),
    .C(_03180_),
    .Y(_02261_));
 sg13g2_nor2_1 _17321_ (.A(net3557),
    .B(net5172),
    .Y(_02262_));
 sg13g2_a21oi_1 _17322_ (.A1(net5443),
    .A2(net5172),
    .Y(_01629_),
    .B1(_02262_));
 sg13g2_nor2_1 _17323_ (.A(net3807),
    .B(net5173),
    .Y(_02263_));
 sg13g2_a21oi_1 _17324_ (.A1(net5502),
    .A2(net5173),
    .Y(_01630_),
    .B1(_02263_));
 sg13g2_nor2_1 _17325_ (.A(net3692),
    .B(net5172),
    .Y(_02264_));
 sg13g2_a21oi_1 _17326_ (.A1(net5546),
    .A2(net5172),
    .Y(_01631_),
    .B1(_02264_));
 sg13g2_nor2_1 _17327_ (.A(net3864),
    .B(net5172),
    .Y(_02265_));
 sg13g2_a21oi_1 _17328_ (.A1(net5589),
    .A2(net5172),
    .Y(_01632_),
    .B1(_02265_));
 sg13g2_nor2_1 _17329_ (.A(net3751),
    .B(net5173),
    .Y(_02266_));
 sg13g2_a21oi_1 _17330_ (.A1(net5635),
    .A2(net5173),
    .Y(_01633_),
    .B1(_02266_));
 sg13g2_nor2_1 _17331_ (.A(net3313),
    .B(net5173),
    .Y(_02267_));
 sg13g2_a21oi_1 _17332_ (.A1(net5680),
    .A2(net5173),
    .Y(_01634_),
    .B1(_02267_));
 sg13g2_nor2_1 _17333_ (.A(net3305),
    .B(net5173),
    .Y(_02268_));
 sg13g2_a21oi_1 _17334_ (.A1(net5725),
    .A2(net5173),
    .Y(_01635_),
    .B1(_02268_));
 sg13g2_nor2_1 _17335_ (.A(net3293),
    .B(net5172),
    .Y(_02269_));
 sg13g2_a21oi_1 _17336_ (.A1(net5772),
    .A2(net5172),
    .Y(_01636_),
    .B1(_02269_));
 sg13g2_nand4_1 _17337_ (.B(net5802),
    .C(net5220),
    .A(net5801),
    .Y(_02270_),
    .D(net5249));
 sg13g2_nand2_1 _17338_ (.Y(_02271_),
    .A(net2214),
    .B(net4871));
 sg13g2_o21ai_1 _17339_ (.B1(_02271_),
    .Y(_01637_),
    .A1(net5443),
    .A2(_02270_));
 sg13g2_nand2_1 _17340_ (.Y(_02272_),
    .A(net2774),
    .B(net4870));
 sg13g2_o21ai_1 _17341_ (.B1(_02272_),
    .Y(_01638_),
    .A1(net5491),
    .A2(net4870));
 sg13g2_nand2_1 _17342_ (.Y(_02273_),
    .A(net2267),
    .B(net4871));
 sg13g2_o21ai_1 _17343_ (.B1(_02273_),
    .Y(_01639_),
    .A1(net5536),
    .A2(net4871));
 sg13g2_nand2_1 _17344_ (.Y(_02274_),
    .A(net3090),
    .B(net4870));
 sg13g2_o21ai_1 _17345_ (.B1(_02274_),
    .Y(_01640_),
    .A1(net5578),
    .A2(net4870));
 sg13g2_nand2_1 _17346_ (.Y(_02275_),
    .A(net2154),
    .B(net4871));
 sg13g2_o21ai_1 _17347_ (.B1(_02275_),
    .Y(_01641_),
    .A1(net5627),
    .A2(net4871));
 sg13g2_nand2_1 _17348_ (.Y(_02276_),
    .A(net2197),
    .B(net4871));
 sg13g2_o21ai_1 _17349_ (.B1(_02276_),
    .Y(_01642_),
    .A1(net5668),
    .A2(net4870));
 sg13g2_nand2_1 _17350_ (.Y(_02277_),
    .A(net2340),
    .B(net4871));
 sg13g2_o21ai_1 _17351_ (.B1(_02277_),
    .Y(_01643_),
    .A1(net5714),
    .A2(net4870));
 sg13g2_nand2_1 _17352_ (.Y(_02278_),
    .A(net3170),
    .B(net4870));
 sg13g2_o21ai_1 _17353_ (.B1(_02278_),
    .Y(_01644_),
    .A1(net5760),
    .A2(net4870));
 sg13g2_nor2_1 _17354_ (.A(net5252),
    .B(net5046),
    .Y(_02279_));
 sg13g2_nor2_1 _17355_ (.A(net4105),
    .B(net4706),
    .Y(_02280_));
 sg13g2_a21oi_1 _17356_ (.A1(net5443),
    .A2(_02279_),
    .Y(_01645_),
    .B1(_02280_));
 sg13g2_nor2_1 _17357_ (.A(net3663),
    .B(net4705),
    .Y(_02281_));
 sg13g2_a21oi_1 _17358_ (.A1(net5491),
    .A2(net4705),
    .Y(_01646_),
    .B1(_02281_));
 sg13g2_nor2_1 _17359_ (.A(net3416),
    .B(net4706),
    .Y(_02282_));
 sg13g2_a21oi_1 _17360_ (.A1(net5536),
    .A2(net4706),
    .Y(_01647_),
    .B1(_02282_));
 sg13g2_nor2_1 _17361_ (.A(net3439),
    .B(net4705),
    .Y(_02283_));
 sg13g2_a21oi_1 _17362_ (.A1(net5578),
    .A2(net4705),
    .Y(_01648_),
    .B1(_02283_));
 sg13g2_nor2_1 _17363_ (.A(net3827),
    .B(net4706),
    .Y(_02284_));
 sg13g2_a21oi_1 _17364_ (.A1(net5627),
    .A2(net4706),
    .Y(_01649_),
    .B1(_02284_));
 sg13g2_nor2_1 _17365_ (.A(net4141),
    .B(net4706),
    .Y(_02285_));
 sg13g2_a21oi_1 _17366_ (.A1(net5678),
    .A2(net4705),
    .Y(_01650_),
    .B1(_02285_));
 sg13g2_nor2_1 _17367_ (.A(net4166),
    .B(net4706),
    .Y(_02286_));
 sg13g2_a21oi_1 _17368_ (.A1(net5714),
    .A2(net4705),
    .Y(_01651_),
    .B1(_02286_));
 sg13g2_nor2_1 _17369_ (.A(net3294),
    .B(net4705),
    .Y(_02287_));
 sg13g2_a21oi_1 _17370_ (.A1(net5759),
    .A2(net4705),
    .Y(_01652_),
    .B1(_02287_));
 sg13g2_nor2_1 _17371_ (.A(net5254),
    .B(net5046),
    .Y(_02288_));
 sg13g2_nor2_1 _17372_ (.A(net3392),
    .B(net4704),
    .Y(_02289_));
 sg13g2_a21oi_1 _17373_ (.A1(net5443),
    .A2(net4704),
    .Y(_01653_),
    .B1(_02289_));
 sg13g2_nor2_1 _17374_ (.A(net3365),
    .B(net4703),
    .Y(_02290_));
 sg13g2_a21oi_1 _17375_ (.A1(net5491),
    .A2(net4703),
    .Y(_01654_),
    .B1(_02290_));
 sg13g2_nor2_1 _17376_ (.A(net3903),
    .B(net4704),
    .Y(_02291_));
 sg13g2_a21oi_1 _17377_ (.A1(net5536),
    .A2(net4704),
    .Y(_01655_),
    .B1(_02291_));
 sg13g2_nor2_1 _17378_ (.A(net3581),
    .B(net4703),
    .Y(_02292_));
 sg13g2_a21oi_1 _17379_ (.A1(net5578),
    .A2(net4703),
    .Y(_01656_),
    .B1(_02292_));
 sg13g2_nor2_1 _17380_ (.A(net3299),
    .B(net4704),
    .Y(_02293_));
 sg13g2_a21oi_1 _17381_ (.A1(net5625),
    .A2(net4704),
    .Y(_01657_),
    .B1(_02293_));
 sg13g2_nor2_1 _17382_ (.A(net2864),
    .B(net4703),
    .Y(_02294_));
 sg13g2_a21oi_1 _17383_ (.A1(net5678),
    .A2(net4703),
    .Y(_01658_),
    .B1(_02294_));
 sg13g2_nor2_1 _17384_ (.A(net4113),
    .B(net4704),
    .Y(_02295_));
 sg13g2_a21oi_1 _17385_ (.A1(net5714),
    .A2(net4704),
    .Y(_01659_),
    .B1(_02295_));
 sg13g2_nor2_1 _17386_ (.A(net3419),
    .B(net4703),
    .Y(_02296_));
 sg13g2_a21oi_1 _17387_ (.A1(net5759),
    .A2(net4703),
    .Y(_01660_),
    .B1(_02296_));
 sg13g2_nor2_1 _17388_ (.A(_03120_),
    .B(net5046),
    .Y(_02297_));
 sg13g2_nor2_1 _17389_ (.A(net4135),
    .B(net4702),
    .Y(_02298_));
 sg13g2_a21oi_1 _17390_ (.A1(net5445),
    .A2(net4702),
    .Y(_01661_),
    .B1(_02298_));
 sg13g2_nor2_1 _17391_ (.A(net3914),
    .B(net4701),
    .Y(_02299_));
 sg13g2_a21oi_1 _17392_ (.A1(net5491),
    .A2(net4701),
    .Y(_01662_),
    .B1(_02299_));
 sg13g2_nor2_1 _17393_ (.A(net4073),
    .B(net4702),
    .Y(_02300_));
 sg13g2_a21oi_1 _17394_ (.A1(net5537),
    .A2(net4702),
    .Y(_01663_),
    .B1(_02300_));
 sg13g2_nor2_1 _17395_ (.A(net3521),
    .B(net4701),
    .Y(_02301_));
 sg13g2_a21oi_1 _17396_ (.A1(net5578),
    .A2(net4701),
    .Y(_01664_),
    .B1(_02301_));
 sg13g2_nor2_1 _17397_ (.A(net4069),
    .B(net4702),
    .Y(_02302_));
 sg13g2_a21oi_1 _17398_ (.A1(net5625),
    .A2(net4702),
    .Y(_01665_),
    .B1(_02302_));
 sg13g2_nor2_1 _17399_ (.A(net3850),
    .B(net4701),
    .Y(_02303_));
 sg13g2_a21oi_1 _17400_ (.A1(net5678),
    .A2(net4701),
    .Y(_01666_),
    .B1(_02303_));
 sg13g2_nor2_1 _17401_ (.A(net4057),
    .B(net4702),
    .Y(_02304_));
 sg13g2_a21oi_1 _17402_ (.A1(net5714),
    .A2(net4702),
    .Y(_01667_),
    .B1(_02304_));
 sg13g2_nor2_1 _17403_ (.A(net3822),
    .B(net4701),
    .Y(_02305_));
 sg13g2_a21oi_1 _17404_ (.A1(net5759),
    .A2(net4701),
    .Y(_01668_),
    .B1(_02305_));
 sg13g2_nor2_1 _17405_ (.A(_03109_),
    .B(net5046),
    .Y(_02306_));
 sg13g2_nor2_1 _17406_ (.A(net3944),
    .B(net4700),
    .Y(_02307_));
 sg13g2_a21oi_1 _17407_ (.A1(net5443),
    .A2(net4700),
    .Y(_01669_),
    .B1(_02307_));
 sg13g2_nor2_1 _17408_ (.A(net4096),
    .B(net4700),
    .Y(_02308_));
 sg13g2_a21oi_1 _17409_ (.A1(net5490),
    .A2(net4700),
    .Y(_01670_),
    .B1(_02308_));
 sg13g2_nor2_1 _17410_ (.A(net3967),
    .B(net4700),
    .Y(_02309_));
 sg13g2_a21oi_1 _17411_ (.A1(net5536),
    .A2(net4700),
    .Y(_01671_),
    .B1(_02309_));
 sg13g2_nor2_1 _17412_ (.A(net3382),
    .B(net4699),
    .Y(_02310_));
 sg13g2_a21oi_1 _17413_ (.A1(net5579),
    .A2(net4699),
    .Y(_01672_),
    .B1(_02310_));
 sg13g2_nor2_1 _17414_ (.A(net3682),
    .B(net4700),
    .Y(_02311_));
 sg13g2_a21oi_1 _17415_ (.A1(net5625),
    .A2(net4700),
    .Y(_01673_),
    .B1(_02311_));
 sg13g2_nor2_1 _17416_ (.A(net3257),
    .B(net4699),
    .Y(_02312_));
 sg13g2_a21oi_1 _17417_ (.A1(net5678),
    .A2(net4699),
    .Y(_01674_),
    .B1(_02312_));
 sg13g2_nor2_1 _17418_ (.A(net2984),
    .B(net4699),
    .Y(_02313_));
 sg13g2_a21oi_1 _17419_ (.A1(net5723),
    .A2(net4699),
    .Y(_01675_),
    .B1(_02313_));
 sg13g2_nor2_1 _17420_ (.A(net3615),
    .B(net4699),
    .Y(_02314_));
 sg13g2_a21oi_1 _17421_ (.A1(net5759),
    .A2(net4699),
    .Y(_01676_),
    .B1(_02314_));
 sg13g2_nor2_1 _17422_ (.A(_03201_),
    .B(net5046),
    .Y(_02315_));
 sg13g2_nor2_1 _17423_ (.A(net3503),
    .B(net4698),
    .Y(_02316_));
 sg13g2_a21oi_1 _17424_ (.A1(net5443),
    .A2(net4698),
    .Y(_01677_),
    .B1(_02316_));
 sg13g2_nor2_1 _17425_ (.A(net3384),
    .B(net4698),
    .Y(_02317_));
 sg13g2_a21oi_1 _17426_ (.A1(net5490),
    .A2(net4698),
    .Y(_01678_),
    .B1(_02317_));
 sg13g2_nor2_1 _17427_ (.A(net3332),
    .B(net4698),
    .Y(_02318_));
 sg13g2_a21oi_1 _17428_ (.A1(net5536),
    .A2(net4698),
    .Y(_01679_),
    .B1(_02318_));
 sg13g2_nor2_1 _17429_ (.A(net3630),
    .B(net4697),
    .Y(_02319_));
 sg13g2_a21oi_1 _17430_ (.A1(net5579),
    .A2(net4697),
    .Y(_01680_),
    .B1(_02319_));
 sg13g2_nor2_1 _17431_ (.A(net3790),
    .B(net4698),
    .Y(_02320_));
 sg13g2_a21oi_1 _17432_ (.A1(net5624),
    .A2(net4698),
    .Y(_01681_),
    .B1(_02320_));
 sg13g2_nor2_1 _17433_ (.A(net3579),
    .B(net4697),
    .Y(_02321_));
 sg13g2_a21oi_1 _17434_ (.A1(net5678),
    .A2(net4697),
    .Y(_01682_),
    .B1(_02321_));
 sg13g2_nor2_1 _17435_ (.A(net4032),
    .B(net4697),
    .Y(_02322_));
 sg13g2_a21oi_1 _17436_ (.A1(net5723),
    .A2(net4697),
    .Y(_01683_),
    .B1(_02322_));
 sg13g2_nor2_1 _17437_ (.A(net3981),
    .B(net4697),
    .Y(_02323_));
 sg13g2_a21oi_1 _17438_ (.A1(net5770),
    .A2(net4697),
    .Y(_01684_),
    .B1(_02323_));
 sg13g2_nor2_1 _17439_ (.A(_03067_),
    .B(net5046),
    .Y(_02324_));
 sg13g2_nor2_1 _17440_ (.A(net3929),
    .B(net4696),
    .Y(_02325_));
 sg13g2_a21oi_1 _17441_ (.A1(net5443),
    .A2(net4696),
    .Y(_01685_),
    .B1(_02325_));
 sg13g2_nor2_1 _17442_ (.A(net4101),
    .B(net4696),
    .Y(_02326_));
 sg13g2_a21oi_1 _17443_ (.A1(net5490),
    .A2(net4696),
    .Y(_01686_),
    .B1(_02326_));
 sg13g2_nor2_1 _17444_ (.A(net4039),
    .B(net4696),
    .Y(_02327_));
 sg13g2_a21oi_1 _17445_ (.A1(net5535),
    .A2(net4696),
    .Y(_01687_),
    .B1(_02327_));
 sg13g2_nor2_1 _17446_ (.A(net3496),
    .B(net4695),
    .Y(_02328_));
 sg13g2_a21oi_1 _17447_ (.A1(net5579),
    .A2(net4695),
    .Y(_01688_),
    .B1(_02328_));
 sg13g2_nor2_1 _17448_ (.A(net3001),
    .B(net4696),
    .Y(_02329_));
 sg13g2_a21oi_1 _17449_ (.A1(net5633),
    .A2(net4696),
    .Y(_01689_),
    .B1(_02329_));
 sg13g2_nor2_1 _17450_ (.A(net3863),
    .B(net4695),
    .Y(_02330_));
 sg13g2_a21oi_1 _17451_ (.A1(net5678),
    .A2(net4695),
    .Y(_01690_),
    .B1(_02330_));
 sg13g2_nor2_1 _17452_ (.A(net3025),
    .B(net4695),
    .Y(_02331_));
 sg13g2_a21oi_1 _17453_ (.A1(net5723),
    .A2(net4695),
    .Y(_01691_),
    .B1(_02331_));
 sg13g2_nor2_1 _17454_ (.A(net3306),
    .B(net4695),
    .Y(_02332_));
 sg13g2_a21oi_1 _17455_ (.A1(net5770),
    .A2(net4695),
    .Y(_01692_),
    .B1(_02332_));
 sg13g2_nor2_1 _17456_ (.A(net5142),
    .B(net5252),
    .Y(_02333_));
 sg13g2_nor2_1 _17457_ (.A(net3792),
    .B(net4694),
    .Y(_02334_));
 sg13g2_a21oi_1 _17458_ (.A1(net5438),
    .A2(net4694),
    .Y(_01693_),
    .B1(_02334_));
 sg13g2_nor2_1 _17459_ (.A(net3668),
    .B(net4694),
    .Y(_02335_));
 sg13g2_a21oi_1 _17460_ (.A1(net5482),
    .A2(net4694),
    .Y(_01694_),
    .B1(_02335_));
 sg13g2_nor2_1 _17461_ (.A(net3998),
    .B(net4694),
    .Y(_02336_));
 sg13g2_a21oi_1 _17462_ (.A1(net5529),
    .A2(net4694),
    .Y(_01695_),
    .B1(_02336_));
 sg13g2_nor2_1 _17463_ (.A(net3818),
    .B(_02333_),
    .Y(_02337_));
 sg13g2_a21oi_1 _17464_ (.A1(net5573),
    .A2(net4694),
    .Y(_01696_),
    .B1(_02337_));
 sg13g2_nor2_1 _17465_ (.A(net3395),
    .B(net4693),
    .Y(_02338_));
 sg13g2_a21oi_1 _17466_ (.A1(net5628),
    .A2(net4693),
    .Y(_01697_),
    .B1(_02338_));
 sg13g2_nor2_1 _17467_ (.A(net3490),
    .B(net4693),
    .Y(_02339_));
 sg13g2_a21oi_1 _17468_ (.A1(net5671),
    .A2(net4693),
    .Y(_01698_),
    .B1(_02339_));
 sg13g2_nor2_1 _17469_ (.A(net4140),
    .B(net4693),
    .Y(_02340_));
 sg13g2_a21oi_1 _17470_ (.A1(net5707),
    .A2(net4693),
    .Y(_01699_),
    .B1(_02340_));
 sg13g2_nor2_1 _17471_ (.A(net3980),
    .B(net4693),
    .Y(_02341_));
 sg13g2_a21oi_1 _17472_ (.A1(net5753),
    .A2(net4693),
    .Y(_01700_),
    .B1(_02341_));
 sg13g2_nor2_1 _17473_ (.A(_02939_),
    .B(net5045),
    .Y(_02342_));
 sg13g2_nor2_1 _17474_ (.A(net3623),
    .B(net4691),
    .Y(_02343_));
 sg13g2_a21oi_1 _17475_ (.A1(net5445),
    .A2(net4691),
    .Y(_01701_),
    .B1(_02343_));
 sg13g2_nor2_1 _17476_ (.A(net3838),
    .B(net4692),
    .Y(_02344_));
 sg13g2_a21oi_1 _17477_ (.A1(net5486),
    .A2(net4692),
    .Y(_01702_),
    .B1(_02344_));
 sg13g2_nor2_1 _17478_ (.A(net3749),
    .B(net4691),
    .Y(_02345_));
 sg13g2_a21oi_1 _17479_ (.A1(net5533),
    .A2(net4691),
    .Y(_01703_),
    .B1(_02345_));
 sg13g2_nor2_1 _17480_ (.A(net3617),
    .B(net4691),
    .Y(_02346_));
 sg13g2_a21oi_1 _17481_ (.A1(net5576),
    .A2(net4691),
    .Y(_01704_),
    .B1(_02346_));
 sg13g2_nor2_1 _17482_ (.A(net3642),
    .B(net4692),
    .Y(_02347_));
 sg13g2_a21oi_1 _17483_ (.A1(net5624),
    .A2(net4692),
    .Y(_01705_),
    .B1(_02347_));
 sg13g2_nor2_1 _17484_ (.A(net3499),
    .B(_02342_),
    .Y(_02348_));
 sg13g2_a21oi_1 _17485_ (.A1(net5667),
    .A2(net4692),
    .Y(_01706_),
    .B1(_02348_));
 sg13g2_nor2_1 _17486_ (.A(net3536),
    .B(net4691),
    .Y(_02349_));
 sg13g2_a21oi_1 _17487_ (.A1(net5715),
    .A2(net4691),
    .Y(_01707_),
    .B1(_02349_));
 sg13g2_nor2_1 _17488_ (.A(net4042),
    .B(net4692),
    .Y(_02350_));
 sg13g2_a21oi_1 _17489_ (.A1(net5760),
    .A2(net4692),
    .Y(_01708_),
    .B1(_02350_));
 sg13g2_nor2_1 _17490_ (.A(_03017_),
    .B(net5045),
    .Y(_02351_));
 sg13g2_nor2_1 _17491_ (.A(net3544),
    .B(net4690),
    .Y(_02352_));
 sg13g2_a21oi_1 _17492_ (.A1(net5445),
    .A2(net4690),
    .Y(_01709_),
    .B1(_02352_));
 sg13g2_nor2_1 _17493_ (.A(net4053),
    .B(net4689),
    .Y(_02353_));
 sg13g2_a21oi_1 _17494_ (.A1(net5486),
    .A2(net4689),
    .Y(_01710_),
    .B1(_02353_));
 sg13g2_nor2_1 _17495_ (.A(net3697),
    .B(net4689),
    .Y(_02354_));
 sg13g2_a21oi_1 _17496_ (.A1(net5533),
    .A2(net4689),
    .Y(_01711_),
    .B1(_02354_));
 sg13g2_nor2_1 _17497_ (.A(net3678),
    .B(net4689),
    .Y(_02355_));
 sg13g2_a21oi_1 _17498_ (.A1(net5575),
    .A2(net4689),
    .Y(_01712_),
    .B1(_02355_));
 sg13g2_nor2_1 _17499_ (.A(net3755),
    .B(net4690),
    .Y(_02356_));
 sg13g2_a21oi_1 _17500_ (.A1(net5624),
    .A2(net4690),
    .Y(_01713_),
    .B1(_02356_));
 sg13g2_nor2_1 _17501_ (.A(net3637),
    .B(net4689),
    .Y(_02357_));
 sg13g2_a21oi_1 _17502_ (.A1(net5667),
    .A2(net4689),
    .Y(_01714_),
    .B1(_02357_));
 sg13g2_nor2_1 _17503_ (.A(net3517),
    .B(net4690),
    .Y(_02358_));
 sg13g2_a21oi_1 _17504_ (.A1(net5715),
    .A2(net4690),
    .Y(_01715_),
    .B1(_02358_));
 sg13g2_nor2_1 _17505_ (.A(net4005),
    .B(net4690),
    .Y(_02359_));
 sg13g2_a21oi_1 _17506_ (.A1(net5760),
    .A2(net4690),
    .Y(_01716_),
    .B1(_02359_));
 sg13g2_nor2_1 _17507_ (.A(_02981_),
    .B(net5045),
    .Y(_02360_));
 sg13g2_nor2_1 _17508_ (.A(net4056),
    .B(net4686),
    .Y(_02361_));
 sg13g2_a21oi_1 _17509_ (.A1(net5445),
    .A2(net4686),
    .Y(_01717_),
    .B1(_02361_));
 sg13g2_nor2_1 _17510_ (.A(net3388),
    .B(net4688),
    .Y(_02362_));
 sg13g2_a21oi_1 _17511_ (.A1(net5486),
    .A2(net4688),
    .Y(_01718_),
    .B1(_02362_));
 sg13g2_nor2_1 _17512_ (.A(net3861),
    .B(net4686),
    .Y(_02363_));
 sg13g2_a21oi_1 _17513_ (.A1(net5533),
    .A2(net4686),
    .Y(_01719_),
    .B1(_02363_));
 sg13g2_nor2_1 _17514_ (.A(net3816),
    .B(net4686),
    .Y(_02364_));
 sg13g2_a21oi_1 _17515_ (.A1(net5575),
    .A2(net4686),
    .Y(_01720_),
    .B1(_02364_));
 sg13g2_nor2_1 _17516_ (.A(net3220),
    .B(net4686),
    .Y(_02365_));
 sg13g2_a21oi_1 _17517_ (.A1(net5624),
    .A2(net4686),
    .Y(_01721_),
    .B1(_02365_));
 sg13g2_nor2_1 _17518_ (.A(net3853),
    .B(net4688),
    .Y(_02366_));
 sg13g2_a21oi_1 _17519_ (.A1(net5667),
    .A2(net4688),
    .Y(_01722_),
    .B1(_02366_));
 sg13g2_nor2_1 _17520_ (.A(net4009),
    .B(net4687),
    .Y(_02367_));
 sg13g2_a21oi_1 _17521_ (.A1(net5714),
    .A2(net4687),
    .Y(_01723_),
    .B1(_02367_));
 sg13g2_nor2_1 _17522_ (.A(net3951),
    .B(net4687),
    .Y(_02368_));
 sg13g2_a21oi_1 _17523_ (.A1(net5760),
    .A2(net4687),
    .Y(_01724_),
    .B1(_02368_));
 sg13g2_nor2_1 _17524_ (.A(_02964_),
    .B(net5045),
    .Y(_02369_));
 sg13g2_nor2_1 _17525_ (.A(net3513),
    .B(net4683),
    .Y(_02370_));
 sg13g2_a21oi_1 _17526_ (.A1(net5445),
    .A2(net4683),
    .Y(_01725_),
    .B1(_02370_));
 sg13g2_nor2_1 _17527_ (.A(net3563),
    .B(net4685),
    .Y(_02371_));
 sg13g2_a21oi_1 _17528_ (.A1(net5486),
    .A2(net4685),
    .Y(_01726_),
    .B1(_02371_));
 sg13g2_nor2_1 _17529_ (.A(net4001),
    .B(net4683),
    .Y(_02372_));
 sg13g2_a21oi_1 _17530_ (.A1(net5533),
    .A2(net4683),
    .Y(_01727_),
    .B1(_02372_));
 sg13g2_nor2_1 _17531_ (.A(net3709),
    .B(net4683),
    .Y(_02373_));
 sg13g2_a21oi_1 _17532_ (.A1(net5575),
    .A2(net4683),
    .Y(_01728_),
    .B1(_02373_));
 sg13g2_nor2_1 _17533_ (.A(net3618),
    .B(net4683),
    .Y(_02374_));
 sg13g2_a21oi_1 _17534_ (.A1(net5625),
    .A2(net4683),
    .Y(_01729_),
    .B1(_02374_));
 sg13g2_nor2_1 _17535_ (.A(net4063),
    .B(net4685),
    .Y(_02375_));
 sg13g2_a21oi_1 _17536_ (.A1(net5667),
    .A2(net4685),
    .Y(_01730_),
    .B1(_02375_));
 sg13g2_nor2_1 _17537_ (.A(net3628),
    .B(net4684),
    .Y(_02376_));
 sg13g2_a21oi_1 _17538_ (.A1(net5714),
    .A2(net4684),
    .Y(_01731_),
    .B1(_02376_));
 sg13g2_nor2_1 _17539_ (.A(net3702),
    .B(net4684),
    .Y(_02377_));
 sg13g2_a21oi_1 _17540_ (.A1(net5760),
    .A2(net4684),
    .Y(_01732_),
    .B1(_02377_));
 sg13g2_nor2_1 _17541_ (.A(_03467_),
    .B(net5045),
    .Y(_02378_));
 sg13g2_nor2_1 _17542_ (.A(net3330),
    .B(net4682),
    .Y(_02379_));
 sg13g2_a21oi_1 _17543_ (.A1(net5444),
    .A2(net4682),
    .Y(_01733_),
    .B1(_02379_));
 sg13g2_nor2_1 _17544_ (.A(net3826),
    .B(net4682),
    .Y(_02380_));
 sg13g2_a21oi_1 _17545_ (.A1(net5489),
    .A2(net4682),
    .Y(_01734_),
    .B1(_02380_));
 sg13g2_nor2_1 _17546_ (.A(net3608),
    .B(net4682),
    .Y(_02381_));
 sg13g2_a21oi_1 _17547_ (.A1(net5535),
    .A2(_02378_),
    .Y(_01735_),
    .B1(_02381_));
 sg13g2_nor2_1 _17548_ (.A(net3273),
    .B(net4681),
    .Y(_02382_));
 sg13g2_a21oi_1 _17549_ (.A1(net5578),
    .A2(net4681),
    .Y(_01736_),
    .B1(_02382_));
 sg13g2_nor2_1 _17550_ (.A(net3537),
    .B(net4681),
    .Y(_02383_));
 sg13g2_a21oi_1 _17551_ (.A1(net5624),
    .A2(net4682),
    .Y(_01737_),
    .B1(_02383_));
 sg13g2_nor2_1 _17552_ (.A(net3450),
    .B(net4681),
    .Y(_02384_));
 sg13g2_a21oi_1 _17553_ (.A1(net5667),
    .A2(net4681),
    .Y(_01738_),
    .B1(_02384_));
 sg13g2_nor2_1 _17554_ (.A(net3235),
    .B(net4681),
    .Y(_02385_));
 sg13g2_a21oi_1 _17555_ (.A1(net5715),
    .A2(net4682),
    .Y(_01739_),
    .B1(_02385_));
 sg13g2_nor2_1 _17556_ (.A(net3619),
    .B(net4681),
    .Y(_02386_));
 sg13g2_a21oi_1 _17557_ (.A1(net5759),
    .A2(net4681),
    .Y(_01740_),
    .B1(_02386_));
 sg13g2_nor2_1 _17558_ (.A(_03212_),
    .B(net5045),
    .Y(_02387_));
 sg13g2_nor2_1 _17559_ (.A(net3669),
    .B(net4680),
    .Y(_02388_));
 sg13g2_a21oi_1 _17560_ (.A1(net5444),
    .A2(net4680),
    .Y(_01741_),
    .B1(_02388_));
 sg13g2_nor2_1 _17561_ (.A(net3687),
    .B(_02387_),
    .Y(_02389_));
 sg13g2_a21oi_1 _17562_ (.A1(net5489),
    .A2(net4680),
    .Y(_01742_),
    .B1(_02389_));
 sg13g2_nor2_1 _17563_ (.A(net3890),
    .B(net4680),
    .Y(_02390_));
 sg13g2_a21oi_1 _17564_ (.A1(net5535),
    .A2(net4680),
    .Y(_01743_),
    .B1(_02390_));
 sg13g2_nor2_1 _17565_ (.A(net3548),
    .B(net4679),
    .Y(_02391_));
 sg13g2_a21oi_1 _17566_ (.A1(net5578),
    .A2(net4679),
    .Y(_01744_),
    .B1(_02391_));
 sg13g2_nor2_1 _17567_ (.A(net4038),
    .B(net4679),
    .Y(_02392_));
 sg13g2_a21oi_1 _17568_ (.A1(net5624),
    .A2(net4679),
    .Y(_01745_),
    .B1(_02392_));
 sg13g2_nor2_1 _17569_ (.A(net3469),
    .B(net4679),
    .Y(_02393_));
 sg13g2_a21oi_1 _17570_ (.A1(net5667),
    .A2(net4679),
    .Y(_01746_),
    .B1(_02393_));
 sg13g2_nor2_1 _17571_ (.A(net3638),
    .B(net4680),
    .Y(_02394_));
 sg13g2_a21oi_1 _17572_ (.A1(net5715),
    .A2(net4680),
    .Y(_01747_),
    .B1(_02394_));
 sg13g2_nor2_1 _17573_ (.A(net4002),
    .B(net4679),
    .Y(_02395_));
 sg13g2_a21oi_1 _17574_ (.A1(net5759),
    .A2(net4679),
    .Y(_01748_),
    .B1(_02395_));
 sg13g2_nor2_1 _17575_ (.A(_03375_),
    .B(net5045),
    .Y(_02396_));
 sg13g2_nor2_1 _17576_ (.A(net3941),
    .B(net4678),
    .Y(_02397_));
 sg13g2_a21oi_1 _17577_ (.A1(net5445),
    .A2(net4678),
    .Y(_01749_),
    .B1(_02397_));
 sg13g2_nor2_1 _17578_ (.A(net4151),
    .B(net4678),
    .Y(_02398_));
 sg13g2_a21oi_1 _17579_ (.A1(net5491),
    .A2(net4678),
    .Y(_01750_),
    .B1(_02398_));
 sg13g2_nor2_1 _17580_ (.A(net3535),
    .B(net4678),
    .Y(_02399_));
 sg13g2_a21oi_1 _17581_ (.A1(net5535),
    .A2(net4678),
    .Y(_01751_),
    .B1(_02399_));
 sg13g2_nor2_1 _17582_ (.A(net3104),
    .B(net4677),
    .Y(_02400_));
 sg13g2_a21oi_1 _17583_ (.A1(net5578),
    .A2(net4677),
    .Y(_01752_),
    .B1(_02400_));
 sg13g2_nor2_1 _17584_ (.A(net3252),
    .B(net4678),
    .Y(_02401_));
 sg13g2_a21oi_1 _17585_ (.A1(net5624),
    .A2(net4678),
    .Y(_01753_),
    .B1(_02401_));
 sg13g2_nor2_1 _17586_ (.A(net3502),
    .B(net4677),
    .Y(_02402_));
 sg13g2_a21oi_1 _17587_ (.A1(net5667),
    .A2(net4677),
    .Y(_01754_),
    .B1(_02402_));
 sg13g2_nor2_1 _17588_ (.A(net4138),
    .B(net4677),
    .Y(_02403_));
 sg13g2_a21oi_1 _17589_ (.A1(net5714),
    .A2(net4677),
    .Y(_01755_),
    .B1(_02403_));
 sg13g2_nor2_1 _17590_ (.A(net3705),
    .B(net4677),
    .Y(_02404_));
 sg13g2_a21oi_1 _17591_ (.A1(net5759),
    .A2(net4677),
    .Y(_01756_),
    .B1(_02404_));
 sg13g2_nor2_1 _17592_ (.A(net5240),
    .B(net5045),
    .Y(_02405_));
 sg13g2_nor2_1 _17593_ (.A(net3997),
    .B(net4676),
    .Y(_02406_));
 sg13g2_a21oi_1 _17594_ (.A1(net5445),
    .A2(net4676),
    .Y(_01757_),
    .B1(_02406_));
 sg13g2_nor2_1 _17595_ (.A(net3776),
    .B(net4676),
    .Y(_02407_));
 sg13g2_a21oi_1 _17596_ (.A1(net5489),
    .A2(net4676),
    .Y(_01758_),
    .B1(_02407_));
 sg13g2_nor2_1 _17597_ (.A(net4085),
    .B(net4676),
    .Y(_02408_));
 sg13g2_a21oi_1 _17598_ (.A1(net5535),
    .A2(net4676),
    .Y(_01759_),
    .B1(_02408_));
 sg13g2_nor2_1 _17599_ (.A(net3707),
    .B(net4675),
    .Y(_02409_));
 sg13g2_a21oi_1 _17600_ (.A1(net5578),
    .A2(net4675),
    .Y(_01760_),
    .B1(_02409_));
 sg13g2_nor2_1 _17601_ (.A(net3479),
    .B(net4676),
    .Y(_02410_));
 sg13g2_a21oi_1 _17602_ (.A1(net5624),
    .A2(net4676),
    .Y(_01761_),
    .B1(_02410_));
 sg13g2_nor2_1 _17603_ (.A(net3402),
    .B(net4675),
    .Y(_02411_));
 sg13g2_a21oi_1 _17604_ (.A1(net5667),
    .A2(net4675),
    .Y(_01762_),
    .B1(_02411_));
 sg13g2_nor2_1 _17605_ (.A(net3358),
    .B(net4675),
    .Y(_02412_));
 sg13g2_a21oi_1 _17606_ (.A1(net5714),
    .A2(net4675),
    .Y(_01763_),
    .B1(_02412_));
 sg13g2_nor2_1 _17607_ (.A(net3856),
    .B(net4675),
    .Y(_02413_));
 sg13g2_a21oi_1 _17608_ (.A1(net5759),
    .A2(net4675),
    .Y(_01764_),
    .B1(_02413_));
 sg13g2_nand2_1 _17609_ (.Y(_02414_),
    .A(net5249),
    .B(net5198));
 sg13g2_nand2_1 _17610_ (.Y(_02415_),
    .A(net2693),
    .B(net4868));
 sg13g2_o21ai_1 _17611_ (.B1(_02415_),
    .Y(_01765_),
    .A1(net5460),
    .A2(net4868));
 sg13g2_nand2_1 _17612_ (.Y(_02416_),
    .A(net3051),
    .B(net4869));
 sg13g2_o21ai_1 _17613_ (.B1(_02416_),
    .Y(_01766_),
    .A1(net5507),
    .A2(net4869));
 sg13g2_nand2_1 _17614_ (.Y(_02417_),
    .A(net2541),
    .B(net4869));
 sg13g2_o21ai_1 _17615_ (.B1(_02417_),
    .Y(_01767_),
    .A1(net5554),
    .A2(net4869));
 sg13g2_nand2_1 _17616_ (.Y(_02418_),
    .A(net2469),
    .B(net4869));
 sg13g2_o21ai_1 _17617_ (.B1(_02418_),
    .Y(_01768_),
    .A1(net5600),
    .A2(net4869));
 sg13g2_nand2_1 _17618_ (.Y(_02419_),
    .A(net3436),
    .B(net4869));
 sg13g2_o21ai_1 _17619_ (.B1(_02419_),
    .Y(_01769_),
    .A1(net5645),
    .A2(net4869));
 sg13g2_nand2_1 _17620_ (.Y(_02420_),
    .A(net2161),
    .B(net4868));
 sg13g2_o21ai_1 _17621_ (.B1(_02420_),
    .Y(_01770_),
    .A1(net5688),
    .A2(net4868));
 sg13g2_nand2_1 _17622_ (.Y(_02421_),
    .A(net2349),
    .B(net4868));
 sg13g2_o21ai_1 _17623_ (.B1(_02421_),
    .Y(_01771_),
    .A1(net5734),
    .A2(net4868));
 sg13g2_nand2_1 _17624_ (.Y(_02422_),
    .A(net2983),
    .B(net4868));
 sg13g2_o21ai_1 _17625_ (.B1(_02422_),
    .Y(_01772_),
    .A1(net5779),
    .A2(net4868));
 sg13g2_nor2_1 _17626_ (.A(_03109_),
    .B(net5210),
    .Y(_02423_));
 sg13g2_nor2_1 _17627_ (.A(net3053),
    .B(net4866),
    .Y(_02424_));
 sg13g2_a21oi_1 _17628_ (.A1(net5452),
    .A2(net4866),
    .Y(_01773_),
    .B1(_02424_));
 sg13g2_nor2_1 _17629_ (.A(net4092),
    .B(net4866),
    .Y(_02425_));
 sg13g2_a21oi_1 _17630_ (.A1(net5497),
    .A2(net4866),
    .Y(_01774_),
    .B1(_02425_));
 sg13g2_nor2_1 _17631_ (.A(net4034),
    .B(net4867),
    .Y(_02426_));
 sg13g2_a21oi_1 _17632_ (.A1(net5552),
    .A2(net4867),
    .Y(_01775_),
    .B1(_02426_));
 sg13g2_nor2_1 _17633_ (.A(net3819),
    .B(net4867),
    .Y(_02427_));
 sg13g2_a21oi_1 _17634_ (.A1(net5596),
    .A2(net4867),
    .Y(_01776_),
    .B1(_02427_));
 sg13g2_nor2_1 _17635_ (.A(net3444),
    .B(net4867),
    .Y(_02428_));
 sg13g2_a21oi_1 _17636_ (.A1(net5642),
    .A2(net4867),
    .Y(_01777_),
    .B1(_02428_));
 sg13g2_nor2_1 _17637_ (.A(net3884),
    .B(net4866),
    .Y(_02429_));
 sg13g2_a21oi_1 _17638_ (.A1(net5687),
    .A2(net4866),
    .Y(_01778_),
    .B1(_02429_));
 sg13g2_nor2_1 _17639_ (.A(net3877),
    .B(net4866),
    .Y(_02430_));
 sg13g2_a21oi_1 _17640_ (.A1(net5732),
    .A2(net4866),
    .Y(_01779_),
    .B1(_02430_));
 sg13g2_nor2_1 _17641_ (.A(net3058),
    .B(net4867),
    .Y(_02431_));
 sg13g2_a21oi_1 _17642_ (.A1(net5783),
    .A2(net4867),
    .Y(_01780_),
    .B1(_02431_));
 sg13g2_nand2_1 _17643_ (.Y(_02432_),
    .A(_03079_),
    .B(net5198));
 sg13g2_nand2_1 _17644_ (.Y(_02433_),
    .A(net2981),
    .B(net4864));
 sg13g2_o21ai_1 _17645_ (.B1(_02433_),
    .Y(_01781_),
    .A1(net5462),
    .A2(net4864));
 sg13g2_nand2_1 _17646_ (.Y(_02434_),
    .A(net2696),
    .B(net4865));
 sg13g2_o21ai_1 _17647_ (.B1(_02434_),
    .Y(_01782_),
    .A1(net5507),
    .A2(net4865));
 sg13g2_nand2_1 _17648_ (.Y(_02435_),
    .A(net3114),
    .B(net4865));
 sg13g2_o21ai_1 _17649_ (.B1(_02435_),
    .Y(_01783_),
    .A1(net5554),
    .A2(net4865));
 sg13g2_nand2_1 _17650_ (.Y(_02436_),
    .A(net2650),
    .B(net4865));
 sg13g2_o21ai_1 _17651_ (.B1(_02436_),
    .Y(_01784_),
    .A1(net5600),
    .A2(net4865));
 sg13g2_nand2_1 _17652_ (.Y(_02437_),
    .A(net2234),
    .B(net4865));
 sg13g2_o21ai_1 _17653_ (.B1(_02437_),
    .Y(_01785_),
    .A1(net5645),
    .A2(net4865));
 sg13g2_nand2_1 _17654_ (.Y(_02438_),
    .A(net2272),
    .B(net4864));
 sg13g2_o21ai_1 _17655_ (.B1(_02438_),
    .Y(_01786_),
    .A1(net5688),
    .A2(net4864));
 sg13g2_nand2_1 _17656_ (.Y(_02439_),
    .A(net2194),
    .B(net4864));
 sg13g2_o21ai_1 _17657_ (.B1(_02439_),
    .Y(_01787_),
    .A1(net5734),
    .A2(net4864));
 sg13g2_nand2_1 _17658_ (.Y(_02440_),
    .A(net2955),
    .B(net4864));
 sg13g2_o21ai_1 _17659_ (.B1(_02440_),
    .Y(_01788_),
    .A1(net5779),
    .A2(net4864));
 sg13g2_nand2_1 _17660_ (.Y(_02441_),
    .A(net5253),
    .B(net5198));
 sg13g2_nand2_1 _17661_ (.Y(_02442_),
    .A(net2656),
    .B(net4862));
 sg13g2_o21ai_1 _17662_ (.B1(_02442_),
    .Y(_01789_),
    .A1(net5462),
    .A2(net4862));
 sg13g2_nand2_1 _17663_ (.Y(_02443_),
    .A(net3233),
    .B(net4863));
 sg13g2_o21ai_1 _17664_ (.B1(_02443_),
    .Y(_01790_),
    .A1(net5507),
    .A2(net4863));
 sg13g2_nand2_1 _17665_ (.Y(_02444_),
    .A(net2748),
    .B(net4863));
 sg13g2_o21ai_1 _17666_ (.B1(_02444_),
    .Y(_01791_),
    .A1(net5554),
    .A2(net4863));
 sg13g2_nand2_1 _17667_ (.Y(_02445_),
    .A(net2247),
    .B(net4863));
 sg13g2_o21ai_1 _17668_ (.B1(_02445_),
    .Y(_01792_),
    .A1(net5600),
    .A2(net4863));
 sg13g2_nand2_1 _17669_ (.Y(_02446_),
    .A(net2952),
    .B(net4863));
 sg13g2_o21ai_1 _17670_ (.B1(_02446_),
    .Y(_01793_),
    .A1(net5645),
    .A2(net4863));
 sg13g2_nand2_1 _17671_ (.Y(_02447_),
    .A(net3376),
    .B(net4862));
 sg13g2_o21ai_1 _17672_ (.B1(_02447_),
    .Y(_01794_),
    .A1(net5688),
    .A2(net4862));
 sg13g2_nand2_1 _17673_ (.Y(_02448_),
    .A(net2843),
    .B(net4862));
 sg13g2_o21ai_1 _17674_ (.B1(_02448_),
    .Y(_01795_),
    .A1(net5734),
    .A2(net4862));
 sg13g2_nand2_1 _17675_ (.Y(_02449_),
    .A(net2780),
    .B(net4862));
 sg13g2_o21ai_1 _17676_ (.B1(_02449_),
    .Y(_01796_),
    .A1(net5779),
    .A2(net4862));
 sg13g2_nand2_2 _17677_ (.Y(_02450_),
    .A(net5235),
    .B(net5199));
 sg13g2_nand2_1 _17678_ (.Y(_02451_),
    .A(net2241),
    .B(net4861));
 sg13g2_o21ai_1 _17679_ (.B1(_02451_),
    .Y(_01797_),
    .A1(net5457),
    .A2(net4861));
 sg13g2_nand2_1 _17680_ (.Y(_02452_),
    .A(net2334),
    .B(_02450_));
 sg13g2_o21ai_1 _17681_ (.B1(_02452_),
    .Y(_01798_),
    .A1(net5505),
    .A2(net4860));
 sg13g2_nand2_1 _17682_ (.Y(_02453_),
    .A(net3179),
    .B(net4861));
 sg13g2_o21ai_1 _17683_ (.B1(_02453_),
    .Y(_01799_),
    .A1(net5549),
    .A2(net4860));
 sg13g2_nand2_1 _17684_ (.Y(_02454_),
    .A(net2593),
    .B(net4860));
 sg13g2_o21ai_1 _17685_ (.B1(_02454_),
    .Y(_01800_),
    .A1(net5592),
    .A2(net4860));
 sg13g2_nand2_1 _17686_ (.Y(_02455_),
    .A(net2229),
    .B(net4860));
 sg13g2_o21ai_1 _17687_ (.B1(_02455_),
    .Y(_01801_),
    .A1(net5638),
    .A2(net4860));
 sg13g2_nand2_1 _17688_ (.Y(_02456_),
    .A(net3295),
    .B(net4861));
 sg13g2_o21ai_1 _17689_ (.B1(_02456_),
    .Y(_01802_),
    .A1(net5684),
    .A2(net4861));
 sg13g2_nand2_1 _17690_ (.Y(_02457_),
    .A(net2538),
    .B(net4861));
 sg13g2_o21ai_1 _17691_ (.B1(_02457_),
    .Y(_01803_),
    .A1(net5728),
    .A2(net4861));
 sg13g2_nand2_1 _17692_ (.Y(_02458_),
    .A(net2686),
    .B(net4860));
 sg13g2_o21ai_1 _17693_ (.B1(_02458_),
    .Y(_01804_),
    .A1(net5775),
    .A2(net4860));
 sg13g2_nand2_1 _17694_ (.Y(_02459_),
    .A(net5234),
    .B(net5198));
 sg13g2_nand2_1 _17695_ (.Y(_02460_),
    .A(net2702),
    .B(net4859));
 sg13g2_o21ai_1 _17696_ (.B1(_02460_),
    .Y(_01805_),
    .A1(net5457),
    .A2(net4859));
 sg13g2_nand2_1 _17697_ (.Y(_02461_),
    .A(net3229),
    .B(net4858));
 sg13g2_o21ai_1 _17698_ (.B1(_02461_),
    .Y(_01806_),
    .A1(net5505),
    .A2(net4858));
 sg13g2_nand2_1 _17699_ (.Y(_02462_),
    .A(net2544),
    .B(_02459_));
 sg13g2_o21ai_1 _17700_ (.B1(_02462_),
    .Y(_01807_),
    .A1(net5548),
    .A2(net4858));
 sg13g2_nand2_1 _17701_ (.Y(_02463_),
    .A(net2490),
    .B(net4858));
 sg13g2_o21ai_1 _17702_ (.B1(_02463_),
    .Y(_01808_),
    .A1(net5592),
    .A2(net4858));
 sg13g2_nand2_1 _17703_ (.Y(_02464_),
    .A(net2975),
    .B(net4858));
 sg13g2_o21ai_1 _17704_ (.B1(_02464_),
    .Y(_01809_),
    .A1(net5638),
    .A2(net4858));
 sg13g2_nand2_1 _17705_ (.Y(_02465_),
    .A(net2346),
    .B(net4859));
 sg13g2_o21ai_1 _17706_ (.B1(_02465_),
    .Y(_01810_),
    .A1(net5683),
    .A2(net4859));
 sg13g2_nand2_1 _17707_ (.Y(_02466_),
    .A(net2479),
    .B(net4858));
 sg13g2_o21ai_1 _17708_ (.B1(_02466_),
    .Y(_01811_),
    .A1(net5728),
    .A2(net4859));
 sg13g2_nand2_1 _17709_ (.Y(_02467_),
    .A(net2509),
    .B(net4859));
 sg13g2_o21ai_1 _17710_ (.B1(_02467_),
    .Y(_01812_),
    .A1(net5775),
    .A2(net4859));
 sg13g2_nand2_1 _17711_ (.Y(_02468_),
    .A(net5236),
    .B(net5199));
 sg13g2_nand2_1 _17712_ (.Y(_02469_),
    .A(net3069),
    .B(net4857));
 sg13g2_o21ai_1 _17713_ (.B1(_02469_),
    .Y(_01813_),
    .A1(net5457),
    .A2(net4857));
 sg13g2_nand2_1 _17714_ (.Y(_02470_),
    .A(net2927),
    .B(net4856));
 sg13g2_o21ai_1 _17715_ (.B1(_02470_),
    .Y(_01814_),
    .A1(net5505),
    .A2(net4856));
 sg13g2_nand2_1 _17716_ (.Y(_02471_),
    .A(net2230),
    .B(net4857));
 sg13g2_o21ai_1 _17717_ (.B1(_02471_),
    .Y(_01815_),
    .A1(net5548),
    .A2(_02468_));
 sg13g2_nand2_1 _17718_ (.Y(_02472_),
    .A(net2282),
    .B(net4856));
 sg13g2_o21ai_1 _17719_ (.B1(_02472_),
    .Y(_01816_),
    .A1(net5591),
    .A2(net4856));
 sg13g2_nand2_1 _17720_ (.Y(_02473_),
    .A(net2814),
    .B(net4856));
 sg13g2_o21ai_1 _17721_ (.B1(_02473_),
    .Y(_01817_),
    .A1(net5638),
    .A2(net4856));
 sg13g2_nand2_1 _17722_ (.Y(_02474_),
    .A(net2968),
    .B(net4857));
 sg13g2_o21ai_1 _17723_ (.B1(_02474_),
    .Y(_01818_),
    .A1(net5683),
    .A2(net4857));
 sg13g2_nand2_1 _17724_ (.Y(_02475_),
    .A(net2884),
    .B(net4857));
 sg13g2_o21ai_1 _17725_ (.B1(_02475_),
    .Y(_01819_),
    .A1(net5728),
    .A2(net4857));
 sg13g2_nand2_1 _17726_ (.Y(_02476_),
    .A(net2869),
    .B(net4856));
 sg13g2_o21ai_1 _17727_ (.B1(_02476_),
    .Y(_01820_),
    .A1(net5775),
    .A2(net4856));
 sg13g2_nand2_1 _17728_ (.Y(_02477_),
    .A(net5238),
    .B(net5199));
 sg13g2_nand2_1 _17729_ (.Y(_02478_),
    .A(net2711),
    .B(net4855));
 sg13g2_o21ai_1 _17730_ (.B1(_02478_),
    .Y(_01821_),
    .A1(net5457),
    .A2(net4855));
 sg13g2_nand2_1 _17731_ (.Y(_02479_),
    .A(net2478),
    .B(net4854));
 sg13g2_o21ai_1 _17732_ (.B1(_02479_),
    .Y(_01822_),
    .A1(net5505),
    .A2(net4854));
 sg13g2_nand2_1 _17733_ (.Y(_02480_),
    .A(net2402),
    .B(net4854));
 sg13g2_o21ai_1 _17734_ (.B1(_02480_),
    .Y(_01823_),
    .A1(net5548),
    .A2(net4854));
 sg13g2_nand2_1 _17735_ (.Y(_02481_),
    .A(net2374),
    .B(net4854));
 sg13g2_o21ai_1 _17736_ (.B1(_02481_),
    .Y(_01824_),
    .A1(net5591),
    .A2(net4854));
 sg13g2_nand2_1 _17737_ (.Y(_02482_),
    .A(net2213),
    .B(net4854));
 sg13g2_o21ai_1 _17738_ (.B1(_02482_),
    .Y(_01825_),
    .A1(net5638),
    .A2(net4854));
 sg13g2_nand2_1 _17739_ (.Y(_02483_),
    .A(net3159),
    .B(net4855));
 sg13g2_o21ai_1 _17740_ (.B1(_02483_),
    .Y(_01826_),
    .A1(net5683),
    .A2(net4855));
 sg13g2_nand2_1 _17741_ (.Y(_02484_),
    .A(net2352),
    .B(net4855));
 sg13g2_o21ai_1 _17742_ (.B1(_02484_),
    .Y(_01827_),
    .A1(net5728),
    .A2(net4855));
 sg13g2_nand2_1 _17743_ (.Y(_02485_),
    .A(net3026),
    .B(_02477_));
 sg13g2_o21ai_1 _17744_ (.B1(_02485_),
    .Y(_01828_),
    .A1(net5775),
    .A2(net4855));
 sg13g2_nand2_1 _17745_ (.Y(_02486_),
    .A(net5244),
    .B(net5199));
 sg13g2_nand2_1 _17746_ (.Y(_02487_),
    .A(net2959),
    .B(net4853));
 sg13g2_o21ai_1 _17747_ (.B1(_02487_),
    .Y(_01829_),
    .A1(net5464),
    .A2(net4853));
 sg13g2_nand2_1 _17748_ (.Y(_02488_),
    .A(net2589),
    .B(net4852));
 sg13g2_o21ai_1 _17749_ (.B1(_02488_),
    .Y(_01830_),
    .A1(net5503),
    .A2(net4852));
 sg13g2_nand2_1 _17750_ (.Y(_02489_),
    .A(net2889),
    .B(net4852));
 sg13g2_o21ai_1 _17751_ (.B1(_02489_),
    .Y(_01831_),
    .A1(net5546),
    .A2(net4852));
 sg13g2_nand2_1 _17752_ (.Y(_02490_),
    .A(net2808),
    .B(net4853));
 sg13g2_o21ai_1 _17753_ (.B1(_02490_),
    .Y(_01832_),
    .A1(net5589),
    .A2(net4853));
 sg13g2_nand2_1 _17754_ (.Y(_02491_),
    .A(net3194),
    .B(net4853));
 sg13g2_o21ai_1 _17755_ (.B1(_02491_),
    .Y(_01833_),
    .A1(net5643),
    .A2(net4853));
 sg13g2_nand2_1 _17756_ (.Y(_02492_),
    .A(net2428),
    .B(net4852));
 sg13g2_o21ai_1 _17757_ (.B1(_02492_),
    .Y(_01834_),
    .A1(net5684),
    .A2(net4852));
 sg13g2_nand2_1 _17758_ (.Y(_02493_),
    .A(net2596),
    .B(net4853));
 sg13g2_o21ai_1 _17759_ (.B1(_02493_),
    .Y(_01835_),
    .A1(net5730),
    .A2(net4853));
 sg13g2_nand2_1 _17760_ (.Y(_02494_),
    .A(net2327),
    .B(net4852));
 sg13g2_o21ai_1 _17761_ (.B1(_02494_),
    .Y(_01836_),
    .A1(net5772),
    .A2(net4852));
 sg13g2_nand2_1 _17762_ (.Y(_02495_),
    .A(net5239),
    .B(net5199));
 sg13g2_nand2_1 _17763_ (.Y(_02496_),
    .A(net3131),
    .B(net4851));
 sg13g2_o21ai_1 _17764_ (.B1(_02496_),
    .Y(_01837_),
    .A1(net5459),
    .A2(net4851));
 sg13g2_nand2_1 _17765_ (.Y(_02497_),
    .A(net2781),
    .B(net4850));
 sg13g2_o21ai_1 _17766_ (.B1(_02497_),
    .Y(_01838_),
    .A1(net5503),
    .A2(net4850));
 sg13g2_nand2_1 _17767_ (.Y(_02498_),
    .A(net2476),
    .B(net4850));
 sg13g2_o21ai_1 _17768_ (.B1(_02498_),
    .Y(_01839_),
    .A1(net5545),
    .A2(net4850));
 sg13g2_nand2_1 _17769_ (.Y(_02499_),
    .A(net3284),
    .B(net4851));
 sg13g2_o21ai_1 _17770_ (.B1(_02499_),
    .Y(_01840_),
    .A1(net5602),
    .A2(net4851));
 sg13g2_nand2_1 _17771_ (.Y(_02500_),
    .A(net3134),
    .B(net4851));
 sg13g2_o21ai_1 _17772_ (.B1(_02500_),
    .Y(_01841_),
    .A1(net5640),
    .A2(net4851));
 sg13g2_nand2_1 _17773_ (.Y(_02501_),
    .A(net2441),
    .B(net4850));
 sg13g2_o21ai_1 _17774_ (.B1(_02501_),
    .Y(_01842_),
    .A1(net5684),
    .A2(net4850));
 sg13g2_nand2_1 _17775_ (.Y(_02502_),
    .A(net2842),
    .B(net4851));
 sg13g2_o21ai_1 _17776_ (.B1(_02502_),
    .Y(_01843_),
    .A1(net5733),
    .A2(net4851));
 sg13g2_nand2_1 _17777_ (.Y(_02503_),
    .A(net2268),
    .B(net4850));
 sg13g2_o21ai_1 _17778_ (.B1(_02503_),
    .Y(_01844_),
    .A1(net5772),
    .A2(net4850));
 sg13g2_nand2_1 _17779_ (.Y(_02504_),
    .A(net5242),
    .B(net5199));
 sg13g2_nand2_1 _17780_ (.Y(_02505_),
    .A(net2769),
    .B(net4848));
 sg13g2_o21ai_1 _17781_ (.B1(_02505_),
    .Y(_01845_),
    .A1(net5459),
    .A2(net4848));
 sg13g2_nand2_1 _17782_ (.Y(_02506_),
    .A(net3030),
    .B(net4849));
 sg13g2_o21ai_1 _17783_ (.B1(_02506_),
    .Y(_01846_),
    .A1(net5503),
    .A2(net4849));
 sg13g2_nand2_1 _17784_ (.Y(_02507_),
    .A(net3217),
    .B(net4849));
 sg13g2_o21ai_1 _17785_ (.B1(_02507_),
    .Y(_01847_),
    .A1(net5545),
    .A2(_02504_));
 sg13g2_nand2_1 _17786_ (.Y(_02508_),
    .A(net3047),
    .B(net4848));
 sg13g2_o21ai_1 _17787_ (.B1(_02508_),
    .Y(_01848_),
    .A1(net5589),
    .A2(net4848));
 sg13g2_nand2_1 _17788_ (.Y(_02509_),
    .A(net2754),
    .B(net4848));
 sg13g2_o21ai_1 _17789_ (.B1(_02509_),
    .Y(_01849_),
    .A1(net5640),
    .A2(net4848));
 sg13g2_nand2_1 _17790_ (.Y(_02510_),
    .A(net3118),
    .B(net4849));
 sg13g2_o21ai_1 _17791_ (.B1(_02510_),
    .Y(_01850_),
    .A1(net5684),
    .A2(net4849));
 sg13g2_nand2_1 _17792_ (.Y(_02511_),
    .A(net2439),
    .B(net4848));
 sg13g2_o21ai_1 _17793_ (.B1(_02511_),
    .Y(_01851_),
    .A1(net5733),
    .A2(net4848));
 sg13g2_nand2_1 _17794_ (.Y(_02512_),
    .A(net3277),
    .B(net4849));
 sg13g2_o21ai_1 _17795_ (.B1(_02512_),
    .Y(_01852_),
    .A1(net5775),
    .A2(net4849));
 sg13g2_nor2_1 _17796_ (.A(_03201_),
    .B(net5210),
    .Y(_02513_));
 sg13g2_nor2_1 _17797_ (.A(net4051),
    .B(net4847),
    .Y(_02514_));
 sg13g2_a21oi_1 _17798_ (.A1(net5452),
    .A2(net4847),
    .Y(_01853_),
    .B1(_02514_));
 sg13g2_nor2_1 _17799_ (.A(net3431),
    .B(net4847),
    .Y(_02515_));
 sg13g2_a21oi_1 _17800_ (.A1(net5497),
    .A2(net4847),
    .Y(_01854_),
    .B1(_02515_));
 sg13g2_nor2_1 _17801_ (.A(net3550),
    .B(net4846),
    .Y(_02516_));
 sg13g2_a21oi_1 _17802_ (.A1(net5552),
    .A2(net4846),
    .Y(_01855_),
    .B1(_02516_));
 sg13g2_nor2_1 _17803_ (.A(net4008),
    .B(net4847),
    .Y(_02517_));
 sg13g2_a21oi_1 _17804_ (.A1(net5595),
    .A2(net4846),
    .Y(_01856_),
    .B1(_02517_));
 sg13g2_nor2_1 _17805_ (.A(net3654),
    .B(net4846),
    .Y(_02518_));
 sg13g2_a21oi_1 _17806_ (.A1(net5642),
    .A2(_02513_),
    .Y(_01857_),
    .B1(_02518_));
 sg13g2_nor2_1 _17807_ (.A(net3728),
    .B(net4846),
    .Y(_02519_));
 sg13g2_a21oi_1 _17808_ (.A1(net5687),
    .A2(net4846),
    .Y(_01858_),
    .B1(_02519_));
 sg13g2_nor2_1 _17809_ (.A(net3378),
    .B(net4847),
    .Y(_02520_));
 sg13g2_a21oi_1 _17810_ (.A1(net5732),
    .A2(net4847),
    .Y(_01859_),
    .B1(_02520_));
 sg13g2_nor2_1 _17811_ (.A(net4054),
    .B(net4846),
    .Y(_02521_));
 sg13g2_a21oi_1 _17812_ (.A1(net5783),
    .A2(net4846),
    .Y(_01860_),
    .B1(_02521_));
 sg13g2_nand2_1 _17813_ (.Y(_02522_),
    .A(net5245),
    .B(net5198));
 sg13g2_nand2_1 _17814_ (.Y(_02523_),
    .A(net2444),
    .B(net4845));
 sg13g2_o21ai_1 _17815_ (.B1(_02523_),
    .Y(_01861_),
    .A1(net5460),
    .A2(net4845));
 sg13g2_nand2_1 _17816_ (.Y(_02524_),
    .A(net2206),
    .B(net4844));
 sg13g2_o21ai_1 _17817_ (.B1(_02524_),
    .Y(_01862_),
    .A1(net5502),
    .A2(net4844));
 sg13g2_nand2_1 _17818_ (.Y(_02525_),
    .A(net3304),
    .B(net4844));
 sg13g2_o21ai_1 _17819_ (.B1(_02525_),
    .Y(_01863_),
    .A1(net5548),
    .A2(net4844));
 sg13g2_nand2_1 _17820_ (.Y(_02526_),
    .A(net2563),
    .B(_02522_));
 sg13g2_o21ai_1 _17821_ (.B1(_02526_),
    .Y(_01864_),
    .A1(net5600),
    .A2(net4845));
 sg13g2_nand2_1 _17822_ (.Y(_02527_),
    .A(net2508),
    .B(net4845));
 sg13g2_o21ai_1 _17823_ (.B1(_02527_),
    .Y(_01865_),
    .A1(net5644),
    .A2(net4845));
 sg13g2_nand2_1 _17824_ (.Y(_02528_),
    .A(net2132),
    .B(net4845));
 sg13g2_o21ai_1 _17825_ (.B1(_02528_),
    .Y(_01866_),
    .A1(net5684),
    .A2(net4845));
 sg13g2_nand2_1 _17826_ (.Y(_02529_),
    .A(net2837),
    .B(net4844));
 sg13g2_o21ai_1 _17827_ (.B1(_02529_),
    .Y(_01867_),
    .A1(net5733),
    .A2(net4844));
 sg13g2_nand2_1 _17828_ (.Y(_02530_),
    .A(net2315),
    .B(net4844));
 sg13g2_o21ai_1 _17829_ (.B1(_02530_),
    .Y(_01868_),
    .A1(net5779),
    .A2(net4844));
 sg13g2_nand2_1 _17830_ (.Y(_02531_),
    .A(net5251),
    .B(net5198));
 sg13g2_nand2_1 _17831_ (.Y(_02532_),
    .A(net2409),
    .B(net4843));
 sg13g2_o21ai_1 _17832_ (.B1(_02532_),
    .Y(_01869_),
    .A1(net5460),
    .A2(net4843));
 sg13g2_nand2_1 _17833_ (.Y(_02533_),
    .A(net3437),
    .B(net4842));
 sg13g2_o21ai_1 _17834_ (.B1(_02533_),
    .Y(_01870_),
    .A1(net5502),
    .A2(net4842));
 sg13g2_nand2_1 _17835_ (.Y(_02534_),
    .A(net2329),
    .B(net4842));
 sg13g2_o21ai_1 _17836_ (.B1(_02534_),
    .Y(_01871_),
    .A1(net5545),
    .A2(net4842));
 sg13g2_nand2_1 _17837_ (.Y(_02535_),
    .A(net2310),
    .B(net4842));
 sg13g2_o21ai_1 _17838_ (.B1(_02535_),
    .Y(_01872_),
    .A1(net5600),
    .A2(net4842));
 sg13g2_nand2_1 _17839_ (.Y(_02536_),
    .A(net2393),
    .B(net4842));
 sg13g2_o21ai_1 _17840_ (.B1(_02536_),
    .Y(_01873_),
    .A1(net5644),
    .A2(net4842));
 sg13g2_nand2_1 _17841_ (.Y(_02537_),
    .A(net2483),
    .B(net4843));
 sg13g2_o21ai_1 _17842_ (.B1(_02537_),
    .Y(_01874_),
    .A1(net5684),
    .A2(_02531_));
 sg13g2_nand2_1 _17843_ (.Y(_02538_),
    .A(net2679),
    .B(net4843));
 sg13g2_o21ai_1 _17844_ (.B1(_02538_),
    .Y(_01875_),
    .A1(net5733),
    .A2(net4843));
 sg13g2_nand2_1 _17845_ (.Y(_02539_),
    .A(net2304),
    .B(net4843));
 sg13g2_o21ai_1 _17846_ (.B1(_02539_),
    .Y(_01876_),
    .A1(net5775),
    .A2(net4843));
 sg13g2_nand2_1 _17847_ (.Y(_02540_),
    .A(net5246),
    .B(net5198));
 sg13g2_nand2_1 _17848_ (.Y(_02541_),
    .A(net3133),
    .B(net4841));
 sg13g2_o21ai_1 _17849_ (.B1(_02541_),
    .Y(_01877_),
    .A1(net5461),
    .A2(_02540_));
 sg13g2_nand2_1 _17850_ (.Y(_02542_),
    .A(net2156),
    .B(net4840));
 sg13g2_o21ai_1 _17851_ (.B1(_02542_),
    .Y(_01878_),
    .A1(net5510),
    .A2(net4840));
 sg13g2_nand2_1 _17852_ (.Y(_02543_),
    .A(net2691),
    .B(net4841));
 sg13g2_o21ai_1 _17853_ (.B1(_02543_),
    .Y(_01879_),
    .A1(net5553),
    .A2(net4840));
 sg13g2_nand2_1 _17854_ (.Y(_02544_),
    .A(net2664),
    .B(net4840));
 sg13g2_o21ai_1 _17855_ (.B1(_02544_),
    .Y(_01880_),
    .A1(net5600),
    .A2(net4840));
 sg13g2_nand2_1 _17856_ (.Y(_02545_),
    .A(net2290),
    .B(net4840));
 sg13g2_o21ai_1 _17857_ (.B1(_02545_),
    .Y(_01881_),
    .A1(net5644),
    .A2(net4840));
 sg13g2_nand2_1 _17858_ (.Y(_02546_),
    .A(net2510),
    .B(net4841));
 sg13g2_o21ai_1 _17859_ (.B1(_02546_),
    .Y(_01882_),
    .A1(net5688),
    .A2(net4841));
 sg13g2_nand2_1 _17860_ (.Y(_02547_),
    .A(net2811),
    .B(net4841));
 sg13g2_o21ai_1 _17861_ (.B1(_02547_),
    .Y(_01883_),
    .A1(net5733),
    .A2(net4840));
 sg13g2_nand2_1 _17862_ (.Y(_02548_),
    .A(net2481),
    .B(net4841));
 sg13g2_o21ai_1 _17863_ (.B1(_02548_),
    .Y(_01884_),
    .A1(net5779),
    .A2(net4841));
 sg13g2_nor3_2 _17864_ (.A(_02940_),
    .B(net5229),
    .C(net5240),
    .Y(_02549_));
 sg13g2_nor2_1 _17865_ (.A(net3564),
    .B(_02549_),
    .Y(_02550_));
 sg13g2_a21oi_1 _17866_ (.A1(net5460),
    .A2(net5171),
    .Y(_01885_),
    .B1(_02550_));
 sg13g2_nor2_1 _17867_ (.A(net3922),
    .B(net5171),
    .Y(_02551_));
 sg13g2_a21oi_1 _17868_ (.A1(net5510),
    .A2(net5171),
    .Y(_01886_),
    .B1(_02551_));
 sg13g2_nor2_1 _17869_ (.A(net4103),
    .B(net5171),
    .Y(_02552_));
 sg13g2_a21oi_1 _17870_ (.A1(net5553),
    .A2(net5171),
    .Y(_01887_),
    .B1(_02552_));
 sg13g2_nor2_1 _17871_ (.A(net3791),
    .B(net5170),
    .Y(_02553_));
 sg13g2_a21oi_1 _17872_ (.A1(net5600),
    .A2(net5170),
    .Y(_01888_),
    .B1(_02553_));
 sg13g2_nor2_1 _17873_ (.A(net3876),
    .B(net5171),
    .Y(_02554_));
 sg13g2_a21oi_1 _17874_ (.A1(net5644),
    .A2(net5171),
    .Y(_01889_),
    .B1(_02554_));
 sg13g2_nor2_1 _17875_ (.A(net3553),
    .B(net5170),
    .Y(_02555_));
 sg13g2_a21oi_1 _17876_ (.A1(net5688),
    .A2(net5170),
    .Y(_01890_),
    .B1(_02555_));
 sg13g2_nor2_1 _17877_ (.A(net3828),
    .B(net5170),
    .Y(_02556_));
 sg13g2_a21oi_1 _17878_ (.A1(net5733),
    .A2(net5170),
    .Y(_01891_),
    .B1(_02556_));
 sg13g2_nor2_1 _17879_ (.A(net3694),
    .B(net5170),
    .Y(_02557_));
 sg13g2_a21oi_1 _17880_ (.A1(net5779),
    .A2(net5170),
    .Y(_01892_),
    .B1(_02557_));
 sg13g2_nand2_1 _17881_ (.Y(_02558_),
    .A(net5249),
    .B(net5203));
 sg13g2_nand2_1 _17882_ (.Y(_02559_),
    .A(net2706),
    .B(net4839));
 sg13g2_o21ai_1 _17883_ (.B1(_02559_),
    .Y(_01893_),
    .A1(net5456),
    .A2(net4839));
 sg13g2_nand2_1 _17884_ (.Y(_02560_),
    .A(net2932),
    .B(net4839));
 sg13g2_o21ai_1 _17885_ (.B1(_02560_),
    .Y(_01894_),
    .A1(net5501),
    .A2(net4839));
 sg13g2_nand2_1 _17886_ (.Y(_02561_),
    .A(net3127),
    .B(net4839));
 sg13g2_o21ai_1 _17887_ (.B1(_02561_),
    .Y(_01895_),
    .A1(net5544),
    .A2(net4839));
 sg13g2_nand2_1 _17888_ (.Y(_02562_),
    .A(net2155),
    .B(net4839));
 sg13g2_o21ai_1 _17889_ (.B1(_02562_),
    .Y(_01896_),
    .A1(net5591),
    .A2(_02558_));
 sg13g2_nand2_1 _17890_ (.Y(_02563_),
    .A(net3130),
    .B(net4838));
 sg13g2_o21ai_1 _17891_ (.B1(_02563_),
    .Y(_01897_),
    .A1(net5636),
    .A2(net4838));
 sg13g2_nand2_1 _17892_ (.Y(_02564_),
    .A(net2379),
    .B(net4838));
 sg13g2_o21ai_1 _17893_ (.B1(_02564_),
    .Y(_01898_),
    .A1(net5681),
    .A2(net4838));
 sg13g2_nand2_1 _17894_ (.Y(_02565_),
    .A(net2250),
    .B(net4838));
 sg13g2_o21ai_1 _17895_ (.B1(_02565_),
    .Y(_01899_),
    .A1(net5727),
    .A2(net4838));
 sg13g2_nand2_1 _17896_ (.Y(_02566_),
    .A(net2598),
    .B(net4838));
 sg13g2_o21ai_1 _17897_ (.B1(_02566_),
    .Y(_01900_),
    .A1(net5773),
    .A2(net4838));
 sg13g2_nand2_1 _17898_ (.Y(_02567_),
    .A(_03139_),
    .B(net5203));
 sg13g2_nand2_1 _17899_ (.Y(_02568_),
    .A(net2306),
    .B(net4837));
 sg13g2_o21ai_1 _17900_ (.B1(_02568_),
    .Y(_01901_),
    .A1(net5456),
    .A2(net4837));
 sg13g2_nand2_1 _17901_ (.Y(_02569_),
    .A(net2356),
    .B(net4837));
 sg13g2_o21ai_1 _17902_ (.B1(_02569_),
    .Y(_01902_),
    .A1(net5501),
    .A2(net4837));
 sg13g2_nand2_1 _17903_ (.Y(_02570_),
    .A(net2432),
    .B(_02567_));
 sg13g2_o21ai_1 _17904_ (.B1(_02570_),
    .Y(_01903_),
    .A1(net5545),
    .A2(net4837));
 sg13g2_nand2_1 _17905_ (.Y(_02571_),
    .A(net3078),
    .B(net4837));
 sg13g2_o21ai_1 _17906_ (.B1(_02571_),
    .Y(_01904_),
    .A1(net5591),
    .A2(net4837));
 sg13g2_nand2_1 _17907_ (.Y(_02572_),
    .A(net2658),
    .B(net4836));
 sg13g2_o21ai_1 _17908_ (.B1(_02572_),
    .Y(_01905_),
    .A1(net5636),
    .A2(net4836));
 sg13g2_nand2_1 _17909_ (.Y(_02573_),
    .A(net2347),
    .B(net4836));
 sg13g2_o21ai_1 _17910_ (.B1(_02573_),
    .Y(_01906_),
    .A1(net5681),
    .A2(net4836));
 sg13g2_nand2_1 _17911_ (.Y(_02574_),
    .A(net2880),
    .B(net4836));
 sg13g2_o21ai_1 _17912_ (.B1(_02574_),
    .Y(_01907_),
    .A1(net5727),
    .A2(net4836));
 sg13g2_nand2_1 _17913_ (.Y(_02575_),
    .A(net3003),
    .B(net4836));
 sg13g2_o21ai_1 _17914_ (.B1(_02575_),
    .Y(_01908_),
    .A1(net5773),
    .A2(net4836));
 sg13g2_nand2_1 _17915_ (.Y(_02576_),
    .A(_03079_),
    .B(net5203));
 sg13g2_nand2_1 _17916_ (.Y(_02577_),
    .A(net2501),
    .B(net4835));
 sg13g2_o21ai_1 _17917_ (.B1(_02577_),
    .Y(_01909_),
    .A1(net5456),
    .A2(net4835));
 sg13g2_nand2_1 _17918_ (.Y(_02578_),
    .A(net2578),
    .B(net4835));
 sg13g2_o21ai_1 _17919_ (.B1(_02578_),
    .Y(_01910_),
    .A1(net5501),
    .A2(net4835));
 sg13g2_nand2_1 _17920_ (.Y(_02579_),
    .A(net3374),
    .B(net4835));
 sg13g2_o21ai_1 _17921_ (.B1(_02579_),
    .Y(_01911_),
    .A1(net5544),
    .A2(net4835));
 sg13g2_nand2_1 _17922_ (.Y(_02580_),
    .A(net2137),
    .B(_02576_));
 sg13g2_o21ai_1 _17923_ (.B1(_02580_),
    .Y(_01912_),
    .A1(net5593),
    .A2(net4835));
 sg13g2_nand2_1 _17924_ (.Y(_02581_),
    .A(net3153),
    .B(net4834));
 sg13g2_o21ai_1 _17925_ (.B1(_02581_),
    .Y(_01913_),
    .A1(net5636),
    .A2(net4834));
 sg13g2_nand2_1 _17926_ (.Y(_02582_),
    .A(net3308),
    .B(net4834));
 sg13g2_o21ai_1 _17927_ (.B1(_02582_),
    .Y(_01914_),
    .A1(net5681),
    .A2(net4834));
 sg13g2_nand2_1 _17928_ (.Y(_02583_),
    .A(net3103),
    .B(net4834));
 sg13g2_o21ai_1 _17929_ (.B1(_02583_),
    .Y(_01915_),
    .A1(net5727),
    .A2(net4834));
 sg13g2_nand2_1 _17930_ (.Y(_02584_),
    .A(net2258),
    .B(net4834));
 sg13g2_o21ai_1 _17931_ (.B1(_02584_),
    .Y(_01916_),
    .A1(net5773),
    .A2(net4834));
 sg13g2_nand2_1 _17932_ (.Y(_02585_),
    .A(net5253),
    .B(net5203));
 sg13g2_nand2_1 _17933_ (.Y(_02586_),
    .A(net2830),
    .B(net4832));
 sg13g2_o21ai_1 _17934_ (.B1(_02586_),
    .Y(_01917_),
    .A1(net5456),
    .A2(net4832));
 sg13g2_nand2_1 _17935_ (.Y(_02587_),
    .A(net2453),
    .B(net4833));
 sg13g2_o21ai_1 _17936_ (.B1(_02587_),
    .Y(_01918_),
    .A1(net5501),
    .A2(net4833));
 sg13g2_nand2_1 _17937_ (.Y(_02588_),
    .A(net3292),
    .B(net4833));
 sg13g2_o21ai_1 _17938_ (.B1(_02588_),
    .Y(_01919_),
    .A1(net5550),
    .A2(net4833));
 sg13g2_nand2_1 _17939_ (.Y(_02589_),
    .A(net2807),
    .B(net4833));
 sg13g2_o21ai_1 _17940_ (.B1(_02589_),
    .Y(_01920_),
    .A1(net5593),
    .A2(net4833));
 sg13g2_nand2_1 _17941_ (.Y(_02590_),
    .A(net2630),
    .B(net4833));
 sg13g2_o21ai_1 _17942_ (.B1(_02590_),
    .Y(_01921_),
    .A1(net5636),
    .A2(net4833));
 sg13g2_nand2_1 _17943_ (.Y(_02591_),
    .A(net2704),
    .B(net4832));
 sg13g2_o21ai_1 _17944_ (.B1(_02591_),
    .Y(_01922_),
    .A1(net5681),
    .A2(net4832));
 sg13g2_nand2_1 _17945_ (.Y(_02592_),
    .A(net2853),
    .B(net4832));
 sg13g2_o21ai_1 _17946_ (.B1(_02592_),
    .Y(_01923_),
    .A1(net5727),
    .A2(net4832));
 sg13g2_nand2_1 _17947_ (.Y(_02593_),
    .A(net2799),
    .B(net4832));
 sg13g2_o21ai_1 _17948_ (.B1(_02593_),
    .Y(_01924_),
    .A1(net5773),
    .A2(net4832));
 sg13g2_nand2_2 _17949_ (.Y(_02594_),
    .A(net5235),
    .B(net5203));
 sg13g2_nand2_1 _17950_ (.Y(_02595_),
    .A(net2360),
    .B(net4831));
 sg13g2_o21ai_1 _17951_ (.B1(_02595_),
    .Y(_01925_),
    .A1(net5457),
    .A2(net4831));
 sg13g2_nand2_1 _17952_ (.Y(_02596_),
    .A(net2826),
    .B(net4831));
 sg13g2_o21ai_1 _17953_ (.B1(_02596_),
    .Y(_01926_),
    .A1(net5504),
    .A2(net4831));
 sg13g2_nand2_1 _17954_ (.Y(_02597_),
    .A(net2505),
    .B(net4831));
 sg13g2_o21ai_1 _17955_ (.B1(_02597_),
    .Y(_01927_),
    .A1(net5548),
    .A2(net4831));
 sg13g2_nand2_1 _17956_ (.Y(_02598_),
    .A(net2177),
    .B(net4831));
 sg13g2_o21ai_1 _17957_ (.B1(_02598_),
    .Y(_01928_),
    .A1(net5593),
    .A2(net4831));
 sg13g2_nand2_1 _17958_ (.Y(_02599_),
    .A(net2587),
    .B(net4830));
 sg13g2_o21ai_1 _17959_ (.B1(_02599_),
    .Y(_01929_),
    .A1(net5636),
    .A2(net4830));
 sg13g2_nand2_1 _17960_ (.Y(_02600_),
    .A(net2276),
    .B(net4830));
 sg13g2_o21ai_1 _17961_ (.B1(_02600_),
    .Y(_01930_),
    .A1(net5682),
    .A2(net4830));
 sg13g2_nand2_1 _17962_ (.Y(_02601_),
    .A(net2179),
    .B(net4830));
 sg13g2_o21ai_1 _17963_ (.B1(_02601_),
    .Y(_01931_),
    .A1(net5726),
    .A2(net4830));
 sg13g2_nand2_1 _17964_ (.Y(_02602_),
    .A(net2931),
    .B(net4830));
 sg13g2_o21ai_1 _17965_ (.B1(_02602_),
    .Y(_01932_),
    .A1(net5773),
    .A2(net4830));
 sg13g2_nor2_1 _17966_ (.A(_03067_),
    .B(net5210),
    .Y(_02603_));
 sg13g2_nor2_1 _17967_ (.A(net4035),
    .B(net4828),
    .Y(_02604_));
 sg13g2_a21oi_1 _17968_ (.A1(net5452),
    .A2(net4828),
    .Y(_01933_),
    .B1(_02604_));
 sg13g2_nor2_1 _17969_ (.A(net2794),
    .B(net4828),
    .Y(_02605_));
 sg13g2_a21oi_1 _17970_ (.A1(net5497),
    .A2(net4828),
    .Y(_01934_),
    .B1(_02605_));
 sg13g2_nor2_1 _17971_ (.A(net3612),
    .B(net4828),
    .Y(_02606_));
 sg13g2_a21oi_1 _17972_ (.A1(net5541),
    .A2(net4828),
    .Y(_01935_),
    .B1(_02606_));
 sg13g2_nor2_1 _17973_ (.A(net3723),
    .B(net4829),
    .Y(_02607_));
 sg13g2_a21oi_1 _17974_ (.A1(net5596),
    .A2(net4829),
    .Y(_01936_),
    .B1(_02607_));
 sg13g2_nor2_1 _17975_ (.A(net3575),
    .B(net4829),
    .Y(_02608_));
 sg13g2_a21oi_1 _17976_ (.A1(net5642),
    .A2(net4829),
    .Y(_01937_),
    .B1(_02608_));
 sg13g2_nor2_1 _17977_ (.A(net3227),
    .B(net4829),
    .Y(_02609_));
 sg13g2_a21oi_1 _17978_ (.A1(net5687),
    .A2(net4829),
    .Y(_01938_),
    .B1(_02609_));
 sg13g2_nor2_1 _17979_ (.A(net2871),
    .B(net4829),
    .Y(_02610_));
 sg13g2_a21oi_1 _17980_ (.A1(net5732),
    .A2(net4829),
    .Y(_01939_),
    .B1(_02610_));
 sg13g2_nor2_1 _17981_ (.A(net3772),
    .B(net4828),
    .Y(_02611_));
 sg13g2_a21oi_1 _17982_ (.A1(net5767),
    .A2(net4828),
    .Y(_01940_),
    .B1(_02611_));
 sg13g2_nand2_1 _17983_ (.Y(_02612_),
    .A(net5236),
    .B(net5203));
 sg13g2_nand2_1 _17984_ (.Y(_02613_),
    .A(net2802),
    .B(net4827));
 sg13g2_o21ai_1 _17985_ (.B1(_02613_),
    .Y(_01941_),
    .A1(net5457),
    .A2(net4827));
 sg13g2_nand2_1 _17986_ (.Y(_02614_),
    .A(net3524),
    .B(net4826));
 sg13g2_o21ai_1 _17987_ (.B1(_02614_),
    .Y(_01942_),
    .A1(net5504),
    .A2(net4826));
 sg13g2_nand2_1 _17988_ (.Y(_02615_),
    .A(net3209),
    .B(_02612_));
 sg13g2_o21ai_1 _17989_ (.B1(_02615_),
    .Y(_01943_),
    .A1(net5548),
    .A2(net4827));
 sg13g2_nand2_1 _17990_ (.Y(_02616_),
    .A(net2897),
    .B(net4827));
 sg13g2_o21ai_1 _17991_ (.B1(_02616_),
    .Y(_01944_),
    .A1(net5591),
    .A2(net4827));
 sg13g2_nand2_1 _17992_ (.Y(_02617_),
    .A(net2753),
    .B(net4826));
 sg13g2_o21ai_1 _17993_ (.B1(_02617_),
    .Y(_01945_),
    .A1(net5636),
    .A2(net4826));
 sg13g2_nand2_1 _17994_ (.Y(_02618_),
    .A(net2568),
    .B(net4826));
 sg13g2_o21ai_1 _17995_ (.B1(_02618_),
    .Y(_01946_),
    .A1(net5682),
    .A2(net4826));
 sg13g2_nand2_1 _17996_ (.Y(_02619_),
    .A(net2433),
    .B(net4826));
 sg13g2_o21ai_1 _17997_ (.B1(_02619_),
    .Y(_01947_),
    .A1(net5726),
    .A2(net4826));
 sg13g2_nand2_1 _17998_ (.Y(_02620_),
    .A(net2398),
    .B(net4827));
 sg13g2_o21ai_1 _17999_ (.B1(_02620_),
    .Y(_01948_),
    .A1(net5774),
    .A2(net4827));
 sg13g2_nand2_2 _18000_ (.Y(_02621_),
    .A(net5238),
    .B(net5202));
 sg13g2_nand2_1 _18001_ (.Y(_02622_),
    .A(net2196),
    .B(net4825));
 sg13g2_o21ai_1 _18002_ (.B1(_02622_),
    .Y(_01949_),
    .A1(net5457),
    .A2(net4825));
 sg13g2_nand2_1 _18003_ (.Y(_02623_),
    .A(net3151),
    .B(net4825));
 sg13g2_o21ai_1 _18004_ (.B1(_02623_),
    .Y(_01950_),
    .A1(net5504),
    .A2(net4825));
 sg13g2_nand2_1 _18005_ (.Y(_02624_),
    .A(net2987),
    .B(net4825));
 sg13g2_o21ai_1 _18006_ (.B1(_02624_),
    .Y(_01951_),
    .A1(net5548),
    .A2(net4825));
 sg13g2_nand2_1 _18007_ (.Y(_02625_),
    .A(net2202),
    .B(net4825));
 sg13g2_o21ai_1 _18008_ (.B1(_02625_),
    .Y(_01952_),
    .A1(net5591),
    .A2(net4825));
 sg13g2_nand2_1 _18009_ (.Y(_02626_),
    .A(net2434),
    .B(net4824));
 sg13g2_o21ai_1 _18010_ (.B1(_02626_),
    .Y(_01953_),
    .A1(net5637),
    .A2(net4824));
 sg13g2_nand2_1 _18011_ (.Y(_02627_),
    .A(net2833),
    .B(net4824));
 sg13g2_o21ai_1 _18012_ (.B1(_02627_),
    .Y(_01954_),
    .A1(net5682),
    .A2(net4824));
 sg13g2_nand2_1 _18013_ (.Y(_02628_),
    .A(net2392),
    .B(net4824));
 sg13g2_o21ai_1 _18014_ (.B1(_02628_),
    .Y(_01955_),
    .A1(net5726),
    .A2(net4824));
 sg13g2_nand2_1 _18015_ (.Y(_02629_),
    .A(net2528),
    .B(net4824));
 sg13g2_o21ai_1 _18016_ (.B1(_02629_),
    .Y(_01956_),
    .A1(net5774),
    .A2(net4824));
 sg13g2_nand2_1 _18017_ (.Y(_02630_),
    .A(net5244),
    .B(net5202));
 sg13g2_nand2_1 _18018_ (.Y(_02631_),
    .A(net2281),
    .B(net4821));
 sg13g2_o21ai_1 _18019_ (.B1(_02631_),
    .Y(_01957_),
    .A1(net5456),
    .A2(net4822));
 sg13g2_nand2_1 _18020_ (.Y(_02632_),
    .A(net2967),
    .B(net4822));
 sg13g2_o21ai_1 _18021_ (.B1(_02632_),
    .Y(_01958_),
    .A1(net5504),
    .A2(net4822));
 sg13g2_nand2_1 _18022_ (.Y(_02633_),
    .A(net2459),
    .B(net4822));
 sg13g2_o21ai_1 _18023_ (.B1(_02633_),
    .Y(_01959_),
    .A1(net5550),
    .A2(net4821));
 sg13g2_nand2_1 _18024_ (.Y(_02634_),
    .A(net3124),
    .B(net4821));
 sg13g2_o21ai_1 _18025_ (.B1(_02634_),
    .Y(_01960_),
    .A1(net5593),
    .A2(net4821));
 sg13g2_nand2_1 _18026_ (.Y(_02635_),
    .A(net2171),
    .B(net4823));
 sg13g2_o21ai_1 _18027_ (.B1(_02635_),
    .Y(_01961_),
    .A1(net5637),
    .A2(net4823));
 sg13g2_nand2_1 _18028_ (.Y(_02636_),
    .A(net3088),
    .B(net4823));
 sg13g2_o21ai_1 _18029_ (.B1(_02636_),
    .Y(_01962_),
    .A1(net5681),
    .A2(net4823));
 sg13g2_nand2_1 _18030_ (.Y(_02637_),
    .A(net2498),
    .B(net4821));
 sg13g2_o21ai_1 _18031_ (.B1(_02637_),
    .Y(_01963_),
    .A1(net5727),
    .A2(net4821));
 sg13g2_nand2_1 _18032_ (.Y(_02638_),
    .A(net3171),
    .B(net4821));
 sg13g2_o21ai_1 _18033_ (.B1(_02638_),
    .Y(_01964_),
    .A1(net5774),
    .A2(net4821));
 sg13g2_nand2_1 _18034_ (.Y(_02639_),
    .A(net5239),
    .B(net5202));
 sg13g2_nand2_1 _18035_ (.Y(_02640_),
    .A(net2601),
    .B(net4818));
 sg13g2_o21ai_1 _18036_ (.B1(_02640_),
    .Y(_01965_),
    .A1(net5456),
    .A2(net4818));
 sg13g2_nand2_1 _18037_ (.Y(_02641_),
    .A(net2189),
    .B(net4819));
 sg13g2_o21ai_1 _18038_ (.B1(_02641_),
    .Y(_01966_),
    .A1(net5504),
    .A2(net4819));
 sg13g2_nand2_1 _18039_ (.Y(_02642_),
    .A(net2252),
    .B(net4819));
 sg13g2_o21ai_1 _18040_ (.B1(_02642_),
    .Y(_01967_),
    .A1(net5550),
    .A2(net4819));
 sg13g2_nand2_1 _18041_ (.Y(_02643_),
    .A(net2571),
    .B(net4818));
 sg13g2_o21ai_1 _18042_ (.B1(_02643_),
    .Y(_01968_),
    .A1(net5593),
    .A2(net4818));
 sg13g2_nand2_1 _18043_ (.Y(_02644_),
    .A(net3160),
    .B(net4820));
 sg13g2_o21ai_1 _18044_ (.B1(_02644_),
    .Y(_01969_),
    .A1(net5637),
    .A2(net4820));
 sg13g2_nand2_1 _18045_ (.Y(_02645_),
    .A(net2926),
    .B(net4820));
 sg13g2_o21ai_1 _18046_ (.B1(_02645_),
    .Y(_01970_),
    .A1(net5681),
    .A2(net4820));
 sg13g2_nand2_1 _18047_ (.Y(_02646_),
    .A(net2342),
    .B(net4818));
 sg13g2_o21ai_1 _18048_ (.B1(_02646_),
    .Y(_01971_),
    .A1(net5727),
    .A2(net4818));
 sg13g2_nand2_1 _18049_ (.Y(_02647_),
    .A(net2920),
    .B(net4818));
 sg13g2_o21ai_1 _18050_ (.B1(_02647_),
    .Y(_01972_),
    .A1(net5774),
    .A2(net4818));
 sg13g2_nand2_1 _18051_ (.Y(_02648_),
    .A(net5242),
    .B(net5202));
 sg13g2_nand2_1 _18052_ (.Y(_02649_),
    .A(net2971),
    .B(net4816));
 sg13g2_o21ai_1 _18053_ (.B1(_02649_),
    .Y(_01973_),
    .A1(net5456),
    .A2(net4816));
 sg13g2_nand2_1 _18054_ (.Y(_02650_),
    .A(net2218),
    .B(net4816));
 sg13g2_o21ai_1 _18055_ (.B1(_02650_),
    .Y(_01974_),
    .A1(net5504),
    .A2(net4816));
 sg13g2_nand2_1 _18056_ (.Y(_02651_),
    .A(net3347),
    .B(_02648_));
 sg13g2_o21ai_1 _18057_ (.B1(_02651_),
    .Y(_01975_),
    .A1(net5550),
    .A2(net4817));
 sg13g2_nand2_1 _18058_ (.Y(_02652_),
    .A(net2974),
    .B(net4816));
 sg13g2_o21ai_1 _18059_ (.B1(_02652_),
    .Y(_01976_),
    .A1(net5593),
    .A2(net4816));
 sg13g2_nand2_1 _18060_ (.Y(_02653_),
    .A(net2475),
    .B(net4817));
 sg13g2_o21ai_1 _18061_ (.B1(_02653_),
    .Y(_01977_),
    .A1(net5637),
    .A2(net4817));
 sg13g2_nand2_1 _18062_ (.Y(_02654_),
    .A(net3154),
    .B(net4817));
 sg13g2_o21ai_1 _18063_ (.B1(_02654_),
    .Y(_01978_),
    .A1(net5681),
    .A2(net4817));
 sg13g2_nand2_1 _18064_ (.Y(_02655_),
    .A(net2933),
    .B(net4817));
 sg13g2_o21ai_1 _18065_ (.B1(_02655_),
    .Y(_01979_),
    .A1(net5726),
    .A2(net4817));
 sg13g2_nand2_1 _18066_ (.Y(_02656_),
    .A(net2531),
    .B(net4816));
 sg13g2_o21ai_1 _18067_ (.B1(_02656_),
    .Y(_01980_),
    .A1(net5773),
    .A2(net4816));
 sg13g2_nand2_1 _18068_ (.Y(_02657_),
    .A(net5243),
    .B(net5202));
 sg13g2_nand2_1 _18069_ (.Y(_02658_),
    .A(net3065),
    .B(net4814));
 sg13g2_o21ai_1 _18070_ (.B1(_02658_),
    .Y(_01981_),
    .A1(net5456),
    .A2(net4814));
 sg13g2_nand2_1 _18071_ (.Y(_02659_),
    .A(net3205),
    .B(net4814));
 sg13g2_o21ai_1 _18072_ (.B1(_02659_),
    .Y(_01982_),
    .A1(net5504),
    .A2(net4814));
 sg13g2_nand2_1 _18073_ (.Y(_02660_),
    .A(net2215),
    .B(net4814));
 sg13g2_o21ai_1 _18074_ (.B1(_02660_),
    .Y(_01983_),
    .A1(net5550),
    .A2(net4814));
 sg13g2_nand2_1 _18075_ (.Y(_02661_),
    .A(net2707),
    .B(net4815));
 sg13g2_o21ai_1 _18076_ (.B1(_02661_),
    .Y(_01984_),
    .A1(net5593),
    .A2(_02657_));
 sg13g2_nand2_1 _18077_ (.Y(_02662_),
    .A(net3275),
    .B(net4815));
 sg13g2_o21ai_1 _18078_ (.B1(_02662_),
    .Y(_01985_),
    .A1(net5636),
    .A2(net4815));
 sg13g2_nand2_1 _18079_ (.Y(_02663_),
    .A(net2894),
    .B(net4815));
 sg13g2_o21ai_1 _18080_ (.B1(_02663_),
    .Y(_01986_),
    .A1(net5681),
    .A2(net4815));
 sg13g2_nand2_1 _18081_ (.Y(_02664_),
    .A(net2251),
    .B(net4815));
 sg13g2_o21ai_1 _18082_ (.B1(_02664_),
    .Y(_01987_),
    .A1(net5726),
    .A2(net4815));
 sg13g2_nand2_1 _18083_ (.Y(_02665_),
    .A(net3071),
    .B(net4814));
 sg13g2_o21ai_1 _18084_ (.B1(_02665_),
    .Y(_01988_),
    .A1(net5773),
    .A2(net4814));
 sg13g2_nand2_1 _18085_ (.Y(_02666_),
    .A(net5245),
    .B(net5202));
 sg13g2_nand2_1 _18086_ (.Y(_02667_),
    .A(net2355),
    .B(net4813));
 sg13g2_o21ai_1 _18087_ (.B1(_02667_),
    .Y(_01989_),
    .A1(net5458),
    .A2(net4813));
 sg13g2_nand2_1 _18088_ (.Y(_02668_),
    .A(net2487),
    .B(net4813));
 sg13g2_o21ai_1 _18089_ (.B1(_02668_),
    .Y(_01990_),
    .A1(net5505),
    .A2(net4813));
 sg13g2_nand2_1 _18090_ (.Y(_02669_),
    .A(net2673),
    .B(net4813));
 sg13g2_o21ai_1 _18091_ (.B1(_02669_),
    .Y(_01991_),
    .A1(net5550),
    .A2(net4813));
 sg13g2_nand2_1 _18092_ (.Y(_02670_),
    .A(net3211),
    .B(net4812));
 sg13g2_o21ai_1 _18093_ (.B1(_02670_),
    .Y(_01992_),
    .A1(net5591),
    .A2(net4812));
 sg13g2_nand2_1 _18094_ (.Y(_02671_),
    .A(net2396),
    .B(net4812));
 sg13g2_o21ai_1 _18095_ (.B1(_02671_),
    .Y(_01993_),
    .A1(net5639),
    .A2(net4812));
 sg13g2_nand2_1 _18096_ (.Y(_02672_),
    .A(net2502),
    .B(net4812));
 sg13g2_o21ai_1 _18097_ (.B1(_02672_),
    .Y(_01994_),
    .A1(net5683),
    .A2(net4812));
 sg13g2_nand2_1 _18098_ (.Y(_02673_),
    .A(net2140),
    .B(net4812));
 sg13g2_o21ai_1 _18099_ (.B1(_02673_),
    .Y(_01995_),
    .A1(net5726),
    .A2(net4812));
 sg13g2_nand2_1 _18100_ (.Y(_02674_),
    .A(net2168),
    .B(net4813));
 sg13g2_o21ai_1 _18101_ (.B1(_02674_),
    .Y(_01996_),
    .A1(net5776),
    .A2(net4813));
 sg13g2_nand2_2 _18102_ (.Y(_02675_),
    .A(net5251),
    .B(net5202));
 sg13g2_nand2_1 _18103_ (.Y(_02676_),
    .A(net2416),
    .B(net4810));
 sg13g2_o21ai_1 _18104_ (.B1(_02676_),
    .Y(_01997_),
    .A1(net5458),
    .A2(net4810));
 sg13g2_nand2_1 _18105_ (.Y(_02677_),
    .A(net2286),
    .B(net4810));
 sg13g2_o21ai_1 _18106_ (.B1(_02677_),
    .Y(_01998_),
    .A1(net5505),
    .A2(net4810));
 sg13g2_nand2_1 _18107_ (.Y(_02678_),
    .A(net2320),
    .B(_02675_));
 sg13g2_o21ai_1 _18108_ (.B1(_02678_),
    .Y(_01999_),
    .A1(net5549),
    .A2(net4810));
 sg13g2_nand2_1 _18109_ (.Y(_02679_),
    .A(net2736),
    .B(net4811));
 sg13g2_o21ai_1 _18110_ (.B1(_02679_),
    .Y(_02000_),
    .A1(net5591),
    .A2(net4811));
 sg13g2_nand2_1 _18111_ (.Y(_02680_),
    .A(net3323),
    .B(net4811));
 sg13g2_o21ai_1 _18112_ (.B1(_02680_),
    .Y(_02001_),
    .A1(net5639),
    .A2(net4811));
 sg13g2_nand2_1 _18113_ (.Y(_02681_),
    .A(net3404),
    .B(net4811));
 sg13g2_o21ai_1 _18114_ (.B1(_02681_),
    .Y(_02002_),
    .A1(net5683),
    .A2(net4811));
 sg13g2_nand2_1 _18115_ (.Y(_02682_),
    .A(net3173),
    .B(net4810));
 sg13g2_o21ai_1 _18116_ (.B1(_02682_),
    .Y(_02003_),
    .A1(net5726),
    .A2(net4811));
 sg13g2_nand2_1 _18117_ (.Y(_02683_),
    .A(net2649),
    .B(net4810));
 sg13g2_o21ai_1 _18118_ (.B1(_02683_),
    .Y(_02004_),
    .A1(net5775),
    .A2(net4810));
 sg13g2_nand2_2 _18119_ (.Y(_02684_),
    .A(net5246),
    .B(net5202));
 sg13g2_nand2_1 _18120_ (.Y(_02685_),
    .A(net2667),
    .B(net4808));
 sg13g2_o21ai_1 _18121_ (.B1(_02685_),
    .Y(_02005_),
    .A1(net5458),
    .A2(net4808));
 sg13g2_nand2_1 _18122_ (.Y(_02686_),
    .A(net2249),
    .B(net4808));
 sg13g2_o21ai_1 _18123_ (.B1(_02686_),
    .Y(_02006_),
    .A1(net5505),
    .A2(net4808));
 sg13g2_nand2_1 _18124_ (.Y(_02687_),
    .A(net3102),
    .B(_02684_));
 sg13g2_o21ai_1 _18125_ (.B1(_02687_),
    .Y(_02007_),
    .A1(net5549),
    .A2(net4808));
 sg13g2_nand2_1 _18126_ (.Y(_02688_),
    .A(net2263),
    .B(net4809));
 sg13g2_o21ai_1 _18127_ (.B1(_02688_),
    .Y(_02008_),
    .A1(net5592),
    .A2(net4809));
 sg13g2_nand2_1 _18128_ (.Y(_02689_),
    .A(net2609),
    .B(net4809));
 sg13g2_o21ai_1 _18129_ (.B1(_02689_),
    .Y(_02009_),
    .A1(net5638),
    .A2(net4809));
 sg13g2_nand2_1 _18130_ (.Y(_02690_),
    .A(net2517),
    .B(net4809));
 sg13g2_o21ai_1 _18131_ (.B1(_02690_),
    .Y(_02010_),
    .A1(net5683),
    .A2(net4809));
 sg13g2_nand2_1 _18132_ (.Y(_02691_),
    .A(net2316),
    .B(net4808));
 sg13g2_o21ai_1 _18133_ (.B1(_02691_),
    .Y(_02011_),
    .A1(net5728),
    .A2(net4809));
 sg13g2_nand2_1 _18134_ (.Y(_02692_),
    .A(net2647),
    .B(net4808));
 sg13g2_o21ai_1 _18135_ (.B1(_02692_),
    .Y(_02012_),
    .A1(net5776),
    .A2(net4808));
 sg13g2_nand2_1 _18136_ (.Y(_02693_),
    .A(net5238),
    .B(_03363_));
 sg13g2_nand2_1 _18137_ (.Y(_02694_),
    .A(net2297),
    .B(net4806));
 sg13g2_o21ai_1 _18138_ (.B1(_02694_),
    .Y(_02013_),
    .A1(net5452),
    .A2(net4806));
 sg13g2_nand2_1 _18139_ (.Y(_02695_),
    .A(net2718),
    .B(net4806));
 sg13g2_o21ai_1 _18140_ (.B1(_02695_),
    .Y(_02014_),
    .A1(net5498),
    .A2(net4806));
 sg13g2_nand2_1 _18141_ (.Y(_02696_),
    .A(net2394),
    .B(net4806));
 sg13g2_o21ai_1 _18142_ (.B1(_02696_),
    .Y(_02015_),
    .A1(net5541),
    .A2(net4806));
 sg13g2_nand2_1 _18143_ (.Y(_02697_),
    .A(net2465),
    .B(net4807));
 sg13g2_o21ai_1 _18144_ (.B1(_02697_),
    .Y(_02016_),
    .A1(net5596),
    .A2(net4807));
 sg13g2_nand2_1 _18145_ (.Y(_02698_),
    .A(net2832),
    .B(net4807));
 sg13g2_o21ai_1 _18146_ (.B1(_02698_),
    .Y(_02017_),
    .A1(net5642),
    .A2(net4807));
 sg13g2_nand2_1 _18147_ (.Y(_02699_),
    .A(net2558),
    .B(net4807));
 sg13g2_o21ai_1 _18148_ (.B1(_02699_),
    .Y(_02018_),
    .A1(net5687),
    .A2(net4807));
 sg13g2_nand2_1 _18149_ (.Y(_02700_),
    .A(net2767),
    .B(net4807));
 sg13g2_o21ai_1 _18150_ (.B1(_02700_),
    .Y(_02019_),
    .A1(net5732),
    .A2(net4807));
 sg13g2_nand2_1 _18151_ (.Y(_02701_),
    .A(net2646),
    .B(net4806));
 sg13g2_o21ai_1 _18152_ (.B1(_02701_),
    .Y(_02020_),
    .A1(net5767),
    .A2(net4806));
 sg13g2_and2_1 _18153_ (.A(net5248),
    .B(_06139_),
    .X(_02702_));
 sg13g2_nor2_1 _18154_ (.A(net3860),
    .B(net4805),
    .Y(_02703_));
 sg13g2_a21oi_1 _18155_ (.A1(net5431),
    .A2(net4805),
    .Y(_02021_),
    .B1(_02703_));
 sg13g2_nor2_1 _18156_ (.A(net3909),
    .B(net4804),
    .Y(_02704_));
 sg13g2_a21oi_1 _18157_ (.A1(net5479),
    .A2(net4804),
    .Y(_02022_),
    .B1(_02704_));
 sg13g2_nor2_1 _18158_ (.A(net3789),
    .B(net4805),
    .Y(_02705_));
 sg13g2_a21oi_1 _18159_ (.A1(net5522),
    .A2(net4805),
    .Y(_02023_),
    .B1(_02705_));
 sg13g2_nor2_1 _18160_ (.A(net3520),
    .B(net4804),
    .Y(_02706_));
 sg13g2_a21oi_1 _18161_ (.A1(net5567),
    .A2(net4804),
    .Y(_02024_),
    .B1(_02706_));
 sg13g2_nor2_1 _18162_ (.A(net3508),
    .B(net4804),
    .Y(_02707_));
 sg13g2_a21oi_1 _18163_ (.A1(net5611),
    .A2(net4804),
    .Y(_02025_),
    .B1(_02707_));
 sg13g2_nor2_1 _18164_ (.A(net3710),
    .B(net4805),
    .Y(_02708_));
 sg13g2_a21oi_1 _18165_ (.A1(net5656),
    .A2(net4805),
    .Y(_02026_),
    .B1(_02708_));
 sg13g2_nor2_1 _18166_ (.A(net3677),
    .B(net4805),
    .Y(_02709_));
 sg13g2_a21oi_1 _18167_ (.A1(net5703),
    .A2(net4805),
    .Y(_02027_),
    .B1(_02709_));
 sg13g2_nor2_1 _18168_ (.A(net3624),
    .B(net4804),
    .Y(_02710_));
 sg13g2_a21oi_1 _18169_ (.A1(net5748),
    .A2(net4804),
    .Y(_02028_),
    .B1(_02710_));
 sg13g2_nand2_1 _18170_ (.Y(_02711_),
    .A(_03139_),
    .B(_06139_));
 sg13g2_nand2_1 _18171_ (.Y(_02712_),
    .A(net3082),
    .B(net4803));
 sg13g2_o21ai_1 _18172_ (.B1(_02712_),
    .Y(_02029_),
    .A1(net5431),
    .A2(net4803));
 sg13g2_nand2_1 _18173_ (.Y(_02713_),
    .A(net2841),
    .B(net4803));
 sg13g2_o21ai_1 _18174_ (.B1(_02713_),
    .Y(_02030_),
    .A1(net5479),
    .A2(net4803));
 sg13g2_nand2_1 _18175_ (.Y(_02714_),
    .A(net2366),
    .B(net4803));
 sg13g2_o21ai_1 _18176_ (.B1(_02714_),
    .Y(_02031_),
    .A1(net5521),
    .A2(net4803));
 sg13g2_nand2_1 _18177_ (.Y(_02715_),
    .A(net2338),
    .B(net4802));
 sg13g2_o21ai_1 _18178_ (.B1(_02715_),
    .Y(_02032_),
    .A1(net5566),
    .A2(net4802));
 sg13g2_nand2_1 _18179_ (.Y(_02716_),
    .A(net2766),
    .B(net4802));
 sg13g2_o21ai_1 _18180_ (.B1(_02716_),
    .Y(_02033_),
    .A1(net5611),
    .A2(net4802));
 sg13g2_nand2_1 _18181_ (.Y(_02717_),
    .A(net2430),
    .B(net4802));
 sg13g2_o21ai_1 _18182_ (.B1(_02717_),
    .Y(_02034_),
    .A1(net5660),
    .A2(net4802));
 sg13g2_nand2_1 _18183_ (.Y(_02718_),
    .A(net2530),
    .B(net4803));
 sg13g2_o21ai_1 _18184_ (.B1(_02718_),
    .Y(_02035_),
    .A1(net5710),
    .A2(_02711_));
 sg13g2_nand2_1 _18185_ (.Y(_02719_),
    .A(net3120),
    .B(net4802));
 sg13g2_o21ai_1 _18186_ (.B1(_02719_),
    .Y(_02036_),
    .A1(net5748),
    .A2(net4802));
 sg13g2_nand2_1 _18187_ (.Y(_02720_),
    .A(_03079_),
    .B(_06139_));
 sg13g2_nand2_1 _18188_ (.Y(_02721_),
    .A(net2580),
    .B(net4801));
 sg13g2_o21ai_1 _18189_ (.B1(_02721_),
    .Y(_02037_),
    .A1(net5431),
    .A2(net4801));
 sg13g2_nand2_1 _18190_ (.Y(_02722_),
    .A(net2397),
    .B(net4800));
 sg13g2_o21ai_1 _18191_ (.B1(_02722_),
    .Y(_02038_),
    .A1(net5479),
    .A2(net4800));
 sg13g2_nand2_1 _18192_ (.Y(_02723_),
    .A(net2422),
    .B(net4801));
 sg13g2_o21ai_1 _18193_ (.B1(_02723_),
    .Y(_02039_),
    .A1(net5521),
    .A2(net4801));
 sg13g2_nand2_1 _18194_ (.Y(_02724_),
    .A(net2990),
    .B(net4800));
 sg13g2_o21ai_1 _18195_ (.B1(_02724_),
    .Y(_02040_),
    .A1(net5566),
    .A2(net4800));
 sg13g2_nand2_1 _18196_ (.Y(_02725_),
    .A(net2666),
    .B(net4800));
 sg13g2_o21ai_1 _18197_ (.B1(_02725_),
    .Y(_02041_),
    .A1(net5611),
    .A2(net4800));
 sg13g2_nand2_1 _18198_ (.Y(_02726_),
    .A(net3022),
    .B(net4801));
 sg13g2_o21ai_1 _18199_ (.B1(_02726_),
    .Y(_02042_),
    .A1(net5666),
    .A2(net4801));
 sg13g2_nand2_1 _18200_ (.Y(_02727_),
    .A(net3357),
    .B(net4801));
 sg13g2_o21ai_1 _18201_ (.B1(_02727_),
    .Y(_02043_),
    .A1(net5710),
    .A2(net4801));
 sg13g2_nand2_1 _18202_ (.Y(_02728_),
    .A(net3240),
    .B(net4800));
 sg13g2_o21ai_1 _18203_ (.B1(_02728_),
    .Y(_02044_),
    .A1(net5748),
    .A2(net4800));
 sg13g2_nor2_1 _18204_ (.A(_03120_),
    .B(_06140_),
    .Y(_02729_));
 sg13g2_nor2_1 _18205_ (.A(net3984),
    .B(net5169),
    .Y(_02730_));
 sg13g2_a21oi_1 _18206_ (.A1(net5431),
    .A2(net5169),
    .Y(_02045_),
    .B1(_02730_));
 sg13g2_nor2_1 _18207_ (.A(net4003),
    .B(net5169),
    .Y(_02731_));
 sg13g2_a21oi_1 _18208_ (.A1(net5479),
    .A2(net5169),
    .Y(_02046_),
    .B1(_02731_));
 sg13g2_nor2_1 _18209_ (.A(net3380),
    .B(net5169),
    .Y(_02732_));
 sg13g2_a21oi_1 _18210_ (.A1(net5521),
    .A2(net5169),
    .Y(_02047_),
    .B1(_02732_));
 sg13g2_nor2_1 _18211_ (.A(net3706),
    .B(net5168),
    .Y(_02733_));
 sg13g2_a21oi_1 _18212_ (.A1(net5566),
    .A2(net5168),
    .Y(_02048_),
    .B1(_02733_));
 sg13g2_nor2_1 _18213_ (.A(net3467),
    .B(net5168),
    .Y(_02734_));
 sg13g2_a21oi_1 _18214_ (.A1(net5623),
    .A2(net5168),
    .Y(_02049_),
    .B1(_02734_));
 sg13g2_nor2_1 _18215_ (.A(net3366),
    .B(net5168),
    .Y(_02735_));
 sg13g2_a21oi_1 _18216_ (.A1(net5666),
    .A2(net5168),
    .Y(_02050_),
    .B1(_02735_));
 sg13g2_nor2_1 _18217_ (.A(net3703),
    .B(net5169),
    .Y(_02736_));
 sg13g2_a21oi_1 _18218_ (.A1(net5710),
    .A2(_02729_),
    .Y(_02051_),
    .B1(_02736_));
 sg13g2_nor2_1 _18219_ (.A(net3841),
    .B(net5168),
    .Y(_02737_));
 sg13g2_a21oi_1 _18220_ (.A1(net5748),
    .A2(net5168),
    .Y(_02052_),
    .B1(_02737_));
 sg13g2_nor2_1 _18221_ (.A(_03109_),
    .B(_06140_),
    .Y(_02738_));
 sg13g2_nor2_1 _18222_ (.A(net3578),
    .B(net5166),
    .Y(_02739_));
 sg13g2_a21oi_1 _18223_ (.A1(net5432),
    .A2(net5166),
    .Y(_02053_),
    .B1(_02739_));
 sg13g2_nor2_1 _18224_ (.A(net2937),
    .B(net5167),
    .Y(_02740_));
 sg13g2_a21oi_1 _18225_ (.A1(net5477),
    .A2(net5167),
    .Y(_02054_),
    .B1(_02740_));
 sg13g2_nor2_1 _18226_ (.A(net3667),
    .B(net5167),
    .Y(_02741_));
 sg13g2_a21oi_1 _18227_ (.A1(net5522),
    .A2(net5167),
    .Y(_02055_),
    .B1(_02741_));
 sg13g2_nor2_1 _18228_ (.A(net3423),
    .B(net5167),
    .Y(_02742_));
 sg13g2_a21oi_1 _18229_ (.A1(net5568),
    .A2(net5167),
    .Y(_02056_),
    .B1(_02742_));
 sg13g2_nor2_1 _18230_ (.A(net3963),
    .B(net5166),
    .Y(_02743_));
 sg13g2_a21oi_1 _18231_ (.A1(net5612),
    .A2(net5166),
    .Y(_02057_),
    .B1(_02743_));
 sg13g2_nor2_1 _18232_ (.A(net3646),
    .B(net5166),
    .Y(_02744_));
 sg13g2_a21oi_1 _18233_ (.A1(net5657),
    .A2(net5166),
    .Y(_02058_),
    .B1(_02744_));
 sg13g2_nor2_1 _18234_ (.A(net3742),
    .B(net5167),
    .Y(_02745_));
 sg13g2_a21oi_1 _18235_ (.A1(net5703),
    .A2(net5167),
    .Y(_02059_),
    .B1(_02745_));
 sg13g2_nor2_1 _18236_ (.A(net3906),
    .B(net5166),
    .Y(_02746_));
 sg13g2_a21oi_1 _18237_ (.A1(net5749),
    .A2(net5166),
    .Y(_02060_),
    .B1(_02746_));
 sg13g2_nand2_1 _18238_ (.Y(_02747_),
    .A(net5234),
    .B(_06139_));
 sg13g2_nand2_1 _18239_ (.Y(_02748_),
    .A(net2815),
    .B(net4798));
 sg13g2_o21ai_1 _18240_ (.B1(_02748_),
    .Y(_02061_),
    .A1(net5432),
    .A2(net4798));
 sg13g2_nand2_1 _18241_ (.Y(_02749_),
    .A(net2870),
    .B(net4799));
 sg13g2_o21ai_1 _18242_ (.B1(_02749_),
    .Y(_02062_),
    .A1(net5477),
    .A2(net4799));
 sg13g2_nand2_1 _18243_ (.Y(_02750_),
    .A(net2369),
    .B(net4799));
 sg13g2_o21ai_1 _18244_ (.B1(_02750_),
    .Y(_02063_),
    .A1(net5522),
    .A2(net4799));
 sg13g2_nand2_1 _18245_ (.Y(_02751_),
    .A(net3010),
    .B(net4799));
 sg13g2_o21ai_1 _18246_ (.B1(_02751_),
    .Y(_02064_),
    .A1(net5567),
    .A2(net4799));
 sg13g2_nand2_1 _18247_ (.Y(_02752_),
    .A(net2525),
    .B(net4798));
 sg13g2_o21ai_1 _18248_ (.B1(_02752_),
    .Y(_02065_),
    .A1(net5612),
    .A2(net4798));
 sg13g2_nand2_1 _18249_ (.Y(_02753_),
    .A(net2403),
    .B(net4798));
 sg13g2_o21ai_1 _18250_ (.B1(_02753_),
    .Y(_02066_),
    .A1(net5659),
    .A2(net4798));
 sg13g2_nand2_1 _18251_ (.Y(_02754_),
    .A(net2557),
    .B(net4799));
 sg13g2_o21ai_1 _18252_ (.B1(_02754_),
    .Y(_02067_),
    .A1(net5703),
    .A2(net4799));
 sg13g2_nand2_1 _18253_ (.Y(_02755_),
    .A(net3189),
    .B(net4798));
 sg13g2_o21ai_1 _18254_ (.B1(_02755_),
    .Y(_02068_),
    .A1(net5749),
    .A2(net4798));
 sg13g2_nand2_1 _18255_ (.Y(_02756_),
    .A(net5236),
    .B(_06139_));
 sg13g2_nand2_1 _18256_ (.Y(_02757_),
    .A(net3286),
    .B(net4796));
 sg13g2_o21ai_1 _18257_ (.B1(_02757_),
    .Y(_02069_),
    .A1(net5432),
    .A2(net4796));
 sg13g2_nand2_1 _18258_ (.Y(_02758_),
    .A(net2223),
    .B(net4797));
 sg13g2_o21ai_1 _18259_ (.B1(_02758_),
    .Y(_02070_),
    .A1(net5477),
    .A2(net4797));
 sg13g2_nand2_1 _18260_ (.Y(_02759_),
    .A(net2389),
    .B(net4797));
 sg13g2_o21ai_1 _18261_ (.B1(_02759_),
    .Y(_02071_),
    .A1(net5522),
    .A2(net4797));
 sg13g2_nand2_1 _18262_ (.Y(_02760_),
    .A(net2729),
    .B(net4797));
 sg13g2_o21ai_1 _18263_ (.B1(_02760_),
    .Y(_02072_),
    .A1(net5567),
    .A2(net4797));
 sg13g2_nand2_1 _18264_ (.Y(_02761_),
    .A(net2634),
    .B(net4796));
 sg13g2_o21ai_1 _18265_ (.B1(_02761_),
    .Y(_02073_),
    .A1(net5612),
    .A2(net4796));
 sg13g2_nand2_1 _18266_ (.Y(_02762_),
    .A(net2220),
    .B(net4796));
 sg13g2_o21ai_1 _18267_ (.B1(_02762_),
    .Y(_02074_),
    .A1(net5660),
    .A2(net4796));
 sg13g2_nand2_1 _18268_ (.Y(_02763_),
    .A(net3555),
    .B(net4797));
 sg13g2_o21ai_1 _18269_ (.B1(_02763_),
    .Y(_02075_),
    .A1(net5712),
    .A2(net4797));
 sg13g2_nand2_1 _18270_ (.Y(_02764_),
    .A(net2298),
    .B(net4796));
 sg13g2_o21ai_1 _18271_ (.B1(_02764_),
    .Y(_02076_),
    .A1(net5749),
    .A2(net4796));
 sg13g2_nand2_1 _18272_ (.Y(_02765_),
    .A(net5237),
    .B(_06139_));
 sg13g2_nand2_1 _18273_ (.Y(_02766_),
    .A(net2818),
    .B(net4794));
 sg13g2_o21ai_1 _18274_ (.B1(_02766_),
    .Y(_02077_),
    .A1(net5432),
    .A2(net4794));
 sg13g2_nand2_1 _18275_ (.Y(_02767_),
    .A(net3070),
    .B(net4795));
 sg13g2_o21ai_1 _18276_ (.B1(_02767_),
    .Y(_02078_),
    .A1(net5477),
    .A2(net4795));
 sg13g2_nand2_1 _18277_ (.Y(_02768_),
    .A(net2555),
    .B(net4795));
 sg13g2_o21ai_1 _18278_ (.B1(_02768_),
    .Y(_02079_),
    .A1(net5522),
    .A2(net4795));
 sg13g2_nand2_1 _18279_ (.Y(_02769_),
    .A(net2564),
    .B(net4795));
 sg13g2_o21ai_1 _18280_ (.B1(_02769_),
    .Y(_02080_),
    .A1(net5567),
    .A2(net4795));
 sg13g2_nand2_1 _18281_ (.Y(_02770_),
    .A(net2561),
    .B(net4794));
 sg13g2_o21ai_1 _18282_ (.B1(_02770_),
    .Y(_02081_),
    .A1(net5612),
    .A2(net4794));
 sg13g2_nand2_1 _18283_ (.Y(_02771_),
    .A(net2477),
    .B(net4794));
 sg13g2_o21ai_1 _18284_ (.B1(_02771_),
    .Y(_02082_),
    .A1(net5659),
    .A2(net4794));
 sg13g2_nand2_1 _18285_ (.Y(_02772_),
    .A(net2785),
    .B(net4795));
 sg13g2_o21ai_1 _18286_ (.B1(_02772_),
    .Y(_02083_),
    .A1(net5712),
    .A2(net4795));
 sg13g2_nand2_1 _18287_ (.Y(_02773_),
    .A(net2742),
    .B(net4794));
 sg13g2_o21ai_1 _18288_ (.B1(_02773_),
    .Y(_02084_),
    .A1(net5749),
    .A2(net4794));
 sg13g2_nor2_1 _18289_ (.A(_02939_),
    .B(_06140_),
    .Y(_02774_));
 sg13g2_nor2_1 _18290_ (.A(net4102),
    .B(net5165),
    .Y(_02775_));
 sg13g2_a21oi_1 _18291_ (.A1(net5431),
    .A2(net5165),
    .Y(_02085_),
    .B1(_02775_));
 sg13g2_nor2_1 _18292_ (.A(net3512),
    .B(net5165),
    .Y(_02776_));
 sg13g2_a21oi_1 _18293_ (.A1(net5478),
    .A2(net5165),
    .Y(_02086_),
    .B1(_02776_));
 sg13g2_nor2_1 _18294_ (.A(net3316),
    .B(net5165),
    .Y(_02777_));
 sg13g2_a21oi_1 _18295_ (.A1(net5521),
    .A2(net5165),
    .Y(_02087_),
    .B1(_02777_));
 sg13g2_nor2_1 _18296_ (.A(net3719),
    .B(net5164),
    .Y(_02778_));
 sg13g2_a21oi_1 _18297_ (.A1(net5566),
    .A2(net5164),
    .Y(_02088_),
    .B1(_02778_));
 sg13g2_nor2_1 _18298_ (.A(net3591),
    .B(net5164),
    .Y(_02779_));
 sg13g2_a21oi_1 _18299_ (.A1(net5611),
    .A2(net5164),
    .Y(_02089_),
    .B1(_02779_));
 sg13g2_nor2_1 _18300_ (.A(net4020),
    .B(net5164),
    .Y(_02780_));
 sg13g2_a21oi_1 _18301_ (.A1(net5656),
    .A2(net5164),
    .Y(_02090_),
    .B1(_02780_));
 sg13g2_nor2_1 _18302_ (.A(net3621),
    .B(net5165),
    .Y(_02781_));
 sg13g2_a21oi_1 _18303_ (.A1(net5703),
    .A2(net5165),
    .Y(_02091_),
    .B1(_02781_));
 sg13g2_nor2_1 _18304_ (.A(net4062),
    .B(net5164),
    .Y(_02782_));
 sg13g2_a21oi_1 _18305_ (.A1(net5748),
    .A2(net5164),
    .Y(_02092_),
    .B1(_02782_));
 sg13g2_nor2_1 _18306_ (.A(_02939_),
    .B(net5210),
    .Y(_02783_));
 sg13g2_nor2_1 _18307_ (.A(net4037),
    .B(net4793),
    .Y(_02784_));
 sg13g2_a21oi_1 _18308_ (.A1(net5449),
    .A2(net4793),
    .Y(_02093_),
    .B1(_02784_));
 sg13g2_nor2_1 _18309_ (.A(net3811),
    .B(net4793),
    .Y(_02785_));
 sg13g2_a21oi_1 _18310_ (.A1(net5495),
    .A2(net4793),
    .Y(_02094_),
    .B1(_02785_));
 sg13g2_nor2_1 _18311_ (.A(net4106),
    .B(net4792),
    .Y(_02786_));
 sg13g2_a21oi_1 _18312_ (.A1(net5552),
    .A2(net4793),
    .Y(_02095_),
    .B1(_02786_));
 sg13g2_nor2_1 _18313_ (.A(net4060),
    .B(_02783_),
    .Y(_02787_));
 sg13g2_a21oi_1 _18314_ (.A1(net5595),
    .A2(net4792),
    .Y(_02096_),
    .B1(_02787_));
 sg13g2_nor2_1 _18315_ (.A(net3875),
    .B(net4792),
    .Y(_02788_));
 sg13g2_a21oi_1 _18316_ (.A1(net5640),
    .A2(net4792),
    .Y(_02097_),
    .B1(_02788_));
 sg13g2_nor2_1 _18317_ (.A(net3859),
    .B(net4792),
    .Y(_02789_));
 sg13g2_a21oi_1 _18318_ (.A1(net5686),
    .A2(net4792),
    .Y(_02098_),
    .B1(_02789_));
 sg13g2_nor2_1 _18319_ (.A(net3349),
    .B(net4792),
    .Y(_02790_));
 sg13g2_a21oi_1 _18320_ (.A1(net5730),
    .A2(net4792),
    .Y(_02099_),
    .B1(_02790_));
 sg13g2_nor2_1 _18321_ (.A(net3532),
    .B(net4793),
    .Y(_02791_));
 sg13g2_a21oi_1 _18322_ (.A1(net5765),
    .A2(net4793),
    .Y(_02100_),
    .B1(_02791_));
 sg13g2_nand2_1 _18323_ (.Y(_02792_),
    .A(net5242),
    .B(_06139_));
 sg13g2_nand2_1 _18324_ (.Y(_02793_),
    .A(net3046),
    .B(net4791));
 sg13g2_o21ai_1 _18325_ (.B1(_02793_),
    .Y(_02101_),
    .A1(net5431),
    .A2(net4791));
 sg13g2_nand2_1 _18326_ (.Y(_02794_),
    .A(net2836),
    .B(net4791));
 sg13g2_o21ai_1 _18327_ (.B1(_02794_),
    .Y(_02102_),
    .A1(net5478),
    .A2(net4791));
 sg13g2_nand2_1 _18328_ (.Y(_02795_),
    .A(net3213),
    .B(net4791));
 sg13g2_o21ai_1 _18329_ (.B1(_02795_),
    .Y(_02103_),
    .A1(net5521),
    .A2(net4791));
 sg13g2_nand2_1 _18330_ (.Y(_02796_),
    .A(net3089),
    .B(net4790));
 sg13g2_o21ai_1 _18331_ (.B1(_02796_),
    .Y(_02104_),
    .A1(net5566),
    .A2(net4790));
 sg13g2_nand2_1 _18332_ (.Y(_02797_),
    .A(net2685),
    .B(net4790));
 sg13g2_o21ai_1 _18333_ (.B1(_02797_),
    .Y(_02105_),
    .A1(net5611),
    .A2(net4790));
 sg13g2_nand2_1 _18334_ (.Y(_02798_),
    .A(net2820),
    .B(net4790));
 sg13g2_o21ai_1 _18335_ (.B1(_02798_),
    .Y(_02106_),
    .A1(net5656),
    .A2(net4790));
 sg13g2_nand2_1 _18336_ (.Y(_02799_),
    .A(net2570),
    .B(net4791));
 sg13g2_o21ai_1 _18337_ (.B1(_02799_),
    .Y(_02107_),
    .A1(net5703),
    .A2(net4791));
 sg13g2_nand2_1 _18338_ (.Y(_02800_),
    .A(net3264),
    .B(net4790));
 sg13g2_o21ai_1 _18339_ (.B1(_02800_),
    .Y(_02108_),
    .A1(net5748),
    .A2(net4790));
 sg13g2_nor2_1 _18340_ (.A(_02964_),
    .B(_06140_),
    .Y(_02801_));
 sg13g2_nor2_1 _18341_ (.A(net3800),
    .B(net5163),
    .Y(_02802_));
 sg13g2_a21oi_1 _18342_ (.A1(net5432),
    .A2(net5163),
    .Y(_02109_),
    .B1(_02802_));
 sg13g2_nor2_1 _18343_ (.A(net3872),
    .B(net5163),
    .Y(_02803_));
 sg13g2_a21oi_1 _18344_ (.A1(net5478),
    .A2(net5163),
    .Y(_02110_),
    .B1(_02803_));
 sg13g2_nor2_1 _18345_ (.A(net3625),
    .B(net5163),
    .Y(_02804_));
 sg13g2_a21oi_1 _18346_ (.A1(net5521),
    .A2(net5163),
    .Y(_02111_),
    .B1(_02804_));
 sg13g2_nor2_1 _18347_ (.A(net3991),
    .B(net5162),
    .Y(_02805_));
 sg13g2_a21oi_1 _18348_ (.A1(net5566),
    .A2(net5162),
    .Y(_02112_),
    .B1(_02805_));
 sg13g2_nor2_1 _18349_ (.A(net3965),
    .B(net5162),
    .Y(_02806_));
 sg13g2_a21oi_1 _18350_ (.A1(net5611),
    .A2(net5162),
    .Y(_02113_),
    .B1(_02806_));
 sg13g2_nor2_1 _18351_ (.A(net3814),
    .B(net5162),
    .Y(_02807_));
 sg13g2_a21oi_1 _18352_ (.A1(net5660),
    .A2(net5162),
    .Y(_02114_),
    .B1(_02807_));
 sg13g2_nor2_1 _18353_ (.A(net3483),
    .B(net5163),
    .Y(_02808_));
 sg13g2_a21oi_1 _18354_ (.A1(net5703),
    .A2(net5163),
    .Y(_02115_),
    .B1(_02808_));
 sg13g2_nor2_1 _18355_ (.A(net3554),
    .B(net5162),
    .Y(_02809_));
 sg13g2_a21oi_1 _18356_ (.A1(net5748),
    .A2(net5162),
    .Y(_02116_),
    .B1(_02809_));
 sg13g2_nor2_1 _18357_ (.A(_03017_),
    .B(net5143),
    .Y(_02810_));
 sg13g2_nor2_1 _18358_ (.A(net4023),
    .B(net4674),
    .Y(_02811_));
 sg13g2_a21oi_1 _18359_ (.A1(net5448),
    .A2(net4674),
    .Y(_02117_),
    .B1(_02811_));
 sg13g2_nor2_1 _18360_ (.A(net3837),
    .B(net4673),
    .Y(_02812_));
 sg13g2_a21oi_1 _18361_ (.A1(net5492),
    .A2(net4673),
    .Y(_02118_),
    .B1(_02812_));
 sg13g2_nor2_1 _18362_ (.A(net3547),
    .B(net4674),
    .Y(_02813_));
 sg13g2_a21oi_1 _18363_ (.A1(net5539),
    .A2(net4674),
    .Y(_02119_),
    .B1(_02813_));
 sg13g2_nor2_1 _18364_ (.A(net3891),
    .B(net4673),
    .Y(_02814_));
 sg13g2_a21oi_1 _18365_ (.A1(net5581),
    .A2(net4673),
    .Y(_02120_),
    .B1(_02814_));
 sg13g2_nor2_1 _18366_ (.A(net3540),
    .B(net4674),
    .Y(_02815_));
 sg13g2_a21oi_1 _18367_ (.A1(net5628),
    .A2(net4674),
    .Y(_02121_),
    .B1(_02815_));
 sg13g2_nor2_1 _18368_ (.A(net3758),
    .B(net4673),
    .Y(_02816_));
 sg13g2_a21oi_1 _18369_ (.A1(net5672),
    .A2(net4673),
    .Y(_02122_),
    .B1(_02816_));
 sg13g2_nor2_1 _18370_ (.A(net4000),
    .B(net4673),
    .Y(_02817_));
 sg13g2_a21oi_1 _18371_ (.A1(net5718),
    .A2(net4673),
    .Y(_02123_),
    .B1(_02817_));
 sg13g2_nor2_1 _18372_ (.A(net4116),
    .B(net4674),
    .Y(_02818_));
 sg13g2_a21oi_1 _18373_ (.A1(net5764),
    .A2(net4674),
    .Y(_02124_),
    .B1(_02818_));
 sg13g2_nand2_1 _18374_ (.Y(_02819_),
    .A(net11),
    .B(net4216));
 sg13g2_a21oi_2 _18375_ (.B1(net6176),
    .Y(_02125_),
    .A2(_02819_),
    .A1(net5261));
 sg13g2_a21oi_1 _18376_ (.A1(net5116),
    .A2(_03299_),
    .Y(_00580_),
    .B1(_03300_));
 sg13g2_a21oi_1 _18377_ (.A1(net5116),
    .A2(_03304_),
    .Y(_00581_),
    .B1(_03305_));
 sg13g2_a221oi_1 _18378_ (.B2(_03310_),
    .C1(net6177),
    .B1(net4237),
    .A1(_02830_),
    .Y(_00582_),
    .A2(_03296_));
 sg13g2_a21oi_1 _18379_ (.A1(_02829_),
    .A2(_03296_),
    .Y(_00583_),
    .B1(_03316_));
 sg13g2_nor2_1 _18380_ (.A(net6177),
    .B(_03322_),
    .Y(_00584_));
 sg13g2_nor2_1 _18381_ (.A(net6177),
    .B(_03330_),
    .Y(_00585_));
 sg13g2_a21oi_1 _18382_ (.A1(_03333_),
    .A2(_03336_),
    .Y(_00586_),
    .B1(_03337_));
 sg13g2_nor2_1 _18383_ (.A(net6177),
    .B(_03343_),
    .Y(_00587_));
 sg13g2_dfrbp_1 _18384_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net689),
    .D(_00027_),
    .Q_N(_09188_),
    .Q(\mem.mem[88][0] ));
 sg13g2_dfrbp_1 _18385_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1365),
    .D(_00028_),
    .Q_N(_09187_),
    .Q(\mem.mem[88][1] ));
 sg13g2_dfrbp_1 _18386_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1364),
    .D(_00029_),
    .Q_N(_09186_),
    .Q(\mem.mem[88][2] ));
 sg13g2_dfrbp_1 _18387_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1363),
    .D(_00030_),
    .Q_N(_09185_),
    .Q(\mem.mem[88][3] ));
 sg13g2_dfrbp_1 _18388_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1362),
    .D(_00031_),
    .Q_N(_09184_),
    .Q(\mem.mem[88][4] ));
 sg13g2_dfrbp_1 _18389_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1361),
    .D(_00032_),
    .Q_N(_09183_),
    .Q(\mem.mem[88][5] ));
 sg13g2_dfrbp_1 _18390_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1360),
    .D(_00033_),
    .Q_N(_09182_),
    .Q(\mem.mem[88][6] ));
 sg13g2_dfrbp_1 _18391_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1359),
    .D(_00034_),
    .Q_N(_09181_),
    .Q(\mem.mem[88][7] ));
 sg13g2_dfrbp_1 _18392_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1358),
    .D(_00035_),
    .Q_N(_09180_),
    .Q(\mem.mem[43][0] ));
 sg13g2_dfrbp_1 _18393_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1357),
    .D(_00036_),
    .Q_N(_09179_),
    .Q(\mem.mem[43][1] ));
 sg13g2_dfrbp_1 _18394_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1356),
    .D(_00037_),
    .Q_N(_09178_),
    .Q(\mem.mem[43][2] ));
 sg13g2_dfrbp_1 _18395_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1355),
    .D(_00038_),
    .Q_N(_09177_),
    .Q(\mem.mem[43][3] ));
 sg13g2_dfrbp_1 _18396_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1354),
    .D(_00039_),
    .Q_N(_09176_),
    .Q(\mem.mem[43][4] ));
 sg13g2_dfrbp_1 _18397_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1353),
    .D(_00040_),
    .Q_N(_09175_),
    .Q(\mem.mem[43][5] ));
 sg13g2_dfrbp_1 _18398_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1352),
    .D(_00041_),
    .Q_N(_09174_),
    .Q(\mem.mem[43][6] ));
 sg13g2_dfrbp_1 _18399_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1351),
    .D(_00042_),
    .Q_N(_09173_),
    .Q(\mem.mem[43][7] ));
 sg13g2_dfrbp_1 _18400_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1350),
    .D(_00043_),
    .Q_N(_09172_),
    .Q(\mem.mem[42][0] ));
 sg13g2_dfrbp_1 _18401_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1349),
    .D(_00044_),
    .Q_N(_09171_),
    .Q(\mem.mem[42][1] ));
 sg13g2_dfrbp_1 _18402_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1348),
    .D(_00045_),
    .Q_N(_09170_),
    .Q(\mem.mem[42][2] ));
 sg13g2_dfrbp_1 _18403_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1347),
    .D(_00046_),
    .Q_N(_09169_),
    .Q(\mem.mem[42][3] ));
 sg13g2_dfrbp_1 _18404_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1346),
    .D(_00047_),
    .Q_N(_09168_),
    .Q(\mem.mem[42][4] ));
 sg13g2_dfrbp_1 _18405_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1345),
    .D(_00048_),
    .Q_N(_09167_),
    .Q(\mem.mem[42][5] ));
 sg13g2_dfrbp_1 _18406_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1344),
    .D(_00049_),
    .Q_N(_09166_),
    .Q(\mem.mem[42][6] ));
 sg13g2_dfrbp_1 _18407_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1343),
    .D(_00050_),
    .Q_N(_09165_),
    .Q(\mem.mem[42][7] ));
 sg13g2_dfrbp_1 _18408_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1342),
    .D(_00051_),
    .Q_N(_09164_),
    .Q(\mem.mem[74][0] ));
 sg13g2_dfrbp_1 _18409_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1341),
    .D(_00052_),
    .Q_N(_09163_),
    .Q(\mem.mem[74][1] ));
 sg13g2_dfrbp_1 _18410_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1340),
    .D(_00053_),
    .Q_N(_09162_),
    .Q(\mem.mem[74][2] ));
 sg13g2_dfrbp_1 _18411_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1339),
    .D(_00054_),
    .Q_N(_09161_),
    .Q(\mem.mem[74][3] ));
 sg13g2_dfrbp_1 _18412_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1338),
    .D(_00055_),
    .Q_N(_09160_),
    .Q(\mem.mem[74][4] ));
 sg13g2_dfrbp_1 _18413_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1337),
    .D(_00056_),
    .Q_N(_09159_),
    .Q(\mem.mem[74][5] ));
 sg13g2_dfrbp_1 _18414_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1336),
    .D(_00057_),
    .Q_N(_09158_),
    .Q(\mem.mem[74][6] ));
 sg13g2_dfrbp_1 _18415_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1335),
    .D(_00058_),
    .Q_N(_09157_),
    .Q(\mem.mem[74][7] ));
 sg13g2_dfrbp_1 _18416_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1334),
    .D(_00059_),
    .Q_N(_09156_),
    .Q(\mem.mem[47][0] ));
 sg13g2_dfrbp_1 _18417_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1333),
    .D(_00060_),
    .Q_N(_09155_),
    .Q(\mem.mem[47][1] ));
 sg13g2_dfrbp_1 _18418_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1332),
    .D(_00061_),
    .Q_N(_09154_),
    .Q(\mem.mem[47][2] ));
 sg13g2_dfrbp_1 _18419_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1331),
    .D(_00062_),
    .Q_N(_09153_),
    .Q(\mem.mem[47][3] ));
 sg13g2_dfrbp_1 _18420_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1330),
    .D(_00063_),
    .Q_N(_09152_),
    .Q(\mem.mem[47][4] ));
 sg13g2_dfrbp_1 _18421_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1329),
    .D(_00064_),
    .Q_N(_09151_),
    .Q(\mem.mem[47][5] ));
 sg13g2_dfrbp_1 _18422_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1328),
    .D(_00065_),
    .Q_N(_09150_),
    .Q(\mem.mem[47][6] ));
 sg13g2_dfrbp_1 _18423_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1327),
    .D(_00066_),
    .Q_N(_09149_),
    .Q(\mem.mem[47][7] ));
 sg13g2_dfrbp_1 _18424_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1326),
    .D(_00067_),
    .Q_N(_09148_),
    .Q(\mem.mem[41][0] ));
 sg13g2_dfrbp_1 _18425_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1325),
    .D(_00068_),
    .Q_N(_09147_),
    .Q(\mem.mem[41][1] ));
 sg13g2_dfrbp_1 _18426_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1324),
    .D(_00069_),
    .Q_N(_09146_),
    .Q(\mem.mem[41][2] ));
 sg13g2_dfrbp_1 _18427_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1323),
    .D(_00070_),
    .Q_N(_09145_),
    .Q(\mem.mem[41][3] ));
 sg13g2_dfrbp_1 _18428_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1322),
    .D(_00071_),
    .Q_N(_09144_),
    .Q(\mem.mem[41][4] ));
 sg13g2_dfrbp_1 _18429_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1321),
    .D(_00072_),
    .Q_N(_09143_),
    .Q(\mem.mem[41][5] ));
 sg13g2_dfrbp_1 _18430_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1320),
    .D(_00073_),
    .Q_N(_09142_),
    .Q(\mem.mem[41][6] ));
 sg13g2_dfrbp_1 _18431_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1319),
    .D(_00074_),
    .Q_N(_09141_),
    .Q(\mem.mem[41][7] ));
 sg13g2_dfrbp_1 _18432_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1318),
    .D(_00075_),
    .Q_N(_09140_),
    .Q(\mem.mem[73][0] ));
 sg13g2_dfrbp_1 _18433_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1317),
    .D(_00076_),
    .Q_N(_09139_),
    .Q(\mem.mem[73][1] ));
 sg13g2_dfrbp_1 _18434_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1316),
    .D(_00077_),
    .Q_N(_09138_),
    .Q(\mem.mem[73][2] ));
 sg13g2_dfrbp_1 _18435_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1315),
    .D(_00078_),
    .Q_N(_09137_),
    .Q(\mem.mem[73][3] ));
 sg13g2_dfrbp_1 _18436_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1314),
    .D(_00079_),
    .Q_N(_09136_),
    .Q(\mem.mem[73][4] ));
 sg13g2_dfrbp_1 _18437_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1313),
    .D(_00080_),
    .Q_N(_09135_),
    .Q(\mem.mem[73][5] ));
 sg13g2_dfrbp_1 _18438_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1312),
    .D(_00081_),
    .Q_N(_09134_),
    .Q(\mem.mem[73][6] ));
 sg13g2_dfrbp_1 _18439_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1311),
    .D(_00082_),
    .Q_N(_09133_),
    .Q(\mem.mem[73][7] ));
 sg13g2_dfrbp_1 _18440_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1310),
    .D(_00083_),
    .Q_N(_09132_),
    .Q(\mem.mem[72][0] ));
 sg13g2_dfrbp_1 _18441_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1309),
    .D(_00084_),
    .Q_N(_09131_),
    .Q(\mem.mem[72][1] ));
 sg13g2_dfrbp_1 _18442_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1308),
    .D(_00085_),
    .Q_N(_09130_),
    .Q(\mem.mem[72][2] ));
 sg13g2_dfrbp_1 _18443_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1307),
    .D(_00086_),
    .Q_N(_09129_),
    .Q(\mem.mem[72][3] ));
 sg13g2_dfrbp_1 _18444_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1306),
    .D(_00087_),
    .Q_N(_09128_),
    .Q(\mem.mem[72][4] ));
 sg13g2_dfrbp_1 _18445_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1305),
    .D(_00088_),
    .Q_N(_09127_),
    .Q(\mem.mem[72][5] ));
 sg13g2_dfrbp_1 _18446_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1304),
    .D(_00089_),
    .Q_N(_09126_),
    .Q(\mem.mem[72][6] ));
 sg13g2_dfrbp_1 _18447_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1303),
    .D(_00090_),
    .Q_N(_09125_),
    .Q(\mem.mem[72][7] ));
 sg13g2_dfrbp_1 _18448_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1302),
    .D(_00091_),
    .Q_N(_09124_),
    .Q(\mem.mem[87][0] ));
 sg13g2_dfrbp_1 _18449_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1301),
    .D(_00092_),
    .Q_N(_09123_),
    .Q(\mem.mem[87][1] ));
 sg13g2_dfrbp_1 _18450_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1300),
    .D(_00093_),
    .Q_N(_09122_),
    .Q(\mem.mem[87][2] ));
 sg13g2_dfrbp_1 _18451_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1299),
    .D(_00094_),
    .Q_N(_09121_),
    .Q(\mem.mem[87][3] ));
 sg13g2_dfrbp_1 _18452_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1298),
    .D(_00095_),
    .Q_N(_09120_),
    .Q(\mem.mem[87][4] ));
 sg13g2_dfrbp_1 _18453_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1297),
    .D(_00096_),
    .Q_N(_09119_),
    .Q(\mem.mem[87][5] ));
 sg13g2_dfrbp_1 _18454_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1296),
    .D(_00097_),
    .Q_N(_09118_),
    .Q(\mem.mem[87][6] ));
 sg13g2_dfrbp_1 _18455_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1295),
    .D(_00098_),
    .Q_N(_09117_),
    .Q(\mem.mem[87][7] ));
 sg13g2_dfrbp_1 _18456_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1294),
    .D(_00099_),
    .Q_N(_09116_),
    .Q(\mem.mem[71][0] ));
 sg13g2_dfrbp_1 _18457_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1293),
    .D(_00100_),
    .Q_N(_09115_),
    .Q(\mem.mem[71][1] ));
 sg13g2_dfrbp_1 _18458_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1292),
    .D(_00101_),
    .Q_N(_09114_),
    .Q(\mem.mem[71][2] ));
 sg13g2_dfrbp_1 _18459_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1291),
    .D(_00102_),
    .Q_N(_09113_),
    .Q(\mem.mem[71][3] ));
 sg13g2_dfrbp_1 _18460_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1290),
    .D(_00103_),
    .Q_N(_09112_),
    .Q(\mem.mem[71][4] ));
 sg13g2_dfrbp_1 _18461_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1289),
    .D(_00104_),
    .Q_N(_09111_),
    .Q(\mem.mem[71][5] ));
 sg13g2_dfrbp_1 _18462_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1288),
    .D(_00105_),
    .Q_N(_09110_),
    .Q(\mem.mem[71][6] ));
 sg13g2_dfrbp_1 _18463_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1287),
    .D(_00106_),
    .Q_N(_09109_),
    .Q(\mem.mem[71][7] ));
 sg13g2_dfrbp_1 _18464_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1286),
    .D(_00107_),
    .Q_N(_09108_),
    .Q(\mem.mem[86][0] ));
 sg13g2_dfrbp_1 _18465_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1285),
    .D(_00108_),
    .Q_N(_09107_),
    .Q(\mem.mem[86][1] ));
 sg13g2_dfrbp_1 _18466_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1284),
    .D(_00109_),
    .Q_N(_09106_),
    .Q(\mem.mem[86][2] ));
 sg13g2_dfrbp_1 _18467_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1283),
    .D(_00110_),
    .Q_N(_09105_),
    .Q(\mem.mem[86][3] ));
 sg13g2_dfrbp_1 _18468_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1282),
    .D(_00111_),
    .Q_N(_09104_),
    .Q(\mem.mem[86][4] ));
 sg13g2_dfrbp_1 _18469_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1281),
    .D(_00112_),
    .Q_N(_09103_),
    .Q(\mem.mem[86][5] ));
 sg13g2_dfrbp_1 _18470_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1280),
    .D(_00113_),
    .Q_N(_09102_),
    .Q(\mem.mem[86][6] ));
 sg13g2_dfrbp_1 _18471_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1279),
    .D(_00114_),
    .Q_N(_09101_),
    .Q(\mem.mem[86][7] ));
 sg13g2_dfrbp_1 _18472_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1278),
    .D(_00115_),
    .Q_N(_09100_),
    .Q(\mem.mem[2][0] ));
 sg13g2_dfrbp_1 _18473_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1277),
    .D(_00116_),
    .Q_N(_09099_),
    .Q(\mem.mem[2][1] ));
 sg13g2_dfrbp_1 _18474_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1276),
    .D(_00117_),
    .Q_N(_09098_),
    .Q(\mem.mem[2][2] ));
 sg13g2_dfrbp_1 _18475_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1275),
    .D(_00118_),
    .Q_N(_09097_),
    .Q(\mem.mem[2][3] ));
 sg13g2_dfrbp_1 _18476_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1274),
    .D(_00119_),
    .Q_N(_09096_),
    .Q(\mem.mem[2][4] ));
 sg13g2_dfrbp_1 _18477_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1273),
    .D(_00120_),
    .Q_N(_09095_),
    .Q(\mem.mem[2][5] ));
 sg13g2_dfrbp_1 _18478_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1272),
    .D(_00121_),
    .Q_N(_09094_),
    .Q(\mem.mem[2][6] ));
 sg13g2_dfrbp_1 _18479_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1271),
    .D(_00122_),
    .Q_N(_09093_),
    .Q(\mem.mem[2][7] ));
 sg13g2_dfrbp_1 _18480_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1270),
    .D(_00123_),
    .Q_N(_09092_),
    .Q(\mem.mem[70][0] ));
 sg13g2_dfrbp_1 _18481_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1269),
    .D(_00124_),
    .Q_N(_09091_),
    .Q(\mem.mem[70][1] ));
 sg13g2_dfrbp_1 _18482_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1268),
    .D(_00125_),
    .Q_N(_09090_),
    .Q(\mem.mem[70][2] ));
 sg13g2_dfrbp_1 _18483_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1267),
    .D(_00126_),
    .Q_N(_09089_),
    .Q(\mem.mem[70][3] ));
 sg13g2_dfrbp_1 _18484_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1266),
    .D(_00127_),
    .Q_N(_09088_),
    .Q(\mem.mem[70][4] ));
 sg13g2_dfrbp_1 _18485_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1265),
    .D(_00128_),
    .Q_N(_09087_),
    .Q(\mem.mem[70][5] ));
 sg13g2_dfrbp_1 _18486_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1264),
    .D(_00129_),
    .Q_N(_09086_),
    .Q(\mem.mem[70][6] ));
 sg13g2_dfrbp_1 _18487_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1263),
    .D(_00130_),
    .Q_N(_09085_),
    .Q(\mem.mem[70][7] ));
 sg13g2_dfrbp_1 _18488_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1262),
    .D(_00131_),
    .Q_N(_09084_),
    .Q(\mem.mem[6][0] ));
 sg13g2_dfrbp_1 _18489_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1261),
    .D(_00132_),
    .Q_N(_09083_),
    .Q(\mem.mem[6][1] ));
 sg13g2_dfrbp_1 _18490_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1260),
    .D(_00133_),
    .Q_N(_09082_),
    .Q(\mem.mem[6][2] ));
 sg13g2_dfrbp_1 _18491_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1259),
    .D(_00134_),
    .Q_N(_09081_),
    .Q(\mem.mem[6][3] ));
 sg13g2_dfrbp_1 _18492_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1258),
    .D(_00135_),
    .Q_N(_09080_),
    .Q(\mem.mem[6][4] ));
 sg13g2_dfrbp_1 _18493_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1257),
    .D(_00136_),
    .Q_N(_09079_),
    .Q(\mem.mem[6][5] ));
 sg13g2_dfrbp_1 _18494_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1256),
    .D(_00137_),
    .Q_N(_09078_),
    .Q(\mem.mem[6][6] ));
 sg13g2_dfrbp_1 _18495_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1255),
    .D(_00138_),
    .Q_N(_09077_),
    .Q(\mem.mem[6][7] ));
 sg13g2_dfrbp_1 _18496_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1254),
    .D(_00139_),
    .Q_N(_09076_),
    .Q(\mem.mem[68][0] ));
 sg13g2_dfrbp_1 _18497_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1253),
    .D(_00140_),
    .Q_N(_09075_),
    .Q(\mem.mem[68][1] ));
 sg13g2_dfrbp_1 _18498_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1252),
    .D(_00141_),
    .Q_N(_09074_),
    .Q(\mem.mem[68][2] ));
 sg13g2_dfrbp_1 _18499_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1251),
    .D(_00142_),
    .Q_N(_09073_),
    .Q(\mem.mem[68][3] ));
 sg13g2_dfrbp_1 _18500_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1250),
    .D(_00143_),
    .Q_N(_09072_),
    .Q(\mem.mem[68][4] ));
 sg13g2_dfrbp_1 _18501_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1249),
    .D(_00144_),
    .Q_N(_09071_),
    .Q(\mem.mem[68][5] ));
 sg13g2_dfrbp_1 _18502_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1248),
    .D(_00145_),
    .Q_N(_09070_),
    .Q(\mem.mem[68][6] ));
 sg13g2_dfrbp_1 _18503_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1247),
    .D(_00146_),
    .Q_N(_09069_),
    .Q(\mem.mem[68][7] ));
 sg13g2_dfrbp_1 _18504_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1246),
    .D(_00147_),
    .Q_N(_09068_),
    .Q(\mem.mem[67][0] ));
 sg13g2_dfrbp_1 _18505_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1245),
    .D(_00148_),
    .Q_N(_09067_),
    .Q(\mem.mem[67][1] ));
 sg13g2_dfrbp_1 _18506_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1244),
    .D(_00149_),
    .Q_N(_09066_),
    .Q(\mem.mem[67][2] ));
 sg13g2_dfrbp_1 _18507_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1243),
    .D(_00150_),
    .Q_N(_09065_),
    .Q(\mem.mem[67][3] ));
 sg13g2_dfrbp_1 _18508_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1242),
    .D(_00151_),
    .Q_N(_09064_),
    .Q(\mem.mem[67][4] ));
 sg13g2_dfrbp_1 _18509_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1241),
    .D(_00152_),
    .Q_N(_09063_),
    .Q(\mem.mem[67][5] ));
 sg13g2_dfrbp_1 _18510_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1240),
    .D(_00153_),
    .Q_N(_09062_),
    .Q(\mem.mem[67][6] ));
 sg13g2_dfrbp_1 _18511_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1239),
    .D(_00154_),
    .Q_N(_09061_),
    .Q(\mem.mem[67][7] ));
 sg13g2_dfrbp_1 _18512_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1238),
    .D(_00155_),
    .Q_N(_09060_),
    .Q(\mem.mem[66][0] ));
 sg13g2_dfrbp_1 _18513_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1237),
    .D(_00156_),
    .Q_N(_09059_),
    .Q(\mem.mem[66][1] ));
 sg13g2_dfrbp_1 _18514_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1236),
    .D(_00157_),
    .Q_N(_09058_),
    .Q(\mem.mem[66][2] ));
 sg13g2_dfrbp_1 _18515_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1235),
    .D(_00158_),
    .Q_N(_09057_),
    .Q(\mem.mem[66][3] ));
 sg13g2_dfrbp_1 _18516_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1234),
    .D(_00159_),
    .Q_N(_09056_),
    .Q(\mem.mem[66][4] ));
 sg13g2_dfrbp_1 _18517_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1233),
    .D(_00160_),
    .Q_N(_09055_),
    .Q(\mem.mem[66][5] ));
 sg13g2_dfrbp_1 _18518_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1232),
    .D(_00161_),
    .Q_N(_09054_),
    .Q(\mem.mem[66][6] ));
 sg13g2_dfrbp_1 _18519_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1231),
    .D(_00162_),
    .Q_N(_09053_),
    .Q(\mem.mem[66][7] ));
 sg13g2_dfrbp_1 _18520_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1230),
    .D(_00163_),
    .Q_N(_09052_),
    .Q(\mem.mem[65][0] ));
 sg13g2_dfrbp_1 _18521_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1229),
    .D(_00164_),
    .Q_N(_09051_),
    .Q(\mem.mem[65][1] ));
 sg13g2_dfrbp_1 _18522_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1228),
    .D(_00165_),
    .Q_N(_09050_),
    .Q(\mem.mem[65][2] ));
 sg13g2_dfrbp_1 _18523_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1227),
    .D(_00166_),
    .Q_N(_09049_),
    .Q(\mem.mem[65][3] ));
 sg13g2_dfrbp_1 _18524_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1226),
    .D(_00167_),
    .Q_N(_09048_),
    .Q(\mem.mem[65][4] ));
 sg13g2_dfrbp_1 _18525_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1225),
    .D(_00168_),
    .Q_N(_09047_),
    .Q(\mem.mem[65][5] ));
 sg13g2_dfrbp_1 _18526_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1224),
    .D(_00169_),
    .Q_N(_09046_),
    .Q(\mem.mem[65][6] ));
 sg13g2_dfrbp_1 _18527_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1223),
    .D(_00170_),
    .Q_N(_09045_),
    .Q(\mem.mem[65][7] ));
 sg13g2_dfrbp_1 _18528_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1222),
    .D(_00171_),
    .Q_N(_09044_),
    .Q(\mem.mem[40][0] ));
 sg13g2_dfrbp_1 _18529_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1221),
    .D(_00172_),
    .Q_N(_09043_),
    .Q(\mem.mem[40][1] ));
 sg13g2_dfrbp_1 _18530_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1220),
    .D(_00173_),
    .Q_N(_09042_),
    .Q(\mem.mem[40][2] ));
 sg13g2_dfrbp_1 _18531_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1219),
    .D(_00174_),
    .Q_N(_09041_),
    .Q(\mem.mem[40][3] ));
 sg13g2_dfrbp_1 _18532_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1218),
    .D(_00175_),
    .Q_N(_09040_),
    .Q(\mem.mem[40][4] ));
 sg13g2_dfrbp_1 _18533_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1217),
    .D(_00176_),
    .Q_N(_09039_),
    .Q(\mem.mem[40][5] ));
 sg13g2_dfrbp_1 _18534_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1216),
    .D(_00177_),
    .Q_N(_09038_),
    .Q(\mem.mem[40][6] ));
 sg13g2_dfrbp_1 _18535_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1215),
    .D(_00178_),
    .Q_N(_09037_),
    .Q(\mem.mem[40][7] ));
 sg13g2_dfrbp_1 _18536_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1214),
    .D(_00179_),
    .Q_N(_09036_),
    .Q(\mem.mem[129][0] ));
 sg13g2_dfrbp_1 _18537_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1213),
    .D(_00180_),
    .Q_N(_09035_),
    .Q(\mem.mem[129][1] ));
 sg13g2_dfrbp_1 _18538_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1212),
    .D(_00181_),
    .Q_N(_09034_),
    .Q(\mem.mem[129][2] ));
 sg13g2_dfrbp_1 _18539_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1211),
    .D(_00182_),
    .Q_N(_09033_),
    .Q(\mem.mem[129][3] ));
 sg13g2_dfrbp_1 _18540_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1210),
    .D(_00183_),
    .Q_N(_09032_),
    .Q(\mem.mem[129][4] ));
 sg13g2_dfrbp_1 _18541_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1209),
    .D(_00184_),
    .Q_N(_09031_),
    .Q(\mem.mem[129][5] ));
 sg13g2_dfrbp_1 _18542_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1208),
    .D(_00185_),
    .Q_N(_09030_),
    .Q(\mem.mem[129][6] ));
 sg13g2_dfrbp_1 _18543_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1207),
    .D(_00186_),
    .Q_N(_09029_),
    .Q(\mem.mem[129][7] ));
 sg13g2_dfrbp_1 _18544_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1206),
    .D(_00187_),
    .Q_N(_09028_),
    .Q(\mem.mem[3][0] ));
 sg13g2_dfrbp_1 _18545_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1205),
    .D(_00188_),
    .Q_N(_09027_),
    .Q(\mem.mem[3][1] ));
 sg13g2_dfrbp_1 _18546_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1204),
    .D(_00189_),
    .Q_N(_09026_),
    .Q(\mem.mem[3][2] ));
 sg13g2_dfrbp_1 _18547_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1203),
    .D(_00190_),
    .Q_N(_09025_),
    .Q(\mem.mem[3][3] ));
 sg13g2_dfrbp_1 _18548_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1202),
    .D(_00191_),
    .Q_N(_09024_),
    .Q(\mem.mem[3][4] ));
 sg13g2_dfrbp_1 _18549_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1201),
    .D(_00192_),
    .Q_N(_09023_),
    .Q(\mem.mem[3][5] ));
 sg13g2_dfrbp_1 _18550_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1200),
    .D(_00193_),
    .Q_N(_09022_),
    .Q(\mem.mem[3][6] ));
 sg13g2_dfrbp_1 _18551_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1199),
    .D(_00194_),
    .Q_N(_09021_),
    .Q(\mem.mem[3][7] ));
 sg13g2_dfrbp_1 _18552_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1198),
    .D(_00195_),
    .Q_N(_09020_),
    .Q(\mem.mem[59][0] ));
 sg13g2_dfrbp_1 _18553_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1197),
    .D(_00196_),
    .Q_N(_09019_),
    .Q(\mem.mem[59][1] ));
 sg13g2_dfrbp_1 _18554_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1196),
    .D(_00197_),
    .Q_N(_09018_),
    .Q(\mem.mem[59][2] ));
 sg13g2_dfrbp_1 _18555_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1195),
    .D(_00198_),
    .Q_N(_09017_),
    .Q(\mem.mem[59][3] ));
 sg13g2_dfrbp_1 _18556_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1194),
    .D(_00199_),
    .Q_N(_09016_),
    .Q(\mem.mem[59][4] ));
 sg13g2_dfrbp_1 _18557_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1193),
    .D(_00200_),
    .Q_N(_09015_),
    .Q(\mem.mem[59][5] ));
 sg13g2_dfrbp_1 _18558_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1192),
    .D(_00201_),
    .Q_N(_09014_),
    .Q(\mem.mem[59][6] ));
 sg13g2_dfrbp_1 _18559_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1191),
    .D(_00202_),
    .Q_N(_09013_),
    .Q(\mem.mem[59][7] ));
 sg13g2_dfrbp_1 _18560_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1190),
    .D(_00203_),
    .Q_N(_09012_),
    .Q(\mem.mem[38][0] ));
 sg13g2_dfrbp_1 _18561_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1189),
    .D(_00204_),
    .Q_N(_09011_),
    .Q(\mem.mem[38][1] ));
 sg13g2_dfrbp_1 _18562_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1188),
    .D(_00205_),
    .Q_N(_09010_),
    .Q(\mem.mem[38][2] ));
 sg13g2_dfrbp_1 _18563_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1187),
    .D(_00206_),
    .Q_N(_09009_),
    .Q(\mem.mem[38][3] ));
 sg13g2_dfrbp_1 _18564_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1186),
    .D(_00207_),
    .Q_N(_09008_),
    .Q(\mem.mem[38][4] ));
 sg13g2_dfrbp_1 _18565_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1185),
    .D(_00208_),
    .Q_N(_09007_),
    .Q(\mem.mem[38][5] ));
 sg13g2_dfrbp_1 _18566_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1184),
    .D(_00209_),
    .Q_N(_09006_),
    .Q(\mem.mem[38][6] ));
 sg13g2_dfrbp_1 _18567_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1183),
    .D(_00210_),
    .Q_N(_09005_),
    .Q(\mem.mem[38][7] ));
 sg13g2_dfrbp_1 _18568_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1182),
    .D(_00211_),
    .Q_N(_09004_),
    .Q(\mem.mem[37][0] ));
 sg13g2_dfrbp_1 _18569_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1181),
    .D(_00212_),
    .Q_N(_09003_),
    .Q(\mem.mem[37][1] ));
 sg13g2_dfrbp_1 _18570_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1180),
    .D(_00213_),
    .Q_N(_09002_),
    .Q(\mem.mem[37][2] ));
 sg13g2_dfrbp_1 _18571_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1179),
    .D(_00214_),
    .Q_N(_09001_),
    .Q(\mem.mem[37][3] ));
 sg13g2_dfrbp_1 _18572_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1178),
    .D(_00215_),
    .Q_N(_09000_),
    .Q(\mem.mem[37][4] ));
 sg13g2_dfrbp_1 _18573_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1177),
    .D(_00216_),
    .Q_N(_08999_),
    .Q(\mem.mem[37][5] ));
 sg13g2_dfrbp_1 _18574_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1176),
    .D(_00217_),
    .Q_N(_08998_),
    .Q(\mem.mem[37][6] ));
 sg13g2_dfrbp_1 _18575_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1175),
    .D(_00218_),
    .Q_N(_08997_),
    .Q(\mem.mem[37][7] ));
 sg13g2_dfrbp_1 _18576_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1174),
    .D(_00219_),
    .Q_N(_08996_),
    .Q(\mem.mem[109][0] ));
 sg13g2_dfrbp_1 _18577_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1173),
    .D(_00220_),
    .Q_N(_08995_),
    .Q(\mem.mem[109][1] ));
 sg13g2_dfrbp_1 _18578_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1172),
    .D(_00221_),
    .Q_N(_08994_),
    .Q(\mem.mem[109][2] ));
 sg13g2_dfrbp_1 _18579_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1171),
    .D(_00222_),
    .Q_N(_08993_),
    .Q(\mem.mem[109][3] ));
 sg13g2_dfrbp_1 _18580_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1170),
    .D(_00223_),
    .Q_N(_08992_),
    .Q(\mem.mem[109][4] ));
 sg13g2_dfrbp_1 _18581_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1169),
    .D(_00224_),
    .Q_N(_08991_),
    .Q(\mem.mem[109][5] ));
 sg13g2_dfrbp_1 _18582_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1168),
    .D(_00225_),
    .Q_N(_08990_),
    .Q(\mem.mem[109][6] ));
 sg13g2_dfrbp_1 _18583_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1167),
    .D(_00226_),
    .Q_N(_08989_),
    .Q(\mem.mem[109][7] ));
 sg13g2_dfrbp_1 _18584_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1166),
    .D(_00227_),
    .Q_N(_08988_),
    .Q(\mem.mem[119][0] ));
 sg13g2_dfrbp_1 _18585_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1165),
    .D(_00228_),
    .Q_N(_08987_),
    .Q(\mem.mem[119][1] ));
 sg13g2_dfrbp_1 _18586_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1164),
    .D(_00229_),
    .Q_N(_08986_),
    .Q(\mem.mem[119][2] ));
 sg13g2_dfrbp_1 _18587_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1163),
    .D(_00230_),
    .Q_N(_08985_),
    .Q(\mem.mem[119][3] ));
 sg13g2_dfrbp_1 _18588_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1162),
    .D(_00231_),
    .Q_N(_08984_),
    .Q(\mem.mem[119][4] ));
 sg13g2_dfrbp_1 _18589_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1161),
    .D(_00232_),
    .Q_N(_08983_),
    .Q(\mem.mem[119][5] ));
 sg13g2_dfrbp_1 _18590_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1160),
    .D(_00233_),
    .Q_N(_08982_),
    .Q(\mem.mem[119][6] ));
 sg13g2_dfrbp_1 _18591_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1159),
    .D(_00234_),
    .Q_N(_08981_),
    .Q(\mem.mem[119][7] ));
 sg13g2_dfrbp_1 _18592_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1158),
    .D(_00235_),
    .Q_N(_08980_),
    .Q(\mem.mem[36][0] ));
 sg13g2_dfrbp_1 _18593_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1157),
    .D(_00236_),
    .Q_N(_08979_),
    .Q(\mem.mem[36][1] ));
 sg13g2_dfrbp_1 _18594_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1156),
    .D(_00237_),
    .Q_N(_08978_),
    .Q(\mem.mem[36][2] ));
 sg13g2_dfrbp_1 _18595_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1155),
    .D(_00238_),
    .Q_N(_08977_),
    .Q(\mem.mem[36][3] ));
 sg13g2_dfrbp_1 _18596_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1154),
    .D(_00239_),
    .Q_N(_08976_),
    .Q(\mem.mem[36][4] ));
 sg13g2_dfrbp_1 _18597_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1153),
    .D(_00240_),
    .Q_N(_08975_),
    .Q(\mem.mem[36][5] ));
 sg13g2_dfrbp_1 _18598_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1152),
    .D(_00241_),
    .Q_N(_08974_),
    .Q(\mem.mem[36][6] ));
 sg13g2_dfrbp_1 _18599_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1151),
    .D(_00242_),
    .Q_N(_08973_),
    .Q(\mem.mem[36][7] ));
 sg13g2_dfrbp_1 _18600_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1150),
    .D(_00243_),
    .Q_N(_08972_),
    .Q(\mem.mem[69][0] ));
 sg13g2_dfrbp_1 _18601_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1149),
    .D(_00244_),
    .Q_N(_08971_),
    .Q(\mem.mem[69][1] ));
 sg13g2_dfrbp_1 _18602_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1148),
    .D(_00245_),
    .Q_N(_08970_),
    .Q(\mem.mem[69][2] ));
 sg13g2_dfrbp_1 _18603_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1147),
    .D(_00246_),
    .Q_N(_08969_),
    .Q(\mem.mem[69][3] ));
 sg13g2_dfrbp_1 _18604_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1146),
    .D(_00247_),
    .Q_N(_08968_),
    .Q(\mem.mem[69][4] ));
 sg13g2_dfrbp_1 _18605_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1145),
    .D(_00248_),
    .Q_N(_08967_),
    .Q(\mem.mem[69][5] ));
 sg13g2_dfrbp_1 _18606_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1144),
    .D(_00249_),
    .Q_N(_08966_),
    .Q(\mem.mem[69][6] ));
 sg13g2_dfrbp_1 _18607_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1143),
    .D(_00250_),
    .Q_N(_08965_),
    .Q(\mem.mem[69][7] ));
 sg13g2_dfrbp_1 _18608_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1142),
    .D(_00251_),
    .Q_N(_08964_),
    .Q(\mem.mem[99][0] ));
 sg13g2_dfrbp_1 _18609_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1141),
    .D(_00252_),
    .Q_N(_08963_),
    .Q(\mem.mem[99][1] ));
 sg13g2_dfrbp_1 _18610_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1140),
    .D(_00253_),
    .Q_N(_08962_),
    .Q(\mem.mem[99][2] ));
 sg13g2_dfrbp_1 _18611_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1139),
    .D(_00254_),
    .Q_N(_08961_),
    .Q(\mem.mem[99][3] ));
 sg13g2_dfrbp_1 _18612_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1138),
    .D(_00255_),
    .Q_N(_08960_),
    .Q(\mem.mem[99][4] ));
 sg13g2_dfrbp_1 _18613_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1137),
    .D(_00256_),
    .Q_N(_08959_),
    .Q(\mem.mem[99][5] ));
 sg13g2_dfrbp_1 _18614_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1136),
    .D(_00257_),
    .Q_N(_08958_),
    .Q(\mem.mem[99][6] ));
 sg13g2_dfrbp_1 _18615_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1135),
    .D(_00258_),
    .Q_N(_08957_),
    .Q(\mem.mem[99][7] ));
 sg13g2_dfrbp_1 _18616_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1134),
    .D(_00259_),
    .Q_N(_08956_),
    .Q(\mem.mem[35][0] ));
 sg13g2_dfrbp_1 _18617_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1133),
    .D(_00260_),
    .Q_N(_08955_),
    .Q(\mem.mem[35][1] ));
 sg13g2_dfrbp_1 _18618_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1132),
    .D(_00261_),
    .Q_N(_08954_),
    .Q(\mem.mem[35][2] ));
 sg13g2_dfrbp_1 _18619_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1131),
    .D(_00262_),
    .Q_N(_08953_),
    .Q(\mem.mem[35][3] ));
 sg13g2_dfrbp_1 _18620_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1130),
    .D(_00263_),
    .Q_N(_08952_),
    .Q(\mem.mem[35][4] ));
 sg13g2_dfrbp_1 _18621_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1129),
    .D(_00264_),
    .Q_N(_08951_),
    .Q(\mem.mem[35][5] ));
 sg13g2_dfrbp_1 _18622_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1128),
    .D(_00265_),
    .Q_N(_08950_),
    .Q(\mem.mem[35][6] ));
 sg13g2_dfrbp_1 _18623_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1127),
    .D(_00266_),
    .Q_N(_08949_),
    .Q(\mem.mem[35][7] ));
 sg13g2_dfrbp_1 _18624_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1126),
    .D(_00267_),
    .Q_N(_08948_),
    .Q(prev_run));
 sg13g2_dfrbp_1 _18625_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1125),
    .D(_00268_),
    .Q_N(_08947_),
    .Q(\mem.mem[34][0] ));
 sg13g2_dfrbp_1 _18626_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1124),
    .D(_00269_),
    .Q_N(_08946_),
    .Q(\mem.mem[34][1] ));
 sg13g2_dfrbp_1 _18627_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1123),
    .D(_00270_),
    .Q_N(_08945_),
    .Q(\mem.mem[34][2] ));
 sg13g2_dfrbp_1 _18628_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1122),
    .D(_00271_),
    .Q_N(_08944_),
    .Q(\mem.mem[34][3] ));
 sg13g2_dfrbp_1 _18629_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1121),
    .D(_00272_),
    .Q_N(_08943_),
    .Q(\mem.mem[34][4] ));
 sg13g2_dfrbp_1 _18630_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1120),
    .D(_00273_),
    .Q_N(_08942_),
    .Q(\mem.mem[34][5] ));
 sg13g2_dfrbp_1 _18631_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1119),
    .D(_00274_),
    .Q_N(_08941_),
    .Q(\mem.mem[34][6] ));
 sg13g2_dfrbp_1 _18632_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1118),
    .D(_00275_),
    .Q_N(_08940_),
    .Q(\mem.mem[34][7] ));
 sg13g2_dfrbp_1 _18633_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1117),
    .D(_00276_),
    .Q_N(_08939_),
    .Q(\mem.mem[149][0] ));
 sg13g2_dfrbp_1 _18634_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1116),
    .D(_00277_),
    .Q_N(_08938_),
    .Q(\mem.mem[149][1] ));
 sg13g2_dfrbp_1 _18635_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1115),
    .D(_00278_),
    .Q_N(_08937_),
    .Q(\mem.mem[149][2] ));
 sg13g2_dfrbp_1 _18636_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1114),
    .D(_00279_),
    .Q_N(_08936_),
    .Q(\mem.mem[149][3] ));
 sg13g2_dfrbp_1 _18637_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1113),
    .D(_00280_),
    .Q_N(_08935_),
    .Q(\mem.mem[149][4] ));
 sg13g2_dfrbp_1 _18638_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1112),
    .D(_00281_),
    .Q_N(_08934_),
    .Q(\mem.mem[149][5] ));
 sg13g2_dfrbp_1 _18639_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1111),
    .D(_00282_),
    .Q_N(_08933_),
    .Q(\mem.mem[149][6] ));
 sg13g2_dfrbp_1 _18640_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1110),
    .D(_00283_),
    .Q_N(_08932_),
    .Q(\mem.mem[149][7] ));
 sg13g2_dfrbp_1 _18641_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1109),
    .D(_00284_),
    .Q_N(_08931_),
    .Q(_00000_));
 sg13g2_dfrbp_1 _18642_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1108),
    .D(_00285_),
    .Q_N(_08930_),
    .Q(_00001_));
 sg13g2_dfrbp_1 _18643_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1107),
    .D(_00286_),
    .Q_N(_08929_),
    .Q(_00002_));
 sg13g2_dfrbp_1 _18644_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1106),
    .D(_00287_),
    .Q_N(_08928_),
    .Q(_00003_));
 sg13g2_dfrbp_1 _18645_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1105),
    .D(_00288_),
    .Q_N(_08927_),
    .Q(_00004_));
 sg13g2_dfrbp_1 _18646_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1104),
    .D(_00289_),
    .Q_N(_08926_),
    .Q(_00005_));
 sg13g2_dfrbp_1 _18647_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1103),
    .D(_00290_),
    .Q_N(_08925_),
    .Q(_00006_));
 sg13g2_dfrbp_1 _18648_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1102),
    .D(_00291_),
    .Q_N(_08924_),
    .Q(_00007_));
 sg13g2_dfrbp_1 _18649_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1101),
    .D(_00292_),
    .Q_N(_08923_),
    .Q(\mem.mem[33][0] ));
 sg13g2_dfrbp_1 _18650_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1100),
    .D(_00293_),
    .Q_N(_08922_),
    .Q(\mem.mem[33][1] ));
 sg13g2_dfrbp_1 _18651_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1099),
    .D(_00294_),
    .Q_N(_08921_),
    .Q(\mem.mem[33][2] ));
 sg13g2_dfrbp_1 _18652_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1098),
    .D(_00295_),
    .Q_N(_08920_),
    .Q(\mem.mem[33][3] ));
 sg13g2_dfrbp_1 _18653_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1097),
    .D(_00296_),
    .Q_N(_08919_),
    .Q(\mem.mem[33][4] ));
 sg13g2_dfrbp_1 _18654_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1096),
    .D(_00297_),
    .Q_N(_08918_),
    .Q(\mem.mem[33][5] ));
 sg13g2_dfrbp_1 _18655_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1095),
    .D(_00298_),
    .Q_N(_08917_),
    .Q(\mem.mem[33][6] ));
 sg13g2_dfrbp_1 _18656_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1094),
    .D(_00299_),
    .Q_N(_08916_),
    .Q(\mem.mem[33][7] ));
 sg13g2_dfrbp_1 _18657_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1093),
    .D(_00300_),
    .Q_N(_08915_),
    .Q(\mem.mem[32][0] ));
 sg13g2_dfrbp_1 _18658_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1092),
    .D(_00301_),
    .Q_N(_08914_),
    .Q(\mem.mem[32][1] ));
 sg13g2_dfrbp_1 _18659_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1091),
    .D(_00302_),
    .Q_N(_08913_),
    .Q(\mem.mem[32][2] ));
 sg13g2_dfrbp_1 _18660_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1090),
    .D(_00303_),
    .Q_N(_08912_),
    .Q(\mem.mem[32][3] ));
 sg13g2_dfrbp_1 _18661_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1089),
    .D(_00304_),
    .Q_N(_08911_),
    .Q(\mem.mem[32][4] ));
 sg13g2_dfrbp_1 _18662_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1088),
    .D(_00305_),
    .Q_N(_08910_),
    .Q(\mem.mem[32][5] ));
 sg13g2_dfrbp_1 _18663_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1087),
    .D(_00306_),
    .Q_N(_08909_),
    .Q(\mem.mem[32][6] ));
 sg13g2_dfrbp_1 _18664_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1086),
    .D(_00307_),
    .Q_N(_08908_),
    .Q(\mem.mem[32][7] ));
 sg13g2_dfrbp_1 _18665_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1085),
    .D(_00308_),
    .Q_N(_08907_),
    .Q(\mem.mem[31][0] ));
 sg13g2_dfrbp_1 _18666_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1084),
    .D(_00309_),
    .Q_N(_08906_),
    .Q(\mem.mem[31][1] ));
 sg13g2_dfrbp_1 _18667_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1083),
    .D(_00310_),
    .Q_N(_08905_),
    .Q(\mem.mem[31][2] ));
 sg13g2_dfrbp_1 _18668_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1082),
    .D(_00311_),
    .Q_N(_08904_),
    .Q(\mem.mem[31][3] ));
 sg13g2_dfrbp_1 _18669_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1081),
    .D(_00312_),
    .Q_N(_08903_),
    .Q(\mem.mem[31][4] ));
 sg13g2_dfrbp_1 _18670_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1080),
    .D(_00313_),
    .Q_N(_08902_),
    .Q(\mem.mem[31][5] ));
 sg13g2_dfrbp_1 _18671_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1079),
    .D(_00314_),
    .Q_N(_08901_),
    .Q(\mem.mem[31][6] ));
 sg13g2_dfrbp_1 _18672_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1078),
    .D(_00315_),
    .Q_N(_08900_),
    .Q(\mem.mem[31][7] ));
 sg13g2_dfrbp_1 _18673_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1077),
    .D(_00316_),
    .Q_N(_08899_),
    .Q(\mem.mem[46][0] ));
 sg13g2_dfrbp_1 _18674_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1076),
    .D(_00317_),
    .Q_N(_08898_),
    .Q(\mem.mem[46][1] ));
 sg13g2_dfrbp_1 _18675_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1075),
    .D(_00318_),
    .Q_N(_08897_),
    .Q(\mem.mem[46][2] ));
 sg13g2_dfrbp_1 _18676_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1074),
    .D(_00319_),
    .Q_N(_08896_),
    .Q(\mem.mem[46][3] ));
 sg13g2_dfrbp_1 _18677_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1073),
    .D(_00320_),
    .Q_N(_08895_),
    .Q(\mem.mem[46][4] ));
 sg13g2_dfrbp_1 _18678_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1072),
    .D(_00321_),
    .Q_N(_08894_),
    .Q(\mem.mem[46][5] ));
 sg13g2_dfrbp_1 _18679_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1071),
    .D(_00322_),
    .Q_N(_08893_),
    .Q(\mem.mem[46][6] ));
 sg13g2_dfrbp_1 _18680_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1070),
    .D(_00323_),
    .Q_N(_08892_),
    .Q(\mem.mem[46][7] ));
 sg13g2_dfrbp_1 _18681_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1069),
    .D(_00324_),
    .Q_N(_08891_),
    .Q(\mem.mem[30][0] ));
 sg13g2_dfrbp_1 _18682_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1068),
    .D(_00325_),
    .Q_N(_08890_),
    .Q(\mem.mem[30][1] ));
 sg13g2_dfrbp_1 _18683_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1067),
    .D(_00326_),
    .Q_N(_08889_),
    .Q(\mem.mem[30][2] ));
 sg13g2_dfrbp_1 _18684_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1066),
    .D(_00327_),
    .Q_N(_08888_),
    .Q(\mem.mem[30][3] ));
 sg13g2_dfrbp_1 _18685_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1065),
    .D(_00328_),
    .Q_N(_08887_),
    .Q(\mem.mem[30][4] ));
 sg13g2_dfrbp_1 _18686_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1064),
    .D(_00329_),
    .Q_N(_08886_),
    .Q(\mem.mem[30][5] ));
 sg13g2_dfrbp_1 _18687_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1063),
    .D(_00330_),
    .Q_N(_08885_),
    .Q(\mem.mem[30][6] ));
 sg13g2_dfrbp_1 _18688_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1062),
    .D(_00331_),
    .Q_N(_08884_),
    .Q(\mem.mem[30][7] ));
 sg13g2_dfrbp_1 _18689_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1061),
    .D(_00332_),
    .Q_N(_08883_),
    .Q(\mem.mem[45][0] ));
 sg13g2_dfrbp_1 _18690_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1060),
    .D(_00333_),
    .Q_N(_08882_),
    .Q(\mem.mem[45][1] ));
 sg13g2_dfrbp_1 _18691_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1059),
    .D(_00334_),
    .Q_N(_08881_),
    .Q(\mem.mem[45][2] ));
 sg13g2_dfrbp_1 _18692_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1058),
    .D(_00335_),
    .Q_N(_08880_),
    .Q(\mem.mem[45][3] ));
 sg13g2_dfrbp_1 _18693_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1057),
    .D(_00336_),
    .Q_N(_08879_),
    .Q(\mem.mem[45][4] ));
 sg13g2_dfrbp_1 _18694_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1056),
    .D(_00337_),
    .Q_N(_08878_),
    .Q(\mem.mem[45][5] ));
 sg13g2_dfrbp_1 _18695_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1055),
    .D(_00338_),
    .Q_N(_08877_),
    .Q(\mem.mem[45][6] ));
 sg13g2_dfrbp_1 _18696_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1054),
    .D(_00339_),
    .Q_N(_08876_),
    .Q(\mem.mem[45][7] ));
 sg13g2_dfrbp_1 _18697_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1053),
    .D(_00340_),
    .Q_N(_08875_),
    .Q(\mem.mem[85][0] ));
 sg13g2_dfrbp_1 _18698_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1052),
    .D(_00341_),
    .Q_N(_08874_),
    .Q(\mem.mem[85][1] ));
 sg13g2_dfrbp_1 _18699_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1051),
    .D(_00342_),
    .Q_N(_08873_),
    .Q(\mem.mem[85][2] ));
 sg13g2_dfrbp_1 _18700_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1050),
    .D(_00343_),
    .Q_N(_08872_),
    .Q(\mem.mem[85][3] ));
 sg13g2_dfrbp_1 _18701_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1049),
    .D(_00344_),
    .Q_N(_08871_),
    .Q(\mem.mem[85][4] ));
 sg13g2_dfrbp_1 _18702_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1048),
    .D(_00345_),
    .Q_N(_08870_),
    .Q(\mem.mem[85][5] ));
 sg13g2_dfrbp_1 _18703_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1047),
    .D(_00346_),
    .Q_N(_08869_),
    .Q(\mem.mem[85][6] ));
 sg13g2_dfrbp_1 _18704_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1046),
    .D(_00347_),
    .Q_N(_08868_),
    .Q(\mem.mem[85][7] ));
 sg13g2_dfrbp_1 _18705_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1045),
    .D(_00348_),
    .Q_N(_08867_),
    .Q(\mem.mem[64][0] ));
 sg13g2_dfrbp_1 _18706_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1044),
    .D(_00349_),
    .Q_N(_08866_),
    .Q(\mem.mem[64][1] ));
 sg13g2_dfrbp_1 _18707_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1043),
    .D(_00350_),
    .Q_N(_08865_),
    .Q(\mem.mem[64][2] ));
 sg13g2_dfrbp_1 _18708_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1042),
    .D(_00351_),
    .Q_N(_08864_),
    .Q(\mem.mem[64][3] ));
 sg13g2_dfrbp_1 _18709_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1041),
    .D(_00352_),
    .Q_N(_08863_),
    .Q(\mem.mem[64][4] ));
 sg13g2_dfrbp_1 _18710_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1040),
    .D(_00353_),
    .Q_N(_08862_),
    .Q(\mem.mem[64][5] ));
 sg13g2_dfrbp_1 _18711_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1039),
    .D(_00354_),
    .Q_N(_08861_),
    .Q(\mem.mem[64][6] ));
 sg13g2_dfrbp_1 _18712_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1038),
    .D(_00355_),
    .Q_N(_08860_),
    .Q(\mem.mem[64][7] ));
 sg13g2_dfrbp_1 _18713_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1037),
    .D(_00356_),
    .Q_N(_08859_),
    .Q(\mem.mem[63][0] ));
 sg13g2_dfrbp_1 _18714_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1036),
    .D(_00357_),
    .Q_N(_08858_),
    .Q(\mem.mem[63][1] ));
 sg13g2_dfrbp_1 _18715_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1035),
    .D(_00358_),
    .Q_N(_08857_),
    .Q(\mem.mem[63][2] ));
 sg13g2_dfrbp_1 _18716_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1034),
    .D(_00359_),
    .Q_N(_08856_),
    .Q(\mem.mem[63][3] ));
 sg13g2_dfrbp_1 _18717_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1033),
    .D(_00360_),
    .Q_N(_08855_),
    .Q(\mem.mem[63][4] ));
 sg13g2_dfrbp_1 _18718_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1032),
    .D(_00361_),
    .Q_N(_08854_),
    .Q(\mem.mem[63][5] ));
 sg13g2_dfrbp_1 _18719_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1031),
    .D(_00362_),
    .Q_N(_08853_),
    .Q(\mem.mem[63][6] ));
 sg13g2_dfrbp_1 _18720_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1030),
    .D(_00363_),
    .Q_N(_08852_),
    .Q(\mem.mem[63][7] ));
 sg13g2_dfrbp_1 _18721_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1029),
    .D(_00364_),
    .Q_N(_08851_),
    .Q(\mem.mem[84][0] ));
 sg13g2_dfrbp_1 _18722_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1028),
    .D(_00365_),
    .Q_N(_08850_),
    .Q(\mem.mem[84][1] ));
 sg13g2_dfrbp_1 _18723_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1027),
    .D(net3713),
    .Q_N(_08849_),
    .Q(\mem.mem[84][2] ));
 sg13g2_dfrbp_1 _18724_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1026),
    .D(_00367_),
    .Q_N(_08848_),
    .Q(\mem.mem[84][3] ));
 sg13g2_dfrbp_1 _18725_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1025),
    .D(_00368_),
    .Q_N(_08847_),
    .Q(\mem.mem[84][4] ));
 sg13g2_dfrbp_1 _18726_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1024),
    .D(_00369_),
    .Q_N(_08846_),
    .Q(\mem.mem[84][5] ));
 sg13g2_dfrbp_1 _18727_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1023),
    .D(_00370_),
    .Q_N(_08845_),
    .Q(\mem.mem[84][6] ));
 sg13g2_dfrbp_1 _18728_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1022),
    .D(_00371_),
    .Q_N(_08844_),
    .Q(\mem.mem[84][7] ));
 sg13g2_dfrbp_1 _18729_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1021),
    .D(_00372_),
    .Q_N(_08843_),
    .Q(\mem.mem[62][0] ));
 sg13g2_dfrbp_1 _18730_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1020),
    .D(_00373_),
    .Q_N(_08842_),
    .Q(\mem.mem[62][1] ));
 sg13g2_dfrbp_1 _18731_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1019),
    .D(_00374_),
    .Q_N(_08841_),
    .Q(\mem.mem[62][2] ));
 sg13g2_dfrbp_1 _18732_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1018),
    .D(_00375_),
    .Q_N(_08840_),
    .Q(\mem.mem[62][3] ));
 sg13g2_dfrbp_1 _18733_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1017),
    .D(_00376_),
    .Q_N(_08839_),
    .Q(\mem.mem[62][4] ));
 sg13g2_dfrbp_1 _18734_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1016),
    .D(_00377_),
    .Q_N(_08838_),
    .Q(\mem.mem[62][5] ));
 sg13g2_dfrbp_1 _18735_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1015),
    .D(_00378_),
    .Q_N(_08837_),
    .Q(\mem.mem[62][6] ));
 sg13g2_dfrbp_1 _18736_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1014),
    .D(net3894),
    .Q_N(_08836_),
    .Q(\mem.mem[62][7] ));
 sg13g2_dfrbp_1 _18737_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1013),
    .D(_00380_),
    .Q_N(_08835_),
    .Q(\mem.mem[61][0] ));
 sg13g2_dfrbp_1 _18738_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1012),
    .D(_00381_),
    .Q_N(_08834_),
    .Q(\mem.mem[61][1] ));
 sg13g2_dfrbp_1 _18739_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1011),
    .D(_00382_),
    .Q_N(_08833_),
    .Q(\mem.mem[61][2] ));
 sg13g2_dfrbp_1 _18740_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1010),
    .D(_00383_),
    .Q_N(_08832_),
    .Q(\mem.mem[61][3] ));
 sg13g2_dfrbp_1 _18741_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1009),
    .D(_00384_),
    .Q_N(_08831_),
    .Q(\mem.mem[61][4] ));
 sg13g2_dfrbp_1 _18742_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1008),
    .D(_00385_),
    .Q_N(_08830_),
    .Q(\mem.mem[61][5] ));
 sg13g2_dfrbp_1 _18743_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1007),
    .D(_00386_),
    .Q_N(_08829_),
    .Q(\mem.mem[61][6] ));
 sg13g2_dfrbp_1 _18744_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1006),
    .D(_00387_),
    .Q_N(_08828_),
    .Q(\mem.mem[61][7] ));
 sg13g2_dfrbp_1 _18745_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1005),
    .D(_00388_),
    .Q_N(_08827_),
    .Q(\mem.mem[83][0] ));
 sg13g2_dfrbp_1 _18746_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1004),
    .D(_00389_),
    .Q_N(_08826_),
    .Q(\mem.mem[83][1] ));
 sg13g2_dfrbp_1 _18747_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1003),
    .D(_00390_),
    .Q_N(_08825_),
    .Q(\mem.mem[83][2] ));
 sg13g2_dfrbp_1 _18748_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1002),
    .D(_00391_),
    .Q_N(_08824_),
    .Q(\mem.mem[83][3] ));
 sg13g2_dfrbp_1 _18749_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1001),
    .D(_00392_),
    .Q_N(_08823_),
    .Q(\mem.mem[83][4] ));
 sg13g2_dfrbp_1 _18750_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1000),
    .D(_00393_),
    .Q_N(_08822_),
    .Q(\mem.mem[83][5] ));
 sg13g2_dfrbp_1 _18751_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net999),
    .D(_00394_),
    .Q_N(_08821_),
    .Q(\mem.mem[83][6] ));
 sg13g2_dfrbp_1 _18752_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net998),
    .D(_00395_),
    .Q_N(_08820_),
    .Q(\mem.mem[83][7] ));
 sg13g2_dfrbp_1 _18753_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net997),
    .D(_00396_),
    .Q_N(_08819_),
    .Q(\mem.mem[60][0] ));
 sg13g2_dfrbp_1 _18754_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net996),
    .D(_00397_),
    .Q_N(_08818_),
    .Q(\mem.mem[60][1] ));
 sg13g2_dfrbp_1 _18755_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net995),
    .D(_00398_),
    .Q_N(_08817_),
    .Q(\mem.mem[60][2] ));
 sg13g2_dfrbp_1 _18756_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net994),
    .D(_00399_),
    .Q_N(_08816_),
    .Q(\mem.mem[60][3] ));
 sg13g2_dfrbp_1 _18757_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net993),
    .D(_00400_),
    .Q_N(_08815_),
    .Q(\mem.mem[60][4] ));
 sg13g2_dfrbp_1 _18758_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net992),
    .D(_00401_),
    .Q_N(_08814_),
    .Q(\mem.mem[60][5] ));
 sg13g2_dfrbp_1 _18759_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net991),
    .D(_00402_),
    .Q_N(_08813_),
    .Q(\mem.mem[60][6] ));
 sg13g2_dfrbp_1 _18760_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net990),
    .D(_00403_),
    .Q_N(_08812_),
    .Q(\mem.mem[60][7] ));
 sg13g2_dfrbp_1 _18761_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net989),
    .D(_00404_),
    .Q_N(_08811_),
    .Q(\mem.mem[5][0] ));
 sg13g2_dfrbp_1 _18762_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net988),
    .D(_00405_),
    .Q_N(_08810_),
    .Q(\mem.mem[5][1] ));
 sg13g2_dfrbp_1 _18763_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net987),
    .D(_00406_),
    .Q_N(_08809_),
    .Q(\mem.mem[5][2] ));
 sg13g2_dfrbp_1 _18764_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net986),
    .D(_00407_),
    .Q_N(_08808_),
    .Q(\mem.mem[5][3] ));
 sg13g2_dfrbp_1 _18765_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net985),
    .D(_00408_),
    .Q_N(_08807_),
    .Q(\mem.mem[5][4] ));
 sg13g2_dfrbp_1 _18766_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net984),
    .D(_00409_),
    .Q_N(_08806_),
    .Q(\mem.mem[5][5] ));
 sg13g2_dfrbp_1 _18767_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net983),
    .D(_00410_),
    .Q_N(_08805_),
    .Q(\mem.mem[5][6] ));
 sg13g2_dfrbp_1 _18768_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net982),
    .D(_00411_),
    .Q_N(_08804_),
    .Q(\mem.mem[5][7] ));
 sg13g2_dfrbp_1 _18769_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net981),
    .D(_00412_),
    .Q_N(_08803_),
    .Q(\mem.mem[82][0] ));
 sg13g2_dfrbp_1 _18770_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net980),
    .D(_00413_),
    .Q_N(_08802_),
    .Q(\mem.mem[82][1] ));
 sg13g2_dfrbp_1 _18771_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net979),
    .D(_00414_),
    .Q_N(_08801_),
    .Q(\mem.mem[82][2] ));
 sg13g2_dfrbp_1 _18772_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net978),
    .D(_00415_),
    .Q_N(_08800_),
    .Q(\mem.mem[82][3] ));
 sg13g2_dfrbp_1 _18773_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net977),
    .D(_00416_),
    .Q_N(_08799_),
    .Q(\mem.mem[82][4] ));
 sg13g2_dfrbp_1 _18774_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net976),
    .D(_00417_),
    .Q_N(_08798_),
    .Q(\mem.mem[82][5] ));
 sg13g2_dfrbp_1 _18775_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net975),
    .D(_00418_),
    .Q_N(_08797_),
    .Q(\mem.mem[82][6] ));
 sg13g2_dfrbp_1 _18776_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net974),
    .D(_00419_),
    .Q_N(_08796_),
    .Q(\mem.mem[82][7] ));
 sg13g2_dfrbp_1 _18777_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net973),
    .D(_00420_),
    .Q_N(_08795_),
    .Q(\mem.mem[58][0] ));
 sg13g2_dfrbp_1 _18778_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net972),
    .D(_00421_),
    .Q_N(_08794_),
    .Q(\mem.mem[58][1] ));
 sg13g2_dfrbp_1 _18779_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net971),
    .D(_00422_),
    .Q_N(_08793_),
    .Q(\mem.mem[58][2] ));
 sg13g2_dfrbp_1 _18780_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net970),
    .D(_00423_),
    .Q_N(_08792_),
    .Q(\mem.mem[58][3] ));
 sg13g2_dfrbp_1 _18781_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net969),
    .D(_00424_),
    .Q_N(_08791_),
    .Q(\mem.mem[58][4] ));
 sg13g2_dfrbp_1 _18782_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net968),
    .D(_00425_),
    .Q_N(_08790_),
    .Q(\mem.mem[58][5] ));
 sg13g2_dfrbp_1 _18783_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net967),
    .D(_00426_),
    .Q_N(_08789_),
    .Q(\mem.mem[58][6] ));
 sg13g2_dfrbp_1 _18784_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net966),
    .D(_00427_),
    .Q_N(_08788_),
    .Q(\mem.mem[58][7] ));
 sg13g2_dfrbp_1 _18785_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net965),
    .D(_00428_),
    .Q_N(_08787_),
    .Q(\mem.mem[57][0] ));
 sg13g2_dfrbp_1 _18786_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net964),
    .D(_00429_),
    .Q_N(_08786_),
    .Q(\mem.mem[57][1] ));
 sg13g2_dfrbp_1 _18787_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net963),
    .D(_00430_),
    .Q_N(_08785_),
    .Q(\mem.mem[57][2] ));
 sg13g2_dfrbp_1 _18788_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net962),
    .D(_00431_),
    .Q_N(_08784_),
    .Q(\mem.mem[57][3] ));
 sg13g2_dfrbp_1 _18789_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net961),
    .D(_00432_),
    .Q_N(_08783_),
    .Q(\mem.mem[57][4] ));
 sg13g2_dfrbp_1 _18790_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net960),
    .D(_00433_),
    .Q_N(_08782_),
    .Q(\mem.mem[57][5] ));
 sg13g2_dfrbp_1 _18791_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net959),
    .D(_00434_),
    .Q_N(_08781_),
    .Q(\mem.mem[57][6] ));
 sg13g2_dfrbp_1 _18792_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net958),
    .D(_00435_),
    .Q_N(_08780_),
    .Q(\mem.mem[57][7] ));
 sg13g2_dfrbp_1 _18793_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net957),
    .D(_00436_),
    .Q_N(_08779_),
    .Q(\mem.mem[81][0] ));
 sg13g2_dfrbp_1 _18794_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net956),
    .D(_00437_),
    .Q_N(_08778_),
    .Q(\mem.mem[81][1] ));
 sg13g2_dfrbp_1 _18795_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net955),
    .D(_00438_),
    .Q_N(_08777_),
    .Q(\mem.mem[81][2] ));
 sg13g2_dfrbp_1 _18796_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net954),
    .D(_00439_),
    .Q_N(_08776_),
    .Q(\mem.mem[81][3] ));
 sg13g2_dfrbp_1 _18797_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net953),
    .D(_00440_),
    .Q_N(_08775_),
    .Q(\mem.mem[81][4] ));
 sg13g2_dfrbp_1 _18798_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net952),
    .D(_00441_),
    .Q_N(_08774_),
    .Q(\mem.mem[81][5] ));
 sg13g2_dfrbp_1 _18799_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net951),
    .D(_00442_),
    .Q_N(_08773_),
    .Q(\mem.mem[81][6] ));
 sg13g2_dfrbp_1 _18800_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net950),
    .D(_00443_),
    .Q_N(_08772_),
    .Q(\mem.mem[81][7] ));
 sg13g2_dfrbp_1 _18801_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net949),
    .D(_00444_),
    .Q_N(_08771_),
    .Q(\mem.mem[56][0] ));
 sg13g2_dfrbp_1 _18802_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net948),
    .D(net3506),
    .Q_N(_08770_),
    .Q(\mem.mem[56][1] ));
 sg13g2_dfrbp_1 _18803_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net947),
    .D(_00446_),
    .Q_N(_08769_),
    .Q(\mem.mem[56][2] ));
 sg13g2_dfrbp_1 _18804_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net946),
    .D(_00447_),
    .Q_N(_08768_),
    .Q(\mem.mem[56][3] ));
 sg13g2_dfrbp_1 _18805_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net945),
    .D(_00448_),
    .Q_N(_08767_),
    .Q(\mem.mem[56][4] ));
 sg13g2_dfrbp_1 _18806_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net944),
    .D(_00449_),
    .Q_N(_08766_),
    .Q(\mem.mem[56][5] ));
 sg13g2_dfrbp_1 _18807_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net943),
    .D(_00450_),
    .Q_N(_08765_),
    .Q(\mem.mem[56][6] ));
 sg13g2_dfrbp_1 _18808_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net942),
    .D(_00451_),
    .Q_N(_08764_),
    .Q(\mem.mem[56][7] ));
 sg13g2_dfrbp_1 _18809_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net941),
    .D(_00452_),
    .Q_N(_08763_),
    .Q(\mem.mem[55][0] ));
 sg13g2_dfrbp_1 _18810_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net940),
    .D(_00453_),
    .Q_N(_08762_),
    .Q(\mem.mem[55][1] ));
 sg13g2_dfrbp_1 _18811_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net939),
    .D(_00454_),
    .Q_N(_08761_),
    .Q(\mem.mem[55][2] ));
 sg13g2_dfrbp_1 _18812_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net938),
    .D(_00455_),
    .Q_N(_08760_),
    .Q(\mem.mem[55][3] ));
 sg13g2_dfrbp_1 _18813_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net937),
    .D(_00456_),
    .Q_N(_08759_),
    .Q(\mem.mem[55][4] ));
 sg13g2_dfrbp_1 _18814_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net936),
    .D(_00457_),
    .Q_N(_08758_),
    .Q(\mem.mem[55][5] ));
 sg13g2_dfrbp_1 _18815_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net935),
    .D(_00458_),
    .Q_N(_08757_),
    .Q(\mem.mem[55][6] ));
 sg13g2_dfrbp_1 _18816_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net934),
    .D(_00459_),
    .Q_N(_08756_),
    .Q(\mem.mem[55][7] ));
 sg13g2_dfrbp_1 _18817_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net933),
    .D(_00460_),
    .Q_N(_08755_),
    .Q(\mem.mem[80][0] ));
 sg13g2_dfrbp_1 _18818_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net932),
    .D(_00461_),
    .Q_N(_08754_),
    .Q(\mem.mem[80][1] ));
 sg13g2_dfrbp_1 _18819_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net931),
    .D(_00462_),
    .Q_N(_08753_),
    .Q(\mem.mem[80][2] ));
 sg13g2_dfrbp_1 _18820_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net930),
    .D(_00463_),
    .Q_N(_08752_),
    .Q(\mem.mem[80][3] ));
 sg13g2_dfrbp_1 _18821_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net929),
    .D(_00464_),
    .Q_N(_08751_),
    .Q(\mem.mem[80][4] ));
 sg13g2_dfrbp_1 _18822_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net928),
    .D(_00465_),
    .Q_N(_08750_),
    .Q(\mem.mem[80][5] ));
 sg13g2_dfrbp_1 _18823_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net927),
    .D(_00466_),
    .Q_N(_08749_),
    .Q(\mem.mem[80][6] ));
 sg13g2_dfrbp_1 _18824_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net926),
    .D(_00467_),
    .Q_N(_08748_),
    .Q(\mem.mem[80][7] ));
 sg13g2_dfrbp_1 _18825_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net925),
    .D(_00468_),
    .Q_N(_08747_),
    .Q(\mem.mem[54][0] ));
 sg13g2_dfrbp_1 _18826_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net924),
    .D(_00469_),
    .Q_N(_08746_),
    .Q(\mem.mem[54][1] ));
 sg13g2_dfrbp_1 _18827_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net923),
    .D(_00470_),
    .Q_N(_08745_),
    .Q(\mem.mem[54][2] ));
 sg13g2_dfrbp_1 _18828_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net922),
    .D(_00471_),
    .Q_N(_08744_),
    .Q(\mem.mem[54][3] ));
 sg13g2_dfrbp_1 _18829_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net921),
    .D(_00472_),
    .Q_N(_08743_),
    .Q(\mem.mem[54][4] ));
 sg13g2_dfrbp_1 _18830_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net920),
    .D(_00473_),
    .Q_N(_08742_),
    .Q(\mem.mem[54][5] ));
 sg13g2_dfrbp_1 _18831_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net919),
    .D(_00474_),
    .Q_N(_08741_),
    .Q(\mem.mem[54][6] ));
 sg13g2_dfrbp_1 _18832_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net918),
    .D(_00475_),
    .Q_N(_08740_),
    .Q(\mem.mem[54][7] ));
 sg13g2_dfrbp_1 _18833_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net917),
    .D(_00476_),
    .Q_N(_08739_),
    .Q(\mem.mem[53][0] ));
 sg13g2_dfrbp_1 _18834_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net916),
    .D(_00477_),
    .Q_N(_08738_),
    .Q(\mem.mem[53][1] ));
 sg13g2_dfrbp_1 _18835_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net915),
    .D(_00478_),
    .Q_N(_08737_),
    .Q(\mem.mem[53][2] ));
 sg13g2_dfrbp_1 _18836_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net914),
    .D(_00479_),
    .Q_N(_08736_),
    .Q(\mem.mem[53][3] ));
 sg13g2_dfrbp_1 _18837_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net913),
    .D(_00480_),
    .Q_N(_08735_),
    .Q(\mem.mem[53][4] ));
 sg13g2_dfrbp_1 _18838_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net912),
    .D(_00481_),
    .Q_N(_08734_),
    .Q(\mem.mem[53][5] ));
 sg13g2_dfrbp_1 _18839_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net911),
    .D(_00482_),
    .Q_N(_08733_),
    .Q(\mem.mem[53][6] ));
 sg13g2_dfrbp_1 _18840_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net910),
    .D(_00483_),
    .Q_N(_08732_),
    .Q(\mem.mem[53][7] ));
 sg13g2_dfrbp_1 _18841_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net909),
    .D(_00484_),
    .Q_N(_08731_),
    .Q(\mem.mem[7][0] ));
 sg13g2_dfrbp_1 _18842_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net908),
    .D(_00485_),
    .Q_N(_08730_),
    .Q(\mem.mem[7][1] ));
 sg13g2_dfrbp_1 _18843_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net907),
    .D(_00486_),
    .Q_N(_08729_),
    .Q(\mem.mem[7][2] ));
 sg13g2_dfrbp_1 _18844_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net906),
    .D(_00487_),
    .Q_N(_08728_),
    .Q(\mem.mem[7][3] ));
 sg13g2_dfrbp_1 _18845_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net905),
    .D(_00488_),
    .Q_N(_08727_),
    .Q(\mem.mem[7][4] ));
 sg13g2_dfrbp_1 _18846_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net904),
    .D(_00489_),
    .Q_N(_08726_),
    .Q(\mem.mem[7][5] ));
 sg13g2_dfrbp_1 _18847_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net903),
    .D(_00490_),
    .Q_N(_08725_),
    .Q(\mem.mem[7][6] ));
 sg13g2_dfrbp_1 _18848_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net902),
    .D(_00491_),
    .Q_N(_08724_),
    .Q(\mem.mem[7][7] ));
 sg13g2_dfrbp_1 _18849_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net901),
    .D(_00492_),
    .Q_N(_08723_),
    .Q(\mem.mem[52][0] ));
 sg13g2_dfrbp_1 _18850_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net900),
    .D(_00493_),
    .Q_N(_08722_),
    .Q(\mem.mem[52][1] ));
 sg13g2_dfrbp_1 _18851_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net899),
    .D(_00494_),
    .Q_N(_08721_),
    .Q(\mem.mem[52][2] ));
 sg13g2_dfrbp_1 _18852_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net898),
    .D(_00495_),
    .Q_N(_08720_),
    .Q(\mem.mem[52][3] ));
 sg13g2_dfrbp_1 _18853_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net897),
    .D(net3970),
    .Q_N(_08719_),
    .Q(\mem.mem[52][4] ));
 sg13g2_dfrbp_1 _18854_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net896),
    .D(_00497_),
    .Q_N(_08718_),
    .Q(\mem.mem[52][5] ));
 sg13g2_dfrbp_1 _18855_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net895),
    .D(net4147),
    .Q_N(_08717_),
    .Q(\mem.mem[52][6] ));
 sg13g2_dfrbp_1 _18856_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net894),
    .D(_00499_),
    .Q_N(_08716_),
    .Q(\mem.mem[52][7] ));
 sg13g2_dfrbp_1 _18857_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net893),
    .D(_00500_),
    .Q_N(_08715_),
    .Q(\mem.mem[51][0] ));
 sg13g2_dfrbp_1 _18858_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net892),
    .D(_00501_),
    .Q_N(_08714_),
    .Q(\mem.mem[51][1] ));
 sg13g2_dfrbp_1 _18859_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net891),
    .D(_00502_),
    .Q_N(_08713_),
    .Q(\mem.mem[51][2] ));
 sg13g2_dfrbp_1 _18860_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net890),
    .D(_00503_),
    .Q_N(_08712_),
    .Q(\mem.mem[51][3] ));
 sg13g2_dfrbp_1 _18861_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net889),
    .D(_00504_),
    .Q_N(_08711_),
    .Q(\mem.mem[51][4] ));
 sg13g2_dfrbp_1 _18862_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net888),
    .D(_00505_),
    .Q_N(_08710_),
    .Q(\mem.mem[51][5] ));
 sg13g2_dfrbp_1 _18863_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net887),
    .D(_00506_),
    .Q_N(_08709_),
    .Q(\mem.mem[51][6] ));
 sg13g2_dfrbp_1 _18864_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net886),
    .D(_00507_),
    .Q_N(_08708_),
    .Q(\mem.mem[51][7] ));
 sg13g2_dfrbp_1 _18865_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net885),
    .D(_00508_),
    .Q_N(_08707_),
    .Q(\mem.mem[78][0] ));
 sg13g2_dfrbp_1 _18866_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net884),
    .D(_00509_),
    .Q_N(_08706_),
    .Q(\mem.mem[78][1] ));
 sg13g2_dfrbp_1 _18867_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net883),
    .D(_00510_),
    .Q_N(_08705_),
    .Q(\mem.mem[78][2] ));
 sg13g2_dfrbp_1 _18868_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net882),
    .D(_00511_),
    .Q_N(_08704_),
    .Q(\mem.mem[78][3] ));
 sg13g2_dfrbp_1 _18869_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net881),
    .D(_00512_),
    .Q_N(_08703_),
    .Q(\mem.mem[78][4] ));
 sg13g2_dfrbp_1 _18870_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net880),
    .D(_00513_),
    .Q_N(_08702_),
    .Q(\mem.mem[78][5] ));
 sg13g2_dfrbp_1 _18871_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net879),
    .D(_00514_),
    .Q_N(_08701_),
    .Q(\mem.mem[78][6] ));
 sg13g2_dfrbp_1 _18872_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net878),
    .D(_00515_),
    .Q_N(_08700_),
    .Q(\mem.mem[78][7] ));
 sg13g2_dfrbp_1 _18873_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net877),
    .D(_00516_),
    .Q_N(_08699_),
    .Q(\mem.mem[50][0] ));
 sg13g2_dfrbp_1 _18874_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net876),
    .D(_00517_),
    .Q_N(_08698_),
    .Q(\mem.mem[50][1] ));
 sg13g2_dfrbp_1 _18875_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net875),
    .D(_00518_),
    .Q_N(_08697_),
    .Q(\mem.mem[50][2] ));
 sg13g2_dfrbp_1 _18876_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net874),
    .D(_00519_),
    .Q_N(_08696_),
    .Q(\mem.mem[50][3] ));
 sg13g2_dfrbp_1 _18877_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net873),
    .D(_00520_),
    .Q_N(_08695_),
    .Q(\mem.mem[50][4] ));
 sg13g2_dfrbp_1 _18878_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net872),
    .D(_00521_),
    .Q_N(_08694_),
    .Q(\mem.mem[50][5] ));
 sg13g2_dfrbp_1 _18879_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net871),
    .D(_00522_),
    .Q_N(_08693_),
    .Q(\mem.mem[50][6] ));
 sg13g2_dfrbp_1 _18880_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net870),
    .D(_00523_),
    .Q_N(_08692_),
    .Q(\mem.mem[50][7] ));
 sg13g2_dfrbp_1 _18881_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net869),
    .D(_00524_),
    .Q_N(_08691_),
    .Q(\mem.mem[4][0] ));
 sg13g2_dfrbp_1 _18882_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net868),
    .D(_00525_),
    .Q_N(_08690_),
    .Q(\mem.mem[4][1] ));
 sg13g2_dfrbp_1 _18883_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net867),
    .D(_00526_),
    .Q_N(_08689_),
    .Q(\mem.mem[4][2] ));
 sg13g2_dfrbp_1 _18884_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net866),
    .D(_00527_),
    .Q_N(_08688_),
    .Q(\mem.mem[4][3] ));
 sg13g2_dfrbp_1 _18885_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net865),
    .D(_00528_),
    .Q_N(_08687_),
    .Q(\mem.mem[4][4] ));
 sg13g2_dfrbp_1 _18886_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net864),
    .D(_00529_),
    .Q_N(_08686_),
    .Q(\mem.mem[4][5] ));
 sg13g2_dfrbp_1 _18887_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net863),
    .D(_00530_),
    .Q_N(_08685_),
    .Q(\mem.mem[4][6] ));
 sg13g2_dfrbp_1 _18888_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net862),
    .D(_00531_),
    .Q_N(_08684_),
    .Q(\mem.mem[4][7] ));
 sg13g2_dfrbp_1 _18889_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net861),
    .D(_00532_),
    .Q_N(_08683_),
    .Q(\mem.mem[77][0] ));
 sg13g2_dfrbp_1 _18890_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net860),
    .D(_00533_),
    .Q_N(_08682_),
    .Q(\mem.mem[77][1] ));
 sg13g2_dfrbp_1 _18891_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net859),
    .D(_00534_),
    .Q_N(_08681_),
    .Q(\mem.mem[77][2] ));
 sg13g2_dfrbp_1 _18892_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net858),
    .D(_00535_),
    .Q_N(_08680_),
    .Q(\mem.mem[77][3] ));
 sg13g2_dfrbp_1 _18893_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net857),
    .D(_00536_),
    .Q_N(_08679_),
    .Q(\mem.mem[77][4] ));
 sg13g2_dfrbp_1 _18894_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net856),
    .D(_00537_),
    .Q_N(_08678_),
    .Q(\mem.mem[77][5] ));
 sg13g2_dfrbp_1 _18895_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net855),
    .D(_00538_),
    .Q_N(_08677_),
    .Q(\mem.mem[77][6] ));
 sg13g2_dfrbp_1 _18896_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net854),
    .D(_00539_),
    .Q_N(_08676_),
    .Q(\mem.mem[77][7] ));
 sg13g2_dfrbp_1 _18897_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net853),
    .D(_00540_),
    .Q_N(_08675_),
    .Q(\mem.mem[48][0] ));
 sg13g2_dfrbp_1 _18898_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net852),
    .D(_00541_),
    .Q_N(_08674_),
    .Q(\mem.mem[48][1] ));
 sg13g2_dfrbp_1 _18899_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net851),
    .D(_00542_),
    .Q_N(_08673_),
    .Q(\mem.mem[48][2] ));
 sg13g2_dfrbp_1 _18900_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net850),
    .D(_00543_),
    .Q_N(_08672_),
    .Q(\mem.mem[48][3] ));
 sg13g2_dfrbp_1 _18901_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net849),
    .D(_00544_),
    .Q_N(_08671_),
    .Q(\mem.mem[48][4] ));
 sg13g2_dfrbp_1 _18902_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net848),
    .D(_00545_),
    .Q_N(_08670_),
    .Q(\mem.mem[48][5] ));
 sg13g2_dfrbp_1 _18903_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net847),
    .D(_00546_),
    .Q_N(_08669_),
    .Q(\mem.mem[48][6] ));
 sg13g2_dfrbp_1 _18904_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net846),
    .D(_00547_),
    .Q_N(_08668_),
    .Q(\mem.mem[48][7] ));
 sg13g2_dfrbp_1 _18905_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net845),
    .D(net4184),
    .Q_N(_08667_),
    .Q(\A[0] ));
 sg13g2_dfrbp_1 _18906_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net843),
    .D(net4196),
    .Q_N(_08666_),
    .Q(\A[1] ));
 sg13g2_dfrbp_1 _18907_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net841),
    .D(net4198),
    .Q_N(_08665_),
    .Q(\A[2] ));
 sg13g2_dfrbp_1 _18908_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net839),
    .D(net4182),
    .Q_N(_08664_),
    .Q(\A[3] ));
 sg13g2_dfrbp_1 _18909_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net837),
    .D(_00552_),
    .Q_N(_08663_),
    .Q(\A[4] ));
 sg13g2_dfrbp_1 _18910_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net835),
    .D(net4179),
    .Q_N(_08662_),
    .Q(\A[5] ));
 sg13g2_dfrbp_1 _18911_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net833),
    .D(_00554_),
    .Q_N(_08661_),
    .Q(\A[6] ));
 sg13g2_dfrbp_1 _18912_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net831),
    .D(_00555_),
    .Q_N(_08660_),
    .Q(\A[7] ));
 sg13g2_dfrbp_1 _18913_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net829),
    .D(_00556_),
    .Q_N(_08659_),
    .Q(\B[0] ));
 sg13g2_dfrbp_1 _18914_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net827),
    .D(_00557_),
    .Q_N(_08658_),
    .Q(\B[1] ));
 sg13g2_dfrbp_1 _18915_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net825),
    .D(_00558_),
    .Q_N(_08657_),
    .Q(\B[2] ));
 sg13g2_dfrbp_1 _18916_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net823),
    .D(_00559_),
    .Q_N(_08656_),
    .Q(\B[3] ));
 sg13g2_dfrbp_1 _18917_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net821),
    .D(_00560_),
    .Q_N(_08655_),
    .Q(\B[4] ));
 sg13g2_dfrbp_1 _18918_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net819),
    .D(_00561_),
    .Q_N(_08654_),
    .Q(\B[5] ));
 sg13g2_dfrbp_1 _18919_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net817),
    .D(net4191),
    .Q_N(_08653_),
    .Q(\B[6] ));
 sg13g2_dfrbp_1 _18920_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net815),
    .D(_00563_),
    .Q_N(_08652_),
    .Q(\B[7] ));
 sg13g2_dfrbp_1 _18921_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net813),
    .D(net4186),
    .Q_N(_08651_),
    .Q(\C[0] ));
 sg13g2_dfrbp_1 _18922_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net811),
    .D(net4172),
    .Q_N(_00026_),
    .Q(\C[1] ));
 sg13g2_dfrbp_1 _18923_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net809),
    .D(net4170),
    .Q_N(_00025_),
    .Q(\C[2] ));
 sg13g2_dfrbp_1 _18924_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net807),
    .D(_00567_),
    .Q_N(_00024_),
    .Q(\C[3] ));
 sg13g2_dfrbp_1 _18925_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net805),
    .D(_00568_),
    .Q_N(_00023_),
    .Q(\C[4] ));
 sg13g2_dfrbp_1 _18926_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net803),
    .D(net3920),
    .Q_N(_00022_),
    .Q(\C[5] ));
 sg13g2_dfrbp_1 _18927_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net801),
    .D(_00570_),
    .Q_N(_00021_),
    .Q(\C[6] ));
 sg13g2_dfrbp_1 _18928_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net799),
    .D(net4176),
    .Q_N(_00020_),
    .Q(\C[7] ));
 sg13g2_dfrbp_1 _18929_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net797),
    .D(net4224),
    .Q_N(_00019_),
    .Q(\PC[0] ));
 sg13g2_dfrbp_1 _18930_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net795),
    .D(_00573_),
    .Q_N(_08650_),
    .Q(\PC[1] ));
 sg13g2_dfrbp_1 _18931_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net793),
    .D(_00574_),
    .Q_N(_08649_),
    .Q(\PC[2] ));
 sg13g2_dfrbp_1 _18932_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net791),
    .D(_00575_),
    .Q_N(_08648_),
    .Q(\PC[3] ));
 sg13g2_dfrbp_1 _18933_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net789),
    .D(_00576_),
    .Q_N(_00018_),
    .Q(\PC[4] ));
 sg13g2_dfrbp_1 _18934_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net787),
    .D(net4220),
    .Q_N(_08647_),
    .Q(\PC[5] ));
 sg13g2_dfrbp_1 _18935_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net785),
    .D(net4222),
    .Q_N(_00017_),
    .Q(\PC[6] ));
 sg13g2_dfrbp_1 _18936_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net783),
    .D(net4235),
    .Q_N(_08646_),
    .Q(\PC[7] ));
 sg13g2_dfrbp_1 _18937_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net781),
    .D(net4256),
    .Q_N(_08645_),
    .Q(\mem.addr[0] ));
 sg13g2_dfrbp_1 _18938_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net779),
    .D(_00581_),
    .Q_N(_08644_),
    .Q(\mem.addr[1] ));
 sg13g2_dfrbp_1 _18939_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net777),
    .D(_00582_),
    .Q_N(_08643_),
    .Q(\mem.addr[2] ));
 sg13g2_dfrbp_1 _18940_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net775),
    .D(_00583_),
    .Q_N(_08642_),
    .Q(\mem.addr[3] ));
 sg13g2_dfrbp_1 _18941_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net773),
    .D(_00584_),
    .Q_N(_08641_),
    .Q(\mem.addr[4] ));
 sg13g2_dfrbp_1 _18942_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net771),
    .D(_00585_),
    .Q_N(_08640_),
    .Q(\mem.addr[5] ));
 sg13g2_dfrbp_1 _18943_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net769),
    .D(_00586_),
    .Q_N(_08639_),
    .Q(\mem.addr[6] ));
 sg13g2_dfrbp_1 _18944_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net767),
    .D(_00587_),
    .Q_N(_08638_),
    .Q(\mem.addr[7] ));
 sg13g2_dfrbp_1 _18945_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net765),
    .D(_00588_),
    .Q_N(_08637_),
    .Q(\mem.mem[139][0] ));
 sg13g2_dfrbp_1 _18946_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net764),
    .D(_00589_),
    .Q_N(_08636_),
    .Q(\mem.mem[139][1] ));
 sg13g2_dfrbp_1 _18947_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net763),
    .D(_00590_),
    .Q_N(_08635_),
    .Q(\mem.mem[139][2] ));
 sg13g2_dfrbp_1 _18948_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net762),
    .D(_00591_),
    .Q_N(_08634_),
    .Q(\mem.mem[139][3] ));
 sg13g2_dfrbp_1 _18949_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net761),
    .D(_00592_),
    .Q_N(_08633_),
    .Q(\mem.mem[139][4] ));
 sg13g2_dfrbp_1 _18950_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net760),
    .D(_00593_),
    .Q_N(_08632_),
    .Q(\mem.mem[139][5] ));
 sg13g2_dfrbp_1 _18951_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net759),
    .D(_00594_),
    .Q_N(_08631_),
    .Q(\mem.mem[139][6] ));
 sg13g2_dfrbp_1 _18952_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net758),
    .D(_00595_),
    .Q_N(_08630_),
    .Q(\mem.mem[139][7] ));
 sg13g2_dfrbp_1 _18953_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net757),
    .D(_00596_),
    .Q_N(_08629_),
    .Q(\mem.data_in[0] ));
 sg13g2_dfrbp_1 _18954_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net755),
    .D(_00597_),
    .Q_N(_08628_),
    .Q(\mem.data_in[1] ));
 sg13g2_dfrbp_1 _18955_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net753),
    .D(_00598_),
    .Q_N(_08627_),
    .Q(\mem.data_in[2] ));
 sg13g2_dfrbp_1 _18956_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net751),
    .D(_00599_),
    .Q_N(_08626_),
    .Q(\mem.data_in[3] ));
 sg13g2_dfrbp_1 _18957_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net749),
    .D(_00600_),
    .Q_N(_08625_),
    .Q(\mem.data_in[4] ));
 sg13g2_dfrbp_1 _18958_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net747),
    .D(_00601_),
    .Q_N(_08624_),
    .Q(\mem.data_in[5] ));
 sg13g2_dfrbp_1 _18959_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net745),
    .D(_00602_),
    .Q_N(_08623_),
    .Q(\mem.data_in[6] ));
 sg13g2_dfrbp_1 _18960_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net743),
    .D(_00603_),
    .Q_N(_08622_),
    .Q(\mem.data_in[7] ));
 sg13g2_dfrbp_1 _18961_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net741),
    .D(_00604_),
    .Q_N(_08621_),
    .Q(\mem_A[0] ));
 sg13g2_dfrbp_1 _18962_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net739),
    .D(_00605_),
    .Q_N(_00016_),
    .Q(\mem_A[1] ));
 sg13g2_dfrbp_1 _18963_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net737),
    .D(_00606_),
    .Q_N(_08620_),
    .Q(\mem_A[2] ));
 sg13g2_dfrbp_1 _18964_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net735),
    .D(_00607_),
    .Q_N(_08619_),
    .Q(\mem_A[3] ));
 sg13g2_dfrbp_1 _18965_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net733),
    .D(_00608_),
    .Q_N(_08618_),
    .Q(\mem_A[4] ));
 sg13g2_dfrbp_1 _18966_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net731),
    .D(_00609_),
    .Q_N(_08617_),
    .Q(\mem_A[5] ));
 sg13g2_dfrbp_1 _18967_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net729),
    .D(_00610_),
    .Q_N(_08616_),
    .Q(\mem_A[6] ));
 sg13g2_dfrbp_1 _18968_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net727),
    .D(_00611_),
    .Q_N(_08615_),
    .Q(\mem_A[7] ));
 sg13g2_dfrbp_1 _18969_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net725),
    .D(_00612_),
    .Q_N(_08614_),
    .Q(\mem.mem[76][0] ));
 sg13g2_dfrbp_1 _18970_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net724),
    .D(_00613_),
    .Q_N(_08613_),
    .Q(\mem.mem[76][1] ));
 sg13g2_dfrbp_1 _18971_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net723),
    .D(_00614_),
    .Q_N(_08612_),
    .Q(\mem.mem[76][2] ));
 sg13g2_dfrbp_1 _18972_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net722),
    .D(_00615_),
    .Q_N(_08611_),
    .Q(\mem.mem[76][3] ));
 sg13g2_dfrbp_1 _18973_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net721),
    .D(_00616_),
    .Q_N(_08610_),
    .Q(\mem.mem[76][4] ));
 sg13g2_dfrbp_1 _18974_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net720),
    .D(_00617_),
    .Q_N(_08609_),
    .Q(\mem.mem[76][5] ));
 sg13g2_dfrbp_1 _18975_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net719),
    .D(_00618_),
    .Q_N(_08608_),
    .Q(\mem.mem[76][6] ));
 sg13g2_dfrbp_1 _18976_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net718),
    .D(_00619_),
    .Q_N(_08607_),
    .Q(\mem.mem[76][7] ));
 sg13g2_dfrbp_1 _18977_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net717),
    .D(_00620_),
    .Q_N(_08606_),
    .Q(\mem.mem[75][0] ));
 sg13g2_dfrbp_1 _18978_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net716),
    .D(_00621_),
    .Q_N(_08605_),
    .Q(\mem.mem[75][1] ));
 sg13g2_dfrbp_1 _18979_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net715),
    .D(_00622_),
    .Q_N(_08604_),
    .Q(\mem.mem[75][2] ));
 sg13g2_dfrbp_1 _18980_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net714),
    .D(_00623_),
    .Q_N(_08603_),
    .Q(\mem.mem[75][3] ));
 sg13g2_dfrbp_1 _18981_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net713),
    .D(_00624_),
    .Q_N(_08602_),
    .Q(\mem.mem[75][4] ));
 sg13g2_dfrbp_1 _18982_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net712),
    .D(_00625_),
    .Q_N(_08601_),
    .Q(\mem.mem[75][5] ));
 sg13g2_dfrbp_1 _18983_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net711),
    .D(_00626_),
    .Q_N(_08600_),
    .Q(\mem.mem[75][6] ));
 sg13g2_dfrbp_1 _18984_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net710),
    .D(_00627_),
    .Q_N(_08599_),
    .Q(\mem.mem[75][7] ));
 sg13g2_dfrbp_1 _18985_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net709),
    .D(_00628_),
    .Q_N(_08598_),
    .Q(\mem.mem[28][0] ));
 sg13g2_dfrbp_1 _18986_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net708),
    .D(_00629_),
    .Q_N(_08597_),
    .Q(\mem.mem[28][1] ));
 sg13g2_dfrbp_1 _18987_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net707),
    .D(_00630_),
    .Q_N(_08596_),
    .Q(\mem.mem[28][2] ));
 sg13g2_dfrbp_1 _18988_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net706),
    .D(_00631_),
    .Q_N(_08595_),
    .Q(\mem.mem[28][3] ));
 sg13g2_dfrbp_1 _18989_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net705),
    .D(_00632_),
    .Q_N(_08594_),
    .Q(\mem.mem[28][4] ));
 sg13g2_dfrbp_1 _18990_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net704),
    .D(_00633_),
    .Q_N(_08593_),
    .Q(\mem.mem[28][5] ));
 sg13g2_dfrbp_1 _18991_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net703),
    .D(_00634_),
    .Q_N(_08592_),
    .Q(\mem.mem[28][6] ));
 sg13g2_dfrbp_1 _18992_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net702),
    .D(_00635_),
    .Q_N(_08591_),
    .Q(\mem.mem[28][7] ));
 sg13g2_dfrbp_1 _18993_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net701),
    .D(_00636_),
    .Q_N(_08590_),
    .Q(\mem.mem[27][0] ));
 sg13g2_dfrbp_1 _18994_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net700),
    .D(_00637_),
    .Q_N(_08589_),
    .Q(\mem.mem[27][1] ));
 sg13g2_dfrbp_1 _18995_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net699),
    .D(_00638_),
    .Q_N(_08588_),
    .Q(\mem.mem[27][2] ));
 sg13g2_dfrbp_1 _18996_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net698),
    .D(_00639_),
    .Q_N(_08587_),
    .Q(\mem.mem[27][3] ));
 sg13g2_dfrbp_1 _18997_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net697),
    .D(_00640_),
    .Q_N(_08586_),
    .Q(\mem.mem[27][4] ));
 sg13g2_dfrbp_1 _18998_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net696),
    .D(_00641_),
    .Q_N(_08585_),
    .Q(\mem.mem[27][5] ));
 sg13g2_dfrbp_1 _18999_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net688),
    .D(_00642_),
    .Q_N(_08584_),
    .Q(\mem.mem[27][6] ));
 sg13g2_dfrbp_1 _19000_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net687),
    .D(_00643_),
    .Q_N(_08583_),
    .Q(\mem.mem[27][7] ));
 sg13g2_dfrbp_1 _19001_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net686),
    .D(_00644_),
    .Q_N(_08582_),
    .Q(\mem.mem[26][0] ));
 sg13g2_dfrbp_1 _19002_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net685),
    .D(_00645_),
    .Q_N(_08581_),
    .Q(\mem.mem[26][1] ));
 sg13g2_dfrbp_1 _19003_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net684),
    .D(_00646_),
    .Q_N(_08580_),
    .Q(\mem.mem[26][2] ));
 sg13g2_dfrbp_1 _19004_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net683),
    .D(_00647_),
    .Q_N(_08579_),
    .Q(\mem.mem[26][3] ));
 sg13g2_dfrbp_1 _19005_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net682),
    .D(_00648_),
    .Q_N(_08578_),
    .Q(\mem.mem[26][4] ));
 sg13g2_dfrbp_1 _19006_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net681),
    .D(_00649_),
    .Q_N(_08577_),
    .Q(\mem.mem[26][5] ));
 sg13g2_dfrbp_1 _19007_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net680),
    .D(_00650_),
    .Q_N(_08576_),
    .Q(\mem.mem[26][6] ));
 sg13g2_dfrbp_1 _19008_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net679),
    .D(_00651_),
    .Q_N(_08575_),
    .Q(\mem.mem[26][7] ));
 sg13g2_dfrbp_1 _19009_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net678),
    .D(_00652_),
    .Q_N(_08574_),
    .Q(\mem.mem[25][0] ));
 sg13g2_dfrbp_1 _19010_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net677),
    .D(_00653_),
    .Q_N(_08573_),
    .Q(\mem.mem[25][1] ));
 sg13g2_dfrbp_1 _19011_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net676),
    .D(_00654_),
    .Q_N(_08572_),
    .Q(\mem.mem[25][2] ));
 sg13g2_dfrbp_1 _19012_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net675),
    .D(_00655_),
    .Q_N(_08571_),
    .Q(\mem.mem[25][3] ));
 sg13g2_dfrbp_1 _19013_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net674),
    .D(_00656_),
    .Q_N(_08570_),
    .Q(\mem.mem[25][4] ));
 sg13g2_dfrbp_1 _19014_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net673),
    .D(_00657_),
    .Q_N(_08569_),
    .Q(\mem.mem[25][5] ));
 sg13g2_dfrbp_1 _19015_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net672),
    .D(_00658_),
    .Q_N(_08568_),
    .Q(\mem.mem[25][6] ));
 sg13g2_dfrbp_1 _19016_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net671),
    .D(_00659_),
    .Q_N(_08567_),
    .Q(\mem.mem[25][7] ));
 sg13g2_dfrbp_1 _19017_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net670),
    .D(_00660_),
    .Q_N(_08566_),
    .Q(\mem.mem[252][0] ));
 sg13g2_dfrbp_1 _19018_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net669),
    .D(_00661_),
    .Q_N(_08565_),
    .Q(\mem.mem[252][1] ));
 sg13g2_dfrbp_1 _19019_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net668),
    .D(_00662_),
    .Q_N(_08564_),
    .Q(\mem.mem[252][2] ));
 sg13g2_dfrbp_1 _19020_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net667),
    .D(_00663_),
    .Q_N(_08563_),
    .Q(\mem.mem[252][3] ));
 sg13g2_dfrbp_1 _19021_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net666),
    .D(_00664_),
    .Q_N(_08562_),
    .Q(\mem.mem[252][4] ));
 sg13g2_dfrbp_1 _19022_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net665),
    .D(_00665_),
    .Q_N(_08561_),
    .Q(\mem.mem[252][5] ));
 sg13g2_dfrbp_1 _19023_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net664),
    .D(_00666_),
    .Q_N(_08560_),
    .Q(\mem.mem[252][6] ));
 sg13g2_dfrbp_1 _19024_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net663),
    .D(_00667_),
    .Q_N(_08559_),
    .Q(\mem.mem[252][7] ));
 sg13g2_dfrbp_1 _19025_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net662),
    .D(_00668_),
    .Q_N(_08558_),
    .Q(\mem.mem[249][0] ));
 sg13g2_dfrbp_1 _19026_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net661),
    .D(_00669_),
    .Q_N(_08557_),
    .Q(\mem.mem[249][1] ));
 sg13g2_dfrbp_1 _19027_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net660),
    .D(_00670_),
    .Q_N(_08556_),
    .Q(\mem.mem[249][2] ));
 sg13g2_dfrbp_1 _19028_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net659),
    .D(_00671_),
    .Q_N(_08555_),
    .Q(\mem.mem[249][3] ));
 sg13g2_dfrbp_1 _19029_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net658),
    .D(_00672_),
    .Q_N(_08554_),
    .Q(\mem.mem[249][4] ));
 sg13g2_dfrbp_1 _19030_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net657),
    .D(_00673_),
    .Q_N(_08553_),
    .Q(\mem.mem[249][5] ));
 sg13g2_dfrbp_1 _19031_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net656),
    .D(_00674_),
    .Q_N(_08552_),
    .Q(\mem.mem[249][6] ));
 sg13g2_dfrbp_1 _19032_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net655),
    .D(_00675_),
    .Q_N(_08551_),
    .Q(\mem.mem[249][7] ));
 sg13g2_dfrbp_1 _19033_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net654),
    .D(_00676_),
    .Q_N(_08550_),
    .Q(\mem.mem[239][0] ));
 sg13g2_dfrbp_1 _19034_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net653),
    .D(_00677_),
    .Q_N(_08549_),
    .Q(\mem.mem[239][1] ));
 sg13g2_dfrbp_1 _19035_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net652),
    .D(_00678_),
    .Q_N(_08548_),
    .Q(\mem.mem[239][2] ));
 sg13g2_dfrbp_1 _19036_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net651),
    .D(_00679_),
    .Q_N(_08547_),
    .Q(\mem.mem[239][3] ));
 sg13g2_dfrbp_1 _19037_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net650),
    .D(_00680_),
    .Q_N(_08546_),
    .Q(\mem.mem[239][4] ));
 sg13g2_dfrbp_1 _19038_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net649),
    .D(_00681_),
    .Q_N(_08545_),
    .Q(\mem.mem[239][5] ));
 sg13g2_dfrbp_1 _19039_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net648),
    .D(_00682_),
    .Q_N(_08544_),
    .Q(\mem.mem[239][6] ));
 sg13g2_dfrbp_1 _19040_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net647),
    .D(_00683_),
    .Q_N(_08543_),
    .Q(\mem.mem[239][7] ));
 sg13g2_dfrbp_1 _19041_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net646),
    .D(_00684_),
    .Q_N(_08542_),
    .Q(\mem.mem[229][0] ));
 sg13g2_dfrbp_1 _19042_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net645),
    .D(_00685_),
    .Q_N(_08541_),
    .Q(\mem.mem[229][1] ));
 sg13g2_dfrbp_1 _19043_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net644),
    .D(_00686_),
    .Q_N(_08540_),
    .Q(\mem.mem[229][2] ));
 sg13g2_dfrbp_1 _19044_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net643),
    .D(_00687_),
    .Q_N(_08539_),
    .Q(\mem.mem[229][3] ));
 sg13g2_dfrbp_1 _19045_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net642),
    .D(_00688_),
    .Q_N(_08538_),
    .Q(\mem.mem[229][4] ));
 sg13g2_dfrbp_1 _19046_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net641),
    .D(_00689_),
    .Q_N(_08537_),
    .Q(\mem.mem[229][5] ));
 sg13g2_dfrbp_1 _19047_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net640),
    .D(_00690_),
    .Q_N(_08536_),
    .Q(\mem.mem[229][6] ));
 sg13g2_dfrbp_1 _19048_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net690),
    .D(_00691_),
    .Q_N(_09189_),
    .Q(\mem.mem[229][7] ));
 sg13g2_dfrbp_1 _19049_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net691),
    .D(_00013_),
    .Q_N(_09190_),
    .Q(halted));
 sg13g2_dfrbp_1 _19050_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net692),
    .D(_00008_),
    .Q_N(_09191_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 _19051_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net693),
    .D(_00009_),
    .Q_N(_09192_),
    .Q(\state[2] ));
 sg13g2_dfrbp_1 _19052_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net694),
    .D(_00010_),
    .Q_N(_09193_),
    .Q(\state[3] ));
 sg13g2_dfrbp_1 _19053_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net695),
    .D(_00014_),
    .Q_N(_09194_),
    .Q(\state[4] ));
 sg13g2_dfrbp_1 _19054_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net509),
    .D(_00011_),
    .Q_N(_09195_),
    .Q(\state[5] ));
 sg13g2_dfrbp_1 _19055_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net639),
    .D(_00012_),
    .Q_N(_08535_),
    .Q(\state[6] ));
 sg13g2_dfrbp_1 _19056_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net638),
    .D(_00692_),
    .Q_N(_08534_),
    .Q(\mem.mem[219][0] ));
 sg13g2_dfrbp_1 _19057_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net637),
    .D(_00693_),
    .Q_N(_08533_),
    .Q(\mem.mem[219][1] ));
 sg13g2_dfrbp_1 _19058_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net636),
    .D(_00694_),
    .Q_N(_08532_),
    .Q(\mem.mem[219][2] ));
 sg13g2_dfrbp_1 _19059_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net635),
    .D(_00695_),
    .Q_N(_08531_),
    .Q(\mem.mem[219][3] ));
 sg13g2_dfrbp_1 _19060_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net634),
    .D(_00696_),
    .Q_N(_08530_),
    .Q(\mem.mem[219][4] ));
 sg13g2_dfrbp_1 _19061_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net633),
    .D(_00697_),
    .Q_N(_08529_),
    .Q(\mem.mem[219][5] ));
 sg13g2_dfrbp_1 _19062_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net632),
    .D(_00698_),
    .Q_N(_08528_),
    .Q(\mem.mem[219][6] ));
 sg13g2_dfrbp_1 _19063_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net631),
    .D(_00699_),
    .Q_N(_08527_),
    .Q(\mem.mem[219][7] ));
 sg13g2_dfrbp_1 _19064_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net630),
    .D(_00700_),
    .Q_N(_08526_),
    .Q(\mem.mem[209][0] ));
 sg13g2_dfrbp_1 _19065_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net629),
    .D(_00701_),
    .Q_N(_08525_),
    .Q(\mem.mem[209][1] ));
 sg13g2_dfrbp_1 _19066_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net628),
    .D(_00702_),
    .Q_N(_08524_),
    .Q(\mem.mem[209][2] ));
 sg13g2_dfrbp_1 _19067_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net627),
    .D(_00703_),
    .Q_N(_08523_),
    .Q(\mem.mem[209][3] ));
 sg13g2_dfrbp_1 _19068_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net626),
    .D(_00704_),
    .Q_N(_08522_),
    .Q(\mem.mem[209][4] ));
 sg13g2_dfrbp_1 _19069_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net625),
    .D(_00705_),
    .Q_N(_08521_),
    .Q(\mem.mem[209][5] ));
 sg13g2_dfrbp_1 _19070_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net624),
    .D(_00706_),
    .Q_N(_08520_),
    .Q(\mem.mem[209][6] ));
 sg13g2_dfrbp_1 _19071_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net623),
    .D(_00707_),
    .Q_N(_08519_),
    .Q(\mem.mem[209][7] ));
 sg13g2_dfrbp_1 _19072_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net622),
    .D(_00708_),
    .Q_N(_08518_),
    .Q(\mem.mem[199][0] ));
 sg13g2_dfrbp_1 _19073_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net621),
    .D(_00709_),
    .Q_N(_08517_),
    .Q(\mem.mem[199][1] ));
 sg13g2_dfrbp_1 _19074_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net620),
    .D(_00710_),
    .Q_N(_08516_),
    .Q(\mem.mem[199][2] ));
 sg13g2_dfrbp_1 _19075_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net619),
    .D(_00711_),
    .Q_N(_08515_),
    .Q(\mem.mem[199][3] ));
 sg13g2_dfrbp_1 _19076_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net618),
    .D(_00712_),
    .Q_N(_08514_),
    .Q(\mem.mem[199][4] ));
 sg13g2_dfrbp_1 _19077_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net617),
    .D(_00713_),
    .Q_N(_08513_),
    .Q(\mem.mem[199][5] ));
 sg13g2_dfrbp_1 _19078_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net616),
    .D(_00714_),
    .Q_N(_08512_),
    .Q(\mem.mem[199][6] ));
 sg13g2_dfrbp_1 _19079_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net615),
    .D(_00715_),
    .Q_N(_08511_),
    .Q(\mem.mem[199][7] ));
 sg13g2_dfrbp_1 _19080_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net614),
    .D(_00716_),
    .Q_N(_08510_),
    .Q(\mem.mem[189][0] ));
 sg13g2_dfrbp_1 _19081_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net613),
    .D(_00717_),
    .Q_N(_08509_),
    .Q(\mem.mem[189][1] ));
 sg13g2_dfrbp_1 _19082_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net612),
    .D(_00718_),
    .Q_N(_08508_),
    .Q(\mem.mem[189][2] ));
 sg13g2_dfrbp_1 _19083_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net611),
    .D(_00719_),
    .Q_N(_08507_),
    .Q(\mem.mem[189][3] ));
 sg13g2_dfrbp_1 _19084_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net610),
    .D(_00720_),
    .Q_N(_08506_),
    .Q(\mem.mem[189][4] ));
 sg13g2_dfrbp_1 _19085_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net609),
    .D(_00721_),
    .Q_N(_08505_),
    .Q(\mem.mem[189][5] ));
 sg13g2_dfrbp_1 _19086_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net608),
    .D(_00722_),
    .Q_N(_08504_),
    .Q(\mem.mem[189][6] ));
 sg13g2_dfrbp_1 _19087_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net607),
    .D(_00723_),
    .Q_N(_08503_),
    .Q(\mem.mem[189][7] ));
 sg13g2_dfrbp_1 _19088_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net606),
    .D(_00724_),
    .Q_N(_08502_),
    .Q(\mem.mem[49][0] ));
 sg13g2_dfrbp_1 _19089_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net605),
    .D(_00725_),
    .Q_N(_08501_),
    .Q(\mem.mem[49][1] ));
 sg13g2_dfrbp_1 _19090_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net604),
    .D(_00726_),
    .Q_N(_08500_),
    .Q(\mem.mem[49][2] ));
 sg13g2_dfrbp_1 _19091_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net603),
    .D(_00727_),
    .Q_N(_08499_),
    .Q(\mem.mem[49][3] ));
 sg13g2_dfrbp_1 _19092_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net602),
    .D(_00728_),
    .Q_N(_08498_),
    .Q(\mem.mem[49][4] ));
 sg13g2_dfrbp_1 _19093_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net601),
    .D(_00729_),
    .Q_N(_08497_),
    .Q(\mem.mem[49][5] ));
 sg13g2_dfrbp_1 _19094_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net600),
    .D(_00730_),
    .Q_N(_08496_),
    .Q(\mem.mem[49][6] ));
 sg13g2_dfrbp_1 _19095_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net599),
    .D(_00731_),
    .Q_N(_08495_),
    .Q(\mem.mem[49][7] ));
 sg13g2_dfrbp_1 _19096_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net598),
    .D(_00732_),
    .Q_N(_08494_),
    .Q(\mem.mem[39][0] ));
 sg13g2_dfrbp_1 _19097_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net597),
    .D(_00733_),
    .Q_N(_08493_),
    .Q(\mem.mem[39][1] ));
 sg13g2_dfrbp_1 _19098_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net596),
    .D(_00734_),
    .Q_N(_08492_),
    .Q(\mem.mem[39][2] ));
 sg13g2_dfrbp_1 _19099_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net595),
    .D(_00735_),
    .Q_N(_08491_),
    .Q(\mem.mem[39][3] ));
 sg13g2_dfrbp_1 _19100_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net594),
    .D(_00736_),
    .Q_N(_08490_),
    .Q(\mem.mem[39][4] ));
 sg13g2_dfrbp_1 _19101_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net593),
    .D(_00737_),
    .Q_N(_08489_),
    .Q(\mem.mem[39][5] ));
 sg13g2_dfrbp_1 _19102_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net592),
    .D(_00738_),
    .Q_N(_08488_),
    .Q(\mem.mem[39][6] ));
 sg13g2_dfrbp_1 _19103_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net591),
    .D(_00739_),
    .Q_N(_08487_),
    .Q(\mem.mem[39][7] ));
 sg13g2_dfrbp_1 _19104_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net590),
    .D(_00740_),
    .Q_N(_08486_),
    .Q(\mem.mem[179][0] ));
 sg13g2_dfrbp_1 _19105_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net589),
    .D(_00741_),
    .Q_N(_08485_),
    .Q(\mem.mem[179][1] ));
 sg13g2_dfrbp_1 _19106_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net588),
    .D(_00742_),
    .Q_N(_08484_),
    .Q(\mem.mem[179][2] ));
 sg13g2_dfrbp_1 _19107_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net587),
    .D(_00743_),
    .Q_N(_08483_),
    .Q(\mem.mem[179][3] ));
 sg13g2_dfrbp_1 _19108_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net586),
    .D(_00744_),
    .Q_N(_08482_),
    .Q(\mem.mem[179][4] ));
 sg13g2_dfrbp_1 _19109_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net585),
    .D(_00745_),
    .Q_N(_08481_),
    .Q(\mem.mem[179][5] ));
 sg13g2_dfrbp_1 _19110_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net584),
    .D(_00746_),
    .Q_N(_08480_),
    .Q(\mem.mem[179][6] ));
 sg13g2_dfrbp_1 _19111_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net583),
    .D(_00747_),
    .Q_N(_08479_),
    .Q(\mem.mem[179][7] ));
 sg13g2_dfrbp_1 _19112_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net582),
    .D(_00748_),
    .Q_N(_08478_),
    .Q(\mem.mem[29][0] ));
 sg13g2_dfrbp_1 _19113_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net581),
    .D(_00749_),
    .Q_N(_08477_),
    .Q(\mem.mem[29][1] ));
 sg13g2_dfrbp_1 _19114_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net580),
    .D(_00750_),
    .Q_N(_08476_),
    .Q(\mem.mem[29][2] ));
 sg13g2_dfrbp_1 _19115_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net579),
    .D(_00751_),
    .Q_N(_08475_),
    .Q(\mem.mem[29][3] ));
 sg13g2_dfrbp_1 _19116_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net578),
    .D(_00752_),
    .Q_N(_08474_),
    .Q(\mem.mem[29][4] ));
 sg13g2_dfrbp_1 _19117_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net577),
    .D(_00753_),
    .Q_N(_08473_),
    .Q(\mem.mem[29][5] ));
 sg13g2_dfrbp_1 _19118_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net576),
    .D(_00754_),
    .Q_N(_08472_),
    .Q(\mem.mem[29][6] ));
 sg13g2_dfrbp_1 _19119_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net575),
    .D(_00755_),
    .Q_N(_08471_),
    .Q(\mem.mem[29][7] ));
 sg13g2_dfrbp_1 _19120_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net574),
    .D(_00756_),
    .Q_N(_08470_),
    .Q(\mem.mem[169][0] ));
 sg13g2_dfrbp_1 _19121_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net573),
    .D(_00757_),
    .Q_N(_08469_),
    .Q(\mem.mem[169][1] ));
 sg13g2_dfrbp_1 _19122_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net572),
    .D(_00758_),
    .Q_N(_08468_),
    .Q(\mem.mem[169][2] ));
 sg13g2_dfrbp_1 _19123_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net571),
    .D(_00759_),
    .Q_N(_08467_),
    .Q(\mem.mem[169][3] ));
 sg13g2_dfrbp_1 _19124_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net570),
    .D(_00760_),
    .Q_N(_08466_),
    .Q(\mem.mem[169][4] ));
 sg13g2_dfrbp_1 _19125_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net569),
    .D(_00761_),
    .Q_N(_08465_),
    .Q(\mem.mem[169][5] ));
 sg13g2_dfrbp_1 _19126_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net568),
    .D(_00762_),
    .Q_N(_08464_),
    .Q(\mem.mem[169][6] ));
 sg13g2_dfrbp_1 _19127_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net567),
    .D(_00763_),
    .Q_N(_08463_),
    .Q(\mem.mem[169][7] ));
 sg13g2_dfrbp_1 _19128_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net566),
    .D(_00764_),
    .Q_N(_08462_),
    .Q(\mem.mem[159][0] ));
 sg13g2_dfrbp_1 _19129_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net565),
    .D(_00765_),
    .Q_N(_08461_),
    .Q(\mem.mem[159][1] ));
 sg13g2_dfrbp_1 _19130_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net564),
    .D(_00766_),
    .Q_N(_08460_),
    .Q(\mem.mem[159][2] ));
 sg13g2_dfrbp_1 _19131_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net563),
    .D(_00767_),
    .Q_N(_08459_),
    .Q(\mem.mem[159][3] ));
 sg13g2_dfrbp_1 _19132_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net562),
    .D(_00768_),
    .Q_N(_08458_),
    .Q(\mem.mem[159][4] ));
 sg13g2_dfrbp_1 _19133_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net561),
    .D(_00769_),
    .Q_N(_08457_),
    .Q(\mem.mem[159][5] ));
 sg13g2_dfrbp_1 _19134_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net560),
    .D(_00770_),
    .Q_N(_08456_),
    .Q(\mem.mem[159][6] ));
 sg13g2_dfrbp_1 _19135_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net559),
    .D(_00771_),
    .Q_N(_08455_),
    .Q(\mem.mem[159][7] ));
 sg13g2_dfrbp_1 _19136_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net558),
    .D(_00772_),
    .Q_N(_08454_),
    .Q(\mem.mem[91][0] ));
 sg13g2_dfrbp_1 _19137_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net557),
    .D(_00773_),
    .Q_N(_08453_),
    .Q(\mem.mem[91][1] ));
 sg13g2_dfrbp_1 _19138_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net556),
    .D(_00774_),
    .Q_N(_08452_),
    .Q(\mem.mem[91][2] ));
 sg13g2_dfrbp_1 _19139_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net555),
    .D(_00775_),
    .Q_N(_08451_),
    .Q(\mem.mem[91][3] ));
 sg13g2_dfrbp_1 _19140_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net554),
    .D(_00776_),
    .Q_N(_08450_),
    .Q(\mem.mem[91][4] ));
 sg13g2_dfrbp_1 _19141_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net553),
    .D(_00777_),
    .Q_N(_08449_),
    .Q(\mem.mem[91][5] ));
 sg13g2_dfrbp_1 _19142_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net552),
    .D(_00778_),
    .Q_N(_08448_),
    .Q(\mem.mem[91][6] ));
 sg13g2_dfrbp_1 _19143_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net551),
    .D(_00779_),
    .Q_N(_08447_),
    .Q(\mem.mem[91][7] ));
 sg13g2_dfrbp_1 _19144_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net550),
    .D(_00780_),
    .Q_N(_08446_),
    .Q(\mem.mem[90][0] ));
 sg13g2_dfrbp_1 _19145_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net549),
    .D(_00781_),
    .Q_N(_08445_),
    .Q(\mem.mem[90][1] ));
 sg13g2_dfrbp_1 _19146_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net548),
    .D(_00782_),
    .Q_N(_08444_),
    .Q(\mem.mem[90][2] ));
 sg13g2_dfrbp_1 _19147_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net547),
    .D(_00783_),
    .Q_N(_08443_),
    .Q(\mem.mem[90][3] ));
 sg13g2_dfrbp_1 _19148_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net546),
    .D(_00784_),
    .Q_N(_08442_),
    .Q(\mem.mem[90][4] ));
 sg13g2_dfrbp_1 _19149_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net545),
    .D(_00785_),
    .Q_N(_08441_),
    .Q(\mem.mem[90][5] ));
 sg13g2_dfrbp_1 _19150_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net544),
    .D(_00786_),
    .Q_N(_08440_),
    .Q(\mem.mem[90][6] ));
 sg13g2_dfrbp_1 _19151_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net543),
    .D(_00787_),
    .Q_N(_08439_),
    .Q(\mem.mem[90][7] ));
 sg13g2_dfrbp_1 _19152_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net542),
    .D(_00788_),
    .Q_N(_08438_),
    .Q(\mem.mem[8][0] ));
 sg13g2_dfrbp_1 _19153_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net541),
    .D(_00789_),
    .Q_N(_08437_),
    .Q(\mem.mem[8][1] ));
 sg13g2_dfrbp_1 _19154_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net540),
    .D(_00790_),
    .Q_N(_08436_),
    .Q(\mem.mem[8][2] ));
 sg13g2_dfrbp_1 _19155_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net539),
    .D(_00791_),
    .Q_N(_08435_),
    .Q(\mem.mem[8][3] ));
 sg13g2_dfrbp_1 _19156_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net538),
    .D(_00792_),
    .Q_N(_08434_),
    .Q(\mem.mem[8][4] ));
 sg13g2_dfrbp_1 _19157_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net537),
    .D(_00793_),
    .Q_N(_08433_),
    .Q(\mem.mem[8][5] ));
 sg13g2_dfrbp_1 _19158_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net536),
    .D(_00794_),
    .Q_N(_08432_),
    .Q(\mem.mem[8][6] ));
 sg13g2_dfrbp_1 _19159_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net535),
    .D(_00795_),
    .Q_N(_08431_),
    .Q(\mem.mem[8][7] ));
 sg13g2_dfrbp_1 _19160_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net534),
    .D(_00796_),
    .Q_N(_08430_),
    .Q(\mem.mem[44][0] ));
 sg13g2_dfrbp_1 _19161_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net533),
    .D(_00797_),
    .Q_N(_08429_),
    .Q(\mem.mem[44][1] ));
 sg13g2_dfrbp_1 _19162_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net532),
    .D(_00798_),
    .Q_N(_08428_),
    .Q(\mem.mem[44][2] ));
 sg13g2_dfrbp_1 _19163_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net531),
    .D(_00799_),
    .Q_N(_08427_),
    .Q(\mem.mem[44][3] ));
 sg13g2_dfrbp_1 _19164_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net530),
    .D(_00800_),
    .Q_N(_08426_),
    .Q(\mem.mem[44][4] ));
 sg13g2_dfrbp_1 _19165_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net529),
    .D(_00801_),
    .Q_N(_08425_),
    .Q(\mem.mem[44][5] ));
 sg13g2_dfrbp_1 _19166_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net528),
    .D(_00802_),
    .Q_N(_08424_),
    .Q(\mem.mem[44][6] ));
 sg13g2_dfrbp_1 _19167_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net527),
    .D(_00803_),
    .Q_N(_08423_),
    .Q(\mem.mem[44][7] ));
 sg13g2_dfrbp_1 _19168_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net526),
    .D(net2139),
    .Q_N(_08422_),
    .Q(\mem.out_strobe ));
 sg13g2_dfrbp_1 _19169_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net524),
    .D(net4249),
    .Q_N(_08421_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _19170_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net522),
    .D(_00806_),
    .Q_N(_08420_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _19171_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net520),
    .D(_00807_),
    .Q_N(_08419_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _19172_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net518),
    .D(_00808_),
    .Q_N(_08418_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _19173_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net516),
    .D(_00809_),
    .Q_N(_08417_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _19174_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net514),
    .D(_00810_),
    .Q_N(_08416_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _19175_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net512),
    .D(_00811_),
    .Q_N(_08415_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _19176_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net510),
    .D(_00812_),
    .Q_N(_08414_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _19177_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net508),
    .D(_00813_),
    .Q_N(_08413_),
    .Q(\mem.mem[19][0] ));
 sg13g2_dfrbp_1 _19178_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net507),
    .D(_00814_),
    .Q_N(_08412_),
    .Q(\mem.mem[19][1] ));
 sg13g2_dfrbp_1 _19179_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net506),
    .D(_00815_),
    .Q_N(_08411_),
    .Q(\mem.mem[19][2] ));
 sg13g2_dfrbp_1 _19180_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net505),
    .D(_00816_),
    .Q_N(_08410_),
    .Q(\mem.mem[19][3] ));
 sg13g2_dfrbp_1 _19181_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net504),
    .D(_00817_),
    .Q_N(_08409_),
    .Q(\mem.mem[19][4] ));
 sg13g2_dfrbp_1 _19182_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net503),
    .D(_00818_),
    .Q_N(_08408_),
    .Q(\mem.mem[19][5] ));
 sg13g2_dfrbp_1 _19183_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net502),
    .D(_00819_),
    .Q_N(_08407_),
    .Q(\mem.mem[19][6] ));
 sg13g2_dfrbp_1 _19184_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net501),
    .D(_00820_),
    .Q_N(_08406_),
    .Q(\mem.mem[19][7] ));
 sg13g2_dfrbp_1 _19185_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net500),
    .D(_00821_),
    .Q_N(_08405_),
    .Q(\mem.mem[89][0] ));
 sg13g2_dfrbp_1 _19186_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net499),
    .D(_00822_),
    .Q_N(_08404_),
    .Q(\mem.mem[89][1] ));
 sg13g2_dfrbp_1 _19187_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net498),
    .D(_00823_),
    .Q_N(_08403_),
    .Q(\mem.mem[89][2] ));
 sg13g2_dfrbp_1 _19188_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net497),
    .D(_00824_),
    .Q_N(_08402_),
    .Q(\mem.mem[89][3] ));
 sg13g2_dfrbp_1 _19189_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net496),
    .D(_00825_),
    .Q_N(_08401_),
    .Q(\mem.mem[89][4] ));
 sg13g2_dfrbp_1 _19190_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net495),
    .D(_00826_),
    .Q_N(_08400_),
    .Q(\mem.mem[89][5] ));
 sg13g2_dfrbp_1 _19191_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net494),
    .D(_00827_),
    .Q_N(_08399_),
    .Q(\mem.mem[89][6] ));
 sg13g2_dfrbp_1 _19192_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net493),
    .D(_00828_),
    .Q_N(_08398_),
    .Q(\mem.mem[89][7] ));
 sg13g2_dfrbp_1 _19193_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net492),
    .D(_00829_),
    .Q_N(_08397_),
    .Q(\mem.mem[79][0] ));
 sg13g2_dfrbp_1 _19194_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net491),
    .D(_00830_),
    .Q_N(_08396_),
    .Q(\mem.mem[79][1] ));
 sg13g2_dfrbp_1 _19195_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net490),
    .D(_00831_),
    .Q_N(_08395_),
    .Q(\mem.mem[79][2] ));
 sg13g2_dfrbp_1 _19196_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net489),
    .D(_00832_),
    .Q_N(_08394_),
    .Q(\mem.mem[79][3] ));
 sg13g2_dfrbp_1 _19197_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net488),
    .D(_00833_),
    .Q_N(_08393_),
    .Q(\mem.mem[79][4] ));
 sg13g2_dfrbp_1 _19198_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net487),
    .D(_00834_),
    .Q_N(_08392_),
    .Q(\mem.mem[79][5] ));
 sg13g2_dfrbp_1 _19199_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net486),
    .D(_00835_),
    .Q_N(_08391_),
    .Q(\mem.mem[79][6] ));
 sg13g2_dfrbp_1 _19200_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net485),
    .D(_00836_),
    .Q_N(_08390_),
    .Q(\mem.mem[79][7] ));
 sg13g2_dfrbp_1 _19201_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net484),
    .D(_00837_),
    .Q_N(_08389_),
    .Q(\mem.mem[92][0] ));
 sg13g2_dfrbp_1 _19202_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net483),
    .D(_00838_),
    .Q_N(_08388_),
    .Q(\mem.mem[92][1] ));
 sg13g2_dfrbp_1 _19203_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net482),
    .D(_00839_),
    .Q_N(_08387_),
    .Q(\mem.mem[92][2] ));
 sg13g2_dfrbp_1 _19204_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net481),
    .D(_00840_),
    .Q_N(_08386_),
    .Q(\mem.mem[92][3] ));
 sg13g2_dfrbp_1 _19205_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net480),
    .D(_00841_),
    .Q_N(_08385_),
    .Q(\mem.mem[92][4] ));
 sg13g2_dfrbp_1 _19206_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net479),
    .D(_00842_),
    .Q_N(_08384_),
    .Q(\mem.mem[92][5] ));
 sg13g2_dfrbp_1 _19207_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net478),
    .D(_00843_),
    .Q_N(_08383_),
    .Q(\mem.mem[92][6] ));
 sg13g2_dfrbp_1 _19208_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net477),
    .D(_00844_),
    .Q_N(_08382_),
    .Q(\mem.mem[92][7] ));
 sg13g2_dfrbp_1 _19209_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net476),
    .D(_00845_),
    .Q_N(_08381_),
    .Q(\mem.mem[93][0] ));
 sg13g2_dfrbp_1 _19210_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net475),
    .D(_00846_),
    .Q_N(_08380_),
    .Q(\mem.mem[93][1] ));
 sg13g2_dfrbp_1 _19211_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net474),
    .D(_00847_),
    .Q_N(_08379_),
    .Q(\mem.mem[93][2] ));
 sg13g2_dfrbp_1 _19212_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net473),
    .D(_00848_),
    .Q_N(_08378_),
    .Q(\mem.mem[93][3] ));
 sg13g2_dfrbp_1 _19213_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net472),
    .D(_00849_),
    .Q_N(_08377_),
    .Q(\mem.mem[93][4] ));
 sg13g2_dfrbp_1 _19214_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net471),
    .D(_00850_),
    .Q_N(_08376_),
    .Q(\mem.mem[93][5] ));
 sg13g2_dfrbp_1 _19215_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net470),
    .D(_00851_),
    .Q_N(_08375_),
    .Q(\mem.mem[93][6] ));
 sg13g2_dfrbp_1 _19216_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net469),
    .D(_00852_),
    .Q_N(_08374_),
    .Q(\mem.mem[93][7] ));
 sg13g2_dfrbp_1 _19217_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net468),
    .D(_00853_),
    .Q_N(_08373_),
    .Q(\mem.mem[94][0] ));
 sg13g2_dfrbp_1 _19218_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net467),
    .D(_00854_),
    .Q_N(_08372_),
    .Q(\mem.mem[94][1] ));
 sg13g2_dfrbp_1 _19219_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net466),
    .D(_00855_),
    .Q_N(_08371_),
    .Q(\mem.mem[94][2] ));
 sg13g2_dfrbp_1 _19220_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net465),
    .D(_00856_),
    .Q_N(_08370_),
    .Q(\mem.mem[94][3] ));
 sg13g2_dfrbp_1 _19221_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net464),
    .D(_00857_),
    .Q_N(_08369_),
    .Q(\mem.mem[94][4] ));
 sg13g2_dfrbp_1 _19222_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net463),
    .D(_00858_),
    .Q_N(_08368_),
    .Q(\mem.mem[94][5] ));
 sg13g2_dfrbp_1 _19223_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net462),
    .D(_00859_),
    .Q_N(_08367_),
    .Q(\mem.mem[94][6] ));
 sg13g2_dfrbp_1 _19224_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net461),
    .D(_00860_),
    .Q_N(_08366_),
    .Q(\mem.mem[94][7] ));
 sg13g2_dfrbp_1 _19225_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net460),
    .D(_00861_),
    .Q_N(_08365_),
    .Q(\mem.mem[95][0] ));
 sg13g2_dfrbp_1 _19226_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net459),
    .D(_00862_),
    .Q_N(_08364_),
    .Q(\mem.mem[95][1] ));
 sg13g2_dfrbp_1 _19227_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net458),
    .D(_00863_),
    .Q_N(_08363_),
    .Q(\mem.mem[95][2] ));
 sg13g2_dfrbp_1 _19228_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net457),
    .D(_00864_),
    .Q_N(_08362_),
    .Q(\mem.mem[95][3] ));
 sg13g2_dfrbp_1 _19229_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net456),
    .D(_00865_),
    .Q_N(_08361_),
    .Q(\mem.mem[95][4] ));
 sg13g2_dfrbp_1 _19230_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net455),
    .D(_00866_),
    .Q_N(_08360_),
    .Q(\mem.mem[95][5] ));
 sg13g2_dfrbp_1 _19231_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net454),
    .D(_00867_),
    .Q_N(_08359_),
    .Q(\mem.mem[95][6] ));
 sg13g2_dfrbp_1 _19232_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net453),
    .D(_00868_),
    .Q_N(_08358_),
    .Q(\mem.mem[95][7] ));
 sg13g2_dfrbp_1 _19233_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net452),
    .D(_00869_),
    .Q_N(_08357_),
    .Q(\mem.mem[96][0] ));
 sg13g2_dfrbp_1 _19234_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net451),
    .D(_00870_),
    .Q_N(_08356_),
    .Q(\mem.mem[96][1] ));
 sg13g2_dfrbp_1 _19235_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net450),
    .D(_00871_),
    .Q_N(_08355_),
    .Q(\mem.mem[96][2] ));
 sg13g2_dfrbp_1 _19236_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net449),
    .D(_00872_),
    .Q_N(_08354_),
    .Q(\mem.mem[96][3] ));
 sg13g2_dfrbp_1 _19237_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net448),
    .D(_00873_),
    .Q_N(_08353_),
    .Q(\mem.mem[96][4] ));
 sg13g2_dfrbp_1 _19238_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net447),
    .D(_00874_),
    .Q_N(_08352_),
    .Q(\mem.mem[96][5] ));
 sg13g2_dfrbp_1 _19239_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net446),
    .D(_00875_),
    .Q_N(_08351_),
    .Q(\mem.mem[96][6] ));
 sg13g2_dfrbp_1 _19240_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net445),
    .D(_00876_),
    .Q_N(_08350_),
    .Q(\mem.mem[96][7] ));
 sg13g2_dfrbp_1 _19241_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net444),
    .D(_00877_),
    .Q_N(_08349_),
    .Q(\mem.mem[97][0] ));
 sg13g2_dfrbp_1 _19242_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net443),
    .D(_00878_),
    .Q_N(_08348_),
    .Q(\mem.mem[97][1] ));
 sg13g2_dfrbp_1 _19243_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net442),
    .D(_00879_),
    .Q_N(_08347_),
    .Q(\mem.mem[97][2] ));
 sg13g2_dfrbp_1 _19244_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net441),
    .D(_00880_),
    .Q_N(_08346_),
    .Q(\mem.mem[97][3] ));
 sg13g2_dfrbp_1 _19245_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net440),
    .D(_00881_),
    .Q_N(_08345_),
    .Q(\mem.mem[97][4] ));
 sg13g2_dfrbp_1 _19246_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net439),
    .D(_00882_),
    .Q_N(_08344_),
    .Q(\mem.mem[97][5] ));
 sg13g2_dfrbp_1 _19247_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net438),
    .D(_00883_),
    .Q_N(_08343_),
    .Q(\mem.mem[97][6] ));
 sg13g2_dfrbp_1 _19248_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net437),
    .D(_00884_),
    .Q_N(_08342_),
    .Q(\mem.mem[97][7] ));
 sg13g2_dfrbp_1 _19249_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net436),
    .D(_00885_),
    .Q_N(_08341_),
    .Q(\mem.mem[98][0] ));
 sg13g2_dfrbp_1 _19250_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net435),
    .D(_00886_),
    .Q_N(_08340_),
    .Q(\mem.mem[98][1] ));
 sg13g2_dfrbp_1 _19251_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net434),
    .D(_00887_),
    .Q_N(_08339_),
    .Q(\mem.mem[98][2] ));
 sg13g2_dfrbp_1 _19252_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net433),
    .D(_00888_),
    .Q_N(_08338_),
    .Q(\mem.mem[98][3] ));
 sg13g2_dfrbp_1 _19253_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net432),
    .D(_00889_),
    .Q_N(_08337_),
    .Q(\mem.mem[98][4] ));
 sg13g2_dfrbp_1 _19254_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net431),
    .D(_00890_),
    .Q_N(_08336_),
    .Q(\mem.mem[98][5] ));
 sg13g2_dfrbp_1 _19255_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net430),
    .D(_00891_),
    .Q_N(_08335_),
    .Q(\mem.mem[98][6] ));
 sg13g2_dfrbp_1 _19256_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net429),
    .D(_00892_),
    .Q_N(_08334_),
    .Q(\mem.mem[98][7] ));
 sg13g2_dfrbp_1 _19257_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net428),
    .D(_00893_),
    .Q_N(_08333_),
    .Q(\mem.mem[0][0] ));
 sg13g2_dfrbp_1 _19258_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net427),
    .D(_00894_),
    .Q_N(_08332_),
    .Q(\mem.mem[0][1] ));
 sg13g2_dfrbp_1 _19259_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net426),
    .D(_00895_),
    .Q_N(_08331_),
    .Q(\mem.mem[0][2] ));
 sg13g2_dfrbp_1 _19260_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net425),
    .D(_00896_),
    .Q_N(_08330_),
    .Q(\mem.mem[0][3] ));
 sg13g2_dfrbp_1 _19261_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net424),
    .D(_00897_),
    .Q_N(_08329_),
    .Q(\mem.mem[0][4] ));
 sg13g2_dfrbp_1 _19262_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net423),
    .D(_00898_),
    .Q_N(_08328_),
    .Q(\mem.mem[0][5] ));
 sg13g2_dfrbp_1 _19263_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net422),
    .D(_00899_),
    .Q_N(_08327_),
    .Q(\mem.mem[0][6] ));
 sg13g2_dfrbp_1 _19264_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net421),
    .D(_00900_),
    .Q_N(_08326_),
    .Q(\mem.mem[0][7] ));
 sg13g2_dfrbp_1 _19265_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net420),
    .D(_00901_),
    .Q_N(_08325_),
    .Q(\mem.mem[100][0] ));
 sg13g2_dfrbp_1 _19266_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net419),
    .D(_00902_),
    .Q_N(_08324_),
    .Q(\mem.mem[100][1] ));
 sg13g2_dfrbp_1 _19267_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net418),
    .D(_00903_),
    .Q_N(_08323_),
    .Q(\mem.mem[100][2] ));
 sg13g2_dfrbp_1 _19268_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net417),
    .D(_00904_),
    .Q_N(_08322_),
    .Q(\mem.mem[100][3] ));
 sg13g2_dfrbp_1 _19269_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net416),
    .D(_00905_),
    .Q_N(_08321_),
    .Q(\mem.mem[100][4] ));
 sg13g2_dfrbp_1 _19270_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net415),
    .D(_00906_),
    .Q_N(_08320_),
    .Q(\mem.mem[100][5] ));
 sg13g2_dfrbp_1 _19271_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net414),
    .D(_00907_),
    .Q_N(_08319_),
    .Q(\mem.mem[100][6] ));
 sg13g2_dfrbp_1 _19272_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net413),
    .D(_00908_),
    .Q_N(_08318_),
    .Q(\mem.mem[100][7] ));
 sg13g2_dfrbp_1 _19273_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net412),
    .D(_00909_),
    .Q_N(_08317_),
    .Q(\mem.mem[101][0] ));
 sg13g2_dfrbp_1 _19274_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net411),
    .D(_00910_),
    .Q_N(_08316_),
    .Q(\mem.mem[101][1] ));
 sg13g2_dfrbp_1 _19275_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net410),
    .D(_00911_),
    .Q_N(_08315_),
    .Q(\mem.mem[101][2] ));
 sg13g2_dfrbp_1 _19276_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net409),
    .D(_00912_),
    .Q_N(_08314_),
    .Q(\mem.mem[101][3] ));
 sg13g2_dfrbp_1 _19277_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net408),
    .D(_00913_),
    .Q_N(_08313_),
    .Q(\mem.mem[101][4] ));
 sg13g2_dfrbp_1 _19278_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net407),
    .D(_00914_),
    .Q_N(_08312_),
    .Q(\mem.mem[101][5] ));
 sg13g2_dfrbp_1 _19279_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net406),
    .D(_00915_),
    .Q_N(_08311_),
    .Q(\mem.mem[101][6] ));
 sg13g2_dfrbp_1 _19280_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net405),
    .D(_00916_),
    .Q_N(_08310_),
    .Q(\mem.mem[101][7] ));
 sg13g2_dfrbp_1 _19281_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net404),
    .D(_00917_),
    .Q_N(_08309_),
    .Q(\mem.mem[102][0] ));
 sg13g2_dfrbp_1 _19282_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net403),
    .D(_00918_),
    .Q_N(_08308_),
    .Q(\mem.mem[102][1] ));
 sg13g2_dfrbp_1 _19283_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net402),
    .D(_00919_),
    .Q_N(_08307_),
    .Q(\mem.mem[102][2] ));
 sg13g2_dfrbp_1 _19284_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net401),
    .D(_00920_),
    .Q_N(_08306_),
    .Q(\mem.mem[102][3] ));
 sg13g2_dfrbp_1 _19285_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net400),
    .D(_00921_),
    .Q_N(_08305_),
    .Q(\mem.mem[102][4] ));
 sg13g2_dfrbp_1 _19286_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net399),
    .D(_00922_),
    .Q_N(_08304_),
    .Q(\mem.mem[102][5] ));
 sg13g2_dfrbp_1 _19287_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net398),
    .D(_00923_),
    .Q_N(_08303_),
    .Q(\mem.mem[102][6] ));
 sg13g2_dfrbp_1 _19288_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net397),
    .D(_00924_),
    .Q_N(_08302_),
    .Q(\mem.mem[102][7] ));
 sg13g2_dfrbp_1 _19289_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net396),
    .D(_00925_),
    .Q_N(_08301_),
    .Q(\mem.mem[103][0] ));
 sg13g2_dfrbp_1 _19290_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net395),
    .D(_00926_),
    .Q_N(_08300_),
    .Q(\mem.mem[103][1] ));
 sg13g2_dfrbp_1 _19291_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net394),
    .D(_00927_),
    .Q_N(_08299_),
    .Q(\mem.mem[103][2] ));
 sg13g2_dfrbp_1 _19292_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net393),
    .D(_00928_),
    .Q_N(_08298_),
    .Q(\mem.mem[103][3] ));
 sg13g2_dfrbp_1 _19293_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net392),
    .D(_00929_),
    .Q_N(_08297_),
    .Q(\mem.mem[103][4] ));
 sg13g2_dfrbp_1 _19294_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net391),
    .D(_00930_),
    .Q_N(_08296_),
    .Q(\mem.mem[103][5] ));
 sg13g2_dfrbp_1 _19295_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net390),
    .D(_00931_),
    .Q_N(_08295_),
    .Q(\mem.mem[103][6] ));
 sg13g2_dfrbp_1 _19296_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net389),
    .D(_00932_),
    .Q_N(_08294_),
    .Q(\mem.mem[103][7] ));
 sg13g2_dfrbp_1 _19297_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net388),
    .D(_00933_),
    .Q_N(_08293_),
    .Q(\mem.mem[104][0] ));
 sg13g2_dfrbp_1 _19298_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net387),
    .D(_00934_),
    .Q_N(_08292_),
    .Q(\mem.mem[104][1] ));
 sg13g2_dfrbp_1 _19299_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net386),
    .D(_00935_),
    .Q_N(_08291_),
    .Q(\mem.mem[104][2] ));
 sg13g2_dfrbp_1 _19300_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net385),
    .D(_00936_),
    .Q_N(_08290_),
    .Q(\mem.mem[104][3] ));
 sg13g2_dfrbp_1 _19301_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net384),
    .D(_00937_),
    .Q_N(_08289_),
    .Q(\mem.mem[104][4] ));
 sg13g2_dfrbp_1 _19302_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net383),
    .D(_00938_),
    .Q_N(_08288_),
    .Q(\mem.mem[104][5] ));
 sg13g2_dfrbp_1 _19303_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net382),
    .D(_00939_),
    .Q_N(_08287_),
    .Q(\mem.mem[104][6] ));
 sg13g2_dfrbp_1 _19304_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net381),
    .D(_00940_),
    .Q_N(_08286_),
    .Q(\mem.mem[104][7] ));
 sg13g2_dfrbp_1 _19305_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net380),
    .D(_00941_),
    .Q_N(_08285_),
    .Q(\mem.mem[105][0] ));
 sg13g2_dfrbp_1 _19306_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net379),
    .D(_00942_),
    .Q_N(_08284_),
    .Q(\mem.mem[105][1] ));
 sg13g2_dfrbp_1 _19307_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net378),
    .D(_00943_),
    .Q_N(_08283_),
    .Q(\mem.mem[105][2] ));
 sg13g2_dfrbp_1 _19308_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net377),
    .D(_00944_),
    .Q_N(_08282_),
    .Q(\mem.mem[105][3] ));
 sg13g2_dfrbp_1 _19309_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net376),
    .D(_00945_),
    .Q_N(_08281_),
    .Q(\mem.mem[105][4] ));
 sg13g2_dfrbp_1 _19310_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net375),
    .D(_00946_),
    .Q_N(_08280_),
    .Q(\mem.mem[105][5] ));
 sg13g2_dfrbp_1 _19311_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net374),
    .D(_00947_),
    .Q_N(_08279_),
    .Q(\mem.mem[105][6] ));
 sg13g2_dfrbp_1 _19312_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net373),
    .D(_00948_),
    .Q_N(_08278_),
    .Q(\mem.mem[105][7] ));
 sg13g2_dfrbp_1 _19313_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net372),
    .D(_00949_),
    .Q_N(_08277_),
    .Q(\mem.mem[106][0] ));
 sg13g2_dfrbp_1 _19314_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net371),
    .D(_00950_),
    .Q_N(_08276_),
    .Q(\mem.mem[106][1] ));
 sg13g2_dfrbp_1 _19315_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net370),
    .D(_00951_),
    .Q_N(_08275_),
    .Q(\mem.mem[106][2] ));
 sg13g2_dfrbp_1 _19316_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net369),
    .D(_00952_),
    .Q_N(_08274_),
    .Q(\mem.mem[106][3] ));
 sg13g2_dfrbp_1 _19317_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net368),
    .D(_00953_),
    .Q_N(_08273_),
    .Q(\mem.mem[106][4] ));
 sg13g2_dfrbp_1 _19318_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net367),
    .D(_00954_),
    .Q_N(_08272_),
    .Q(\mem.mem[106][5] ));
 sg13g2_dfrbp_1 _19319_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net366),
    .D(_00955_),
    .Q_N(_08271_),
    .Q(\mem.mem[106][6] ));
 sg13g2_dfrbp_1 _19320_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net365),
    .D(_00956_),
    .Q_N(_08270_),
    .Q(\mem.mem[106][7] ));
 sg13g2_dfrbp_1 _19321_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net364),
    .D(_00957_),
    .Q_N(_08269_),
    .Q(\mem.mem[107][0] ));
 sg13g2_dfrbp_1 _19322_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net363),
    .D(_00958_),
    .Q_N(_08268_),
    .Q(\mem.mem[107][1] ));
 sg13g2_dfrbp_1 _19323_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net362),
    .D(_00959_),
    .Q_N(_08267_),
    .Q(\mem.mem[107][2] ));
 sg13g2_dfrbp_1 _19324_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net361),
    .D(_00960_),
    .Q_N(_08266_),
    .Q(\mem.mem[107][3] ));
 sg13g2_dfrbp_1 _19325_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net360),
    .D(_00961_),
    .Q_N(_08265_),
    .Q(\mem.mem[107][4] ));
 sg13g2_dfrbp_1 _19326_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net359),
    .D(_00962_),
    .Q_N(_08264_),
    .Q(\mem.mem[107][5] ));
 sg13g2_dfrbp_1 _19327_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net358),
    .D(_00963_),
    .Q_N(_08263_),
    .Q(\mem.mem[107][6] ));
 sg13g2_dfrbp_1 _19328_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net357),
    .D(_00964_),
    .Q_N(_08262_),
    .Q(\mem.mem[107][7] ));
 sg13g2_dfrbp_1 _19329_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net356),
    .D(_00965_),
    .Q_N(_08261_),
    .Q(\mem.mem[108][0] ));
 sg13g2_dfrbp_1 _19330_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net355),
    .D(_00966_),
    .Q_N(_08260_),
    .Q(\mem.mem[108][1] ));
 sg13g2_dfrbp_1 _19331_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net354),
    .D(_00967_),
    .Q_N(_08259_),
    .Q(\mem.mem[108][2] ));
 sg13g2_dfrbp_1 _19332_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net353),
    .D(_00968_),
    .Q_N(_08258_),
    .Q(\mem.mem[108][3] ));
 sg13g2_dfrbp_1 _19333_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net352),
    .D(_00969_),
    .Q_N(_08257_),
    .Q(\mem.mem[108][4] ));
 sg13g2_dfrbp_1 _19334_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net351),
    .D(_00970_),
    .Q_N(_08256_),
    .Q(\mem.mem[108][5] ));
 sg13g2_dfrbp_1 _19335_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net350),
    .D(_00971_),
    .Q_N(_08255_),
    .Q(\mem.mem[108][6] ));
 sg13g2_dfrbp_1 _19336_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net349),
    .D(_00972_),
    .Q_N(_08254_),
    .Q(\mem.mem[108][7] ));
 sg13g2_dfrbp_1 _19337_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net348),
    .D(_00973_),
    .Q_N(_08253_),
    .Q(\mem.mem[10][0] ));
 sg13g2_dfrbp_1 _19338_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net347),
    .D(_00974_),
    .Q_N(_08252_),
    .Q(\mem.mem[10][1] ));
 sg13g2_dfrbp_1 _19339_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net346),
    .D(_00975_),
    .Q_N(_08251_),
    .Q(\mem.mem[10][2] ));
 sg13g2_dfrbp_1 _19340_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net345),
    .D(_00976_),
    .Q_N(_08250_),
    .Q(\mem.mem[10][3] ));
 sg13g2_dfrbp_1 _19341_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net344),
    .D(_00977_),
    .Q_N(_08249_),
    .Q(\mem.mem[10][4] ));
 sg13g2_dfrbp_1 _19342_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net343),
    .D(_00978_),
    .Q_N(_08248_),
    .Q(\mem.mem[10][5] ));
 sg13g2_dfrbp_1 _19343_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net342),
    .D(_00979_),
    .Q_N(_08247_),
    .Q(\mem.mem[10][6] ));
 sg13g2_dfrbp_1 _19344_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net341),
    .D(_00980_),
    .Q_N(_08246_),
    .Q(\mem.mem[10][7] ));
 sg13g2_dfrbp_1 _19345_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net340),
    .D(_00981_),
    .Q_N(_08245_),
    .Q(\mem.mem[110][0] ));
 sg13g2_dfrbp_1 _19346_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net339),
    .D(_00982_),
    .Q_N(_08244_),
    .Q(\mem.mem[110][1] ));
 sg13g2_dfrbp_1 _19347_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net338),
    .D(_00983_),
    .Q_N(_08243_),
    .Q(\mem.mem[110][2] ));
 sg13g2_dfrbp_1 _19348_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net337),
    .D(_00984_),
    .Q_N(_08242_),
    .Q(\mem.mem[110][3] ));
 sg13g2_dfrbp_1 _19349_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net336),
    .D(_00985_),
    .Q_N(_08241_),
    .Q(\mem.mem[110][4] ));
 sg13g2_dfrbp_1 _19350_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net335),
    .D(_00986_),
    .Q_N(_08240_),
    .Q(\mem.mem[110][5] ));
 sg13g2_dfrbp_1 _19351_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net334),
    .D(_00987_),
    .Q_N(_08239_),
    .Q(\mem.mem[110][6] ));
 sg13g2_dfrbp_1 _19352_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net333),
    .D(_00988_),
    .Q_N(_08238_),
    .Q(\mem.mem[110][7] ));
 sg13g2_dfrbp_1 _19353_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net332),
    .D(_00989_),
    .Q_N(_08237_),
    .Q(\mem.mem[111][0] ));
 sg13g2_dfrbp_1 _19354_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net331),
    .D(_00990_),
    .Q_N(_08236_),
    .Q(\mem.mem[111][1] ));
 sg13g2_dfrbp_1 _19355_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net330),
    .D(_00991_),
    .Q_N(_08235_),
    .Q(\mem.mem[111][2] ));
 sg13g2_dfrbp_1 _19356_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net329),
    .D(_00992_),
    .Q_N(_08234_),
    .Q(\mem.mem[111][3] ));
 sg13g2_dfrbp_1 _19357_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net328),
    .D(_00993_),
    .Q_N(_08233_),
    .Q(\mem.mem[111][4] ));
 sg13g2_dfrbp_1 _19358_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net327),
    .D(_00994_),
    .Q_N(_08232_),
    .Q(\mem.mem[111][5] ));
 sg13g2_dfrbp_1 _19359_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net326),
    .D(_00995_),
    .Q_N(_08231_),
    .Q(\mem.mem[111][6] ));
 sg13g2_dfrbp_1 _19360_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net325),
    .D(_00996_),
    .Q_N(_08230_),
    .Q(\mem.mem[111][7] ));
 sg13g2_dfrbp_1 _19361_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net324),
    .D(_00997_),
    .Q_N(_08229_),
    .Q(\mem.mem[112][0] ));
 sg13g2_dfrbp_1 _19362_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net323),
    .D(_00998_),
    .Q_N(_08228_),
    .Q(\mem.mem[112][1] ));
 sg13g2_dfrbp_1 _19363_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net322),
    .D(_00999_),
    .Q_N(_08227_),
    .Q(\mem.mem[112][2] ));
 sg13g2_dfrbp_1 _19364_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net321),
    .D(_01000_),
    .Q_N(_08226_),
    .Q(\mem.mem[112][3] ));
 sg13g2_dfrbp_1 _19365_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net320),
    .D(_01001_),
    .Q_N(_08225_),
    .Q(\mem.mem[112][4] ));
 sg13g2_dfrbp_1 _19366_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net319),
    .D(_01002_),
    .Q_N(_08224_),
    .Q(\mem.mem[112][5] ));
 sg13g2_dfrbp_1 _19367_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net318),
    .D(_01003_),
    .Q_N(_08223_),
    .Q(\mem.mem[112][6] ));
 sg13g2_dfrbp_1 _19368_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net317),
    .D(_01004_),
    .Q_N(_08222_),
    .Q(\mem.mem[112][7] ));
 sg13g2_dfrbp_1 _19369_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net316),
    .D(_01005_),
    .Q_N(_08221_),
    .Q(\mem.mem[113][0] ));
 sg13g2_dfrbp_1 _19370_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net315),
    .D(_01006_),
    .Q_N(_08220_),
    .Q(\mem.mem[113][1] ));
 sg13g2_dfrbp_1 _19371_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net314),
    .D(_01007_),
    .Q_N(_08219_),
    .Q(\mem.mem[113][2] ));
 sg13g2_dfrbp_1 _19372_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net313),
    .D(_01008_),
    .Q_N(_08218_),
    .Q(\mem.mem[113][3] ));
 sg13g2_dfrbp_1 _19373_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net312),
    .D(_01009_),
    .Q_N(_08217_),
    .Q(\mem.mem[113][4] ));
 sg13g2_dfrbp_1 _19374_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net311),
    .D(_01010_),
    .Q_N(_08216_),
    .Q(\mem.mem[113][5] ));
 sg13g2_dfrbp_1 _19375_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net310),
    .D(_01011_),
    .Q_N(_08215_),
    .Q(\mem.mem[113][6] ));
 sg13g2_dfrbp_1 _19376_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net309),
    .D(_01012_),
    .Q_N(_08214_),
    .Q(\mem.mem[113][7] ));
 sg13g2_dfrbp_1 _19377_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net308),
    .D(_01013_),
    .Q_N(_08213_),
    .Q(\mem.mem[114][0] ));
 sg13g2_dfrbp_1 _19378_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net307),
    .D(_01014_),
    .Q_N(_08212_),
    .Q(\mem.mem[114][1] ));
 sg13g2_dfrbp_1 _19379_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net306),
    .D(_01015_),
    .Q_N(_08211_),
    .Q(\mem.mem[114][2] ));
 sg13g2_dfrbp_1 _19380_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net305),
    .D(_01016_),
    .Q_N(_08210_),
    .Q(\mem.mem[114][3] ));
 sg13g2_dfrbp_1 _19381_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net304),
    .D(_01017_),
    .Q_N(_08209_),
    .Q(\mem.mem[114][4] ));
 sg13g2_dfrbp_1 _19382_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net303),
    .D(_01018_),
    .Q_N(_08208_),
    .Q(\mem.mem[114][5] ));
 sg13g2_dfrbp_1 _19383_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net302),
    .D(_01019_),
    .Q_N(_08207_),
    .Q(\mem.mem[114][6] ));
 sg13g2_dfrbp_1 _19384_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net301),
    .D(_01020_),
    .Q_N(_08206_),
    .Q(\mem.mem[114][7] ));
 sg13g2_dfrbp_1 _19385_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net300),
    .D(_01021_),
    .Q_N(_08205_),
    .Q(\mem.mem[115][0] ));
 sg13g2_dfrbp_1 _19386_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net299),
    .D(_01022_),
    .Q_N(_08204_),
    .Q(\mem.mem[115][1] ));
 sg13g2_dfrbp_1 _19387_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net298),
    .D(_01023_),
    .Q_N(_08203_),
    .Q(\mem.mem[115][2] ));
 sg13g2_dfrbp_1 _19388_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net297),
    .D(_01024_),
    .Q_N(_08202_),
    .Q(\mem.mem[115][3] ));
 sg13g2_dfrbp_1 _19389_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net296),
    .D(_01025_),
    .Q_N(_08201_),
    .Q(\mem.mem[115][4] ));
 sg13g2_dfrbp_1 _19390_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net295),
    .D(_01026_),
    .Q_N(_08200_),
    .Q(\mem.mem[115][5] ));
 sg13g2_dfrbp_1 _19391_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net294),
    .D(_01027_),
    .Q_N(_08199_),
    .Q(\mem.mem[115][6] ));
 sg13g2_dfrbp_1 _19392_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net293),
    .D(_01028_),
    .Q_N(_08198_),
    .Q(\mem.mem[115][7] ));
 sg13g2_dfrbp_1 _19393_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net292),
    .D(_01029_),
    .Q_N(_08197_),
    .Q(\mem.mem[116][0] ));
 sg13g2_dfrbp_1 _19394_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net291),
    .D(_01030_),
    .Q_N(_08196_),
    .Q(\mem.mem[116][1] ));
 sg13g2_dfrbp_1 _19395_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net290),
    .D(_01031_),
    .Q_N(_08195_),
    .Q(\mem.mem[116][2] ));
 sg13g2_dfrbp_1 _19396_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net289),
    .D(_01032_),
    .Q_N(_08194_),
    .Q(\mem.mem[116][3] ));
 sg13g2_dfrbp_1 _19397_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net288),
    .D(_01033_),
    .Q_N(_08193_),
    .Q(\mem.mem[116][4] ));
 sg13g2_dfrbp_1 _19398_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net287),
    .D(_01034_),
    .Q_N(_08192_),
    .Q(\mem.mem[116][5] ));
 sg13g2_dfrbp_1 _19399_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net286),
    .D(_01035_),
    .Q_N(_08191_),
    .Q(\mem.mem[116][6] ));
 sg13g2_dfrbp_1 _19400_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net285),
    .D(_01036_),
    .Q_N(_08190_),
    .Q(\mem.mem[116][7] ));
 sg13g2_dfrbp_1 _19401_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net284),
    .D(_01037_),
    .Q_N(_08189_),
    .Q(\mem.mem[117][0] ));
 sg13g2_dfrbp_1 _19402_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net283),
    .D(_01038_),
    .Q_N(_08188_),
    .Q(\mem.mem[117][1] ));
 sg13g2_dfrbp_1 _19403_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net282),
    .D(_01039_),
    .Q_N(_08187_),
    .Q(\mem.mem[117][2] ));
 sg13g2_dfrbp_1 _19404_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net281),
    .D(_01040_),
    .Q_N(_08186_),
    .Q(\mem.mem[117][3] ));
 sg13g2_dfrbp_1 _19405_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net280),
    .D(_01041_),
    .Q_N(_08185_),
    .Q(\mem.mem[117][4] ));
 sg13g2_dfrbp_1 _19406_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net279),
    .D(_01042_),
    .Q_N(_08184_),
    .Q(\mem.mem[117][5] ));
 sg13g2_dfrbp_1 _19407_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net278),
    .D(_01043_),
    .Q_N(_08183_),
    .Q(\mem.mem[117][6] ));
 sg13g2_dfrbp_1 _19408_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net277),
    .D(_01044_),
    .Q_N(_08182_),
    .Q(\mem.mem[117][7] ));
 sg13g2_dfrbp_1 _19409_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net276),
    .D(net3092),
    .Q_N(_08181_),
    .Q(\mem.mem[118][0] ));
 sg13g2_dfrbp_1 _19410_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net275),
    .D(_01046_),
    .Q_N(_08180_),
    .Q(\mem.mem[118][1] ));
 sg13g2_dfrbp_1 _19411_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net274),
    .D(_01047_),
    .Q_N(_08179_),
    .Q(\mem.mem[118][2] ));
 sg13g2_dfrbp_1 _19412_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net273),
    .D(_01048_),
    .Q_N(_08178_),
    .Q(\mem.mem[118][3] ));
 sg13g2_dfrbp_1 _19413_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net272),
    .D(_01049_),
    .Q_N(_08177_),
    .Q(\mem.mem[118][4] ));
 sg13g2_dfrbp_1 _19414_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net271),
    .D(_01050_),
    .Q_N(_08176_),
    .Q(\mem.mem[118][5] ));
 sg13g2_dfrbp_1 _19415_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net270),
    .D(_01051_),
    .Q_N(_08175_),
    .Q(\mem.mem[118][6] ));
 sg13g2_dfrbp_1 _19416_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net269),
    .D(_01052_),
    .Q_N(_08174_),
    .Q(\mem.mem[118][7] ));
 sg13g2_dfrbp_1 _19417_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net268),
    .D(_01053_),
    .Q_N(_08173_),
    .Q(\mem.mem[11][0] ));
 sg13g2_dfrbp_1 _19418_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net267),
    .D(_01054_),
    .Q_N(_08172_),
    .Q(\mem.mem[11][1] ));
 sg13g2_dfrbp_1 _19419_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net266),
    .D(_01055_),
    .Q_N(_08171_),
    .Q(\mem.mem[11][2] ));
 sg13g2_dfrbp_1 _19420_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net265),
    .D(_01056_),
    .Q_N(_08170_),
    .Q(\mem.mem[11][3] ));
 sg13g2_dfrbp_1 _19421_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net264),
    .D(_01057_),
    .Q_N(_08169_),
    .Q(\mem.mem[11][4] ));
 sg13g2_dfrbp_1 _19422_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net263),
    .D(_01058_),
    .Q_N(_08168_),
    .Q(\mem.mem[11][5] ));
 sg13g2_dfrbp_1 _19423_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net262),
    .D(_01059_),
    .Q_N(_08167_),
    .Q(\mem.mem[11][6] ));
 sg13g2_dfrbp_1 _19424_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net261),
    .D(_01060_),
    .Q_N(_08166_),
    .Q(\mem.mem[11][7] ));
 sg13g2_dfrbp_1 _19425_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net260),
    .D(_01061_),
    .Q_N(_08165_),
    .Q(\mem.mem[120][0] ));
 sg13g2_dfrbp_1 _19426_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net259),
    .D(_01062_),
    .Q_N(_08164_),
    .Q(\mem.mem[120][1] ));
 sg13g2_dfrbp_1 _19427_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net258),
    .D(_01063_),
    .Q_N(_08163_),
    .Q(\mem.mem[120][2] ));
 sg13g2_dfrbp_1 _19428_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net257),
    .D(_01064_),
    .Q_N(_08162_),
    .Q(\mem.mem[120][3] ));
 sg13g2_dfrbp_1 _19429_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net256),
    .D(_01065_),
    .Q_N(_08161_),
    .Q(\mem.mem[120][4] ));
 sg13g2_dfrbp_1 _19430_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net255),
    .D(_01066_),
    .Q_N(_08160_),
    .Q(\mem.mem[120][5] ));
 sg13g2_dfrbp_1 _19431_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net254),
    .D(_01067_),
    .Q_N(_08159_),
    .Q(\mem.mem[120][6] ));
 sg13g2_dfrbp_1 _19432_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net253),
    .D(_01068_),
    .Q_N(_08158_),
    .Q(\mem.mem[120][7] ));
 sg13g2_dfrbp_1 _19433_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net252),
    .D(_01069_),
    .Q_N(_08157_),
    .Q(\mem.mem[121][0] ));
 sg13g2_dfrbp_1 _19434_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net251),
    .D(_01070_),
    .Q_N(_08156_),
    .Q(\mem.mem[121][1] ));
 sg13g2_dfrbp_1 _19435_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net250),
    .D(_01071_),
    .Q_N(_08155_),
    .Q(\mem.mem[121][2] ));
 sg13g2_dfrbp_1 _19436_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net249),
    .D(_01072_),
    .Q_N(_08154_),
    .Q(\mem.mem[121][3] ));
 sg13g2_dfrbp_1 _19437_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net248),
    .D(_01073_),
    .Q_N(_08153_),
    .Q(\mem.mem[121][4] ));
 sg13g2_dfrbp_1 _19438_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net247),
    .D(_01074_),
    .Q_N(_08152_),
    .Q(\mem.mem[121][5] ));
 sg13g2_dfrbp_1 _19439_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net246),
    .D(_01075_),
    .Q_N(_08151_),
    .Q(\mem.mem[121][6] ));
 sg13g2_dfrbp_1 _19440_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net245),
    .D(_01076_),
    .Q_N(_08150_),
    .Q(\mem.mem[121][7] ));
 sg13g2_dfrbp_1 _19441_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net244),
    .D(_01077_),
    .Q_N(_08149_),
    .Q(\mem.mem[122][0] ));
 sg13g2_dfrbp_1 _19442_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net243),
    .D(_01078_),
    .Q_N(_08148_),
    .Q(\mem.mem[122][1] ));
 sg13g2_dfrbp_1 _19443_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net242),
    .D(_01079_),
    .Q_N(_08147_),
    .Q(\mem.mem[122][2] ));
 sg13g2_dfrbp_1 _19444_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net241),
    .D(_01080_),
    .Q_N(_08146_),
    .Q(\mem.mem[122][3] ));
 sg13g2_dfrbp_1 _19445_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net240),
    .D(_01081_),
    .Q_N(_08145_),
    .Q(\mem.mem[122][4] ));
 sg13g2_dfrbp_1 _19446_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net239),
    .D(_01082_),
    .Q_N(_08144_),
    .Q(\mem.mem[122][5] ));
 sg13g2_dfrbp_1 _19447_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net238),
    .D(_01083_),
    .Q_N(_08143_),
    .Q(\mem.mem[122][6] ));
 sg13g2_dfrbp_1 _19448_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net237),
    .D(_01084_),
    .Q_N(_08142_),
    .Q(\mem.mem[122][7] ));
 sg13g2_dfrbp_1 _19449_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net236),
    .D(_01085_),
    .Q_N(_08141_),
    .Q(\mem.mem[123][0] ));
 sg13g2_dfrbp_1 _19450_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net235),
    .D(_01086_),
    .Q_N(_08140_),
    .Q(\mem.mem[123][1] ));
 sg13g2_dfrbp_1 _19451_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net234),
    .D(_01087_),
    .Q_N(_08139_),
    .Q(\mem.mem[123][2] ));
 sg13g2_dfrbp_1 _19452_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net233),
    .D(_01088_),
    .Q_N(_08138_),
    .Q(\mem.mem[123][3] ));
 sg13g2_dfrbp_1 _19453_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net232),
    .D(_01089_),
    .Q_N(_08137_),
    .Q(\mem.mem[123][4] ));
 sg13g2_dfrbp_1 _19454_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net231),
    .D(_01090_),
    .Q_N(_08136_),
    .Q(\mem.mem[123][5] ));
 sg13g2_dfrbp_1 _19455_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net230),
    .D(_01091_),
    .Q_N(_08135_),
    .Q(\mem.mem[123][6] ));
 sg13g2_dfrbp_1 _19456_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net229),
    .D(_01092_),
    .Q_N(_08134_),
    .Q(\mem.mem[123][7] ));
 sg13g2_dfrbp_1 _19457_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net228),
    .D(_01093_),
    .Q_N(_08133_),
    .Q(\mem.mem[124][0] ));
 sg13g2_dfrbp_1 _19458_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net227),
    .D(_01094_),
    .Q_N(_08132_),
    .Q(\mem.mem[124][1] ));
 sg13g2_dfrbp_1 _19459_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net226),
    .D(_01095_),
    .Q_N(_08131_),
    .Q(\mem.mem[124][2] ));
 sg13g2_dfrbp_1 _19460_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net225),
    .D(_01096_),
    .Q_N(_08130_),
    .Q(\mem.mem[124][3] ));
 sg13g2_dfrbp_1 _19461_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net224),
    .D(_01097_),
    .Q_N(_08129_),
    .Q(\mem.mem[124][4] ));
 sg13g2_dfrbp_1 _19462_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net223),
    .D(_01098_),
    .Q_N(_08128_),
    .Q(\mem.mem[124][5] ));
 sg13g2_dfrbp_1 _19463_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net222),
    .D(_01099_),
    .Q_N(_08127_),
    .Q(\mem.mem[124][6] ));
 sg13g2_dfrbp_1 _19464_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net221),
    .D(_01100_),
    .Q_N(_08126_),
    .Q(\mem.mem[124][7] ));
 sg13g2_dfrbp_1 _19465_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net220),
    .D(_01101_),
    .Q_N(_08125_),
    .Q(\mem.mem[125][0] ));
 sg13g2_dfrbp_1 _19466_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net219),
    .D(_01102_),
    .Q_N(_08124_),
    .Q(\mem.mem[125][1] ));
 sg13g2_dfrbp_1 _19467_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net218),
    .D(_01103_),
    .Q_N(_08123_),
    .Q(\mem.mem[125][2] ));
 sg13g2_dfrbp_1 _19468_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net217),
    .D(_01104_),
    .Q_N(_08122_),
    .Q(\mem.mem[125][3] ));
 sg13g2_dfrbp_1 _19469_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net216),
    .D(_01105_),
    .Q_N(_08121_),
    .Q(\mem.mem[125][4] ));
 sg13g2_dfrbp_1 _19470_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net215),
    .D(_01106_),
    .Q_N(_08120_),
    .Q(\mem.mem[125][5] ));
 sg13g2_dfrbp_1 _19471_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net214),
    .D(_01107_),
    .Q_N(_08119_),
    .Q(\mem.mem[125][6] ));
 sg13g2_dfrbp_1 _19472_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net213),
    .D(_01108_),
    .Q_N(_08118_),
    .Q(\mem.mem[125][7] ));
 sg13g2_dfrbp_1 _19473_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net212),
    .D(_01109_),
    .Q_N(_08117_),
    .Q(\mem.mem[126][0] ));
 sg13g2_dfrbp_1 _19474_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net211),
    .D(_01110_),
    .Q_N(_08116_),
    .Q(\mem.mem[126][1] ));
 sg13g2_dfrbp_1 _19475_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net210),
    .D(_01111_),
    .Q_N(_08115_),
    .Q(\mem.mem[126][2] ));
 sg13g2_dfrbp_1 _19476_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net209),
    .D(_01112_),
    .Q_N(_08114_),
    .Q(\mem.mem[126][3] ));
 sg13g2_dfrbp_1 _19477_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net208),
    .D(_01113_),
    .Q_N(_08113_),
    .Q(\mem.mem[126][4] ));
 sg13g2_dfrbp_1 _19478_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net207),
    .D(_01114_),
    .Q_N(_08112_),
    .Q(\mem.mem[126][5] ));
 sg13g2_dfrbp_1 _19479_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net206),
    .D(_01115_),
    .Q_N(_08111_),
    .Q(\mem.mem[126][6] ));
 sg13g2_dfrbp_1 _19480_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net205),
    .D(_01116_),
    .Q_N(_08110_),
    .Q(\mem.mem[126][7] ));
 sg13g2_dfrbp_1 _19481_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net204),
    .D(_01117_),
    .Q_N(_08109_),
    .Q(\mem.mem[127][0] ));
 sg13g2_dfrbp_1 _19482_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net203),
    .D(_01118_),
    .Q_N(_08108_),
    .Q(\mem.mem[127][1] ));
 sg13g2_dfrbp_1 _19483_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net202),
    .D(_01119_),
    .Q_N(_08107_),
    .Q(\mem.mem[127][2] ));
 sg13g2_dfrbp_1 _19484_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net201),
    .D(_01120_),
    .Q_N(_08106_),
    .Q(\mem.mem[127][3] ));
 sg13g2_dfrbp_1 _19485_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net200),
    .D(_01121_),
    .Q_N(_08105_),
    .Q(\mem.mem[127][4] ));
 sg13g2_dfrbp_1 _19486_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net199),
    .D(_01122_),
    .Q_N(_08104_),
    .Q(\mem.mem[127][5] ));
 sg13g2_dfrbp_1 _19487_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net198),
    .D(_01123_),
    .Q_N(_08103_),
    .Q(\mem.mem[127][6] ));
 sg13g2_dfrbp_1 _19488_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net197),
    .D(_01124_),
    .Q_N(_08102_),
    .Q(\mem.mem[127][7] ));
 sg13g2_dfrbp_1 _19489_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net196),
    .D(_01125_),
    .Q_N(_08101_),
    .Q(\mem.mem[128][0] ));
 sg13g2_dfrbp_1 _19490_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net195),
    .D(_01126_),
    .Q_N(_08100_),
    .Q(\mem.mem[128][1] ));
 sg13g2_dfrbp_1 _19491_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net194),
    .D(_01127_),
    .Q_N(_08099_),
    .Q(\mem.mem[128][2] ));
 sg13g2_dfrbp_1 _19492_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net193),
    .D(_01128_),
    .Q_N(_08098_),
    .Q(\mem.mem[128][3] ));
 sg13g2_dfrbp_1 _19493_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net192),
    .D(_01129_),
    .Q_N(_08097_),
    .Q(\mem.mem[128][4] ));
 sg13g2_dfrbp_1 _19494_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net191),
    .D(_01130_),
    .Q_N(_08096_),
    .Q(\mem.mem[128][5] ));
 sg13g2_dfrbp_1 _19495_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net190),
    .D(_01131_),
    .Q_N(_08095_),
    .Q(\mem.mem[128][6] ));
 sg13g2_dfrbp_1 _19496_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net189),
    .D(_01132_),
    .Q_N(_08094_),
    .Q(\mem.mem[128][7] ));
 sg13g2_dfrbp_1 _19497_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net188),
    .D(_01133_),
    .Q_N(_08093_),
    .Q(\mem.mem[12][0] ));
 sg13g2_dfrbp_1 _19498_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net187),
    .D(_01134_),
    .Q_N(_08092_),
    .Q(\mem.mem[12][1] ));
 sg13g2_dfrbp_1 _19499_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net186),
    .D(_01135_),
    .Q_N(_08091_),
    .Q(\mem.mem[12][2] ));
 sg13g2_dfrbp_1 _19500_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net185),
    .D(_01136_),
    .Q_N(_08090_),
    .Q(\mem.mem[12][3] ));
 sg13g2_dfrbp_1 _19501_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net184),
    .D(_01137_),
    .Q_N(_08089_),
    .Q(\mem.mem[12][4] ));
 sg13g2_dfrbp_1 _19502_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net183),
    .D(_01138_),
    .Q_N(_08088_),
    .Q(\mem.mem[12][5] ));
 sg13g2_dfrbp_1 _19503_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net182),
    .D(_01139_),
    .Q_N(_08087_),
    .Q(\mem.mem[12][6] ));
 sg13g2_dfrbp_1 _19504_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net181),
    .D(_01140_),
    .Q_N(_08086_),
    .Q(\mem.mem[12][7] ));
 sg13g2_dfrbp_1 _19505_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net180),
    .D(_01141_),
    .Q_N(_08085_),
    .Q(\mem.mem[130][0] ));
 sg13g2_dfrbp_1 _19506_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net179),
    .D(_01142_),
    .Q_N(_08084_),
    .Q(\mem.mem[130][1] ));
 sg13g2_dfrbp_1 _19507_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net178),
    .D(_01143_),
    .Q_N(_08083_),
    .Q(\mem.mem[130][2] ));
 sg13g2_dfrbp_1 _19508_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net177),
    .D(_01144_),
    .Q_N(_08082_),
    .Q(\mem.mem[130][3] ));
 sg13g2_dfrbp_1 _19509_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net176),
    .D(_01145_),
    .Q_N(_08081_),
    .Q(\mem.mem[130][4] ));
 sg13g2_dfrbp_1 _19510_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net175),
    .D(_01146_),
    .Q_N(_08080_),
    .Q(\mem.mem[130][5] ));
 sg13g2_dfrbp_1 _19511_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net174),
    .D(_01147_),
    .Q_N(_08079_),
    .Q(\mem.mem[130][6] ));
 sg13g2_dfrbp_1 _19512_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net173),
    .D(_01148_),
    .Q_N(_08078_),
    .Q(\mem.mem[130][7] ));
 sg13g2_dfrbp_1 _19513_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net172),
    .D(_01149_),
    .Q_N(_08077_),
    .Q(\mem.mem[131][0] ));
 sg13g2_dfrbp_1 _19514_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net171),
    .D(_01150_),
    .Q_N(_08076_),
    .Q(\mem.mem[131][1] ));
 sg13g2_dfrbp_1 _19515_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net170),
    .D(_01151_),
    .Q_N(_08075_),
    .Q(\mem.mem[131][2] ));
 sg13g2_dfrbp_1 _19516_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net169),
    .D(_01152_),
    .Q_N(_08074_),
    .Q(\mem.mem[131][3] ));
 sg13g2_dfrbp_1 _19517_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net168),
    .D(_01153_),
    .Q_N(_08073_),
    .Q(\mem.mem[131][4] ));
 sg13g2_dfrbp_1 _19518_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net167),
    .D(_01154_),
    .Q_N(_08072_),
    .Q(\mem.mem[131][5] ));
 sg13g2_dfrbp_1 _19519_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net166),
    .D(_01155_),
    .Q_N(_08071_),
    .Q(\mem.mem[131][6] ));
 sg13g2_dfrbp_1 _19520_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net165),
    .D(_01156_),
    .Q_N(_08070_),
    .Q(\mem.mem[131][7] ));
 sg13g2_dfrbp_1 _19521_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net164),
    .D(_01157_),
    .Q_N(_08069_),
    .Q(\mem.mem[132][0] ));
 sg13g2_dfrbp_1 _19522_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net163),
    .D(_01158_),
    .Q_N(_08068_),
    .Q(\mem.mem[132][1] ));
 sg13g2_dfrbp_1 _19523_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net162),
    .D(_01159_),
    .Q_N(_08067_),
    .Q(\mem.mem[132][2] ));
 sg13g2_dfrbp_1 _19524_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net161),
    .D(_01160_),
    .Q_N(_08066_),
    .Q(\mem.mem[132][3] ));
 sg13g2_dfrbp_1 _19525_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net160),
    .D(_01161_),
    .Q_N(_08065_),
    .Q(\mem.mem[132][4] ));
 sg13g2_dfrbp_1 _19526_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net159),
    .D(_01162_),
    .Q_N(_08064_),
    .Q(\mem.mem[132][5] ));
 sg13g2_dfrbp_1 _19527_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net158),
    .D(_01163_),
    .Q_N(_08063_),
    .Q(\mem.mem[132][6] ));
 sg13g2_dfrbp_1 _19528_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net157),
    .D(_01164_),
    .Q_N(_08062_),
    .Q(\mem.mem[132][7] ));
 sg13g2_dfrbp_1 _19529_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net156),
    .D(_01165_),
    .Q_N(_08061_),
    .Q(\mem.mem[133][0] ));
 sg13g2_dfrbp_1 _19530_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net155),
    .D(_01166_),
    .Q_N(_08060_),
    .Q(\mem.mem[133][1] ));
 sg13g2_dfrbp_1 _19531_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net154),
    .D(_01167_),
    .Q_N(_08059_),
    .Q(\mem.mem[133][2] ));
 sg13g2_dfrbp_1 _19532_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net153),
    .D(_01168_),
    .Q_N(_08058_),
    .Q(\mem.mem[133][3] ));
 sg13g2_dfrbp_1 _19533_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net152),
    .D(_01169_),
    .Q_N(_08057_),
    .Q(\mem.mem[133][4] ));
 sg13g2_dfrbp_1 _19534_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net151),
    .D(_01170_),
    .Q_N(_08056_),
    .Q(\mem.mem[133][5] ));
 sg13g2_dfrbp_1 _19535_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net150),
    .D(_01171_),
    .Q_N(_08055_),
    .Q(\mem.mem[133][6] ));
 sg13g2_dfrbp_1 _19536_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net149),
    .D(_01172_),
    .Q_N(_08054_),
    .Q(\mem.mem[133][7] ));
 sg13g2_dfrbp_1 _19537_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net148),
    .D(_01173_),
    .Q_N(_08053_),
    .Q(\mem.mem[134][0] ));
 sg13g2_dfrbp_1 _19538_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net147),
    .D(_01174_),
    .Q_N(_08052_),
    .Q(\mem.mem[134][1] ));
 sg13g2_dfrbp_1 _19539_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net146),
    .D(_01175_),
    .Q_N(_08051_),
    .Q(\mem.mem[134][2] ));
 sg13g2_dfrbp_1 _19540_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net145),
    .D(_01176_),
    .Q_N(_08050_),
    .Q(\mem.mem[134][3] ));
 sg13g2_dfrbp_1 _19541_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net144),
    .D(_01177_),
    .Q_N(_08049_),
    .Q(\mem.mem[134][4] ));
 sg13g2_dfrbp_1 _19542_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net143),
    .D(_01178_),
    .Q_N(_08048_),
    .Q(\mem.mem[134][5] ));
 sg13g2_dfrbp_1 _19543_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net142),
    .D(_01179_),
    .Q_N(_08047_),
    .Q(\mem.mem[134][6] ));
 sg13g2_dfrbp_1 _19544_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net141),
    .D(_01180_),
    .Q_N(_08046_),
    .Q(\mem.mem[134][7] ));
 sg13g2_dfrbp_1 _19545_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net140),
    .D(_01181_),
    .Q_N(_08045_),
    .Q(\mem.mem[135][0] ));
 sg13g2_dfrbp_1 _19546_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net139),
    .D(_01182_),
    .Q_N(_08044_),
    .Q(\mem.mem[135][1] ));
 sg13g2_dfrbp_1 _19547_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net138),
    .D(_01183_),
    .Q_N(_08043_),
    .Q(\mem.mem[135][2] ));
 sg13g2_dfrbp_1 _19548_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net137),
    .D(_01184_),
    .Q_N(_08042_),
    .Q(\mem.mem[135][3] ));
 sg13g2_dfrbp_1 _19549_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net136),
    .D(_01185_),
    .Q_N(_08041_),
    .Q(\mem.mem[135][4] ));
 sg13g2_dfrbp_1 _19550_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net135),
    .D(_01186_),
    .Q_N(_08040_),
    .Q(\mem.mem[135][5] ));
 sg13g2_dfrbp_1 _19551_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net134),
    .D(_01187_),
    .Q_N(_08039_),
    .Q(\mem.mem[135][6] ));
 sg13g2_dfrbp_1 _19552_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net133),
    .D(_01188_),
    .Q_N(_08038_),
    .Q(\mem.mem[135][7] ));
 sg13g2_dfrbp_1 _19553_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net132),
    .D(_01189_),
    .Q_N(_08037_),
    .Q(\mem.mem[136][0] ));
 sg13g2_dfrbp_1 _19554_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net131),
    .D(_01190_),
    .Q_N(_08036_),
    .Q(\mem.mem[136][1] ));
 sg13g2_dfrbp_1 _19555_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net130),
    .D(_01191_),
    .Q_N(_08035_),
    .Q(\mem.mem[136][2] ));
 sg13g2_dfrbp_1 _19556_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net129),
    .D(_01192_),
    .Q_N(_08034_),
    .Q(\mem.mem[136][3] ));
 sg13g2_dfrbp_1 _19557_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net128),
    .D(_01193_),
    .Q_N(_08033_),
    .Q(\mem.mem[136][4] ));
 sg13g2_dfrbp_1 _19558_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net127),
    .D(_01194_),
    .Q_N(_08032_),
    .Q(\mem.mem[136][5] ));
 sg13g2_dfrbp_1 _19559_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net126),
    .D(_01195_),
    .Q_N(_08031_),
    .Q(\mem.mem[136][6] ));
 sg13g2_dfrbp_1 _19560_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net125),
    .D(_01196_),
    .Q_N(_08030_),
    .Q(\mem.mem[136][7] ));
 sg13g2_dfrbp_1 _19561_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net124),
    .D(_01197_),
    .Q_N(_08029_),
    .Q(\mem.mem[137][0] ));
 sg13g2_dfrbp_1 _19562_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net123),
    .D(_01198_),
    .Q_N(_08028_),
    .Q(\mem.mem[137][1] ));
 sg13g2_dfrbp_1 _19563_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net122),
    .D(_01199_),
    .Q_N(_08027_),
    .Q(\mem.mem[137][2] ));
 sg13g2_dfrbp_1 _19564_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net121),
    .D(_01200_),
    .Q_N(_08026_),
    .Q(\mem.mem[137][3] ));
 sg13g2_dfrbp_1 _19565_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net120),
    .D(_01201_),
    .Q_N(_08025_),
    .Q(\mem.mem[137][4] ));
 sg13g2_dfrbp_1 _19566_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net119),
    .D(_01202_),
    .Q_N(_08024_),
    .Q(\mem.mem[137][5] ));
 sg13g2_dfrbp_1 _19567_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net118),
    .D(_01203_),
    .Q_N(_08023_),
    .Q(\mem.mem[137][6] ));
 sg13g2_dfrbp_1 _19568_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net117),
    .D(_01204_),
    .Q_N(_08022_),
    .Q(\mem.mem[137][7] ));
 sg13g2_dfrbp_1 _19569_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net116),
    .D(_01205_),
    .Q_N(_08021_),
    .Q(\mem.mem[138][0] ));
 sg13g2_dfrbp_1 _19570_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net115),
    .D(_01206_),
    .Q_N(_08020_),
    .Q(\mem.mem[138][1] ));
 sg13g2_dfrbp_1 _19571_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net114),
    .D(_01207_),
    .Q_N(_08019_),
    .Q(\mem.mem[138][2] ));
 sg13g2_dfrbp_1 _19572_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net113),
    .D(_01208_),
    .Q_N(_08018_),
    .Q(\mem.mem[138][3] ));
 sg13g2_dfrbp_1 _19573_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net112),
    .D(_01209_),
    .Q_N(_08017_),
    .Q(\mem.mem[138][4] ));
 sg13g2_dfrbp_1 _19574_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net111),
    .D(_01210_),
    .Q_N(_08016_),
    .Q(\mem.mem[138][5] ));
 sg13g2_dfrbp_1 _19575_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net110),
    .D(_01211_),
    .Q_N(_08015_),
    .Q(\mem.mem[138][6] ));
 sg13g2_dfrbp_1 _19576_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net109),
    .D(_01212_),
    .Q_N(_08014_),
    .Q(\mem.mem[138][7] ));
 sg13g2_dfrbp_1 _19577_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net108),
    .D(_01213_),
    .Q_N(_08013_),
    .Q(\mem.mem[13][0] ));
 sg13g2_dfrbp_1 _19578_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net107),
    .D(_01214_),
    .Q_N(_08012_),
    .Q(\mem.mem[13][1] ));
 sg13g2_dfrbp_1 _19579_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net106),
    .D(_01215_),
    .Q_N(_08011_),
    .Q(\mem.mem[13][2] ));
 sg13g2_dfrbp_1 _19580_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net105),
    .D(_01216_),
    .Q_N(_08010_),
    .Q(\mem.mem[13][3] ));
 sg13g2_dfrbp_1 _19581_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net104),
    .D(_01217_),
    .Q_N(_08009_),
    .Q(\mem.mem[13][4] ));
 sg13g2_dfrbp_1 _19582_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net103),
    .D(_01218_),
    .Q_N(_08008_),
    .Q(\mem.mem[13][5] ));
 sg13g2_dfrbp_1 _19583_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net102),
    .D(_01219_),
    .Q_N(_08007_),
    .Q(\mem.mem[13][6] ));
 sg13g2_dfrbp_1 _19584_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net101),
    .D(_01220_),
    .Q_N(_08006_),
    .Q(\mem.mem[13][7] ));
 sg13g2_dfrbp_1 _19585_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net100),
    .D(_01221_),
    .Q_N(_08005_),
    .Q(\mem.mem[140][0] ));
 sg13g2_dfrbp_1 _19586_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net99),
    .D(_01222_),
    .Q_N(_08004_),
    .Q(\mem.mem[140][1] ));
 sg13g2_dfrbp_1 _19587_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net98),
    .D(_01223_),
    .Q_N(_08003_),
    .Q(\mem.mem[140][2] ));
 sg13g2_dfrbp_1 _19588_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net97),
    .D(_01224_),
    .Q_N(_08002_),
    .Q(\mem.mem[140][3] ));
 sg13g2_dfrbp_1 _19589_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net96),
    .D(_01225_),
    .Q_N(_08001_),
    .Q(\mem.mem[140][4] ));
 sg13g2_dfrbp_1 _19590_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net95),
    .D(_01226_),
    .Q_N(_08000_),
    .Q(\mem.mem[140][5] ));
 sg13g2_dfrbp_1 _19591_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net94),
    .D(_01227_),
    .Q_N(_07999_),
    .Q(\mem.mem[140][6] ));
 sg13g2_dfrbp_1 _19592_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net93),
    .D(_01228_),
    .Q_N(_07998_),
    .Q(\mem.mem[140][7] ));
 sg13g2_dfrbp_1 _19593_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net92),
    .D(_01229_),
    .Q_N(_07997_),
    .Q(\mem.mem[141][0] ));
 sg13g2_dfrbp_1 _19594_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net91),
    .D(_01230_),
    .Q_N(_07996_),
    .Q(\mem.mem[141][1] ));
 sg13g2_dfrbp_1 _19595_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net90),
    .D(_01231_),
    .Q_N(_07995_),
    .Q(\mem.mem[141][2] ));
 sg13g2_dfrbp_1 _19596_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net89),
    .D(_01232_),
    .Q_N(_07994_),
    .Q(\mem.mem[141][3] ));
 sg13g2_dfrbp_1 _19597_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net88),
    .D(_01233_),
    .Q_N(_07993_),
    .Q(\mem.mem[141][4] ));
 sg13g2_dfrbp_1 _19598_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net87),
    .D(_01234_),
    .Q_N(_07992_),
    .Q(\mem.mem[141][5] ));
 sg13g2_dfrbp_1 _19599_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net86),
    .D(_01235_),
    .Q_N(_07991_),
    .Q(\mem.mem[141][6] ));
 sg13g2_dfrbp_1 _19600_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net85),
    .D(_01236_),
    .Q_N(_07990_),
    .Q(\mem.mem[141][7] ));
 sg13g2_dfrbp_1 _19601_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net84),
    .D(_01237_),
    .Q_N(_07989_),
    .Q(\mem.mem[142][0] ));
 sg13g2_dfrbp_1 _19602_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net83),
    .D(_01238_),
    .Q_N(_07988_),
    .Q(\mem.mem[142][1] ));
 sg13g2_dfrbp_1 _19603_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net82),
    .D(_01239_),
    .Q_N(_07987_),
    .Q(\mem.mem[142][2] ));
 sg13g2_dfrbp_1 _19604_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net81),
    .D(_01240_),
    .Q_N(_07986_),
    .Q(\mem.mem[142][3] ));
 sg13g2_dfrbp_1 _19605_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net80),
    .D(_01241_),
    .Q_N(_07985_),
    .Q(\mem.mem[142][4] ));
 sg13g2_dfrbp_1 _19606_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net79),
    .D(_01242_),
    .Q_N(_07984_),
    .Q(\mem.mem[142][5] ));
 sg13g2_dfrbp_1 _19607_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net78),
    .D(_01243_),
    .Q_N(_07983_),
    .Q(\mem.mem[142][6] ));
 sg13g2_dfrbp_1 _19608_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net77),
    .D(_01244_),
    .Q_N(_07982_),
    .Q(\mem.mem[142][7] ));
 sg13g2_dfrbp_1 _19609_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net76),
    .D(_01245_),
    .Q_N(_07981_),
    .Q(\mem.mem[143][0] ));
 sg13g2_dfrbp_1 _19610_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net75),
    .D(_01246_),
    .Q_N(_07980_),
    .Q(\mem.mem[143][1] ));
 sg13g2_dfrbp_1 _19611_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net74),
    .D(_01247_),
    .Q_N(_07979_),
    .Q(\mem.mem[143][2] ));
 sg13g2_dfrbp_1 _19612_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net73),
    .D(_01248_),
    .Q_N(_07978_),
    .Q(\mem.mem[143][3] ));
 sg13g2_dfrbp_1 _19613_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net72),
    .D(_01249_),
    .Q_N(_07977_),
    .Q(\mem.mem[143][4] ));
 sg13g2_dfrbp_1 _19614_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net71),
    .D(_01250_),
    .Q_N(_07976_),
    .Q(\mem.mem[143][5] ));
 sg13g2_dfrbp_1 _19615_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net70),
    .D(_01251_),
    .Q_N(_07975_),
    .Q(\mem.mem[143][6] ));
 sg13g2_dfrbp_1 _19616_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net69),
    .D(_01252_),
    .Q_N(_07974_),
    .Q(\mem.mem[143][7] ));
 sg13g2_dfrbp_1 _19617_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net68),
    .D(_01253_),
    .Q_N(_07973_),
    .Q(\mem.mem[144][0] ));
 sg13g2_dfrbp_1 _19618_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net67),
    .D(_01254_),
    .Q_N(_07972_),
    .Q(\mem.mem[144][1] ));
 sg13g2_dfrbp_1 _19619_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net66),
    .D(_01255_),
    .Q_N(_07971_),
    .Q(\mem.mem[144][2] ));
 sg13g2_dfrbp_1 _19620_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net65),
    .D(net3905),
    .Q_N(_07970_),
    .Q(\mem.mem[144][3] ));
 sg13g2_dfrbp_1 _19621_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net64),
    .D(_01257_),
    .Q_N(_07969_),
    .Q(\mem.mem[144][4] ));
 sg13g2_dfrbp_1 _19622_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net63),
    .D(_01258_),
    .Q_N(_07968_),
    .Q(\mem.mem[144][5] ));
 sg13g2_dfrbp_1 _19623_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net62),
    .D(_01259_),
    .Q_N(_07967_),
    .Q(\mem.mem[144][6] ));
 sg13g2_dfrbp_1 _19624_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net61),
    .D(_01260_),
    .Q_N(_07966_),
    .Q(\mem.mem[144][7] ));
 sg13g2_dfrbp_1 _19625_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net60),
    .D(_01261_),
    .Q_N(_07965_),
    .Q(\mem.mem[145][0] ));
 sg13g2_dfrbp_1 _19626_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net59),
    .D(_01262_),
    .Q_N(_07964_),
    .Q(\mem.mem[145][1] ));
 sg13g2_dfrbp_1 _19627_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net58),
    .D(_01263_),
    .Q_N(_07963_),
    .Q(\mem.mem[145][2] ));
 sg13g2_dfrbp_1 _19628_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net57),
    .D(_01264_),
    .Q_N(_07962_),
    .Q(\mem.mem[145][3] ));
 sg13g2_dfrbp_1 _19629_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net56),
    .D(_01265_),
    .Q_N(_07961_),
    .Q(\mem.mem[145][4] ));
 sg13g2_dfrbp_1 _19630_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net55),
    .D(_01266_),
    .Q_N(_07960_),
    .Q(\mem.mem[145][5] ));
 sg13g2_dfrbp_1 _19631_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net54),
    .D(_01267_),
    .Q_N(_07959_),
    .Q(\mem.mem[145][6] ));
 sg13g2_dfrbp_1 _19632_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net53),
    .D(_01268_),
    .Q_N(_07958_),
    .Q(\mem.mem[145][7] ));
 sg13g2_dfrbp_1 _19633_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net52),
    .D(_01269_),
    .Q_N(_07957_),
    .Q(\mem.mem[146][0] ));
 sg13g2_dfrbp_1 _19634_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net51),
    .D(_01270_),
    .Q_N(_07956_),
    .Q(\mem.mem[146][1] ));
 sg13g2_dfrbp_1 _19635_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net50),
    .D(_01271_),
    .Q_N(_07955_),
    .Q(\mem.mem[146][2] ));
 sg13g2_dfrbp_1 _19636_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net49),
    .D(_01272_),
    .Q_N(_07954_),
    .Q(\mem.mem[146][3] ));
 sg13g2_dfrbp_1 _19637_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net48),
    .D(_01273_),
    .Q_N(_07953_),
    .Q(\mem.mem[146][4] ));
 sg13g2_dfrbp_1 _19638_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net47),
    .D(_01274_),
    .Q_N(_07952_),
    .Q(\mem.mem[146][5] ));
 sg13g2_dfrbp_1 _19639_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net46),
    .D(_01275_),
    .Q_N(_07951_),
    .Q(\mem.mem[146][6] ));
 sg13g2_dfrbp_1 _19640_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net45),
    .D(_01276_),
    .Q_N(_07950_),
    .Q(\mem.mem[146][7] ));
 sg13g2_dfrbp_1 _19641_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net44),
    .D(_01277_),
    .Q_N(_07949_),
    .Q(\mem.mem[147][0] ));
 sg13g2_dfrbp_1 _19642_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net43),
    .D(_01278_),
    .Q_N(_07948_),
    .Q(\mem.mem[147][1] ));
 sg13g2_dfrbp_1 _19643_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net42),
    .D(_01279_),
    .Q_N(_07947_),
    .Q(\mem.mem[147][2] ));
 sg13g2_dfrbp_1 _19644_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net41),
    .D(_01280_),
    .Q_N(_07946_),
    .Q(\mem.mem[147][3] ));
 sg13g2_dfrbp_1 _19645_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net40),
    .D(_01281_),
    .Q_N(_07945_),
    .Q(\mem.mem[147][4] ));
 sg13g2_dfrbp_1 _19646_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net39),
    .D(_01282_),
    .Q_N(_07944_),
    .Q(\mem.mem[147][5] ));
 sg13g2_dfrbp_1 _19647_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net38),
    .D(_01283_),
    .Q_N(_07943_),
    .Q(\mem.mem[147][6] ));
 sg13g2_dfrbp_1 _19648_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net37),
    .D(_01284_),
    .Q_N(_07942_),
    .Q(\mem.mem[147][7] ));
 sg13g2_dfrbp_1 _19649_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net36),
    .D(_01285_),
    .Q_N(_07941_),
    .Q(\mem.mem[148][0] ));
 sg13g2_dfrbp_1 _19650_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net35),
    .D(_01286_),
    .Q_N(_07940_),
    .Q(\mem.mem[148][1] ));
 sg13g2_dfrbp_1 _19651_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net34),
    .D(_01287_),
    .Q_N(_07939_),
    .Q(\mem.mem[148][2] ));
 sg13g2_dfrbp_1 _19652_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net33),
    .D(_01288_),
    .Q_N(_07938_),
    .Q(\mem.mem[148][3] ));
 sg13g2_dfrbp_1 _19653_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net32),
    .D(_01289_),
    .Q_N(_07937_),
    .Q(\mem.mem[148][4] ));
 sg13g2_dfrbp_1 _19654_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net31),
    .D(_01290_),
    .Q_N(_07936_),
    .Q(\mem.mem[148][5] ));
 sg13g2_dfrbp_1 _19655_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net30),
    .D(_01291_),
    .Q_N(_07935_),
    .Q(\mem.mem[148][6] ));
 sg13g2_dfrbp_1 _19656_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net29),
    .D(_01292_),
    .Q_N(_07934_),
    .Q(\mem.mem[148][7] ));
 sg13g2_dfrbp_1 _19657_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net28),
    .D(_01293_),
    .Q_N(_07933_),
    .Q(\mem.mem[14][0] ));
 sg13g2_dfrbp_1 _19658_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net27),
    .D(_01294_),
    .Q_N(_07932_),
    .Q(\mem.mem[14][1] ));
 sg13g2_dfrbp_1 _19659_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net26),
    .D(_01295_),
    .Q_N(_07931_),
    .Q(\mem.mem[14][2] ));
 sg13g2_dfrbp_1 _19660_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net25),
    .D(_01296_),
    .Q_N(_07930_),
    .Q(\mem.mem[14][3] ));
 sg13g2_dfrbp_1 _19661_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net24),
    .D(_01297_),
    .Q_N(_07929_),
    .Q(\mem.mem[14][4] ));
 sg13g2_dfrbp_1 _19662_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2129),
    .D(_01298_),
    .Q_N(_07928_),
    .Q(\mem.mem[14][5] ));
 sg13g2_dfrbp_1 _19663_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2128),
    .D(_01299_),
    .Q_N(_07927_),
    .Q(\mem.mem[14][6] ));
 sg13g2_dfrbp_1 _19664_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2127),
    .D(_01300_),
    .Q_N(_07926_),
    .Q(\mem.mem[14][7] ));
 sg13g2_dfrbp_1 _19665_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2126),
    .D(_01301_),
    .Q_N(_07925_),
    .Q(\mem.mem[150][0] ));
 sg13g2_dfrbp_1 _19666_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2125),
    .D(_01302_),
    .Q_N(_07924_),
    .Q(\mem.mem[150][1] ));
 sg13g2_dfrbp_1 _19667_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2124),
    .D(_01303_),
    .Q_N(_07923_),
    .Q(\mem.mem[150][2] ));
 sg13g2_dfrbp_1 _19668_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2123),
    .D(_01304_),
    .Q_N(_07922_),
    .Q(\mem.mem[150][3] ));
 sg13g2_dfrbp_1 _19669_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2122),
    .D(_01305_),
    .Q_N(_07921_),
    .Q(\mem.mem[150][4] ));
 sg13g2_dfrbp_1 _19670_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2121),
    .D(_01306_),
    .Q_N(_07920_),
    .Q(\mem.mem[150][5] ));
 sg13g2_dfrbp_1 _19671_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2120),
    .D(_01307_),
    .Q_N(_07919_),
    .Q(\mem.mem[150][6] ));
 sg13g2_dfrbp_1 _19672_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2119),
    .D(_01308_),
    .Q_N(_07918_),
    .Q(\mem.mem[150][7] ));
 sg13g2_dfrbp_1 _19673_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net2118),
    .D(_01309_),
    .Q_N(_07917_),
    .Q(\mem.mem[151][0] ));
 sg13g2_dfrbp_1 _19674_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2117),
    .D(_01310_),
    .Q_N(_07916_),
    .Q(\mem.mem[151][1] ));
 sg13g2_dfrbp_1 _19675_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net2116),
    .D(_01311_),
    .Q_N(_07915_),
    .Q(\mem.mem[151][2] ));
 sg13g2_dfrbp_1 _19676_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2115),
    .D(_01312_),
    .Q_N(_07914_),
    .Q(\mem.mem[151][3] ));
 sg13g2_dfrbp_1 _19677_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2114),
    .D(_01313_),
    .Q_N(_07913_),
    .Q(\mem.mem[151][4] ));
 sg13g2_dfrbp_1 _19678_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2113),
    .D(_01314_),
    .Q_N(_07912_),
    .Q(\mem.mem[151][5] ));
 sg13g2_dfrbp_1 _19679_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2112),
    .D(_01315_),
    .Q_N(_07911_),
    .Q(\mem.mem[151][6] ));
 sg13g2_dfrbp_1 _19680_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2111),
    .D(_01316_),
    .Q_N(_07910_),
    .Q(\mem.mem[151][7] ));
 sg13g2_dfrbp_1 _19681_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2110),
    .D(_01317_),
    .Q_N(_07909_),
    .Q(\mem.mem[152][0] ));
 sg13g2_dfrbp_1 _19682_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2109),
    .D(_01318_),
    .Q_N(_07908_),
    .Q(\mem.mem[152][1] ));
 sg13g2_dfrbp_1 _19683_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2108),
    .D(_01319_),
    .Q_N(_07907_),
    .Q(\mem.mem[152][2] ));
 sg13g2_dfrbp_1 _19684_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2107),
    .D(_01320_),
    .Q_N(_07906_),
    .Q(\mem.mem[152][3] ));
 sg13g2_dfrbp_1 _19685_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2106),
    .D(_01321_),
    .Q_N(_07905_),
    .Q(\mem.mem[152][4] ));
 sg13g2_dfrbp_1 _19686_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2105),
    .D(_01322_),
    .Q_N(_07904_),
    .Q(\mem.mem[152][5] ));
 sg13g2_dfrbp_1 _19687_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2104),
    .D(_01323_),
    .Q_N(_07903_),
    .Q(\mem.mem[152][6] ));
 sg13g2_dfrbp_1 _19688_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2103),
    .D(_01324_),
    .Q_N(_07902_),
    .Q(\mem.mem[152][7] ));
 sg13g2_dfrbp_1 _19689_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2102),
    .D(_01325_),
    .Q_N(_07901_),
    .Q(\mem.mem[153][0] ));
 sg13g2_dfrbp_1 _19690_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2101),
    .D(_01326_),
    .Q_N(_07900_),
    .Q(\mem.mem[153][1] ));
 sg13g2_dfrbp_1 _19691_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2100),
    .D(_01327_),
    .Q_N(_07899_),
    .Q(\mem.mem[153][2] ));
 sg13g2_dfrbp_1 _19692_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2099),
    .D(_01328_),
    .Q_N(_07898_),
    .Q(\mem.mem[153][3] ));
 sg13g2_dfrbp_1 _19693_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2098),
    .D(_01329_),
    .Q_N(_07897_),
    .Q(\mem.mem[153][4] ));
 sg13g2_dfrbp_1 _19694_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2097),
    .D(_01330_),
    .Q_N(_07896_),
    .Q(\mem.mem[153][5] ));
 sg13g2_dfrbp_1 _19695_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2096),
    .D(_01331_),
    .Q_N(_07895_),
    .Q(\mem.mem[153][6] ));
 sg13g2_dfrbp_1 _19696_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2095),
    .D(_01332_),
    .Q_N(_07894_),
    .Q(\mem.mem[153][7] ));
 sg13g2_dfrbp_1 _19697_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2094),
    .D(_01333_),
    .Q_N(_07893_),
    .Q(\mem.mem[154][0] ));
 sg13g2_dfrbp_1 _19698_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2093),
    .D(_01334_),
    .Q_N(_07892_),
    .Q(\mem.mem[154][1] ));
 sg13g2_dfrbp_1 _19699_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2092),
    .D(_01335_),
    .Q_N(_07891_),
    .Q(\mem.mem[154][2] ));
 sg13g2_dfrbp_1 _19700_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2091),
    .D(_01336_),
    .Q_N(_07890_),
    .Q(\mem.mem[154][3] ));
 sg13g2_dfrbp_1 _19701_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2090),
    .D(_01337_),
    .Q_N(_07889_),
    .Q(\mem.mem[154][4] ));
 sg13g2_dfrbp_1 _19702_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2089),
    .D(_01338_),
    .Q_N(_07888_),
    .Q(\mem.mem[154][5] ));
 sg13g2_dfrbp_1 _19703_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2088),
    .D(_01339_),
    .Q_N(_07887_),
    .Q(\mem.mem[154][6] ));
 sg13g2_dfrbp_1 _19704_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2087),
    .D(_01340_),
    .Q_N(_07886_),
    .Q(\mem.mem[154][7] ));
 sg13g2_dfrbp_1 _19705_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2086),
    .D(_01341_),
    .Q_N(_07885_),
    .Q(\mem.mem[155][0] ));
 sg13g2_dfrbp_1 _19706_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2085),
    .D(_01342_),
    .Q_N(_07884_),
    .Q(\mem.mem[155][1] ));
 sg13g2_dfrbp_1 _19707_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2084),
    .D(_01343_),
    .Q_N(_07883_),
    .Q(\mem.mem[155][2] ));
 sg13g2_dfrbp_1 _19708_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2083),
    .D(_01344_),
    .Q_N(_07882_),
    .Q(\mem.mem[155][3] ));
 sg13g2_dfrbp_1 _19709_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2082),
    .D(_01345_),
    .Q_N(_07881_),
    .Q(\mem.mem[155][4] ));
 sg13g2_dfrbp_1 _19710_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2081),
    .D(_01346_),
    .Q_N(_07880_),
    .Q(\mem.mem[155][5] ));
 sg13g2_dfrbp_1 _19711_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2080),
    .D(_01347_),
    .Q_N(_07879_),
    .Q(\mem.mem[155][6] ));
 sg13g2_dfrbp_1 _19712_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2079),
    .D(_01348_),
    .Q_N(_07878_),
    .Q(\mem.mem[155][7] ));
 sg13g2_dfrbp_1 _19713_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2078),
    .D(_01349_),
    .Q_N(_07877_),
    .Q(\mem.mem[156][0] ));
 sg13g2_dfrbp_1 _19714_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2077),
    .D(_01350_),
    .Q_N(_07876_),
    .Q(\mem.mem[156][1] ));
 sg13g2_dfrbp_1 _19715_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2076),
    .D(_01351_),
    .Q_N(_07875_),
    .Q(\mem.mem[156][2] ));
 sg13g2_dfrbp_1 _19716_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2075),
    .D(_01352_),
    .Q_N(_07874_),
    .Q(\mem.mem[156][3] ));
 sg13g2_dfrbp_1 _19717_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2074),
    .D(_01353_),
    .Q_N(_07873_),
    .Q(\mem.mem[156][4] ));
 sg13g2_dfrbp_1 _19718_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2073),
    .D(_01354_),
    .Q_N(_07872_),
    .Q(\mem.mem[156][5] ));
 sg13g2_dfrbp_1 _19719_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2072),
    .D(_01355_),
    .Q_N(_07871_),
    .Q(\mem.mem[156][6] ));
 sg13g2_dfrbp_1 _19720_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2071),
    .D(_01356_),
    .Q_N(_07870_),
    .Q(\mem.mem[156][7] ));
 sg13g2_dfrbp_1 _19721_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2070),
    .D(_01357_),
    .Q_N(_07869_),
    .Q(\mem.mem[157][0] ));
 sg13g2_dfrbp_1 _19722_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2069),
    .D(_01358_),
    .Q_N(_07868_),
    .Q(\mem.mem[157][1] ));
 sg13g2_dfrbp_1 _19723_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2068),
    .D(_01359_),
    .Q_N(_07867_),
    .Q(\mem.mem[157][2] ));
 sg13g2_dfrbp_1 _19724_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2067),
    .D(_01360_),
    .Q_N(_07866_),
    .Q(\mem.mem[157][3] ));
 sg13g2_dfrbp_1 _19725_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2066),
    .D(_01361_),
    .Q_N(_07865_),
    .Q(\mem.mem[157][4] ));
 sg13g2_dfrbp_1 _19726_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2065),
    .D(_01362_),
    .Q_N(_07864_),
    .Q(\mem.mem[157][5] ));
 sg13g2_dfrbp_1 _19727_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2064),
    .D(_01363_),
    .Q_N(_07863_),
    .Q(\mem.mem[157][6] ));
 sg13g2_dfrbp_1 _19728_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2063),
    .D(_01364_),
    .Q_N(_07862_),
    .Q(\mem.mem[157][7] ));
 sg13g2_dfrbp_1 _19729_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2062),
    .D(_01365_),
    .Q_N(_07861_),
    .Q(\mem.mem[158][0] ));
 sg13g2_dfrbp_1 _19730_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2061),
    .D(_01366_),
    .Q_N(_07860_),
    .Q(\mem.mem[158][1] ));
 sg13g2_dfrbp_1 _19731_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2060),
    .D(_01367_),
    .Q_N(_07859_),
    .Q(\mem.mem[158][2] ));
 sg13g2_dfrbp_1 _19732_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2059),
    .D(_01368_),
    .Q_N(_07858_),
    .Q(\mem.mem[158][3] ));
 sg13g2_dfrbp_1 _19733_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2058),
    .D(_01369_),
    .Q_N(_07857_),
    .Q(\mem.mem[158][4] ));
 sg13g2_dfrbp_1 _19734_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2057),
    .D(_01370_),
    .Q_N(_07856_),
    .Q(\mem.mem[158][5] ));
 sg13g2_dfrbp_1 _19735_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2056),
    .D(_01371_),
    .Q_N(_07855_),
    .Q(\mem.mem[158][6] ));
 sg13g2_dfrbp_1 _19736_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2055),
    .D(_01372_),
    .Q_N(_07854_),
    .Q(\mem.mem[158][7] ));
 sg13g2_dfrbp_1 _19737_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2054),
    .D(_01373_),
    .Q_N(_07853_),
    .Q(\mem.mem[15][0] ));
 sg13g2_dfrbp_1 _19738_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2053),
    .D(_01374_),
    .Q_N(_07852_),
    .Q(\mem.mem[15][1] ));
 sg13g2_dfrbp_1 _19739_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2052),
    .D(_01375_),
    .Q_N(_07851_),
    .Q(\mem.mem[15][2] ));
 sg13g2_dfrbp_1 _19740_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2051),
    .D(_01376_),
    .Q_N(_07850_),
    .Q(\mem.mem[15][3] ));
 sg13g2_dfrbp_1 _19741_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2050),
    .D(_01377_),
    .Q_N(_07849_),
    .Q(\mem.mem[15][4] ));
 sg13g2_dfrbp_1 _19742_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2049),
    .D(_01378_),
    .Q_N(_07848_),
    .Q(\mem.mem[15][5] ));
 sg13g2_dfrbp_1 _19743_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net2048),
    .D(_01379_),
    .Q_N(_07847_),
    .Q(\mem.mem[15][6] ));
 sg13g2_dfrbp_1 _19744_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2047),
    .D(_01380_),
    .Q_N(_07846_),
    .Q(\mem.mem[15][7] ));
 sg13g2_dfrbp_1 _19745_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2046),
    .D(_01381_),
    .Q_N(_07845_),
    .Q(\mem.mem[160][0] ));
 sg13g2_dfrbp_1 _19746_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2045),
    .D(_01382_),
    .Q_N(_07844_),
    .Q(\mem.mem[160][1] ));
 sg13g2_dfrbp_1 _19747_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2044),
    .D(_01383_),
    .Q_N(_07843_),
    .Q(\mem.mem[160][2] ));
 sg13g2_dfrbp_1 _19748_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2043),
    .D(_01384_),
    .Q_N(_07842_),
    .Q(\mem.mem[160][3] ));
 sg13g2_dfrbp_1 _19749_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2042),
    .D(_01385_),
    .Q_N(_07841_),
    .Q(\mem.mem[160][4] ));
 sg13g2_dfrbp_1 _19750_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2041),
    .D(_01386_),
    .Q_N(_07840_),
    .Q(\mem.mem[160][5] ));
 sg13g2_dfrbp_1 _19751_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2040),
    .D(_01387_),
    .Q_N(_07839_),
    .Q(\mem.mem[160][6] ));
 sg13g2_dfrbp_1 _19752_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2039),
    .D(_01388_),
    .Q_N(_07838_),
    .Q(\mem.mem[160][7] ));
 sg13g2_dfrbp_1 _19753_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2038),
    .D(_01389_),
    .Q_N(_07837_),
    .Q(\mem.mem[161][0] ));
 sg13g2_dfrbp_1 _19754_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2037),
    .D(_01390_),
    .Q_N(_07836_),
    .Q(\mem.mem[161][1] ));
 sg13g2_dfrbp_1 _19755_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2036),
    .D(_01391_),
    .Q_N(_07835_),
    .Q(\mem.mem[161][2] ));
 sg13g2_dfrbp_1 _19756_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2035),
    .D(_01392_),
    .Q_N(_07834_),
    .Q(\mem.mem[161][3] ));
 sg13g2_dfrbp_1 _19757_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2034),
    .D(_01393_),
    .Q_N(_07833_),
    .Q(\mem.mem[161][4] ));
 sg13g2_dfrbp_1 _19758_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2033),
    .D(_01394_),
    .Q_N(_07832_),
    .Q(\mem.mem[161][5] ));
 sg13g2_dfrbp_1 _19759_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2032),
    .D(_01395_),
    .Q_N(_07831_),
    .Q(\mem.mem[161][6] ));
 sg13g2_dfrbp_1 _19760_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2031),
    .D(_01396_),
    .Q_N(_07830_),
    .Q(\mem.mem[161][7] ));
 sg13g2_dfrbp_1 _19761_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2030),
    .D(_01397_),
    .Q_N(_07829_),
    .Q(\mem.mem[162][0] ));
 sg13g2_dfrbp_1 _19762_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2029),
    .D(_01398_),
    .Q_N(_07828_),
    .Q(\mem.mem[162][1] ));
 sg13g2_dfrbp_1 _19763_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2028),
    .D(_01399_),
    .Q_N(_07827_),
    .Q(\mem.mem[162][2] ));
 sg13g2_dfrbp_1 _19764_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2027),
    .D(_01400_),
    .Q_N(_07826_),
    .Q(\mem.mem[162][3] ));
 sg13g2_dfrbp_1 _19765_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2026),
    .D(_01401_),
    .Q_N(_07825_),
    .Q(\mem.mem[162][4] ));
 sg13g2_dfrbp_1 _19766_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2025),
    .D(_01402_),
    .Q_N(_07824_),
    .Q(\mem.mem[162][5] ));
 sg13g2_dfrbp_1 _19767_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2024),
    .D(_01403_),
    .Q_N(_07823_),
    .Q(\mem.mem[162][6] ));
 sg13g2_dfrbp_1 _19768_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2023),
    .D(_01404_),
    .Q_N(_07822_),
    .Q(\mem.mem[162][7] ));
 sg13g2_dfrbp_1 _19769_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2022),
    .D(_01405_),
    .Q_N(_07821_),
    .Q(\mem.mem[163][0] ));
 sg13g2_dfrbp_1 _19770_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2021),
    .D(_01406_),
    .Q_N(_07820_),
    .Q(\mem.mem[163][1] ));
 sg13g2_dfrbp_1 _19771_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2020),
    .D(_01407_),
    .Q_N(_07819_),
    .Q(\mem.mem[163][2] ));
 sg13g2_dfrbp_1 _19772_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2019),
    .D(_01408_),
    .Q_N(_07818_),
    .Q(\mem.mem[163][3] ));
 sg13g2_dfrbp_1 _19773_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2018),
    .D(_01409_),
    .Q_N(_07817_),
    .Q(\mem.mem[163][4] ));
 sg13g2_dfrbp_1 _19774_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2017),
    .D(_01410_),
    .Q_N(_07816_),
    .Q(\mem.mem[163][5] ));
 sg13g2_dfrbp_1 _19775_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2016),
    .D(_01411_),
    .Q_N(_07815_),
    .Q(\mem.mem[163][6] ));
 sg13g2_dfrbp_1 _19776_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2015),
    .D(_01412_),
    .Q_N(_07814_),
    .Q(\mem.mem[163][7] ));
 sg13g2_dfrbp_1 _19777_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2014),
    .D(_01413_),
    .Q_N(_07813_),
    .Q(\mem.mem[164][0] ));
 sg13g2_dfrbp_1 _19778_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2013),
    .D(_01414_),
    .Q_N(_07812_),
    .Q(\mem.mem[164][1] ));
 sg13g2_dfrbp_1 _19779_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2012),
    .D(_01415_),
    .Q_N(_07811_),
    .Q(\mem.mem[164][2] ));
 sg13g2_dfrbp_1 _19780_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2011),
    .D(_01416_),
    .Q_N(_07810_),
    .Q(\mem.mem[164][3] ));
 sg13g2_dfrbp_1 _19781_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2010),
    .D(_01417_),
    .Q_N(_07809_),
    .Q(\mem.mem[164][4] ));
 sg13g2_dfrbp_1 _19782_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2009),
    .D(_01418_),
    .Q_N(_07808_),
    .Q(\mem.mem[164][5] ));
 sg13g2_dfrbp_1 _19783_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2008),
    .D(_01419_),
    .Q_N(_07807_),
    .Q(\mem.mem[164][6] ));
 sg13g2_dfrbp_1 _19784_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2007),
    .D(_01420_),
    .Q_N(_07806_),
    .Q(\mem.mem[164][7] ));
 sg13g2_dfrbp_1 _19785_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2006),
    .D(_01421_),
    .Q_N(_07805_),
    .Q(\mem.mem[165][0] ));
 sg13g2_dfrbp_1 _19786_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2005),
    .D(_01422_),
    .Q_N(_07804_),
    .Q(\mem.mem[165][1] ));
 sg13g2_dfrbp_1 _19787_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2004),
    .D(_01423_),
    .Q_N(_07803_),
    .Q(\mem.mem[165][2] ));
 sg13g2_dfrbp_1 _19788_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2003),
    .D(_01424_),
    .Q_N(_07802_),
    .Q(\mem.mem[165][3] ));
 sg13g2_dfrbp_1 _19789_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2002),
    .D(_01425_),
    .Q_N(_07801_),
    .Q(\mem.mem[165][4] ));
 sg13g2_dfrbp_1 _19790_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2001),
    .D(_01426_),
    .Q_N(_07800_),
    .Q(\mem.mem[165][5] ));
 sg13g2_dfrbp_1 _19791_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2000),
    .D(_01427_),
    .Q_N(_07799_),
    .Q(\mem.mem[165][6] ));
 sg13g2_dfrbp_1 _19792_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1999),
    .D(_01428_),
    .Q_N(_07798_),
    .Q(\mem.mem[165][7] ));
 sg13g2_dfrbp_1 _19793_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1998),
    .D(_01429_),
    .Q_N(_07797_),
    .Q(\mem.mem[166][0] ));
 sg13g2_dfrbp_1 _19794_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1997),
    .D(_01430_),
    .Q_N(_07796_),
    .Q(\mem.mem[166][1] ));
 sg13g2_dfrbp_1 _19795_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1996),
    .D(_01431_),
    .Q_N(_07795_),
    .Q(\mem.mem[166][2] ));
 sg13g2_dfrbp_1 _19796_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1995),
    .D(_01432_),
    .Q_N(_07794_),
    .Q(\mem.mem[166][3] ));
 sg13g2_dfrbp_1 _19797_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1994),
    .D(_01433_),
    .Q_N(_07793_),
    .Q(\mem.mem[166][4] ));
 sg13g2_dfrbp_1 _19798_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1993),
    .D(_01434_),
    .Q_N(_07792_),
    .Q(\mem.mem[166][5] ));
 sg13g2_dfrbp_1 _19799_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1992),
    .D(_01435_),
    .Q_N(_07791_),
    .Q(\mem.mem[166][6] ));
 sg13g2_dfrbp_1 _19800_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1991),
    .D(net3386),
    .Q_N(_07790_),
    .Q(\mem.mem[166][7] ));
 sg13g2_dfrbp_1 _19801_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1990),
    .D(_01437_),
    .Q_N(_07789_),
    .Q(\mem.mem[167][0] ));
 sg13g2_dfrbp_1 _19802_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1989),
    .D(_01438_),
    .Q_N(_07788_),
    .Q(\mem.mem[167][1] ));
 sg13g2_dfrbp_1 _19803_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1988),
    .D(_01439_),
    .Q_N(_07787_),
    .Q(\mem.mem[167][2] ));
 sg13g2_dfrbp_1 _19804_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1987),
    .D(_01440_),
    .Q_N(_07786_),
    .Q(\mem.mem[167][3] ));
 sg13g2_dfrbp_1 _19805_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1986),
    .D(_01441_),
    .Q_N(_07785_),
    .Q(\mem.mem[167][4] ));
 sg13g2_dfrbp_1 _19806_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1985),
    .D(_01442_),
    .Q_N(_07784_),
    .Q(\mem.mem[167][5] ));
 sg13g2_dfrbp_1 _19807_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1984),
    .D(_01443_),
    .Q_N(_07783_),
    .Q(\mem.mem[167][6] ));
 sg13g2_dfrbp_1 _19808_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1983),
    .D(_01444_),
    .Q_N(_07782_),
    .Q(\mem.mem[167][7] ));
 sg13g2_dfrbp_1 _19809_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1982),
    .D(_01445_),
    .Q_N(_07781_),
    .Q(\mem.mem[168][0] ));
 sg13g2_dfrbp_1 _19810_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1981),
    .D(_01446_),
    .Q_N(_07780_),
    .Q(\mem.mem[168][1] ));
 sg13g2_dfrbp_1 _19811_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1980),
    .D(_01447_),
    .Q_N(_07779_),
    .Q(\mem.mem[168][2] ));
 sg13g2_dfrbp_1 _19812_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1979),
    .D(_01448_),
    .Q_N(_07778_),
    .Q(\mem.mem[168][3] ));
 sg13g2_dfrbp_1 _19813_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1978),
    .D(_01449_),
    .Q_N(_07777_),
    .Q(\mem.mem[168][4] ));
 sg13g2_dfrbp_1 _19814_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1977),
    .D(_01450_),
    .Q_N(_07776_),
    .Q(\mem.mem[168][5] ));
 sg13g2_dfrbp_1 _19815_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1976),
    .D(_01451_),
    .Q_N(_07775_),
    .Q(\mem.mem[168][6] ));
 sg13g2_dfrbp_1 _19816_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1975),
    .D(_01452_),
    .Q_N(_07774_),
    .Q(\mem.mem[168][7] ));
 sg13g2_dfrbp_1 _19817_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1974),
    .D(_01453_),
    .Q_N(_07773_),
    .Q(\mem.mem[16][0] ));
 sg13g2_dfrbp_1 _19818_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1973),
    .D(_01454_),
    .Q_N(_07772_),
    .Q(\mem.mem[16][1] ));
 sg13g2_dfrbp_1 _19819_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1972),
    .D(_01455_),
    .Q_N(_07771_),
    .Q(\mem.mem[16][2] ));
 sg13g2_dfrbp_1 _19820_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1971),
    .D(_01456_),
    .Q_N(_07770_),
    .Q(\mem.mem[16][3] ));
 sg13g2_dfrbp_1 _19821_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1970),
    .D(_01457_),
    .Q_N(_07769_),
    .Q(\mem.mem[16][4] ));
 sg13g2_dfrbp_1 _19822_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1969),
    .D(_01458_),
    .Q_N(_07768_),
    .Q(\mem.mem[16][5] ));
 sg13g2_dfrbp_1 _19823_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1968),
    .D(_01459_),
    .Q_N(_07767_),
    .Q(\mem.mem[16][6] ));
 sg13g2_dfrbp_1 _19824_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1967),
    .D(_01460_),
    .Q_N(_07766_),
    .Q(\mem.mem[16][7] ));
 sg13g2_dfrbp_1 _19825_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1966),
    .D(_01461_),
    .Q_N(_07765_),
    .Q(\mem.mem[170][0] ));
 sg13g2_dfrbp_1 _19826_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1965),
    .D(_01462_),
    .Q_N(_07764_),
    .Q(\mem.mem[170][1] ));
 sg13g2_dfrbp_1 _19827_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1964),
    .D(_01463_),
    .Q_N(_07763_),
    .Q(\mem.mem[170][2] ));
 sg13g2_dfrbp_1 _19828_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1963),
    .D(_01464_),
    .Q_N(_07762_),
    .Q(\mem.mem[170][3] ));
 sg13g2_dfrbp_1 _19829_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1962),
    .D(_01465_),
    .Q_N(_07761_),
    .Q(\mem.mem[170][4] ));
 sg13g2_dfrbp_1 _19830_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1961),
    .D(_01466_),
    .Q_N(_07760_),
    .Q(\mem.mem[170][5] ));
 sg13g2_dfrbp_1 _19831_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1960),
    .D(_01467_),
    .Q_N(_07759_),
    .Q(\mem.mem[170][6] ));
 sg13g2_dfrbp_1 _19832_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1959),
    .D(_01468_),
    .Q_N(_07758_),
    .Q(\mem.mem[170][7] ));
 sg13g2_dfrbp_1 _19833_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1958),
    .D(_01469_),
    .Q_N(_07757_),
    .Q(\mem.mem[171][0] ));
 sg13g2_dfrbp_1 _19834_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1957),
    .D(_01470_),
    .Q_N(_07756_),
    .Q(\mem.mem[171][1] ));
 sg13g2_dfrbp_1 _19835_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1956),
    .D(_01471_),
    .Q_N(_07755_),
    .Q(\mem.mem[171][2] ));
 sg13g2_dfrbp_1 _19836_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1955),
    .D(_01472_),
    .Q_N(_07754_),
    .Q(\mem.mem[171][3] ));
 sg13g2_dfrbp_1 _19837_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1954),
    .D(_01473_),
    .Q_N(_07753_),
    .Q(\mem.mem[171][4] ));
 sg13g2_dfrbp_1 _19838_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1953),
    .D(_01474_),
    .Q_N(_07752_),
    .Q(\mem.mem[171][5] ));
 sg13g2_dfrbp_1 _19839_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1952),
    .D(_01475_),
    .Q_N(_07751_),
    .Q(\mem.mem[171][6] ));
 sg13g2_dfrbp_1 _19840_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1951),
    .D(_01476_),
    .Q_N(_07750_),
    .Q(\mem.mem[171][7] ));
 sg13g2_dfrbp_1 _19841_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1950),
    .D(_01477_),
    .Q_N(_07749_),
    .Q(\mem.mem[172][0] ));
 sg13g2_dfrbp_1 _19842_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1949),
    .D(_01478_),
    .Q_N(_07748_),
    .Q(\mem.mem[172][1] ));
 sg13g2_dfrbp_1 _19843_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1948),
    .D(_01479_),
    .Q_N(_07747_),
    .Q(\mem.mem[172][2] ));
 sg13g2_dfrbp_1 _19844_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1947),
    .D(_01480_),
    .Q_N(_07746_),
    .Q(\mem.mem[172][3] ));
 sg13g2_dfrbp_1 _19845_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1946),
    .D(_01481_),
    .Q_N(_07745_),
    .Q(\mem.mem[172][4] ));
 sg13g2_dfrbp_1 _19846_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1945),
    .D(_01482_),
    .Q_N(_07744_),
    .Q(\mem.mem[172][5] ));
 sg13g2_dfrbp_1 _19847_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1944),
    .D(_01483_),
    .Q_N(_07743_),
    .Q(\mem.mem[172][6] ));
 sg13g2_dfrbp_1 _19848_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1943),
    .D(_01484_),
    .Q_N(_07742_),
    .Q(\mem.mem[172][7] ));
 sg13g2_dfrbp_1 _19849_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1942),
    .D(_01485_),
    .Q_N(_07741_),
    .Q(\mem.mem[173][0] ));
 sg13g2_dfrbp_1 _19850_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1941),
    .D(_01486_),
    .Q_N(_07740_),
    .Q(\mem.mem[173][1] ));
 sg13g2_dfrbp_1 _19851_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1940),
    .D(_01487_),
    .Q_N(_07739_),
    .Q(\mem.mem[173][2] ));
 sg13g2_dfrbp_1 _19852_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1939),
    .D(_01488_),
    .Q_N(_07738_),
    .Q(\mem.mem[173][3] ));
 sg13g2_dfrbp_1 _19853_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1938),
    .D(_01489_),
    .Q_N(_07737_),
    .Q(\mem.mem[173][4] ));
 sg13g2_dfrbp_1 _19854_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1937),
    .D(_01490_),
    .Q_N(_07736_),
    .Q(\mem.mem[173][5] ));
 sg13g2_dfrbp_1 _19855_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1936),
    .D(_01491_),
    .Q_N(_07735_),
    .Q(\mem.mem[173][6] ));
 sg13g2_dfrbp_1 _19856_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1935),
    .D(_01492_),
    .Q_N(_07734_),
    .Q(\mem.mem[173][7] ));
 sg13g2_dfrbp_1 _19857_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1934),
    .D(_01493_),
    .Q_N(_07733_),
    .Q(\mem.mem[174][0] ));
 sg13g2_dfrbp_1 _19858_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1933),
    .D(_01494_),
    .Q_N(_07732_),
    .Q(\mem.mem[174][1] ));
 sg13g2_dfrbp_1 _19859_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1932),
    .D(_01495_),
    .Q_N(_07731_),
    .Q(\mem.mem[174][2] ));
 sg13g2_dfrbp_1 _19860_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1931),
    .D(_01496_),
    .Q_N(_07730_),
    .Q(\mem.mem[174][3] ));
 sg13g2_dfrbp_1 _19861_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1930),
    .D(_01497_),
    .Q_N(_07729_),
    .Q(\mem.mem[174][4] ));
 sg13g2_dfrbp_1 _19862_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1929),
    .D(_01498_),
    .Q_N(_07728_),
    .Q(\mem.mem[174][5] ));
 sg13g2_dfrbp_1 _19863_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1928),
    .D(_01499_),
    .Q_N(_07727_),
    .Q(\mem.mem[174][6] ));
 sg13g2_dfrbp_1 _19864_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1927),
    .D(_01500_),
    .Q_N(_07726_),
    .Q(\mem.mem[174][7] ));
 sg13g2_dfrbp_1 _19865_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1926),
    .D(_01501_),
    .Q_N(_07725_),
    .Q(\mem.mem[175][0] ));
 sg13g2_dfrbp_1 _19866_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1925),
    .D(_01502_),
    .Q_N(_07724_),
    .Q(\mem.mem[175][1] ));
 sg13g2_dfrbp_1 _19867_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1924),
    .D(_01503_),
    .Q_N(_07723_),
    .Q(\mem.mem[175][2] ));
 sg13g2_dfrbp_1 _19868_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1923),
    .D(_01504_),
    .Q_N(_07722_),
    .Q(\mem.mem[175][3] ));
 sg13g2_dfrbp_1 _19869_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1922),
    .D(_01505_),
    .Q_N(_07721_),
    .Q(\mem.mem[175][4] ));
 sg13g2_dfrbp_1 _19870_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1921),
    .D(_01506_),
    .Q_N(_07720_),
    .Q(\mem.mem[175][5] ));
 sg13g2_dfrbp_1 _19871_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1920),
    .D(_01507_),
    .Q_N(_07719_),
    .Q(\mem.mem[175][6] ));
 sg13g2_dfrbp_1 _19872_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1919),
    .D(_01508_),
    .Q_N(_07718_),
    .Q(\mem.mem[175][7] ));
 sg13g2_dfrbp_1 _19873_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1918),
    .D(_01509_),
    .Q_N(_07717_),
    .Q(\mem.mem[176][0] ));
 sg13g2_dfrbp_1 _19874_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1917),
    .D(_01510_),
    .Q_N(_07716_),
    .Q(\mem.mem[176][1] ));
 sg13g2_dfrbp_1 _19875_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1916),
    .D(_01511_),
    .Q_N(_07715_),
    .Q(\mem.mem[176][2] ));
 sg13g2_dfrbp_1 _19876_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1915),
    .D(_01512_),
    .Q_N(_07714_),
    .Q(\mem.mem[176][3] ));
 sg13g2_dfrbp_1 _19877_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1914),
    .D(_01513_),
    .Q_N(_07713_),
    .Q(\mem.mem[176][4] ));
 sg13g2_dfrbp_1 _19878_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1913),
    .D(_01514_),
    .Q_N(_07712_),
    .Q(\mem.mem[176][5] ));
 sg13g2_dfrbp_1 _19879_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1912),
    .D(_01515_),
    .Q_N(_07711_),
    .Q(\mem.mem[176][6] ));
 sg13g2_dfrbp_1 _19880_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1911),
    .D(_01516_),
    .Q_N(_07710_),
    .Q(\mem.mem[176][7] ));
 sg13g2_dfrbp_1 _19881_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1910),
    .D(_01517_),
    .Q_N(_07709_),
    .Q(\mem.mem[177][0] ));
 sg13g2_dfrbp_1 _19882_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1909),
    .D(_01518_),
    .Q_N(_07708_),
    .Q(\mem.mem[177][1] ));
 sg13g2_dfrbp_1 _19883_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1908),
    .D(_01519_),
    .Q_N(_07707_),
    .Q(\mem.mem[177][2] ));
 sg13g2_dfrbp_1 _19884_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1907),
    .D(_01520_),
    .Q_N(_07706_),
    .Q(\mem.mem[177][3] ));
 sg13g2_dfrbp_1 _19885_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1906),
    .D(_01521_),
    .Q_N(_07705_),
    .Q(\mem.mem[177][4] ));
 sg13g2_dfrbp_1 _19886_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1905),
    .D(_01522_),
    .Q_N(_07704_),
    .Q(\mem.mem[177][5] ));
 sg13g2_dfrbp_1 _19887_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1904),
    .D(_01523_),
    .Q_N(_07703_),
    .Q(\mem.mem[177][6] ));
 sg13g2_dfrbp_1 _19888_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1903),
    .D(_01524_),
    .Q_N(_07702_),
    .Q(\mem.mem[177][7] ));
 sg13g2_dfrbp_1 _19889_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1902),
    .D(_01525_),
    .Q_N(_07701_),
    .Q(\mem.mem[178][0] ));
 sg13g2_dfrbp_1 _19890_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1901),
    .D(_01526_),
    .Q_N(_07700_),
    .Q(\mem.mem[178][1] ));
 sg13g2_dfrbp_1 _19891_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1900),
    .D(_01527_),
    .Q_N(_07699_),
    .Q(\mem.mem[178][2] ));
 sg13g2_dfrbp_1 _19892_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1899),
    .D(_01528_),
    .Q_N(_07698_),
    .Q(\mem.mem[178][3] ));
 sg13g2_dfrbp_1 _19893_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1898),
    .D(_01529_),
    .Q_N(_07697_),
    .Q(\mem.mem[178][4] ));
 sg13g2_dfrbp_1 _19894_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1897),
    .D(_01530_),
    .Q_N(_07696_),
    .Q(\mem.mem[178][5] ));
 sg13g2_dfrbp_1 _19895_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1896),
    .D(_01531_),
    .Q_N(_07695_),
    .Q(\mem.mem[178][6] ));
 sg13g2_dfrbp_1 _19896_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1895),
    .D(_01532_),
    .Q_N(_07694_),
    .Q(\mem.mem[178][7] ));
 sg13g2_dfrbp_1 _19897_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1894),
    .D(_01533_),
    .Q_N(_07693_),
    .Q(\mem.mem[17][0] ));
 sg13g2_dfrbp_1 _19898_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1893),
    .D(_01534_),
    .Q_N(_07692_),
    .Q(\mem.mem[17][1] ));
 sg13g2_dfrbp_1 _19899_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1892),
    .D(_01535_),
    .Q_N(_07691_),
    .Q(\mem.mem[17][2] ));
 sg13g2_dfrbp_1 _19900_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1891),
    .D(_01536_),
    .Q_N(_07690_),
    .Q(\mem.mem[17][3] ));
 sg13g2_dfrbp_1 _19901_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1890),
    .D(_01537_),
    .Q_N(_07689_),
    .Q(\mem.mem[17][4] ));
 sg13g2_dfrbp_1 _19902_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1889),
    .D(_01538_),
    .Q_N(_07688_),
    .Q(\mem.mem[17][5] ));
 sg13g2_dfrbp_1 _19903_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1888),
    .D(_01539_),
    .Q_N(_07687_),
    .Q(\mem.mem[17][6] ));
 sg13g2_dfrbp_1 _19904_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1887),
    .D(_01540_),
    .Q_N(_07686_),
    .Q(\mem.mem[17][7] ));
 sg13g2_dfrbp_1 _19905_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1886),
    .D(_01541_),
    .Q_N(_07685_),
    .Q(\mem.mem[180][0] ));
 sg13g2_dfrbp_1 _19906_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1885),
    .D(_01542_),
    .Q_N(_07684_),
    .Q(\mem.mem[180][1] ));
 sg13g2_dfrbp_1 _19907_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1884),
    .D(_01543_),
    .Q_N(_07683_),
    .Q(\mem.mem[180][2] ));
 sg13g2_dfrbp_1 _19908_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1883),
    .D(_01544_),
    .Q_N(_07682_),
    .Q(\mem.mem[180][3] ));
 sg13g2_dfrbp_1 _19909_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1882),
    .D(_01545_),
    .Q_N(_07681_),
    .Q(\mem.mem[180][4] ));
 sg13g2_dfrbp_1 _19910_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1881),
    .D(_01546_),
    .Q_N(_07680_),
    .Q(\mem.mem[180][5] ));
 sg13g2_dfrbp_1 _19911_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1880),
    .D(_01547_),
    .Q_N(_07679_),
    .Q(\mem.mem[180][6] ));
 sg13g2_dfrbp_1 _19912_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1879),
    .D(_01548_),
    .Q_N(_07678_),
    .Q(\mem.mem[180][7] ));
 sg13g2_dfrbp_1 _19913_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1878),
    .D(_01549_),
    .Q_N(_07677_),
    .Q(\mem.mem[181][0] ));
 sg13g2_dfrbp_1 _19914_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1877),
    .D(_01550_),
    .Q_N(_07676_),
    .Q(\mem.mem[181][1] ));
 sg13g2_dfrbp_1 _19915_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1876),
    .D(_01551_),
    .Q_N(_07675_),
    .Q(\mem.mem[181][2] ));
 sg13g2_dfrbp_1 _19916_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1875),
    .D(_01552_),
    .Q_N(_07674_),
    .Q(\mem.mem[181][3] ));
 sg13g2_dfrbp_1 _19917_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1874),
    .D(_01553_),
    .Q_N(_07673_),
    .Q(\mem.mem[181][4] ));
 sg13g2_dfrbp_1 _19918_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1873),
    .D(_01554_),
    .Q_N(_07672_),
    .Q(\mem.mem[181][5] ));
 sg13g2_dfrbp_1 _19919_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1872),
    .D(_01555_),
    .Q_N(_07671_),
    .Q(\mem.mem[181][6] ));
 sg13g2_dfrbp_1 _19920_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1871),
    .D(_01556_),
    .Q_N(_07670_),
    .Q(\mem.mem[181][7] ));
 sg13g2_dfrbp_1 _19921_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1870),
    .D(_01557_),
    .Q_N(_07669_),
    .Q(\mem.mem[182][0] ));
 sg13g2_dfrbp_1 _19922_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1869),
    .D(_01558_),
    .Q_N(_07668_),
    .Q(\mem.mem[182][1] ));
 sg13g2_dfrbp_1 _19923_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1868),
    .D(_01559_),
    .Q_N(_07667_),
    .Q(\mem.mem[182][2] ));
 sg13g2_dfrbp_1 _19924_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1867),
    .D(_01560_),
    .Q_N(_07666_),
    .Q(\mem.mem[182][3] ));
 sg13g2_dfrbp_1 _19925_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1866),
    .D(_01561_),
    .Q_N(_07665_),
    .Q(\mem.mem[182][4] ));
 sg13g2_dfrbp_1 _19926_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1865),
    .D(_01562_),
    .Q_N(_07664_),
    .Q(\mem.mem[182][5] ));
 sg13g2_dfrbp_1 _19927_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1864),
    .D(_01563_),
    .Q_N(_07663_),
    .Q(\mem.mem[182][6] ));
 sg13g2_dfrbp_1 _19928_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1863),
    .D(_01564_),
    .Q_N(_07662_),
    .Q(\mem.mem[182][7] ));
 sg13g2_dfrbp_1 _19929_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1862),
    .D(_01565_),
    .Q_N(_07661_),
    .Q(\mem.mem[183][0] ));
 sg13g2_dfrbp_1 _19930_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1861),
    .D(_01566_),
    .Q_N(_07660_),
    .Q(\mem.mem[183][1] ));
 sg13g2_dfrbp_1 _19931_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1860),
    .D(_01567_),
    .Q_N(_07659_),
    .Q(\mem.mem[183][2] ));
 sg13g2_dfrbp_1 _19932_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1859),
    .D(_01568_),
    .Q_N(_07658_),
    .Q(\mem.mem[183][3] ));
 sg13g2_dfrbp_1 _19933_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1858),
    .D(_01569_),
    .Q_N(_07657_),
    .Q(\mem.mem[183][4] ));
 sg13g2_dfrbp_1 _19934_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1857),
    .D(_01570_),
    .Q_N(_07656_),
    .Q(\mem.mem[183][5] ));
 sg13g2_dfrbp_1 _19935_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1856),
    .D(_01571_),
    .Q_N(_07655_),
    .Q(\mem.mem[183][6] ));
 sg13g2_dfrbp_1 _19936_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1855),
    .D(_01572_),
    .Q_N(_07654_),
    .Q(\mem.mem[183][7] ));
 sg13g2_dfrbp_1 _19937_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1854),
    .D(_01573_),
    .Q_N(_07653_),
    .Q(\mem.mem[184][0] ));
 sg13g2_dfrbp_1 _19938_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1853),
    .D(_01574_),
    .Q_N(_07652_),
    .Q(\mem.mem[184][1] ));
 sg13g2_dfrbp_1 _19939_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1852),
    .D(_01575_),
    .Q_N(_07651_),
    .Q(\mem.mem[184][2] ));
 sg13g2_dfrbp_1 _19940_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1851),
    .D(_01576_),
    .Q_N(_07650_),
    .Q(\mem.mem[184][3] ));
 sg13g2_dfrbp_1 _19941_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1850),
    .D(_01577_),
    .Q_N(_07649_),
    .Q(\mem.mem[184][4] ));
 sg13g2_dfrbp_1 _19942_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1849),
    .D(_01578_),
    .Q_N(_07648_),
    .Q(\mem.mem[184][5] ));
 sg13g2_dfrbp_1 _19943_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1848),
    .D(_01579_),
    .Q_N(_07647_),
    .Q(\mem.mem[184][6] ));
 sg13g2_dfrbp_1 _19944_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1847),
    .D(_01580_),
    .Q_N(_07646_),
    .Q(\mem.mem[184][7] ));
 sg13g2_dfrbp_1 _19945_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1846),
    .D(_01581_),
    .Q_N(_07645_),
    .Q(\mem.mem[185][0] ));
 sg13g2_dfrbp_1 _19946_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1845),
    .D(_01582_),
    .Q_N(_07644_),
    .Q(\mem.mem[185][1] ));
 sg13g2_dfrbp_1 _19947_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1844),
    .D(_01583_),
    .Q_N(_07643_),
    .Q(\mem.mem[185][2] ));
 sg13g2_dfrbp_1 _19948_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1843),
    .D(_01584_),
    .Q_N(_07642_),
    .Q(\mem.mem[185][3] ));
 sg13g2_dfrbp_1 _19949_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1842),
    .D(_01585_),
    .Q_N(_07641_),
    .Q(\mem.mem[185][4] ));
 sg13g2_dfrbp_1 _19950_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1841),
    .D(_01586_),
    .Q_N(_07640_),
    .Q(\mem.mem[185][5] ));
 sg13g2_dfrbp_1 _19951_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1840),
    .D(_01587_),
    .Q_N(_07639_),
    .Q(\mem.mem[185][6] ));
 sg13g2_dfrbp_1 _19952_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1839),
    .D(_01588_),
    .Q_N(_07638_),
    .Q(\mem.mem[185][7] ));
 sg13g2_dfrbp_1 _19953_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1838),
    .D(_01589_),
    .Q_N(_07637_),
    .Q(\mem.mem[186][0] ));
 sg13g2_dfrbp_1 _19954_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1837),
    .D(_01590_),
    .Q_N(_07636_),
    .Q(\mem.mem[186][1] ));
 sg13g2_dfrbp_1 _19955_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1836),
    .D(_01591_),
    .Q_N(_07635_),
    .Q(\mem.mem[186][2] ));
 sg13g2_dfrbp_1 _19956_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1835),
    .D(_01592_),
    .Q_N(_07634_),
    .Q(\mem.mem[186][3] ));
 sg13g2_dfrbp_1 _19957_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1834),
    .D(_01593_),
    .Q_N(_07633_),
    .Q(\mem.mem[186][4] ));
 sg13g2_dfrbp_1 _19958_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1833),
    .D(_01594_),
    .Q_N(_07632_),
    .Q(\mem.mem[186][5] ));
 sg13g2_dfrbp_1 _19959_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1832),
    .D(_01595_),
    .Q_N(_07631_),
    .Q(\mem.mem[186][6] ));
 sg13g2_dfrbp_1 _19960_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1831),
    .D(_01596_),
    .Q_N(_07630_),
    .Q(\mem.mem[186][7] ));
 sg13g2_dfrbp_1 _19961_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1830),
    .D(_01597_),
    .Q_N(_07629_),
    .Q(\mem.mem[187][0] ));
 sg13g2_dfrbp_1 _19962_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1829),
    .D(_01598_),
    .Q_N(_07628_),
    .Q(\mem.mem[187][1] ));
 sg13g2_dfrbp_1 _19963_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1828),
    .D(_01599_),
    .Q_N(_07627_),
    .Q(\mem.mem[187][2] ));
 sg13g2_dfrbp_1 _19964_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1827),
    .D(_01600_),
    .Q_N(_07626_),
    .Q(\mem.mem[187][3] ));
 sg13g2_dfrbp_1 _19965_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1826),
    .D(_01601_),
    .Q_N(_07625_),
    .Q(\mem.mem[187][4] ));
 sg13g2_dfrbp_1 _19966_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1825),
    .D(_01602_),
    .Q_N(_07624_),
    .Q(\mem.mem[187][5] ));
 sg13g2_dfrbp_1 _19967_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1824),
    .D(_01603_),
    .Q_N(_07623_),
    .Q(\mem.mem[187][6] ));
 sg13g2_dfrbp_1 _19968_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1823),
    .D(_01604_),
    .Q_N(_07622_),
    .Q(\mem.mem[187][7] ));
 sg13g2_dfrbp_1 _19969_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1822),
    .D(_01605_),
    .Q_N(_07621_),
    .Q(\mem.mem[188][0] ));
 sg13g2_dfrbp_1 _19970_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1821),
    .D(_01606_),
    .Q_N(_07620_),
    .Q(\mem.mem[188][1] ));
 sg13g2_dfrbp_1 _19971_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1820),
    .D(_01607_),
    .Q_N(_07619_),
    .Q(\mem.mem[188][2] ));
 sg13g2_dfrbp_1 _19972_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1819),
    .D(_01608_),
    .Q_N(_07618_),
    .Q(\mem.mem[188][3] ));
 sg13g2_dfrbp_1 _19973_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1818),
    .D(_01609_),
    .Q_N(_07617_),
    .Q(\mem.mem[188][4] ));
 sg13g2_dfrbp_1 _19974_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1817),
    .D(_01610_),
    .Q_N(_07616_),
    .Q(\mem.mem[188][5] ));
 sg13g2_dfrbp_1 _19975_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1816),
    .D(_01611_),
    .Q_N(_07615_),
    .Q(\mem.mem[188][6] ));
 sg13g2_dfrbp_1 _19976_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1815),
    .D(_01612_),
    .Q_N(_07614_),
    .Q(\mem.mem[188][7] ));
 sg13g2_dfrbp_1 _19977_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1814),
    .D(_01613_),
    .Q_N(_07613_),
    .Q(\mem.mem[18][0] ));
 sg13g2_dfrbp_1 _19978_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1813),
    .D(_01614_),
    .Q_N(_07612_),
    .Q(\mem.mem[18][1] ));
 sg13g2_dfrbp_1 _19979_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1812),
    .D(_01615_),
    .Q_N(_07611_),
    .Q(\mem.mem[18][2] ));
 sg13g2_dfrbp_1 _19980_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1811),
    .D(_01616_),
    .Q_N(_07610_),
    .Q(\mem.mem[18][3] ));
 sg13g2_dfrbp_1 _19981_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1810),
    .D(_01617_),
    .Q_N(_07609_),
    .Q(\mem.mem[18][4] ));
 sg13g2_dfrbp_1 _19982_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1809),
    .D(_01618_),
    .Q_N(_07608_),
    .Q(\mem.mem[18][5] ));
 sg13g2_dfrbp_1 _19983_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1808),
    .D(_01619_),
    .Q_N(_07607_),
    .Q(\mem.mem[18][6] ));
 sg13g2_dfrbp_1 _19984_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1807),
    .D(_01620_),
    .Q_N(_07606_),
    .Q(\mem.mem[18][7] ));
 sg13g2_dfrbp_1 _19985_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1806),
    .D(_01621_),
    .Q_N(_07605_),
    .Q(\mem.mem[190][0] ));
 sg13g2_dfrbp_1 _19986_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1805),
    .D(_01622_),
    .Q_N(_07604_),
    .Q(\mem.mem[190][1] ));
 sg13g2_dfrbp_1 _19987_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1804),
    .D(_01623_),
    .Q_N(_07603_),
    .Q(\mem.mem[190][2] ));
 sg13g2_dfrbp_1 _19988_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1803),
    .D(_01624_),
    .Q_N(_07602_),
    .Q(\mem.mem[190][3] ));
 sg13g2_dfrbp_1 _19989_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1802),
    .D(_01625_),
    .Q_N(_07601_),
    .Q(\mem.mem[190][4] ));
 sg13g2_dfrbp_1 _19990_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1801),
    .D(_01626_),
    .Q_N(_07600_),
    .Q(\mem.mem[190][5] ));
 sg13g2_dfrbp_1 _19991_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1800),
    .D(_01627_),
    .Q_N(_07599_),
    .Q(\mem.mem[190][6] ));
 sg13g2_dfrbp_1 _19992_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1799),
    .D(_01628_),
    .Q_N(_07598_),
    .Q(\mem.mem[190][7] ));
 sg13g2_dfrbp_1 _19993_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1798),
    .D(_01629_),
    .Q_N(_07597_),
    .Q(\mem.mem[191][0] ));
 sg13g2_dfrbp_1 _19994_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1797),
    .D(_01630_),
    .Q_N(_07596_),
    .Q(\mem.mem[191][1] ));
 sg13g2_dfrbp_1 _19995_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1796),
    .D(_01631_),
    .Q_N(_07595_),
    .Q(\mem.mem[191][2] ));
 sg13g2_dfrbp_1 _19996_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1795),
    .D(_01632_),
    .Q_N(_07594_),
    .Q(\mem.mem[191][3] ));
 sg13g2_dfrbp_1 _19997_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1794),
    .D(_01633_),
    .Q_N(_07593_),
    .Q(\mem.mem[191][4] ));
 sg13g2_dfrbp_1 _19998_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1793),
    .D(_01634_),
    .Q_N(_07592_),
    .Q(\mem.mem[191][5] ));
 sg13g2_dfrbp_1 _19999_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1792),
    .D(_01635_),
    .Q_N(_07591_),
    .Q(\mem.mem[191][6] ));
 sg13g2_dfrbp_1 _20000_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1791),
    .D(_01636_),
    .Q_N(_07590_),
    .Q(\mem.mem[191][7] ));
 sg13g2_dfrbp_1 _20001_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1790),
    .D(_01637_),
    .Q_N(_07589_),
    .Q(\mem.mem[192][0] ));
 sg13g2_dfrbp_1 _20002_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1789),
    .D(_01638_),
    .Q_N(_07588_),
    .Q(\mem.mem[192][1] ));
 sg13g2_dfrbp_1 _20003_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1788),
    .D(_01639_),
    .Q_N(_07587_),
    .Q(\mem.mem[192][2] ));
 sg13g2_dfrbp_1 _20004_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1787),
    .D(_01640_),
    .Q_N(_07586_),
    .Q(\mem.mem[192][3] ));
 sg13g2_dfrbp_1 _20005_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1786),
    .D(_01641_),
    .Q_N(_07585_),
    .Q(\mem.mem[192][4] ));
 sg13g2_dfrbp_1 _20006_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1785),
    .D(_01642_),
    .Q_N(_07584_),
    .Q(\mem.mem[192][5] ));
 sg13g2_dfrbp_1 _20007_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1784),
    .D(_01643_),
    .Q_N(_07583_),
    .Q(\mem.mem[192][6] ));
 sg13g2_dfrbp_1 _20008_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1783),
    .D(_01644_),
    .Q_N(_07582_),
    .Q(\mem.mem[192][7] ));
 sg13g2_dfrbp_1 _20009_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1782),
    .D(_01645_),
    .Q_N(_07581_),
    .Q(\mem.mem[193][0] ));
 sg13g2_dfrbp_1 _20010_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1781),
    .D(_01646_),
    .Q_N(_07580_),
    .Q(\mem.mem[193][1] ));
 sg13g2_dfrbp_1 _20011_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1780),
    .D(_01647_),
    .Q_N(_07579_),
    .Q(\mem.mem[193][2] ));
 sg13g2_dfrbp_1 _20012_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1779),
    .D(_01648_),
    .Q_N(_07578_),
    .Q(\mem.mem[193][3] ));
 sg13g2_dfrbp_1 _20013_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1778),
    .D(_01649_),
    .Q_N(_07577_),
    .Q(\mem.mem[193][4] ));
 sg13g2_dfrbp_1 _20014_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1777),
    .D(_01650_),
    .Q_N(_07576_),
    .Q(\mem.mem[193][5] ));
 sg13g2_dfrbp_1 _20015_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1776),
    .D(_01651_),
    .Q_N(_07575_),
    .Q(\mem.mem[193][6] ));
 sg13g2_dfrbp_1 _20016_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1775),
    .D(_01652_),
    .Q_N(_07574_),
    .Q(\mem.mem[193][7] ));
 sg13g2_dfrbp_1 _20017_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1774),
    .D(_01653_),
    .Q_N(_07573_),
    .Q(\mem.mem[194][0] ));
 sg13g2_dfrbp_1 _20018_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1773),
    .D(_01654_),
    .Q_N(_07572_),
    .Q(\mem.mem[194][1] ));
 sg13g2_dfrbp_1 _20019_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1772),
    .D(_01655_),
    .Q_N(_07571_),
    .Q(\mem.mem[194][2] ));
 sg13g2_dfrbp_1 _20020_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1771),
    .D(_01656_),
    .Q_N(_07570_),
    .Q(\mem.mem[194][3] ));
 sg13g2_dfrbp_1 _20021_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1770),
    .D(_01657_),
    .Q_N(_07569_),
    .Q(\mem.mem[194][4] ));
 sg13g2_dfrbp_1 _20022_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1769),
    .D(_01658_),
    .Q_N(_07568_),
    .Q(\mem.mem[194][5] ));
 sg13g2_dfrbp_1 _20023_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1768),
    .D(_01659_),
    .Q_N(_07567_),
    .Q(\mem.mem[194][6] ));
 sg13g2_dfrbp_1 _20024_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1767),
    .D(_01660_),
    .Q_N(_07566_),
    .Q(\mem.mem[194][7] ));
 sg13g2_dfrbp_1 _20025_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1766),
    .D(_01661_),
    .Q_N(_07565_),
    .Q(\mem.mem[195][0] ));
 sg13g2_dfrbp_1 _20026_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1765),
    .D(_01662_),
    .Q_N(_07564_),
    .Q(\mem.mem[195][1] ));
 sg13g2_dfrbp_1 _20027_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1764),
    .D(_01663_),
    .Q_N(_07563_),
    .Q(\mem.mem[195][2] ));
 sg13g2_dfrbp_1 _20028_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1763),
    .D(_01664_),
    .Q_N(_07562_),
    .Q(\mem.mem[195][3] ));
 sg13g2_dfrbp_1 _20029_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1762),
    .D(_01665_),
    .Q_N(_07561_),
    .Q(\mem.mem[195][4] ));
 sg13g2_dfrbp_1 _20030_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1761),
    .D(_01666_),
    .Q_N(_07560_),
    .Q(\mem.mem[195][5] ));
 sg13g2_dfrbp_1 _20031_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1760),
    .D(_01667_),
    .Q_N(_07559_),
    .Q(\mem.mem[195][6] ));
 sg13g2_dfrbp_1 _20032_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1759),
    .D(_01668_),
    .Q_N(_07558_),
    .Q(\mem.mem[195][7] ));
 sg13g2_dfrbp_1 _20033_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1758),
    .D(_01669_),
    .Q_N(_07557_),
    .Q(\mem.mem[196][0] ));
 sg13g2_dfrbp_1 _20034_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1757),
    .D(_01670_),
    .Q_N(_07556_),
    .Q(\mem.mem[196][1] ));
 sg13g2_dfrbp_1 _20035_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1756),
    .D(_01671_),
    .Q_N(_07555_),
    .Q(\mem.mem[196][2] ));
 sg13g2_dfrbp_1 _20036_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1755),
    .D(_01672_),
    .Q_N(_07554_),
    .Q(\mem.mem[196][3] ));
 sg13g2_dfrbp_1 _20037_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1754),
    .D(_01673_),
    .Q_N(_07553_),
    .Q(\mem.mem[196][4] ));
 sg13g2_dfrbp_1 _20038_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1753),
    .D(_01674_),
    .Q_N(_07552_),
    .Q(\mem.mem[196][5] ));
 sg13g2_dfrbp_1 _20039_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1752),
    .D(_01675_),
    .Q_N(_07551_),
    .Q(\mem.mem[196][6] ));
 sg13g2_dfrbp_1 _20040_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1751),
    .D(_01676_),
    .Q_N(_07550_),
    .Q(\mem.mem[196][7] ));
 sg13g2_dfrbp_1 _20041_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1750),
    .D(_01677_),
    .Q_N(_07549_),
    .Q(\mem.mem[197][0] ));
 sg13g2_dfrbp_1 _20042_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1749),
    .D(_01678_),
    .Q_N(_07548_),
    .Q(\mem.mem[197][1] ));
 sg13g2_dfrbp_1 _20043_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1748),
    .D(_01679_),
    .Q_N(_07547_),
    .Q(\mem.mem[197][2] ));
 sg13g2_dfrbp_1 _20044_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1747),
    .D(_01680_),
    .Q_N(_07546_),
    .Q(\mem.mem[197][3] ));
 sg13g2_dfrbp_1 _20045_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1746),
    .D(_01681_),
    .Q_N(_07545_),
    .Q(\mem.mem[197][4] ));
 sg13g2_dfrbp_1 _20046_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1745),
    .D(_01682_),
    .Q_N(_07544_),
    .Q(\mem.mem[197][5] ));
 sg13g2_dfrbp_1 _20047_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1744),
    .D(_01683_),
    .Q_N(_07543_),
    .Q(\mem.mem[197][6] ));
 sg13g2_dfrbp_1 _20048_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1743),
    .D(_01684_),
    .Q_N(_07542_),
    .Q(\mem.mem[197][7] ));
 sg13g2_dfrbp_1 _20049_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1742),
    .D(_01685_),
    .Q_N(_07541_),
    .Q(\mem.mem[198][0] ));
 sg13g2_dfrbp_1 _20050_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1741),
    .D(_01686_),
    .Q_N(_07540_),
    .Q(\mem.mem[198][1] ));
 sg13g2_dfrbp_1 _20051_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1740),
    .D(_01687_),
    .Q_N(_07539_),
    .Q(\mem.mem[198][2] ));
 sg13g2_dfrbp_1 _20052_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1739),
    .D(_01688_),
    .Q_N(_07538_),
    .Q(\mem.mem[198][3] ));
 sg13g2_dfrbp_1 _20053_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1738),
    .D(_01689_),
    .Q_N(_07537_),
    .Q(\mem.mem[198][4] ));
 sg13g2_dfrbp_1 _20054_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1737),
    .D(_01690_),
    .Q_N(_07536_),
    .Q(\mem.mem[198][5] ));
 sg13g2_dfrbp_1 _20055_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1736),
    .D(_01691_),
    .Q_N(_07535_),
    .Q(\mem.mem[198][6] ));
 sg13g2_dfrbp_1 _20056_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1735),
    .D(_01692_),
    .Q_N(_07534_),
    .Q(\mem.mem[198][7] ));
 sg13g2_dfrbp_1 _20057_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1734),
    .D(_01693_),
    .Q_N(_07533_),
    .Q(\mem.mem[1][0] ));
 sg13g2_dfrbp_1 _20058_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1733),
    .D(_01694_),
    .Q_N(_07532_),
    .Q(\mem.mem[1][1] ));
 sg13g2_dfrbp_1 _20059_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1732),
    .D(_01695_),
    .Q_N(_07531_),
    .Q(\mem.mem[1][2] ));
 sg13g2_dfrbp_1 _20060_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1731),
    .D(_01696_),
    .Q_N(_07530_),
    .Q(\mem.mem[1][3] ));
 sg13g2_dfrbp_1 _20061_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1730),
    .D(_01697_),
    .Q_N(_07529_),
    .Q(\mem.mem[1][4] ));
 sg13g2_dfrbp_1 _20062_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1729),
    .D(_01698_),
    .Q_N(_07528_),
    .Q(\mem.mem[1][5] ));
 sg13g2_dfrbp_1 _20063_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1728),
    .D(_01699_),
    .Q_N(_07527_),
    .Q(\mem.mem[1][6] ));
 sg13g2_dfrbp_1 _20064_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1727),
    .D(_01700_),
    .Q_N(_07526_),
    .Q(\mem.mem[1][7] ));
 sg13g2_dfrbp_1 _20065_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1726),
    .D(_01701_),
    .Q_N(_07525_),
    .Q(\mem.mem[200][0] ));
 sg13g2_dfrbp_1 _20066_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1725),
    .D(_01702_),
    .Q_N(_07524_),
    .Q(\mem.mem[200][1] ));
 sg13g2_dfrbp_1 _20067_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1724),
    .D(_01703_),
    .Q_N(_07523_),
    .Q(\mem.mem[200][2] ));
 sg13g2_dfrbp_1 _20068_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1723),
    .D(_01704_),
    .Q_N(_07522_),
    .Q(\mem.mem[200][3] ));
 sg13g2_dfrbp_1 _20069_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1722),
    .D(_01705_),
    .Q_N(_07521_),
    .Q(\mem.mem[200][4] ));
 sg13g2_dfrbp_1 _20070_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1721),
    .D(_01706_),
    .Q_N(_07520_),
    .Q(\mem.mem[200][5] ));
 sg13g2_dfrbp_1 _20071_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1720),
    .D(_01707_),
    .Q_N(_07519_),
    .Q(\mem.mem[200][6] ));
 sg13g2_dfrbp_1 _20072_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1719),
    .D(_01708_),
    .Q_N(_07518_),
    .Q(\mem.mem[200][7] ));
 sg13g2_dfrbp_1 _20073_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1718),
    .D(_01709_),
    .Q_N(_07517_),
    .Q(\mem.mem[201][0] ));
 sg13g2_dfrbp_1 _20074_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1717),
    .D(_01710_),
    .Q_N(_07516_),
    .Q(\mem.mem[201][1] ));
 sg13g2_dfrbp_1 _20075_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1716),
    .D(_01711_),
    .Q_N(_07515_),
    .Q(\mem.mem[201][2] ));
 sg13g2_dfrbp_1 _20076_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1715),
    .D(_01712_),
    .Q_N(_07514_),
    .Q(\mem.mem[201][3] ));
 sg13g2_dfrbp_1 _20077_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1714),
    .D(_01713_),
    .Q_N(_07513_),
    .Q(\mem.mem[201][4] ));
 sg13g2_dfrbp_1 _20078_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1713),
    .D(_01714_),
    .Q_N(_07512_),
    .Q(\mem.mem[201][5] ));
 sg13g2_dfrbp_1 _20079_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1712),
    .D(_01715_),
    .Q_N(_07511_),
    .Q(\mem.mem[201][6] ));
 sg13g2_dfrbp_1 _20080_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1711),
    .D(_01716_),
    .Q_N(_07510_),
    .Q(\mem.mem[201][7] ));
 sg13g2_dfrbp_1 _20081_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1710),
    .D(_01717_),
    .Q_N(_07509_),
    .Q(\mem.mem[202][0] ));
 sg13g2_dfrbp_1 _20082_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1709),
    .D(_01718_),
    .Q_N(_07508_),
    .Q(\mem.mem[202][1] ));
 sg13g2_dfrbp_1 _20083_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1708),
    .D(_01719_),
    .Q_N(_07507_),
    .Q(\mem.mem[202][2] ));
 sg13g2_dfrbp_1 _20084_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1707),
    .D(_01720_),
    .Q_N(_07506_),
    .Q(\mem.mem[202][3] ));
 sg13g2_dfrbp_1 _20085_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1706),
    .D(_01721_),
    .Q_N(_07505_),
    .Q(\mem.mem[202][4] ));
 sg13g2_dfrbp_1 _20086_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1705),
    .D(_01722_),
    .Q_N(_07504_),
    .Q(\mem.mem[202][5] ));
 sg13g2_dfrbp_1 _20087_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1704),
    .D(_01723_),
    .Q_N(_07503_),
    .Q(\mem.mem[202][6] ));
 sg13g2_dfrbp_1 _20088_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1703),
    .D(_01724_),
    .Q_N(_07502_),
    .Q(\mem.mem[202][7] ));
 sg13g2_dfrbp_1 _20089_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1702),
    .D(_01725_),
    .Q_N(_07501_),
    .Q(\mem.mem[203][0] ));
 sg13g2_dfrbp_1 _20090_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1701),
    .D(_01726_),
    .Q_N(_07500_),
    .Q(\mem.mem[203][1] ));
 sg13g2_dfrbp_1 _20091_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1700),
    .D(_01727_),
    .Q_N(_07499_),
    .Q(\mem.mem[203][2] ));
 sg13g2_dfrbp_1 _20092_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1699),
    .D(_01728_),
    .Q_N(_07498_),
    .Q(\mem.mem[203][3] ));
 sg13g2_dfrbp_1 _20093_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1698),
    .D(_01729_),
    .Q_N(_07497_),
    .Q(\mem.mem[203][4] ));
 sg13g2_dfrbp_1 _20094_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1697),
    .D(_01730_),
    .Q_N(_07496_),
    .Q(\mem.mem[203][5] ));
 sg13g2_dfrbp_1 _20095_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1696),
    .D(_01731_),
    .Q_N(_07495_),
    .Q(\mem.mem[203][6] ));
 sg13g2_dfrbp_1 _20096_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1695),
    .D(_01732_),
    .Q_N(_07494_),
    .Q(\mem.mem[203][7] ));
 sg13g2_dfrbp_1 _20097_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1694),
    .D(_01733_),
    .Q_N(_07493_),
    .Q(\mem.mem[204][0] ));
 sg13g2_dfrbp_1 _20098_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1693),
    .D(_01734_),
    .Q_N(_07492_),
    .Q(\mem.mem[204][1] ));
 sg13g2_dfrbp_1 _20099_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1692),
    .D(_01735_),
    .Q_N(_07491_),
    .Q(\mem.mem[204][2] ));
 sg13g2_dfrbp_1 _20100_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1691),
    .D(_01736_),
    .Q_N(_07490_),
    .Q(\mem.mem[204][3] ));
 sg13g2_dfrbp_1 _20101_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1690),
    .D(_01737_),
    .Q_N(_07489_),
    .Q(\mem.mem[204][4] ));
 sg13g2_dfrbp_1 _20102_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1689),
    .D(_01738_),
    .Q_N(_07488_),
    .Q(\mem.mem[204][5] ));
 sg13g2_dfrbp_1 _20103_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1688),
    .D(_01739_),
    .Q_N(_07487_),
    .Q(\mem.mem[204][6] ));
 sg13g2_dfrbp_1 _20104_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1687),
    .D(_01740_),
    .Q_N(_07486_),
    .Q(\mem.mem[204][7] ));
 sg13g2_dfrbp_1 _20105_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1686),
    .D(_01741_),
    .Q_N(_07485_),
    .Q(\mem.mem[205][0] ));
 sg13g2_dfrbp_1 _20106_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1685),
    .D(_01742_),
    .Q_N(_07484_),
    .Q(\mem.mem[205][1] ));
 sg13g2_dfrbp_1 _20107_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1684),
    .D(_01743_),
    .Q_N(_07483_),
    .Q(\mem.mem[205][2] ));
 sg13g2_dfrbp_1 _20108_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1683),
    .D(_01744_),
    .Q_N(_07482_),
    .Q(\mem.mem[205][3] ));
 sg13g2_dfrbp_1 _20109_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1682),
    .D(_01745_),
    .Q_N(_07481_),
    .Q(\mem.mem[205][4] ));
 sg13g2_dfrbp_1 _20110_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1681),
    .D(_01746_),
    .Q_N(_07480_),
    .Q(\mem.mem[205][5] ));
 sg13g2_dfrbp_1 _20111_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1680),
    .D(_01747_),
    .Q_N(_07479_),
    .Q(\mem.mem[205][6] ));
 sg13g2_dfrbp_1 _20112_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1679),
    .D(_01748_),
    .Q_N(_07478_),
    .Q(\mem.mem[205][7] ));
 sg13g2_dfrbp_1 _20113_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1678),
    .D(_01749_),
    .Q_N(_07477_),
    .Q(\mem.mem[206][0] ));
 sg13g2_dfrbp_1 _20114_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1677),
    .D(_01750_),
    .Q_N(_07476_),
    .Q(\mem.mem[206][1] ));
 sg13g2_dfrbp_1 _20115_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1676),
    .D(_01751_),
    .Q_N(_07475_),
    .Q(\mem.mem[206][2] ));
 sg13g2_dfrbp_1 _20116_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1675),
    .D(_01752_),
    .Q_N(_07474_),
    .Q(\mem.mem[206][3] ));
 sg13g2_dfrbp_1 _20117_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1674),
    .D(_01753_),
    .Q_N(_07473_),
    .Q(\mem.mem[206][4] ));
 sg13g2_dfrbp_1 _20118_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1673),
    .D(_01754_),
    .Q_N(_07472_),
    .Q(\mem.mem[206][5] ));
 sg13g2_dfrbp_1 _20119_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1672),
    .D(_01755_),
    .Q_N(_07471_),
    .Q(\mem.mem[206][6] ));
 sg13g2_dfrbp_1 _20120_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1671),
    .D(_01756_),
    .Q_N(_07470_),
    .Q(\mem.mem[206][7] ));
 sg13g2_dfrbp_1 _20121_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1670),
    .D(_01757_),
    .Q_N(_07469_),
    .Q(\mem.mem[207][0] ));
 sg13g2_dfrbp_1 _20122_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1669),
    .D(_01758_),
    .Q_N(_07468_),
    .Q(\mem.mem[207][1] ));
 sg13g2_dfrbp_1 _20123_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1668),
    .D(_01759_),
    .Q_N(_07467_),
    .Q(\mem.mem[207][2] ));
 sg13g2_dfrbp_1 _20124_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1667),
    .D(_01760_),
    .Q_N(_07466_),
    .Q(\mem.mem[207][3] ));
 sg13g2_dfrbp_1 _20125_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1666),
    .D(_01761_),
    .Q_N(_07465_),
    .Q(\mem.mem[207][4] ));
 sg13g2_dfrbp_1 _20126_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1665),
    .D(_01762_),
    .Q_N(_07464_),
    .Q(\mem.mem[207][5] ));
 sg13g2_dfrbp_1 _20127_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1664),
    .D(_01763_),
    .Q_N(_07463_),
    .Q(\mem.mem[207][6] ));
 sg13g2_dfrbp_1 _20128_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1663),
    .D(_01764_),
    .Q_N(_07462_),
    .Q(\mem.mem[207][7] ));
 sg13g2_dfrbp_1 _20129_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1662),
    .D(_01765_),
    .Q_N(_07461_),
    .Q(\mem.mem[208][0] ));
 sg13g2_dfrbp_1 _20130_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1661),
    .D(_01766_),
    .Q_N(_07460_),
    .Q(\mem.mem[208][1] ));
 sg13g2_dfrbp_1 _20131_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1660),
    .D(_01767_),
    .Q_N(_07459_),
    .Q(\mem.mem[208][2] ));
 sg13g2_dfrbp_1 _20132_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1659),
    .D(_01768_),
    .Q_N(_07458_),
    .Q(\mem.mem[208][3] ));
 sg13g2_dfrbp_1 _20133_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1658),
    .D(_01769_),
    .Q_N(_07457_),
    .Q(\mem.mem[208][4] ));
 sg13g2_dfrbp_1 _20134_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1657),
    .D(_01770_),
    .Q_N(_07456_),
    .Q(\mem.mem[208][5] ));
 sg13g2_dfrbp_1 _20135_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1656),
    .D(_01771_),
    .Q_N(_07455_),
    .Q(\mem.mem[208][6] ));
 sg13g2_dfrbp_1 _20136_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1655),
    .D(_01772_),
    .Q_N(_07454_),
    .Q(\mem.mem[208][7] ));
 sg13g2_dfrbp_1 _20137_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1654),
    .D(_01773_),
    .Q_N(_07453_),
    .Q(\mem.mem[20][0] ));
 sg13g2_dfrbp_1 _20138_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1653),
    .D(_01774_),
    .Q_N(_07452_),
    .Q(\mem.mem[20][1] ));
 sg13g2_dfrbp_1 _20139_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1652),
    .D(_01775_),
    .Q_N(_07451_),
    .Q(\mem.mem[20][2] ));
 sg13g2_dfrbp_1 _20140_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1651),
    .D(_01776_),
    .Q_N(_07450_),
    .Q(\mem.mem[20][3] ));
 sg13g2_dfrbp_1 _20141_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1650),
    .D(_01777_),
    .Q_N(_07449_),
    .Q(\mem.mem[20][4] ));
 sg13g2_dfrbp_1 _20142_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1649),
    .D(_01778_),
    .Q_N(_07448_),
    .Q(\mem.mem[20][5] ));
 sg13g2_dfrbp_1 _20143_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1648),
    .D(_01779_),
    .Q_N(_07447_),
    .Q(\mem.mem[20][6] ));
 sg13g2_dfrbp_1 _20144_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1647),
    .D(_01780_),
    .Q_N(_07446_),
    .Q(\mem.mem[20][7] ));
 sg13g2_dfrbp_1 _20145_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1646),
    .D(_01781_),
    .Q_N(_07445_),
    .Q(\mem.mem[210][0] ));
 sg13g2_dfrbp_1 _20146_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1645),
    .D(_01782_),
    .Q_N(_07444_),
    .Q(\mem.mem[210][1] ));
 sg13g2_dfrbp_1 _20147_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1644),
    .D(_01783_),
    .Q_N(_07443_),
    .Q(\mem.mem[210][2] ));
 sg13g2_dfrbp_1 _20148_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1643),
    .D(_01784_),
    .Q_N(_07442_),
    .Q(\mem.mem[210][3] ));
 sg13g2_dfrbp_1 _20149_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1642),
    .D(_01785_),
    .Q_N(_07441_),
    .Q(\mem.mem[210][4] ));
 sg13g2_dfrbp_1 _20150_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1641),
    .D(_01786_),
    .Q_N(_07440_),
    .Q(\mem.mem[210][5] ));
 sg13g2_dfrbp_1 _20151_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1640),
    .D(_01787_),
    .Q_N(_07439_),
    .Q(\mem.mem[210][6] ));
 sg13g2_dfrbp_1 _20152_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1639),
    .D(_01788_),
    .Q_N(_07438_),
    .Q(\mem.mem[210][7] ));
 sg13g2_dfrbp_1 _20153_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1638),
    .D(_01789_),
    .Q_N(_07437_),
    .Q(\mem.mem[211][0] ));
 sg13g2_dfrbp_1 _20154_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1637),
    .D(_01790_),
    .Q_N(_07436_),
    .Q(\mem.mem[211][1] ));
 sg13g2_dfrbp_1 _20155_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1636),
    .D(_01791_),
    .Q_N(_07435_),
    .Q(\mem.mem[211][2] ));
 sg13g2_dfrbp_1 _20156_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1635),
    .D(_01792_),
    .Q_N(_07434_),
    .Q(\mem.mem[211][3] ));
 sg13g2_dfrbp_1 _20157_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1634),
    .D(_01793_),
    .Q_N(_07433_),
    .Q(\mem.mem[211][4] ));
 sg13g2_dfrbp_1 _20158_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1633),
    .D(_01794_),
    .Q_N(_07432_),
    .Q(\mem.mem[211][5] ));
 sg13g2_dfrbp_1 _20159_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1632),
    .D(_01795_),
    .Q_N(_07431_),
    .Q(\mem.mem[211][6] ));
 sg13g2_dfrbp_1 _20160_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1631),
    .D(_01796_),
    .Q_N(_07430_),
    .Q(\mem.mem[211][7] ));
 sg13g2_dfrbp_1 _20161_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1630),
    .D(_01797_),
    .Q_N(_07429_),
    .Q(\mem.mem[212][0] ));
 sg13g2_dfrbp_1 _20162_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1629),
    .D(_01798_),
    .Q_N(_07428_),
    .Q(\mem.mem[212][1] ));
 sg13g2_dfrbp_1 _20163_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1628),
    .D(_01799_),
    .Q_N(_07427_),
    .Q(\mem.mem[212][2] ));
 sg13g2_dfrbp_1 _20164_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1627),
    .D(_01800_),
    .Q_N(_07426_),
    .Q(\mem.mem[212][3] ));
 sg13g2_dfrbp_1 _20165_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1626),
    .D(_01801_),
    .Q_N(_07425_),
    .Q(\mem.mem[212][4] ));
 sg13g2_dfrbp_1 _20166_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1625),
    .D(_01802_),
    .Q_N(_07424_),
    .Q(\mem.mem[212][5] ));
 sg13g2_dfrbp_1 _20167_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1624),
    .D(_01803_),
    .Q_N(_07423_),
    .Q(\mem.mem[212][6] ));
 sg13g2_dfrbp_1 _20168_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1623),
    .D(_01804_),
    .Q_N(_07422_),
    .Q(\mem.mem[212][7] ));
 sg13g2_dfrbp_1 _20169_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1622),
    .D(_01805_),
    .Q_N(_07421_),
    .Q(\mem.mem[213][0] ));
 sg13g2_dfrbp_1 _20170_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1621),
    .D(_01806_),
    .Q_N(_07420_),
    .Q(\mem.mem[213][1] ));
 sg13g2_dfrbp_1 _20171_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1620),
    .D(_01807_),
    .Q_N(_07419_),
    .Q(\mem.mem[213][2] ));
 sg13g2_dfrbp_1 _20172_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1619),
    .D(_01808_),
    .Q_N(_07418_),
    .Q(\mem.mem[213][3] ));
 sg13g2_dfrbp_1 _20173_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1618),
    .D(_01809_),
    .Q_N(_07417_),
    .Q(\mem.mem[213][4] ));
 sg13g2_dfrbp_1 _20174_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1617),
    .D(_01810_),
    .Q_N(_07416_),
    .Q(\mem.mem[213][5] ));
 sg13g2_dfrbp_1 _20175_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1616),
    .D(_01811_),
    .Q_N(_07415_),
    .Q(\mem.mem[213][6] ));
 sg13g2_dfrbp_1 _20176_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1615),
    .D(_01812_),
    .Q_N(_07414_),
    .Q(\mem.mem[213][7] ));
 sg13g2_dfrbp_1 _20177_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1614),
    .D(_01813_),
    .Q_N(_07413_),
    .Q(\mem.mem[214][0] ));
 sg13g2_dfrbp_1 _20178_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1613),
    .D(_01814_),
    .Q_N(_07412_),
    .Q(\mem.mem[214][1] ));
 sg13g2_dfrbp_1 _20179_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1612),
    .D(_01815_),
    .Q_N(_07411_),
    .Q(\mem.mem[214][2] ));
 sg13g2_dfrbp_1 _20180_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1611),
    .D(_01816_),
    .Q_N(_07410_),
    .Q(\mem.mem[214][3] ));
 sg13g2_dfrbp_1 _20181_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1610),
    .D(_01817_),
    .Q_N(_07409_),
    .Q(\mem.mem[214][4] ));
 sg13g2_dfrbp_1 _20182_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1609),
    .D(_01818_),
    .Q_N(_07408_),
    .Q(\mem.mem[214][5] ));
 sg13g2_dfrbp_1 _20183_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1608),
    .D(_01819_),
    .Q_N(_07407_),
    .Q(\mem.mem[214][6] ));
 sg13g2_dfrbp_1 _20184_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1607),
    .D(_01820_),
    .Q_N(_07406_),
    .Q(\mem.mem[214][7] ));
 sg13g2_dfrbp_1 _20185_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1606),
    .D(_01821_),
    .Q_N(_07405_),
    .Q(\mem.mem[215][0] ));
 sg13g2_dfrbp_1 _20186_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1605),
    .D(_01822_),
    .Q_N(_07404_),
    .Q(\mem.mem[215][1] ));
 sg13g2_dfrbp_1 _20187_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1604),
    .D(_01823_),
    .Q_N(_07403_),
    .Q(\mem.mem[215][2] ));
 sg13g2_dfrbp_1 _20188_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1603),
    .D(_01824_),
    .Q_N(_07402_),
    .Q(\mem.mem[215][3] ));
 sg13g2_dfrbp_1 _20189_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1602),
    .D(_01825_),
    .Q_N(_07401_),
    .Q(\mem.mem[215][4] ));
 sg13g2_dfrbp_1 _20190_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1601),
    .D(_01826_),
    .Q_N(_07400_),
    .Q(\mem.mem[215][5] ));
 sg13g2_dfrbp_1 _20191_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1600),
    .D(_01827_),
    .Q_N(_07399_),
    .Q(\mem.mem[215][6] ));
 sg13g2_dfrbp_1 _20192_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1599),
    .D(_01828_),
    .Q_N(_07398_),
    .Q(\mem.mem[215][7] ));
 sg13g2_dfrbp_1 _20193_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1598),
    .D(_01829_),
    .Q_N(_07397_),
    .Q(\mem.mem[216][0] ));
 sg13g2_dfrbp_1 _20194_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1597),
    .D(_01830_),
    .Q_N(_07396_),
    .Q(\mem.mem[216][1] ));
 sg13g2_dfrbp_1 _20195_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1596),
    .D(_01831_),
    .Q_N(_07395_),
    .Q(\mem.mem[216][2] ));
 sg13g2_dfrbp_1 _20196_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1595),
    .D(_01832_),
    .Q_N(_07394_),
    .Q(\mem.mem[216][3] ));
 sg13g2_dfrbp_1 _20197_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1594),
    .D(_01833_),
    .Q_N(_07393_),
    .Q(\mem.mem[216][4] ));
 sg13g2_dfrbp_1 _20198_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1593),
    .D(_01834_),
    .Q_N(_07392_),
    .Q(\mem.mem[216][5] ));
 sg13g2_dfrbp_1 _20199_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1592),
    .D(_01835_),
    .Q_N(_07391_),
    .Q(\mem.mem[216][6] ));
 sg13g2_dfrbp_1 _20200_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1591),
    .D(_01836_),
    .Q_N(_07390_),
    .Q(\mem.mem[216][7] ));
 sg13g2_dfrbp_1 _20201_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1590),
    .D(_01837_),
    .Q_N(_07389_),
    .Q(\mem.mem[217][0] ));
 sg13g2_dfrbp_1 _20202_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1589),
    .D(_01838_),
    .Q_N(_07388_),
    .Q(\mem.mem[217][1] ));
 sg13g2_dfrbp_1 _20203_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1588),
    .D(_01839_),
    .Q_N(_07387_),
    .Q(\mem.mem[217][2] ));
 sg13g2_dfrbp_1 _20204_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1587),
    .D(_01840_),
    .Q_N(_07386_),
    .Q(\mem.mem[217][3] ));
 sg13g2_dfrbp_1 _20205_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1586),
    .D(_01841_),
    .Q_N(_07385_),
    .Q(\mem.mem[217][4] ));
 sg13g2_dfrbp_1 _20206_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1585),
    .D(_01842_),
    .Q_N(_07384_),
    .Q(\mem.mem[217][5] ));
 sg13g2_dfrbp_1 _20207_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1584),
    .D(_01843_),
    .Q_N(_07383_),
    .Q(\mem.mem[217][6] ));
 sg13g2_dfrbp_1 _20208_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1583),
    .D(_01844_),
    .Q_N(_07382_),
    .Q(\mem.mem[217][7] ));
 sg13g2_dfrbp_1 _20209_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1582),
    .D(_01845_),
    .Q_N(_07381_),
    .Q(\mem.mem[218][0] ));
 sg13g2_dfrbp_1 _20210_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1581),
    .D(_01846_),
    .Q_N(_07380_),
    .Q(\mem.mem[218][1] ));
 sg13g2_dfrbp_1 _20211_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1580),
    .D(_01847_),
    .Q_N(_07379_),
    .Q(\mem.mem[218][2] ));
 sg13g2_dfrbp_1 _20212_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1579),
    .D(_01848_),
    .Q_N(_07378_),
    .Q(\mem.mem[218][3] ));
 sg13g2_dfrbp_1 _20213_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1578),
    .D(_01849_),
    .Q_N(_07377_),
    .Q(\mem.mem[218][4] ));
 sg13g2_dfrbp_1 _20214_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1577),
    .D(_01850_),
    .Q_N(_07376_),
    .Q(\mem.mem[218][5] ));
 sg13g2_dfrbp_1 _20215_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1576),
    .D(_01851_),
    .Q_N(_07375_),
    .Q(\mem.mem[218][6] ));
 sg13g2_dfrbp_1 _20216_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1575),
    .D(_01852_),
    .Q_N(_07374_),
    .Q(\mem.mem[218][7] ));
 sg13g2_dfrbp_1 _20217_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1574),
    .D(_01853_),
    .Q_N(_07373_),
    .Q(\mem.mem[21][0] ));
 sg13g2_dfrbp_1 _20218_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1573),
    .D(_01854_),
    .Q_N(_07372_),
    .Q(\mem.mem[21][1] ));
 sg13g2_dfrbp_1 _20219_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1572),
    .D(_01855_),
    .Q_N(_07371_),
    .Q(\mem.mem[21][2] ));
 sg13g2_dfrbp_1 _20220_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1571),
    .D(_01856_),
    .Q_N(_07370_),
    .Q(\mem.mem[21][3] ));
 sg13g2_dfrbp_1 _20221_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1570),
    .D(_01857_),
    .Q_N(_07369_),
    .Q(\mem.mem[21][4] ));
 sg13g2_dfrbp_1 _20222_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1569),
    .D(_01858_),
    .Q_N(_07368_),
    .Q(\mem.mem[21][5] ));
 sg13g2_dfrbp_1 _20223_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1568),
    .D(_01859_),
    .Q_N(_07367_),
    .Q(\mem.mem[21][6] ));
 sg13g2_dfrbp_1 _20224_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1567),
    .D(_01860_),
    .Q_N(_07366_),
    .Q(\mem.mem[21][7] ));
 sg13g2_dfrbp_1 _20225_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1566),
    .D(_01861_),
    .Q_N(_07365_),
    .Q(\mem.mem[220][0] ));
 sg13g2_dfrbp_1 _20226_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1565),
    .D(_01862_),
    .Q_N(_07364_),
    .Q(\mem.mem[220][1] ));
 sg13g2_dfrbp_1 _20227_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1564),
    .D(_01863_),
    .Q_N(_07363_),
    .Q(\mem.mem[220][2] ));
 sg13g2_dfrbp_1 _20228_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1563),
    .D(_01864_),
    .Q_N(_07362_),
    .Q(\mem.mem[220][3] ));
 sg13g2_dfrbp_1 _20229_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1562),
    .D(_01865_),
    .Q_N(_07361_),
    .Q(\mem.mem[220][4] ));
 sg13g2_dfrbp_1 _20230_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1561),
    .D(_01866_),
    .Q_N(_07360_),
    .Q(\mem.mem[220][5] ));
 sg13g2_dfrbp_1 _20231_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1560),
    .D(_01867_),
    .Q_N(_07359_),
    .Q(\mem.mem[220][6] ));
 sg13g2_dfrbp_1 _20232_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1559),
    .D(_01868_),
    .Q_N(_07358_),
    .Q(\mem.mem[220][7] ));
 sg13g2_dfrbp_1 _20233_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1558),
    .D(_01869_),
    .Q_N(_07357_),
    .Q(\mem.mem[221][0] ));
 sg13g2_dfrbp_1 _20234_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1557),
    .D(_01870_),
    .Q_N(_07356_),
    .Q(\mem.mem[221][1] ));
 sg13g2_dfrbp_1 _20235_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1556),
    .D(_01871_),
    .Q_N(_07355_),
    .Q(\mem.mem[221][2] ));
 sg13g2_dfrbp_1 _20236_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1555),
    .D(_01872_),
    .Q_N(_07354_),
    .Q(\mem.mem[221][3] ));
 sg13g2_dfrbp_1 _20237_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1554),
    .D(_01873_),
    .Q_N(_07353_),
    .Q(\mem.mem[221][4] ));
 sg13g2_dfrbp_1 _20238_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1553),
    .D(_01874_),
    .Q_N(_07352_),
    .Q(\mem.mem[221][5] ));
 sg13g2_dfrbp_1 _20239_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1552),
    .D(_01875_),
    .Q_N(_07351_),
    .Q(\mem.mem[221][6] ));
 sg13g2_dfrbp_1 _20240_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1551),
    .D(_01876_),
    .Q_N(_07350_),
    .Q(\mem.mem[221][7] ));
 sg13g2_dfrbp_1 _20241_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1550),
    .D(_01877_),
    .Q_N(_07349_),
    .Q(\mem.mem[222][0] ));
 sg13g2_dfrbp_1 _20242_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1549),
    .D(_01878_),
    .Q_N(_07348_),
    .Q(\mem.mem[222][1] ));
 sg13g2_dfrbp_1 _20243_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1548),
    .D(_01879_),
    .Q_N(_07347_),
    .Q(\mem.mem[222][2] ));
 sg13g2_dfrbp_1 _20244_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1547),
    .D(_01880_),
    .Q_N(_07346_),
    .Q(\mem.mem[222][3] ));
 sg13g2_dfrbp_1 _20245_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1546),
    .D(_01881_),
    .Q_N(_07345_),
    .Q(\mem.mem[222][4] ));
 sg13g2_dfrbp_1 _20246_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1545),
    .D(_01882_),
    .Q_N(_07344_),
    .Q(\mem.mem[222][5] ));
 sg13g2_dfrbp_1 _20247_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1544),
    .D(_01883_),
    .Q_N(_07343_),
    .Q(\mem.mem[222][6] ));
 sg13g2_dfrbp_1 _20248_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1543),
    .D(_01884_),
    .Q_N(_07342_),
    .Q(\mem.mem[222][7] ));
 sg13g2_dfrbp_1 _20249_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1542),
    .D(_01885_),
    .Q_N(_07341_),
    .Q(\mem.mem[223][0] ));
 sg13g2_dfrbp_1 _20250_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1541),
    .D(_01886_),
    .Q_N(_07340_),
    .Q(\mem.mem[223][1] ));
 sg13g2_dfrbp_1 _20251_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1540),
    .D(_01887_),
    .Q_N(_07339_),
    .Q(\mem.mem[223][2] ));
 sg13g2_dfrbp_1 _20252_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1539),
    .D(_01888_),
    .Q_N(_07338_),
    .Q(\mem.mem[223][3] ));
 sg13g2_dfrbp_1 _20253_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1538),
    .D(_01889_),
    .Q_N(_07337_),
    .Q(\mem.mem[223][4] ));
 sg13g2_dfrbp_1 _20254_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1537),
    .D(_01890_),
    .Q_N(_07336_),
    .Q(\mem.mem[223][5] ));
 sg13g2_dfrbp_1 _20255_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1536),
    .D(_01891_),
    .Q_N(_07335_),
    .Q(\mem.mem[223][6] ));
 sg13g2_dfrbp_1 _20256_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1535),
    .D(_01892_),
    .Q_N(_07334_),
    .Q(\mem.mem[223][7] ));
 sg13g2_dfrbp_1 _20257_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1534),
    .D(_01893_),
    .Q_N(_07333_),
    .Q(\mem.mem[224][0] ));
 sg13g2_dfrbp_1 _20258_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1533),
    .D(_01894_),
    .Q_N(_07332_),
    .Q(\mem.mem[224][1] ));
 sg13g2_dfrbp_1 _20259_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1532),
    .D(_01895_),
    .Q_N(_07331_),
    .Q(\mem.mem[224][2] ));
 sg13g2_dfrbp_1 _20260_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1531),
    .D(_01896_),
    .Q_N(_07330_),
    .Q(\mem.mem[224][3] ));
 sg13g2_dfrbp_1 _20261_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1530),
    .D(_01897_),
    .Q_N(_07329_),
    .Q(\mem.mem[224][4] ));
 sg13g2_dfrbp_1 _20262_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1529),
    .D(_01898_),
    .Q_N(_07328_),
    .Q(\mem.mem[224][5] ));
 sg13g2_dfrbp_1 _20263_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1528),
    .D(_01899_),
    .Q_N(_07327_),
    .Q(\mem.mem[224][6] ));
 sg13g2_dfrbp_1 _20264_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1527),
    .D(_01900_),
    .Q_N(_07326_),
    .Q(\mem.mem[224][7] ));
 sg13g2_dfrbp_1 _20265_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1526),
    .D(_01901_),
    .Q_N(_07325_),
    .Q(\mem.mem[225][0] ));
 sg13g2_dfrbp_1 _20266_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1525),
    .D(_01902_),
    .Q_N(_07324_),
    .Q(\mem.mem[225][1] ));
 sg13g2_dfrbp_1 _20267_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1524),
    .D(_01903_),
    .Q_N(_07323_),
    .Q(\mem.mem[225][2] ));
 sg13g2_dfrbp_1 _20268_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1523),
    .D(_01904_),
    .Q_N(_07322_),
    .Q(\mem.mem[225][3] ));
 sg13g2_dfrbp_1 _20269_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1522),
    .D(_01905_),
    .Q_N(_07321_),
    .Q(\mem.mem[225][4] ));
 sg13g2_dfrbp_1 _20270_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1521),
    .D(_01906_),
    .Q_N(_07320_),
    .Q(\mem.mem[225][5] ));
 sg13g2_dfrbp_1 _20271_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1520),
    .D(_01907_),
    .Q_N(_07319_),
    .Q(\mem.mem[225][6] ));
 sg13g2_dfrbp_1 _20272_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1519),
    .D(_01908_),
    .Q_N(_07318_),
    .Q(\mem.mem[225][7] ));
 sg13g2_dfrbp_1 _20273_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1518),
    .D(_01909_),
    .Q_N(_07317_),
    .Q(\mem.mem[226][0] ));
 sg13g2_dfrbp_1 _20274_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1517),
    .D(_01910_),
    .Q_N(_07316_),
    .Q(\mem.mem[226][1] ));
 sg13g2_dfrbp_1 _20275_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1516),
    .D(_01911_),
    .Q_N(_07315_),
    .Q(\mem.mem[226][2] ));
 sg13g2_dfrbp_1 _20276_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1515),
    .D(_01912_),
    .Q_N(_07314_),
    .Q(\mem.mem[226][3] ));
 sg13g2_dfrbp_1 _20277_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1514),
    .D(_01913_),
    .Q_N(_07313_),
    .Q(\mem.mem[226][4] ));
 sg13g2_dfrbp_1 _20278_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1513),
    .D(_01914_),
    .Q_N(_07312_),
    .Q(\mem.mem[226][5] ));
 sg13g2_dfrbp_1 _20279_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1512),
    .D(_01915_),
    .Q_N(_07311_),
    .Q(\mem.mem[226][6] ));
 sg13g2_dfrbp_1 _20280_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1511),
    .D(_01916_),
    .Q_N(_07310_),
    .Q(\mem.mem[226][7] ));
 sg13g2_dfrbp_1 _20281_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1510),
    .D(_01917_),
    .Q_N(_07309_),
    .Q(\mem.mem[227][0] ));
 sg13g2_dfrbp_1 _20282_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1509),
    .D(_01918_),
    .Q_N(_07308_),
    .Q(\mem.mem[227][1] ));
 sg13g2_dfrbp_1 _20283_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1508),
    .D(_01919_),
    .Q_N(_07307_),
    .Q(\mem.mem[227][2] ));
 sg13g2_dfrbp_1 _20284_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1507),
    .D(_01920_),
    .Q_N(_07306_),
    .Q(\mem.mem[227][3] ));
 sg13g2_dfrbp_1 _20285_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1506),
    .D(_01921_),
    .Q_N(_07305_),
    .Q(\mem.mem[227][4] ));
 sg13g2_dfrbp_1 _20286_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1505),
    .D(_01922_),
    .Q_N(_07304_),
    .Q(\mem.mem[227][5] ));
 sg13g2_dfrbp_1 _20287_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1504),
    .D(_01923_),
    .Q_N(_07303_),
    .Q(\mem.mem[227][6] ));
 sg13g2_dfrbp_1 _20288_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1503),
    .D(_01924_),
    .Q_N(_07302_),
    .Q(\mem.mem[227][7] ));
 sg13g2_dfrbp_1 _20289_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1502),
    .D(_01925_),
    .Q_N(_07301_),
    .Q(\mem.mem[228][0] ));
 sg13g2_dfrbp_1 _20290_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1501),
    .D(_01926_),
    .Q_N(_07300_),
    .Q(\mem.mem[228][1] ));
 sg13g2_dfrbp_1 _20291_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1500),
    .D(_01927_),
    .Q_N(_07299_),
    .Q(\mem.mem[228][2] ));
 sg13g2_dfrbp_1 _20292_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1499),
    .D(_01928_),
    .Q_N(_07298_),
    .Q(\mem.mem[228][3] ));
 sg13g2_dfrbp_1 _20293_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1498),
    .D(_01929_),
    .Q_N(_07297_),
    .Q(\mem.mem[228][4] ));
 sg13g2_dfrbp_1 _20294_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1497),
    .D(_01930_),
    .Q_N(_07296_),
    .Q(\mem.mem[228][5] ));
 sg13g2_dfrbp_1 _20295_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1496),
    .D(_01931_),
    .Q_N(_07295_),
    .Q(\mem.mem[228][6] ));
 sg13g2_dfrbp_1 _20296_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1495),
    .D(_01932_),
    .Q_N(_07294_),
    .Q(\mem.mem[228][7] ));
 sg13g2_dfrbp_1 _20297_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1494),
    .D(_01933_),
    .Q_N(_07293_),
    .Q(\mem.mem[22][0] ));
 sg13g2_dfrbp_1 _20298_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1493),
    .D(_01934_),
    .Q_N(_07292_),
    .Q(\mem.mem[22][1] ));
 sg13g2_dfrbp_1 _20299_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1492),
    .D(_01935_),
    .Q_N(_07291_),
    .Q(\mem.mem[22][2] ));
 sg13g2_dfrbp_1 _20300_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1491),
    .D(_01936_),
    .Q_N(_07290_),
    .Q(\mem.mem[22][3] ));
 sg13g2_dfrbp_1 _20301_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1490),
    .D(_01937_),
    .Q_N(_07289_),
    .Q(\mem.mem[22][4] ));
 sg13g2_dfrbp_1 _20302_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1489),
    .D(_01938_),
    .Q_N(_07288_),
    .Q(\mem.mem[22][5] ));
 sg13g2_dfrbp_1 _20303_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1488),
    .D(_01939_),
    .Q_N(_07287_),
    .Q(\mem.mem[22][6] ));
 sg13g2_dfrbp_1 _20304_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1487),
    .D(_01940_),
    .Q_N(_07286_),
    .Q(\mem.mem[22][7] ));
 sg13g2_dfrbp_1 _20305_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1486),
    .D(_01941_),
    .Q_N(_07285_),
    .Q(\mem.mem[230][0] ));
 sg13g2_dfrbp_1 _20306_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1485),
    .D(_01942_),
    .Q_N(_07284_),
    .Q(\mem.mem[230][1] ));
 sg13g2_dfrbp_1 _20307_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1484),
    .D(_01943_),
    .Q_N(_07283_),
    .Q(\mem.mem[230][2] ));
 sg13g2_dfrbp_1 _20308_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1483),
    .D(_01944_),
    .Q_N(_07282_),
    .Q(\mem.mem[230][3] ));
 sg13g2_dfrbp_1 _20309_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1482),
    .D(_01945_),
    .Q_N(_07281_),
    .Q(\mem.mem[230][4] ));
 sg13g2_dfrbp_1 _20310_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1481),
    .D(_01946_),
    .Q_N(_07280_),
    .Q(\mem.mem[230][5] ));
 sg13g2_dfrbp_1 _20311_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1480),
    .D(_01947_),
    .Q_N(_07279_),
    .Q(\mem.mem[230][6] ));
 sg13g2_dfrbp_1 _20312_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1479),
    .D(_01948_),
    .Q_N(_07278_),
    .Q(\mem.mem[230][7] ));
 sg13g2_dfrbp_1 _20313_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1478),
    .D(_01949_),
    .Q_N(_07277_),
    .Q(\mem.mem[231][0] ));
 sg13g2_dfrbp_1 _20314_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1477),
    .D(_01950_),
    .Q_N(_07276_),
    .Q(\mem.mem[231][1] ));
 sg13g2_dfrbp_1 _20315_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1476),
    .D(_01951_),
    .Q_N(_07275_),
    .Q(\mem.mem[231][2] ));
 sg13g2_dfrbp_1 _20316_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1475),
    .D(_01952_),
    .Q_N(_07274_),
    .Q(\mem.mem[231][3] ));
 sg13g2_dfrbp_1 _20317_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1474),
    .D(_01953_),
    .Q_N(_07273_),
    .Q(\mem.mem[231][4] ));
 sg13g2_dfrbp_1 _20318_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1473),
    .D(_01954_),
    .Q_N(_07272_),
    .Q(\mem.mem[231][5] ));
 sg13g2_dfrbp_1 _20319_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1472),
    .D(_01955_),
    .Q_N(_07271_),
    .Q(\mem.mem[231][6] ));
 sg13g2_dfrbp_1 _20320_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1471),
    .D(_01956_),
    .Q_N(_07270_),
    .Q(\mem.mem[231][7] ));
 sg13g2_dfrbp_1 _20321_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1470),
    .D(_01957_),
    .Q_N(_07269_),
    .Q(\mem.mem[232][0] ));
 sg13g2_dfrbp_1 _20322_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1469),
    .D(_01958_),
    .Q_N(_07268_),
    .Q(\mem.mem[232][1] ));
 sg13g2_dfrbp_1 _20323_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1468),
    .D(_01959_),
    .Q_N(_07267_),
    .Q(\mem.mem[232][2] ));
 sg13g2_dfrbp_1 _20324_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1467),
    .D(_01960_),
    .Q_N(_07266_),
    .Q(\mem.mem[232][3] ));
 sg13g2_dfrbp_1 _20325_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1466),
    .D(_01961_),
    .Q_N(_07265_),
    .Q(\mem.mem[232][4] ));
 sg13g2_dfrbp_1 _20326_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1465),
    .D(_01962_),
    .Q_N(_07264_),
    .Q(\mem.mem[232][5] ));
 sg13g2_dfrbp_1 _20327_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1464),
    .D(_01963_),
    .Q_N(_07263_),
    .Q(\mem.mem[232][6] ));
 sg13g2_dfrbp_1 _20328_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1463),
    .D(_01964_),
    .Q_N(_07262_),
    .Q(\mem.mem[232][7] ));
 sg13g2_dfrbp_1 _20329_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1462),
    .D(_01965_),
    .Q_N(_07261_),
    .Q(\mem.mem[233][0] ));
 sg13g2_dfrbp_1 _20330_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1461),
    .D(_01966_),
    .Q_N(_07260_),
    .Q(\mem.mem[233][1] ));
 sg13g2_dfrbp_1 _20331_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1460),
    .D(_01967_),
    .Q_N(_07259_),
    .Q(\mem.mem[233][2] ));
 sg13g2_dfrbp_1 _20332_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1459),
    .D(_01968_),
    .Q_N(_07258_),
    .Q(\mem.mem[233][3] ));
 sg13g2_dfrbp_1 _20333_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1458),
    .D(_01969_),
    .Q_N(_07257_),
    .Q(\mem.mem[233][4] ));
 sg13g2_dfrbp_1 _20334_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1457),
    .D(_01970_),
    .Q_N(_07256_),
    .Q(\mem.mem[233][5] ));
 sg13g2_dfrbp_1 _20335_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1456),
    .D(_01971_),
    .Q_N(_07255_),
    .Q(\mem.mem[233][6] ));
 sg13g2_dfrbp_1 _20336_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1455),
    .D(_01972_),
    .Q_N(_07254_),
    .Q(\mem.mem[233][7] ));
 sg13g2_dfrbp_1 _20337_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1454),
    .D(_01973_),
    .Q_N(_07253_),
    .Q(\mem.mem[234][0] ));
 sg13g2_dfrbp_1 _20338_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1453),
    .D(_01974_),
    .Q_N(_07252_),
    .Q(\mem.mem[234][1] ));
 sg13g2_dfrbp_1 _20339_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1452),
    .D(_01975_),
    .Q_N(_07251_),
    .Q(\mem.mem[234][2] ));
 sg13g2_dfrbp_1 _20340_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1451),
    .D(_01976_),
    .Q_N(_07250_),
    .Q(\mem.mem[234][3] ));
 sg13g2_dfrbp_1 _20341_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1450),
    .D(_01977_),
    .Q_N(_07249_),
    .Q(\mem.mem[234][4] ));
 sg13g2_dfrbp_1 _20342_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1449),
    .D(_01978_),
    .Q_N(_07248_),
    .Q(\mem.mem[234][5] ));
 sg13g2_dfrbp_1 _20343_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1448),
    .D(_01979_),
    .Q_N(_07247_),
    .Q(\mem.mem[234][6] ));
 sg13g2_dfrbp_1 _20344_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1447),
    .D(_01980_),
    .Q_N(_07246_),
    .Q(\mem.mem[234][7] ));
 sg13g2_dfrbp_1 _20345_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1446),
    .D(_01981_),
    .Q_N(_07245_),
    .Q(\mem.mem[235][0] ));
 sg13g2_dfrbp_1 _20346_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1445),
    .D(_01982_),
    .Q_N(_07244_),
    .Q(\mem.mem[235][1] ));
 sg13g2_dfrbp_1 _20347_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1444),
    .D(_01983_),
    .Q_N(_07243_),
    .Q(\mem.mem[235][2] ));
 sg13g2_dfrbp_1 _20348_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1443),
    .D(_01984_),
    .Q_N(_07242_),
    .Q(\mem.mem[235][3] ));
 sg13g2_dfrbp_1 _20349_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1442),
    .D(_01985_),
    .Q_N(_07241_),
    .Q(\mem.mem[235][4] ));
 sg13g2_dfrbp_1 _20350_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1441),
    .D(_01986_),
    .Q_N(_07240_),
    .Q(\mem.mem[235][5] ));
 sg13g2_dfrbp_1 _20351_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1440),
    .D(_01987_),
    .Q_N(_07239_),
    .Q(\mem.mem[235][6] ));
 sg13g2_dfrbp_1 _20352_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1439),
    .D(_01988_),
    .Q_N(_07238_),
    .Q(\mem.mem[235][7] ));
 sg13g2_dfrbp_1 _20353_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1438),
    .D(_01989_),
    .Q_N(_07237_),
    .Q(\mem.mem[236][0] ));
 sg13g2_dfrbp_1 _20354_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1437),
    .D(_01990_),
    .Q_N(_07236_),
    .Q(\mem.mem[236][1] ));
 sg13g2_dfrbp_1 _20355_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1436),
    .D(_01991_),
    .Q_N(_07235_),
    .Q(\mem.mem[236][2] ));
 sg13g2_dfrbp_1 _20356_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1435),
    .D(_01992_),
    .Q_N(_07234_),
    .Q(\mem.mem[236][3] ));
 sg13g2_dfrbp_1 _20357_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1434),
    .D(_01993_),
    .Q_N(_07233_),
    .Q(\mem.mem[236][4] ));
 sg13g2_dfrbp_1 _20358_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1433),
    .D(_01994_),
    .Q_N(_07232_),
    .Q(\mem.mem[236][5] ));
 sg13g2_dfrbp_1 _20359_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1432),
    .D(_01995_),
    .Q_N(_07231_),
    .Q(\mem.mem[236][6] ));
 sg13g2_dfrbp_1 _20360_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1431),
    .D(_01996_),
    .Q_N(_07230_),
    .Q(\mem.mem[236][7] ));
 sg13g2_dfrbp_1 _20361_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1430),
    .D(_01997_),
    .Q_N(_07229_),
    .Q(\mem.mem[237][0] ));
 sg13g2_dfrbp_1 _20362_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1429),
    .D(_01998_),
    .Q_N(_07228_),
    .Q(\mem.mem[237][1] ));
 sg13g2_dfrbp_1 _20363_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1428),
    .D(_01999_),
    .Q_N(_07227_),
    .Q(\mem.mem[237][2] ));
 sg13g2_dfrbp_1 _20364_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1427),
    .D(_02000_),
    .Q_N(_07226_),
    .Q(\mem.mem[237][3] ));
 sg13g2_dfrbp_1 _20365_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1426),
    .D(_02001_),
    .Q_N(_07225_),
    .Q(\mem.mem[237][4] ));
 sg13g2_dfrbp_1 _20366_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1425),
    .D(_02002_),
    .Q_N(_07224_),
    .Q(\mem.mem[237][5] ));
 sg13g2_dfrbp_1 _20367_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1424),
    .D(_02003_),
    .Q_N(_07223_),
    .Q(\mem.mem[237][6] ));
 sg13g2_dfrbp_1 _20368_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1423),
    .D(_02004_),
    .Q_N(_07222_),
    .Q(\mem.mem[237][7] ));
 sg13g2_dfrbp_1 _20369_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1422),
    .D(_02005_),
    .Q_N(_07221_),
    .Q(\mem.mem[238][0] ));
 sg13g2_dfrbp_1 _20370_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1421),
    .D(_02006_),
    .Q_N(_07220_),
    .Q(\mem.mem[238][1] ));
 sg13g2_dfrbp_1 _20371_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1420),
    .D(_02007_),
    .Q_N(_07219_),
    .Q(\mem.mem[238][2] ));
 sg13g2_dfrbp_1 _20372_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1419),
    .D(_02008_),
    .Q_N(_07218_),
    .Q(\mem.mem[238][3] ));
 sg13g2_dfrbp_1 _20373_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1418),
    .D(_02009_),
    .Q_N(_07217_),
    .Q(\mem.mem[238][4] ));
 sg13g2_dfrbp_1 _20374_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1417),
    .D(_02010_),
    .Q_N(_07216_),
    .Q(\mem.mem[238][5] ));
 sg13g2_dfrbp_1 _20375_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1416),
    .D(_02011_),
    .Q_N(_07215_),
    .Q(\mem.mem[238][6] ));
 sg13g2_dfrbp_1 _20376_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1415),
    .D(_02012_),
    .Q_N(_07214_),
    .Q(\mem.mem[238][7] ));
 sg13g2_dfrbp_1 _20377_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1414),
    .D(_02013_),
    .Q_N(_07213_),
    .Q(\mem.mem[23][0] ));
 sg13g2_dfrbp_1 _20378_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1413),
    .D(_02014_),
    .Q_N(_07212_),
    .Q(\mem.mem[23][1] ));
 sg13g2_dfrbp_1 _20379_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1412),
    .D(_02015_),
    .Q_N(_07211_),
    .Q(\mem.mem[23][2] ));
 sg13g2_dfrbp_1 _20380_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1411),
    .D(_02016_),
    .Q_N(_07210_),
    .Q(\mem.mem[23][3] ));
 sg13g2_dfrbp_1 _20381_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1410),
    .D(_02017_),
    .Q_N(_07209_),
    .Q(\mem.mem[23][4] ));
 sg13g2_dfrbp_1 _20382_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1409),
    .D(_02018_),
    .Q_N(_07208_),
    .Q(\mem.mem[23][5] ));
 sg13g2_dfrbp_1 _20383_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1408),
    .D(_02019_),
    .Q_N(_07207_),
    .Q(\mem.mem[23][6] ));
 sg13g2_dfrbp_1 _20384_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1407),
    .D(_02020_),
    .Q_N(_07206_),
    .Q(\mem.mem[23][7] ));
 sg13g2_dfrbp_1 _20385_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1406),
    .D(_02021_),
    .Q_N(_07205_),
    .Q(\mem.mem[240][0] ));
 sg13g2_dfrbp_1 _20386_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1405),
    .D(_02022_),
    .Q_N(_07204_),
    .Q(\mem.mem[240][1] ));
 sg13g2_dfrbp_1 _20387_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1404),
    .D(_02023_),
    .Q_N(_07203_),
    .Q(\mem.mem[240][2] ));
 sg13g2_dfrbp_1 _20388_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1403),
    .D(_02024_),
    .Q_N(_07202_),
    .Q(\mem.mem[240][3] ));
 sg13g2_dfrbp_1 _20389_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1402),
    .D(_02025_),
    .Q_N(_07201_),
    .Q(\mem.mem[240][4] ));
 sg13g2_dfrbp_1 _20390_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1401),
    .D(_02026_),
    .Q_N(_07200_),
    .Q(\mem.mem[240][5] ));
 sg13g2_dfrbp_1 _20391_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1400),
    .D(_02027_),
    .Q_N(_07199_),
    .Q(\mem.mem[240][6] ));
 sg13g2_dfrbp_1 _20392_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1399),
    .D(_02028_),
    .Q_N(_07198_),
    .Q(\mem.mem[240][7] ));
 sg13g2_dfrbp_1 _20393_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1398),
    .D(_02029_),
    .Q_N(_07197_),
    .Q(\mem.mem[241][0] ));
 sg13g2_dfrbp_1 _20394_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1397),
    .D(_02030_),
    .Q_N(_07196_),
    .Q(\mem.mem[241][1] ));
 sg13g2_dfrbp_1 _20395_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1396),
    .D(_02031_),
    .Q_N(_07195_),
    .Q(\mem.mem[241][2] ));
 sg13g2_dfrbp_1 _20396_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1395),
    .D(_02032_),
    .Q_N(_07194_),
    .Q(\mem.mem[241][3] ));
 sg13g2_dfrbp_1 _20397_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1394),
    .D(_02033_),
    .Q_N(_07193_),
    .Q(\mem.mem[241][4] ));
 sg13g2_dfrbp_1 _20398_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1393),
    .D(_02034_),
    .Q_N(_07192_),
    .Q(\mem.mem[241][5] ));
 sg13g2_dfrbp_1 _20399_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1392),
    .D(_02035_),
    .Q_N(_07191_),
    .Q(\mem.mem[241][6] ));
 sg13g2_dfrbp_1 _20400_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1391),
    .D(_02036_),
    .Q_N(_07190_),
    .Q(\mem.mem[241][7] ));
 sg13g2_dfrbp_1 _20401_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1390),
    .D(_02037_),
    .Q_N(_07189_),
    .Q(\mem.mem[242][0] ));
 sg13g2_dfrbp_1 _20402_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1389),
    .D(_02038_),
    .Q_N(_07188_),
    .Q(\mem.mem[242][1] ));
 sg13g2_dfrbp_1 _20403_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1388),
    .D(_02039_),
    .Q_N(_07187_),
    .Q(\mem.mem[242][2] ));
 sg13g2_dfrbp_1 _20404_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1387),
    .D(_02040_),
    .Q_N(_07186_),
    .Q(\mem.mem[242][3] ));
 sg13g2_dfrbp_1 _20405_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1386),
    .D(_02041_),
    .Q_N(_07185_),
    .Q(\mem.mem[242][4] ));
 sg13g2_dfrbp_1 _20406_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1385),
    .D(_02042_),
    .Q_N(_07184_),
    .Q(\mem.mem[242][5] ));
 sg13g2_dfrbp_1 _20407_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1384),
    .D(_02043_),
    .Q_N(_07183_),
    .Q(\mem.mem[242][6] ));
 sg13g2_dfrbp_1 _20408_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1383),
    .D(_02044_),
    .Q_N(_07182_),
    .Q(\mem.mem[242][7] ));
 sg13g2_dfrbp_1 _20409_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1382),
    .D(_02045_),
    .Q_N(_07181_),
    .Q(\mem.mem[243][0] ));
 sg13g2_dfrbp_1 _20410_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1381),
    .D(_02046_),
    .Q_N(_07180_),
    .Q(\mem.mem[243][1] ));
 sg13g2_dfrbp_1 _20411_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1380),
    .D(_02047_),
    .Q_N(_07179_),
    .Q(\mem.mem[243][2] ));
 sg13g2_dfrbp_1 _20412_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1379),
    .D(_02048_),
    .Q_N(_07178_),
    .Q(\mem.mem[243][3] ));
 sg13g2_dfrbp_1 _20413_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1378),
    .D(_02049_),
    .Q_N(_07177_),
    .Q(\mem.mem[243][4] ));
 sg13g2_dfrbp_1 _20414_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1377),
    .D(_02050_),
    .Q_N(_07176_),
    .Q(\mem.mem[243][5] ));
 sg13g2_dfrbp_1 _20415_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1376),
    .D(_02051_),
    .Q_N(_07175_),
    .Q(\mem.mem[243][6] ));
 sg13g2_dfrbp_1 _20416_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1375),
    .D(_02052_),
    .Q_N(_07174_),
    .Q(\mem.mem[243][7] ));
 sg13g2_dfrbp_1 _20417_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1374),
    .D(_02053_),
    .Q_N(_07173_),
    .Q(\mem.mem[244][0] ));
 sg13g2_dfrbp_1 _20418_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1373),
    .D(_02054_),
    .Q_N(_07172_),
    .Q(\mem.mem[244][1] ));
 sg13g2_dfrbp_1 _20419_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1372),
    .D(_02055_),
    .Q_N(_07171_),
    .Q(\mem.mem[244][2] ));
 sg13g2_dfrbp_1 _20420_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1371),
    .D(_02056_),
    .Q_N(_07170_),
    .Q(\mem.mem[244][3] ));
 sg13g2_dfrbp_1 _20421_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1370),
    .D(_02057_),
    .Q_N(_07169_),
    .Q(\mem.mem[244][4] ));
 sg13g2_dfrbp_1 _20422_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1369),
    .D(_02058_),
    .Q_N(_07168_),
    .Q(\mem.mem[244][5] ));
 sg13g2_dfrbp_1 _20423_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1368),
    .D(_02059_),
    .Q_N(_07167_),
    .Q(\mem.mem[244][6] ));
 sg13g2_dfrbp_1 _20424_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1367),
    .D(_02060_),
    .Q_N(_07166_),
    .Q(\mem.mem[244][7] ));
 sg13g2_dfrbp_1 _20425_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1366),
    .D(_02061_),
    .Q_N(_07165_),
    .Q(\mem.mem[245][0] ));
 sg13g2_dfrbp_1 _20426_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net844),
    .D(_02062_),
    .Q_N(_07164_),
    .Q(\mem.mem[245][1] ));
 sg13g2_dfrbp_1 _20427_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net842),
    .D(_02063_),
    .Q_N(_07163_),
    .Q(\mem.mem[245][2] ));
 sg13g2_dfrbp_1 _20428_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net840),
    .D(_02064_),
    .Q_N(_07162_),
    .Q(\mem.mem[245][3] ));
 sg13g2_dfrbp_1 _20429_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net838),
    .D(_02065_),
    .Q_N(_07161_),
    .Q(\mem.mem[245][4] ));
 sg13g2_dfrbp_1 _20430_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net836),
    .D(_02066_),
    .Q_N(_07160_),
    .Q(\mem.mem[245][5] ));
 sg13g2_dfrbp_1 _20431_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net834),
    .D(_02067_),
    .Q_N(_07159_),
    .Q(\mem.mem[245][6] ));
 sg13g2_dfrbp_1 _20432_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net832),
    .D(_02068_),
    .Q_N(_07158_),
    .Q(\mem.mem[245][7] ));
 sg13g2_dfrbp_1 _20433_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net830),
    .D(_02069_),
    .Q_N(_07157_),
    .Q(\mem.mem[246][0] ));
 sg13g2_dfrbp_1 _20434_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net828),
    .D(_02070_),
    .Q_N(_07156_),
    .Q(\mem.mem[246][1] ));
 sg13g2_dfrbp_1 _20435_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net826),
    .D(_02071_),
    .Q_N(_07155_),
    .Q(\mem.mem[246][2] ));
 sg13g2_dfrbp_1 _20436_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net824),
    .D(_02072_),
    .Q_N(_07154_),
    .Q(\mem.mem[246][3] ));
 sg13g2_dfrbp_1 _20437_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net822),
    .D(_02073_),
    .Q_N(_07153_),
    .Q(\mem.mem[246][4] ));
 sg13g2_dfrbp_1 _20438_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net820),
    .D(_02074_),
    .Q_N(_07152_),
    .Q(\mem.mem[246][5] ));
 sg13g2_dfrbp_1 _20439_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net818),
    .D(_02075_),
    .Q_N(_07151_),
    .Q(\mem.mem[246][6] ));
 sg13g2_dfrbp_1 _20440_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net816),
    .D(_02076_),
    .Q_N(_07150_),
    .Q(\mem.mem[246][7] ));
 sg13g2_dfrbp_1 _20441_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net814),
    .D(_02077_),
    .Q_N(_07149_),
    .Q(\mem.mem[247][0] ));
 sg13g2_dfrbp_1 _20442_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net812),
    .D(_02078_),
    .Q_N(_07148_),
    .Q(\mem.mem[247][1] ));
 sg13g2_dfrbp_1 _20443_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net810),
    .D(_02079_),
    .Q_N(_07147_),
    .Q(\mem.mem[247][2] ));
 sg13g2_dfrbp_1 _20444_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net808),
    .D(_02080_),
    .Q_N(_07146_),
    .Q(\mem.mem[247][3] ));
 sg13g2_dfrbp_1 _20445_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net806),
    .D(_02081_),
    .Q_N(_07145_),
    .Q(\mem.mem[247][4] ));
 sg13g2_dfrbp_1 _20446_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net804),
    .D(_02082_),
    .Q_N(_07144_),
    .Q(\mem.mem[247][5] ));
 sg13g2_dfrbp_1 _20447_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net802),
    .D(_02083_),
    .Q_N(_07143_),
    .Q(\mem.mem[247][6] ));
 sg13g2_dfrbp_1 _20448_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net800),
    .D(_02084_),
    .Q_N(_07142_),
    .Q(\mem.mem[247][7] ));
 sg13g2_dfrbp_1 _20449_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net798),
    .D(_02085_),
    .Q_N(_07141_),
    .Q(\mem.mem[248][0] ));
 sg13g2_dfrbp_1 _20450_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net796),
    .D(_02086_),
    .Q_N(_07140_),
    .Q(\mem.mem[248][1] ));
 sg13g2_dfrbp_1 _20451_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net794),
    .D(_02087_),
    .Q_N(_07139_),
    .Q(\mem.mem[248][2] ));
 sg13g2_dfrbp_1 _20452_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net792),
    .D(_02088_),
    .Q_N(_07138_),
    .Q(\mem.mem[248][3] ));
 sg13g2_dfrbp_1 _20453_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net790),
    .D(_02089_),
    .Q_N(_07137_),
    .Q(\mem.mem[248][4] ));
 sg13g2_dfrbp_1 _20454_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net788),
    .D(_02090_),
    .Q_N(_07136_),
    .Q(\mem.mem[248][5] ));
 sg13g2_dfrbp_1 _20455_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net786),
    .D(_02091_),
    .Q_N(_07135_),
    .Q(\mem.mem[248][6] ));
 sg13g2_dfrbp_1 _20456_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net784),
    .D(_02092_),
    .Q_N(_07134_),
    .Q(\mem.mem[248][7] ));
 sg13g2_dfrbp_1 _20457_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net782),
    .D(_02093_),
    .Q_N(_07133_),
    .Q(\mem.mem[24][0] ));
 sg13g2_dfrbp_1 _20458_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net780),
    .D(_02094_),
    .Q_N(_07132_),
    .Q(\mem.mem[24][1] ));
 sg13g2_dfrbp_1 _20459_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net778),
    .D(_02095_),
    .Q_N(_07131_),
    .Q(\mem.mem[24][2] ));
 sg13g2_dfrbp_1 _20460_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net776),
    .D(_02096_),
    .Q_N(_07130_),
    .Q(\mem.mem[24][3] ));
 sg13g2_dfrbp_1 _20461_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net774),
    .D(_02097_),
    .Q_N(_07129_),
    .Q(\mem.mem[24][4] ));
 sg13g2_dfrbp_1 _20462_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net772),
    .D(_02098_),
    .Q_N(_07128_),
    .Q(\mem.mem[24][5] ));
 sg13g2_dfrbp_1 _20463_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net770),
    .D(_02099_),
    .Q_N(_07127_),
    .Q(\mem.mem[24][6] ));
 sg13g2_dfrbp_1 _20464_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net768),
    .D(_02100_),
    .Q_N(_07126_),
    .Q(\mem.mem[24][7] ));
 sg13g2_dfrbp_1 _20465_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net766),
    .D(_02101_),
    .Q_N(_07125_),
    .Q(\mem.mem[250][0] ));
 sg13g2_dfrbp_1 _20466_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net756),
    .D(_02102_),
    .Q_N(_07124_),
    .Q(\mem.mem[250][1] ));
 sg13g2_dfrbp_1 _20467_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net754),
    .D(_02103_),
    .Q_N(_07123_),
    .Q(\mem.mem[250][2] ));
 sg13g2_dfrbp_1 _20468_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net752),
    .D(_02104_),
    .Q_N(_07122_),
    .Q(\mem.mem[250][3] ));
 sg13g2_dfrbp_1 _20469_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net750),
    .D(_02105_),
    .Q_N(_07121_),
    .Q(\mem.mem[250][4] ));
 sg13g2_dfrbp_1 _20470_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net748),
    .D(_02106_),
    .Q_N(_07120_),
    .Q(\mem.mem[250][5] ));
 sg13g2_dfrbp_1 _20471_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net746),
    .D(_02107_),
    .Q_N(_07119_),
    .Q(\mem.mem[250][6] ));
 sg13g2_dfrbp_1 _20472_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net744),
    .D(_02108_),
    .Q_N(_07118_),
    .Q(\mem.mem[250][7] ));
 sg13g2_dfrbp_1 _20473_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net742),
    .D(_02109_),
    .Q_N(_07117_),
    .Q(\mem.mem[251][0] ));
 sg13g2_dfrbp_1 _20474_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net740),
    .D(_02110_),
    .Q_N(_07116_),
    .Q(\mem.mem[251][1] ));
 sg13g2_dfrbp_1 _20475_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net738),
    .D(_02111_),
    .Q_N(_07115_),
    .Q(\mem.mem[251][2] ));
 sg13g2_dfrbp_1 _20476_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net736),
    .D(_02112_),
    .Q_N(_07114_),
    .Q(\mem.mem[251][3] ));
 sg13g2_dfrbp_1 _20477_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net734),
    .D(_02113_),
    .Q_N(_07113_),
    .Q(\mem.mem[251][4] ));
 sg13g2_dfrbp_1 _20478_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net732),
    .D(_02114_),
    .Q_N(_07112_),
    .Q(\mem.mem[251][5] ));
 sg13g2_dfrbp_1 _20479_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net730),
    .D(_02115_),
    .Q_N(_07111_),
    .Q(\mem.mem[251][6] ));
 sg13g2_dfrbp_1 _20480_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net728),
    .D(_02116_),
    .Q_N(_07110_),
    .Q(\mem.mem[251][7] ));
 sg13g2_dfrbp_1 _20481_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net726),
    .D(_02117_),
    .Q_N(_07109_),
    .Q(\mem.mem[9][0] ));
 sg13g2_dfrbp_1 _20482_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net525),
    .D(_02118_),
    .Q_N(_07108_),
    .Q(\mem.mem[9][1] ));
 sg13g2_dfrbp_1 _20483_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net523),
    .D(_02119_),
    .Q_N(_07107_),
    .Q(\mem.mem[9][2] ));
 sg13g2_dfrbp_1 _20484_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net521),
    .D(_02120_),
    .Q_N(_07106_),
    .Q(\mem.mem[9][3] ));
 sg13g2_dfrbp_1 _20485_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net519),
    .D(_02121_),
    .Q_N(_07105_),
    .Q(\mem.mem[9][4] ));
 sg13g2_dfrbp_1 _20486_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net517),
    .D(_02122_),
    .Q_N(_07104_),
    .Q(\mem.mem[9][5] ));
 sg13g2_dfrbp_1 _20487_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net515),
    .D(_02123_),
    .Q_N(_07103_),
    .Q(\mem.mem[9][6] ));
 sg13g2_dfrbp_1 _20488_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net513),
    .D(_02124_),
    .Q_N(_07102_),
    .Q(\mem.mem[9][7] ));
 sg13g2_dfrbp_1 _20489_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net511),
    .D(_02125_),
    .Q_N(_00015_),
    .Q(\mem.wr_en ));
 sg13g2_tiehi _19660__25 (.L_HI(net25));
 sg13g2_tiehi _19659__26 (.L_HI(net26));
 sg13g2_tiehi _19658__27 (.L_HI(net27));
 sg13g2_tiehi _19657__28 (.L_HI(net28));
 sg13g2_tiehi _19656__29 (.L_HI(net29));
 sg13g2_tiehi _19655__30 (.L_HI(net30));
 sg13g2_tiehi _19654__31 (.L_HI(net31));
 sg13g2_tiehi _19653__32 (.L_HI(net32));
 sg13g2_tiehi _19652__33 (.L_HI(net33));
 sg13g2_tiehi _19651__34 (.L_HI(net34));
 sg13g2_tiehi _19650__35 (.L_HI(net35));
 sg13g2_tiehi _19649__36 (.L_HI(net36));
 sg13g2_tiehi _19648__37 (.L_HI(net37));
 sg13g2_tiehi _19647__38 (.L_HI(net38));
 sg13g2_tiehi _19646__39 (.L_HI(net39));
 sg13g2_tiehi _19645__40 (.L_HI(net40));
 sg13g2_tiehi _19644__41 (.L_HI(net41));
 sg13g2_tiehi _19643__42 (.L_HI(net42));
 sg13g2_tiehi _19642__43 (.L_HI(net43));
 sg13g2_tiehi _19641__44 (.L_HI(net44));
 sg13g2_tiehi _19640__45 (.L_HI(net45));
 sg13g2_tiehi _19639__46 (.L_HI(net46));
 sg13g2_tiehi _19638__47 (.L_HI(net47));
 sg13g2_tiehi _19637__48 (.L_HI(net48));
 sg13g2_tiehi _19636__49 (.L_HI(net49));
 sg13g2_tiehi _19635__50 (.L_HI(net50));
 sg13g2_tiehi _19634__51 (.L_HI(net51));
 sg13g2_tiehi _19633__52 (.L_HI(net52));
 sg13g2_tiehi _19632__53 (.L_HI(net53));
 sg13g2_tiehi _19631__54 (.L_HI(net54));
 sg13g2_tiehi _19630__55 (.L_HI(net55));
 sg13g2_tiehi _19629__56 (.L_HI(net56));
 sg13g2_tiehi _19628__57 (.L_HI(net57));
 sg13g2_tiehi _19627__58 (.L_HI(net58));
 sg13g2_tiehi _19626__59 (.L_HI(net59));
 sg13g2_tiehi _19625__60 (.L_HI(net60));
 sg13g2_tiehi _19624__61 (.L_HI(net61));
 sg13g2_tiehi _19623__62 (.L_HI(net62));
 sg13g2_tiehi _19622__63 (.L_HI(net63));
 sg13g2_tiehi _19621__64 (.L_HI(net64));
 sg13g2_tiehi _19620__65 (.L_HI(net65));
 sg13g2_tiehi _19619__66 (.L_HI(net66));
 sg13g2_tiehi _19618__67 (.L_HI(net67));
 sg13g2_tiehi _19617__68 (.L_HI(net68));
 sg13g2_tiehi _19616__69 (.L_HI(net69));
 sg13g2_tiehi _19615__70 (.L_HI(net70));
 sg13g2_tiehi _19614__71 (.L_HI(net71));
 sg13g2_tiehi _19613__72 (.L_HI(net72));
 sg13g2_tiehi _19612__73 (.L_HI(net73));
 sg13g2_tiehi _19611__74 (.L_HI(net74));
 sg13g2_tiehi _19610__75 (.L_HI(net75));
 sg13g2_tiehi _19609__76 (.L_HI(net76));
 sg13g2_tiehi _19608__77 (.L_HI(net77));
 sg13g2_tiehi _19607__78 (.L_HI(net78));
 sg13g2_tiehi _19606__79 (.L_HI(net79));
 sg13g2_tiehi _19605__80 (.L_HI(net80));
 sg13g2_tiehi _19604__81 (.L_HI(net81));
 sg13g2_tiehi _19603__82 (.L_HI(net82));
 sg13g2_tiehi _19602__83 (.L_HI(net83));
 sg13g2_tiehi _19601__84 (.L_HI(net84));
 sg13g2_tiehi _19600__85 (.L_HI(net85));
 sg13g2_tiehi _19599__86 (.L_HI(net86));
 sg13g2_tiehi _19598__87 (.L_HI(net87));
 sg13g2_tiehi _19597__88 (.L_HI(net88));
 sg13g2_tiehi _19596__89 (.L_HI(net89));
 sg13g2_tiehi _19595__90 (.L_HI(net90));
 sg13g2_tiehi _19594__91 (.L_HI(net91));
 sg13g2_tiehi _19593__92 (.L_HI(net92));
 sg13g2_tiehi _19592__93 (.L_HI(net93));
 sg13g2_tiehi _19591__94 (.L_HI(net94));
 sg13g2_tiehi _19590__95 (.L_HI(net95));
 sg13g2_tiehi _19589__96 (.L_HI(net96));
 sg13g2_tiehi _19588__97 (.L_HI(net97));
 sg13g2_tiehi _19587__98 (.L_HI(net98));
 sg13g2_tiehi _19586__99 (.L_HI(net99));
 sg13g2_tiehi _19585__100 (.L_HI(net100));
 sg13g2_tiehi _19584__101 (.L_HI(net101));
 sg13g2_tiehi _19583__102 (.L_HI(net102));
 sg13g2_tiehi _19582__103 (.L_HI(net103));
 sg13g2_tiehi _19581__104 (.L_HI(net104));
 sg13g2_tiehi _19580__105 (.L_HI(net105));
 sg13g2_tiehi _19579__106 (.L_HI(net106));
 sg13g2_tiehi _19578__107 (.L_HI(net107));
 sg13g2_tiehi _19577__108 (.L_HI(net108));
 sg13g2_tiehi _19576__109 (.L_HI(net109));
 sg13g2_tiehi _19575__110 (.L_HI(net110));
 sg13g2_tiehi _19574__111 (.L_HI(net111));
 sg13g2_tiehi _19573__112 (.L_HI(net112));
 sg13g2_tiehi _19572__113 (.L_HI(net113));
 sg13g2_tiehi _19571__114 (.L_HI(net114));
 sg13g2_tiehi _19570__115 (.L_HI(net115));
 sg13g2_tiehi _19569__116 (.L_HI(net116));
 sg13g2_tiehi _19568__117 (.L_HI(net117));
 sg13g2_tiehi _19567__118 (.L_HI(net118));
 sg13g2_tiehi _19566__119 (.L_HI(net119));
 sg13g2_tiehi _19565__120 (.L_HI(net120));
 sg13g2_tiehi _19564__121 (.L_HI(net121));
 sg13g2_tiehi _19563__122 (.L_HI(net122));
 sg13g2_tiehi _19562__123 (.L_HI(net123));
 sg13g2_tiehi _19561__124 (.L_HI(net124));
 sg13g2_tiehi _19560__125 (.L_HI(net125));
 sg13g2_tiehi _19559__126 (.L_HI(net126));
 sg13g2_tiehi _19558__127 (.L_HI(net127));
 sg13g2_tiehi _19557__128 (.L_HI(net128));
 sg13g2_tiehi _19556__129 (.L_HI(net129));
 sg13g2_tiehi _19555__130 (.L_HI(net130));
 sg13g2_tiehi _19554__131 (.L_HI(net131));
 sg13g2_tiehi _19553__132 (.L_HI(net132));
 sg13g2_tiehi _19552__133 (.L_HI(net133));
 sg13g2_tiehi _19551__134 (.L_HI(net134));
 sg13g2_tiehi _19550__135 (.L_HI(net135));
 sg13g2_tiehi _19549__136 (.L_HI(net136));
 sg13g2_tiehi _19548__137 (.L_HI(net137));
 sg13g2_tiehi _19547__138 (.L_HI(net138));
 sg13g2_tiehi _19546__139 (.L_HI(net139));
 sg13g2_tiehi _19545__140 (.L_HI(net140));
 sg13g2_tiehi _19544__141 (.L_HI(net141));
 sg13g2_tiehi _19543__142 (.L_HI(net142));
 sg13g2_tiehi _19542__143 (.L_HI(net143));
 sg13g2_tiehi _19541__144 (.L_HI(net144));
 sg13g2_tiehi _19540__145 (.L_HI(net145));
 sg13g2_tiehi _19539__146 (.L_HI(net146));
 sg13g2_tiehi _19538__147 (.L_HI(net147));
 sg13g2_tiehi _19537__148 (.L_HI(net148));
 sg13g2_tiehi _19536__149 (.L_HI(net149));
 sg13g2_tiehi _19535__150 (.L_HI(net150));
 sg13g2_tiehi _19534__151 (.L_HI(net151));
 sg13g2_tiehi _19533__152 (.L_HI(net152));
 sg13g2_tiehi _19532__153 (.L_HI(net153));
 sg13g2_tiehi _19531__154 (.L_HI(net154));
 sg13g2_tiehi _19530__155 (.L_HI(net155));
 sg13g2_tiehi _19529__156 (.L_HI(net156));
 sg13g2_tiehi _19528__157 (.L_HI(net157));
 sg13g2_tiehi _19527__158 (.L_HI(net158));
 sg13g2_tiehi _19526__159 (.L_HI(net159));
 sg13g2_tiehi _19525__160 (.L_HI(net160));
 sg13g2_tiehi _19524__161 (.L_HI(net161));
 sg13g2_tiehi _19523__162 (.L_HI(net162));
 sg13g2_tiehi _19522__163 (.L_HI(net163));
 sg13g2_tiehi _19521__164 (.L_HI(net164));
 sg13g2_tiehi _19520__165 (.L_HI(net165));
 sg13g2_tiehi _19519__166 (.L_HI(net166));
 sg13g2_tiehi _19518__167 (.L_HI(net167));
 sg13g2_tiehi _19517__168 (.L_HI(net168));
 sg13g2_tiehi _19516__169 (.L_HI(net169));
 sg13g2_tiehi _19515__170 (.L_HI(net170));
 sg13g2_tiehi _19514__171 (.L_HI(net171));
 sg13g2_tiehi _19513__172 (.L_HI(net172));
 sg13g2_tiehi _19512__173 (.L_HI(net173));
 sg13g2_tiehi _19511__174 (.L_HI(net174));
 sg13g2_tiehi _19510__175 (.L_HI(net175));
 sg13g2_tiehi _19509__176 (.L_HI(net176));
 sg13g2_tiehi _19508__177 (.L_HI(net177));
 sg13g2_tiehi _19507__178 (.L_HI(net178));
 sg13g2_tiehi _19506__179 (.L_HI(net179));
 sg13g2_tiehi _19505__180 (.L_HI(net180));
 sg13g2_tiehi _19504__181 (.L_HI(net181));
 sg13g2_tiehi _19503__182 (.L_HI(net182));
 sg13g2_tiehi _19502__183 (.L_HI(net183));
 sg13g2_tiehi _19501__184 (.L_HI(net184));
 sg13g2_tiehi _19500__185 (.L_HI(net185));
 sg13g2_tiehi _19499__186 (.L_HI(net186));
 sg13g2_tiehi _19498__187 (.L_HI(net187));
 sg13g2_tiehi _19497__188 (.L_HI(net188));
 sg13g2_tiehi _19496__189 (.L_HI(net189));
 sg13g2_tiehi _19495__190 (.L_HI(net190));
 sg13g2_tiehi _19494__191 (.L_HI(net191));
 sg13g2_tiehi _19493__192 (.L_HI(net192));
 sg13g2_tiehi _19492__193 (.L_HI(net193));
 sg13g2_tiehi _19491__194 (.L_HI(net194));
 sg13g2_tiehi _19490__195 (.L_HI(net195));
 sg13g2_tiehi _19489__196 (.L_HI(net196));
 sg13g2_tiehi _19488__197 (.L_HI(net197));
 sg13g2_tiehi _19487__198 (.L_HI(net198));
 sg13g2_tiehi _19486__199 (.L_HI(net199));
 sg13g2_tiehi _19485__200 (.L_HI(net200));
 sg13g2_tiehi _19484__201 (.L_HI(net201));
 sg13g2_tiehi _19483__202 (.L_HI(net202));
 sg13g2_tiehi _19482__203 (.L_HI(net203));
 sg13g2_tiehi _19481__204 (.L_HI(net204));
 sg13g2_tiehi _19480__205 (.L_HI(net205));
 sg13g2_tiehi _19479__206 (.L_HI(net206));
 sg13g2_tiehi _19478__207 (.L_HI(net207));
 sg13g2_tiehi _19477__208 (.L_HI(net208));
 sg13g2_tiehi _19476__209 (.L_HI(net209));
 sg13g2_tiehi _19475__210 (.L_HI(net210));
 sg13g2_tiehi _19474__211 (.L_HI(net211));
 sg13g2_tiehi _19473__212 (.L_HI(net212));
 sg13g2_tiehi _19472__213 (.L_HI(net213));
 sg13g2_tiehi _19471__214 (.L_HI(net214));
 sg13g2_tiehi _19470__215 (.L_HI(net215));
 sg13g2_tiehi _19469__216 (.L_HI(net216));
 sg13g2_tiehi _19468__217 (.L_HI(net217));
 sg13g2_tiehi _19467__218 (.L_HI(net218));
 sg13g2_tiehi _19466__219 (.L_HI(net219));
 sg13g2_tiehi _19465__220 (.L_HI(net220));
 sg13g2_tiehi _19464__221 (.L_HI(net221));
 sg13g2_tiehi _19463__222 (.L_HI(net222));
 sg13g2_tiehi _19462__223 (.L_HI(net223));
 sg13g2_tiehi _19461__224 (.L_HI(net224));
 sg13g2_tiehi _19460__225 (.L_HI(net225));
 sg13g2_tiehi _19459__226 (.L_HI(net226));
 sg13g2_tiehi _19458__227 (.L_HI(net227));
 sg13g2_tiehi _19457__228 (.L_HI(net228));
 sg13g2_tiehi _19456__229 (.L_HI(net229));
 sg13g2_tiehi _19455__230 (.L_HI(net230));
 sg13g2_tiehi _19454__231 (.L_HI(net231));
 sg13g2_tiehi _19453__232 (.L_HI(net232));
 sg13g2_tiehi _19452__233 (.L_HI(net233));
 sg13g2_tiehi _19451__234 (.L_HI(net234));
 sg13g2_tiehi _19450__235 (.L_HI(net235));
 sg13g2_tiehi _19449__236 (.L_HI(net236));
 sg13g2_tiehi _19448__237 (.L_HI(net237));
 sg13g2_tiehi _19447__238 (.L_HI(net238));
 sg13g2_tiehi _19446__239 (.L_HI(net239));
 sg13g2_tiehi _19445__240 (.L_HI(net240));
 sg13g2_tiehi _19444__241 (.L_HI(net241));
 sg13g2_tiehi _19443__242 (.L_HI(net242));
 sg13g2_tiehi _19442__243 (.L_HI(net243));
 sg13g2_tiehi _19441__244 (.L_HI(net244));
 sg13g2_tiehi _19440__245 (.L_HI(net245));
 sg13g2_tiehi _19439__246 (.L_HI(net246));
 sg13g2_tiehi _19438__247 (.L_HI(net247));
 sg13g2_tiehi _19437__248 (.L_HI(net248));
 sg13g2_tiehi _19436__249 (.L_HI(net249));
 sg13g2_tiehi _19435__250 (.L_HI(net250));
 sg13g2_tiehi _19434__251 (.L_HI(net251));
 sg13g2_tiehi _19433__252 (.L_HI(net252));
 sg13g2_tiehi _19432__253 (.L_HI(net253));
 sg13g2_tiehi _19431__254 (.L_HI(net254));
 sg13g2_tiehi _19430__255 (.L_HI(net255));
 sg13g2_tiehi _19429__256 (.L_HI(net256));
 sg13g2_tiehi _19428__257 (.L_HI(net257));
 sg13g2_tiehi _19427__258 (.L_HI(net258));
 sg13g2_tiehi _19426__259 (.L_HI(net259));
 sg13g2_tiehi _19425__260 (.L_HI(net260));
 sg13g2_tiehi _19424__261 (.L_HI(net261));
 sg13g2_tiehi _19423__262 (.L_HI(net262));
 sg13g2_tiehi _19422__263 (.L_HI(net263));
 sg13g2_tiehi _19421__264 (.L_HI(net264));
 sg13g2_tiehi _19420__265 (.L_HI(net265));
 sg13g2_tiehi _19419__266 (.L_HI(net266));
 sg13g2_tiehi _19418__267 (.L_HI(net267));
 sg13g2_tiehi _19417__268 (.L_HI(net268));
 sg13g2_tiehi _19416__269 (.L_HI(net269));
 sg13g2_tiehi _19415__270 (.L_HI(net270));
 sg13g2_tiehi _19414__271 (.L_HI(net271));
 sg13g2_tiehi _19413__272 (.L_HI(net272));
 sg13g2_tiehi _19412__273 (.L_HI(net273));
 sg13g2_tiehi _19411__274 (.L_HI(net274));
 sg13g2_tiehi _19410__275 (.L_HI(net275));
 sg13g2_tiehi _19409__276 (.L_HI(net276));
 sg13g2_tiehi _19408__277 (.L_HI(net277));
 sg13g2_tiehi _19407__278 (.L_HI(net278));
 sg13g2_tiehi _19406__279 (.L_HI(net279));
 sg13g2_tiehi _19405__280 (.L_HI(net280));
 sg13g2_tiehi _19404__281 (.L_HI(net281));
 sg13g2_tiehi _19403__282 (.L_HI(net282));
 sg13g2_tiehi _19402__283 (.L_HI(net283));
 sg13g2_tiehi _19401__284 (.L_HI(net284));
 sg13g2_tiehi _19400__285 (.L_HI(net285));
 sg13g2_tiehi _19399__286 (.L_HI(net286));
 sg13g2_tiehi _19398__287 (.L_HI(net287));
 sg13g2_tiehi _19397__288 (.L_HI(net288));
 sg13g2_tiehi _19396__289 (.L_HI(net289));
 sg13g2_tiehi _19395__290 (.L_HI(net290));
 sg13g2_tiehi _19394__291 (.L_HI(net291));
 sg13g2_tiehi _19393__292 (.L_HI(net292));
 sg13g2_tiehi _19392__293 (.L_HI(net293));
 sg13g2_tiehi _19391__294 (.L_HI(net294));
 sg13g2_tiehi _19390__295 (.L_HI(net295));
 sg13g2_tiehi _19389__296 (.L_HI(net296));
 sg13g2_tiehi _19388__297 (.L_HI(net297));
 sg13g2_tiehi _19387__298 (.L_HI(net298));
 sg13g2_tiehi _19386__299 (.L_HI(net299));
 sg13g2_tiehi _19385__300 (.L_HI(net300));
 sg13g2_tiehi _19384__301 (.L_HI(net301));
 sg13g2_tiehi _19383__302 (.L_HI(net302));
 sg13g2_tiehi _19382__303 (.L_HI(net303));
 sg13g2_tiehi _19381__304 (.L_HI(net304));
 sg13g2_tiehi _19380__305 (.L_HI(net305));
 sg13g2_tiehi _19379__306 (.L_HI(net306));
 sg13g2_tiehi _19378__307 (.L_HI(net307));
 sg13g2_tiehi _19377__308 (.L_HI(net308));
 sg13g2_tiehi _19376__309 (.L_HI(net309));
 sg13g2_tiehi _19375__310 (.L_HI(net310));
 sg13g2_tiehi _19374__311 (.L_HI(net311));
 sg13g2_tiehi _19373__312 (.L_HI(net312));
 sg13g2_tiehi _19372__313 (.L_HI(net313));
 sg13g2_tiehi _19371__314 (.L_HI(net314));
 sg13g2_tiehi _19370__315 (.L_HI(net315));
 sg13g2_tiehi _19369__316 (.L_HI(net316));
 sg13g2_tiehi _19368__317 (.L_HI(net317));
 sg13g2_tiehi _19367__318 (.L_HI(net318));
 sg13g2_tiehi _19366__319 (.L_HI(net319));
 sg13g2_tiehi _19365__320 (.L_HI(net320));
 sg13g2_tiehi _19364__321 (.L_HI(net321));
 sg13g2_tiehi _19363__322 (.L_HI(net322));
 sg13g2_tiehi _19362__323 (.L_HI(net323));
 sg13g2_tiehi _19361__324 (.L_HI(net324));
 sg13g2_tiehi _19360__325 (.L_HI(net325));
 sg13g2_tiehi _19359__326 (.L_HI(net326));
 sg13g2_tiehi _19358__327 (.L_HI(net327));
 sg13g2_tiehi _19357__328 (.L_HI(net328));
 sg13g2_tiehi _19356__329 (.L_HI(net329));
 sg13g2_tiehi _19355__330 (.L_HI(net330));
 sg13g2_tiehi _19354__331 (.L_HI(net331));
 sg13g2_tiehi _19353__332 (.L_HI(net332));
 sg13g2_tiehi _19352__333 (.L_HI(net333));
 sg13g2_tiehi _19351__334 (.L_HI(net334));
 sg13g2_tiehi _19350__335 (.L_HI(net335));
 sg13g2_tiehi _19349__336 (.L_HI(net336));
 sg13g2_tiehi _19348__337 (.L_HI(net337));
 sg13g2_tiehi _19347__338 (.L_HI(net338));
 sg13g2_tiehi _19346__339 (.L_HI(net339));
 sg13g2_tiehi _19345__340 (.L_HI(net340));
 sg13g2_tiehi _19344__341 (.L_HI(net341));
 sg13g2_tiehi _19343__342 (.L_HI(net342));
 sg13g2_tiehi _19342__343 (.L_HI(net343));
 sg13g2_tiehi _19341__344 (.L_HI(net344));
 sg13g2_tiehi _19340__345 (.L_HI(net345));
 sg13g2_tiehi _19339__346 (.L_HI(net346));
 sg13g2_tiehi _19338__347 (.L_HI(net347));
 sg13g2_tiehi _19337__348 (.L_HI(net348));
 sg13g2_tiehi _19336__349 (.L_HI(net349));
 sg13g2_tiehi _19335__350 (.L_HI(net350));
 sg13g2_tiehi _19334__351 (.L_HI(net351));
 sg13g2_tiehi _19333__352 (.L_HI(net352));
 sg13g2_tiehi _19332__353 (.L_HI(net353));
 sg13g2_tiehi _19331__354 (.L_HI(net354));
 sg13g2_tiehi _19330__355 (.L_HI(net355));
 sg13g2_tiehi _19329__356 (.L_HI(net356));
 sg13g2_tiehi _19328__357 (.L_HI(net357));
 sg13g2_tiehi _19327__358 (.L_HI(net358));
 sg13g2_tiehi _19326__359 (.L_HI(net359));
 sg13g2_tiehi _19325__360 (.L_HI(net360));
 sg13g2_tiehi _19324__361 (.L_HI(net361));
 sg13g2_tiehi _19323__362 (.L_HI(net362));
 sg13g2_tiehi _19322__363 (.L_HI(net363));
 sg13g2_tiehi _19321__364 (.L_HI(net364));
 sg13g2_tiehi _19320__365 (.L_HI(net365));
 sg13g2_tiehi _19319__366 (.L_HI(net366));
 sg13g2_tiehi _19318__367 (.L_HI(net367));
 sg13g2_tiehi _19317__368 (.L_HI(net368));
 sg13g2_tiehi _19316__369 (.L_HI(net369));
 sg13g2_tiehi _19315__370 (.L_HI(net370));
 sg13g2_tiehi _19314__371 (.L_HI(net371));
 sg13g2_tiehi _19313__372 (.L_HI(net372));
 sg13g2_tiehi _19312__373 (.L_HI(net373));
 sg13g2_tiehi _19311__374 (.L_HI(net374));
 sg13g2_tiehi _19310__375 (.L_HI(net375));
 sg13g2_tiehi _19309__376 (.L_HI(net376));
 sg13g2_tiehi _19308__377 (.L_HI(net377));
 sg13g2_tiehi _19307__378 (.L_HI(net378));
 sg13g2_tiehi _19306__379 (.L_HI(net379));
 sg13g2_tiehi _19305__380 (.L_HI(net380));
 sg13g2_tiehi _19304__381 (.L_HI(net381));
 sg13g2_tiehi _19303__382 (.L_HI(net382));
 sg13g2_tiehi _19302__383 (.L_HI(net383));
 sg13g2_tiehi _19301__384 (.L_HI(net384));
 sg13g2_tiehi _19300__385 (.L_HI(net385));
 sg13g2_tiehi _19299__386 (.L_HI(net386));
 sg13g2_tiehi _19298__387 (.L_HI(net387));
 sg13g2_tiehi _19297__388 (.L_HI(net388));
 sg13g2_tiehi _19296__389 (.L_HI(net389));
 sg13g2_tiehi _19295__390 (.L_HI(net390));
 sg13g2_tiehi _19294__391 (.L_HI(net391));
 sg13g2_tiehi _19293__392 (.L_HI(net392));
 sg13g2_tiehi _19292__393 (.L_HI(net393));
 sg13g2_tiehi _19291__394 (.L_HI(net394));
 sg13g2_tiehi _19290__395 (.L_HI(net395));
 sg13g2_tiehi _19289__396 (.L_HI(net396));
 sg13g2_tiehi _19288__397 (.L_HI(net397));
 sg13g2_tiehi _19287__398 (.L_HI(net398));
 sg13g2_tiehi _19286__399 (.L_HI(net399));
 sg13g2_tiehi _19285__400 (.L_HI(net400));
 sg13g2_tiehi _19284__401 (.L_HI(net401));
 sg13g2_tiehi _19283__402 (.L_HI(net402));
 sg13g2_tiehi _19282__403 (.L_HI(net403));
 sg13g2_tiehi _19281__404 (.L_HI(net404));
 sg13g2_tiehi _19280__405 (.L_HI(net405));
 sg13g2_tiehi _19279__406 (.L_HI(net406));
 sg13g2_tiehi _19278__407 (.L_HI(net407));
 sg13g2_tiehi _19277__408 (.L_HI(net408));
 sg13g2_tiehi _19276__409 (.L_HI(net409));
 sg13g2_tiehi _19275__410 (.L_HI(net410));
 sg13g2_tiehi _19274__411 (.L_HI(net411));
 sg13g2_tiehi _19273__412 (.L_HI(net412));
 sg13g2_tiehi _19272__413 (.L_HI(net413));
 sg13g2_tiehi _19271__414 (.L_HI(net414));
 sg13g2_tiehi _19270__415 (.L_HI(net415));
 sg13g2_tiehi _19269__416 (.L_HI(net416));
 sg13g2_tiehi _19268__417 (.L_HI(net417));
 sg13g2_tiehi _19267__418 (.L_HI(net418));
 sg13g2_tiehi _19266__419 (.L_HI(net419));
 sg13g2_tiehi _19265__420 (.L_HI(net420));
 sg13g2_tiehi _19264__421 (.L_HI(net421));
 sg13g2_tiehi _19263__422 (.L_HI(net422));
 sg13g2_tiehi _19262__423 (.L_HI(net423));
 sg13g2_tiehi _19261__424 (.L_HI(net424));
 sg13g2_tiehi _19260__425 (.L_HI(net425));
 sg13g2_tiehi _19259__426 (.L_HI(net426));
 sg13g2_tiehi _19258__427 (.L_HI(net427));
 sg13g2_tiehi _19257__428 (.L_HI(net428));
 sg13g2_tiehi _19256__429 (.L_HI(net429));
 sg13g2_tiehi _19255__430 (.L_HI(net430));
 sg13g2_tiehi _19254__431 (.L_HI(net431));
 sg13g2_tiehi _19253__432 (.L_HI(net432));
 sg13g2_tiehi _19252__433 (.L_HI(net433));
 sg13g2_tiehi _19251__434 (.L_HI(net434));
 sg13g2_tiehi _19250__435 (.L_HI(net435));
 sg13g2_tiehi _19249__436 (.L_HI(net436));
 sg13g2_tiehi _19248__437 (.L_HI(net437));
 sg13g2_tiehi _19247__438 (.L_HI(net438));
 sg13g2_tiehi _19246__439 (.L_HI(net439));
 sg13g2_tiehi _19245__440 (.L_HI(net440));
 sg13g2_tiehi _19244__441 (.L_HI(net441));
 sg13g2_tiehi _19243__442 (.L_HI(net442));
 sg13g2_tiehi _19242__443 (.L_HI(net443));
 sg13g2_tiehi _19241__444 (.L_HI(net444));
 sg13g2_tiehi _19240__445 (.L_HI(net445));
 sg13g2_tiehi _19239__446 (.L_HI(net446));
 sg13g2_tiehi _19238__447 (.L_HI(net447));
 sg13g2_tiehi _19237__448 (.L_HI(net448));
 sg13g2_tiehi _19236__449 (.L_HI(net449));
 sg13g2_tiehi _19235__450 (.L_HI(net450));
 sg13g2_tiehi _19234__451 (.L_HI(net451));
 sg13g2_tiehi _19233__452 (.L_HI(net452));
 sg13g2_tiehi _19232__453 (.L_HI(net453));
 sg13g2_tiehi _19231__454 (.L_HI(net454));
 sg13g2_tiehi _19230__455 (.L_HI(net455));
 sg13g2_tiehi _19229__456 (.L_HI(net456));
 sg13g2_tiehi _19228__457 (.L_HI(net457));
 sg13g2_tiehi _19227__458 (.L_HI(net458));
 sg13g2_tiehi _19226__459 (.L_HI(net459));
 sg13g2_tiehi _19225__460 (.L_HI(net460));
 sg13g2_tiehi _19224__461 (.L_HI(net461));
 sg13g2_tiehi _19223__462 (.L_HI(net462));
 sg13g2_tiehi _19222__463 (.L_HI(net463));
 sg13g2_tiehi _19221__464 (.L_HI(net464));
 sg13g2_tiehi _19220__465 (.L_HI(net465));
 sg13g2_tiehi _19219__466 (.L_HI(net466));
 sg13g2_tiehi _19218__467 (.L_HI(net467));
 sg13g2_tiehi _19217__468 (.L_HI(net468));
 sg13g2_tiehi _19216__469 (.L_HI(net469));
 sg13g2_tiehi _19215__470 (.L_HI(net470));
 sg13g2_tiehi _19214__471 (.L_HI(net471));
 sg13g2_tiehi _19213__472 (.L_HI(net472));
 sg13g2_tiehi _19212__473 (.L_HI(net473));
 sg13g2_tiehi _19211__474 (.L_HI(net474));
 sg13g2_tiehi _19210__475 (.L_HI(net475));
 sg13g2_tiehi _19209__476 (.L_HI(net476));
 sg13g2_tiehi _19208__477 (.L_HI(net477));
 sg13g2_tiehi _19207__478 (.L_HI(net478));
 sg13g2_tiehi _19206__479 (.L_HI(net479));
 sg13g2_tiehi _19205__480 (.L_HI(net480));
 sg13g2_tiehi _19204__481 (.L_HI(net481));
 sg13g2_tiehi _19203__482 (.L_HI(net482));
 sg13g2_tiehi _19202__483 (.L_HI(net483));
 sg13g2_tiehi _19201__484 (.L_HI(net484));
 sg13g2_tiehi _19200__485 (.L_HI(net485));
 sg13g2_tiehi _19199__486 (.L_HI(net486));
 sg13g2_tiehi _19198__487 (.L_HI(net487));
 sg13g2_tiehi _19197__488 (.L_HI(net488));
 sg13g2_tiehi _19196__489 (.L_HI(net489));
 sg13g2_tiehi _19195__490 (.L_HI(net490));
 sg13g2_tiehi _19194__491 (.L_HI(net491));
 sg13g2_tiehi _19193__492 (.L_HI(net492));
 sg13g2_tiehi _19192__493 (.L_HI(net493));
 sg13g2_tiehi _19191__494 (.L_HI(net494));
 sg13g2_tiehi _19190__495 (.L_HI(net495));
 sg13g2_tiehi _19189__496 (.L_HI(net496));
 sg13g2_tiehi _19188__497 (.L_HI(net497));
 sg13g2_tiehi _19187__498 (.L_HI(net498));
 sg13g2_tiehi _19186__499 (.L_HI(net499));
 sg13g2_tiehi _19185__500 (.L_HI(net500));
 sg13g2_tiehi _19184__501 (.L_HI(net501));
 sg13g2_tiehi _19183__502 (.L_HI(net502));
 sg13g2_tiehi _19182__503 (.L_HI(net503));
 sg13g2_tiehi _19181__504 (.L_HI(net504));
 sg13g2_tiehi _19180__505 (.L_HI(net505));
 sg13g2_tiehi _19179__506 (.L_HI(net506));
 sg13g2_tiehi _19178__507 (.L_HI(net507));
 sg13g2_tiehi _19177__508 (.L_HI(net508));
 sg13g2_tiehi _19054__509 (.L_HI(net509));
 sg13g2_tiehi _19176__510 (.L_HI(net510));
 sg13g2_tiehi _20489__511 (.L_HI(net511));
 sg13g2_tiehi _19175__512 (.L_HI(net512));
 sg13g2_tiehi _20488__513 (.L_HI(net513));
 sg13g2_tiehi _19174__514 (.L_HI(net514));
 sg13g2_tiehi _20487__515 (.L_HI(net515));
 sg13g2_tiehi _19173__516 (.L_HI(net516));
 sg13g2_tiehi _20486__517 (.L_HI(net517));
 sg13g2_tiehi _19172__518 (.L_HI(net518));
 sg13g2_tiehi _20485__519 (.L_HI(net519));
 sg13g2_tiehi _19171__520 (.L_HI(net520));
 sg13g2_tiehi _20484__521 (.L_HI(net521));
 sg13g2_tiehi _19170__522 (.L_HI(net522));
 sg13g2_tiehi _20483__523 (.L_HI(net523));
 sg13g2_tiehi _19169__524 (.L_HI(net524));
 sg13g2_tiehi _20482__525 (.L_HI(net525));
 sg13g2_tiehi _19168__526 (.L_HI(net526));
 sg13g2_tiehi _19167__527 (.L_HI(net527));
 sg13g2_tiehi _19166__528 (.L_HI(net528));
 sg13g2_tiehi _19165__529 (.L_HI(net529));
 sg13g2_tiehi _19164__530 (.L_HI(net530));
 sg13g2_tiehi _19163__531 (.L_HI(net531));
 sg13g2_tiehi _19162__532 (.L_HI(net532));
 sg13g2_tiehi _19161__533 (.L_HI(net533));
 sg13g2_tiehi _19160__534 (.L_HI(net534));
 sg13g2_tiehi _19159__535 (.L_HI(net535));
 sg13g2_tiehi _19158__536 (.L_HI(net536));
 sg13g2_tiehi _19157__537 (.L_HI(net537));
 sg13g2_tiehi _19156__538 (.L_HI(net538));
 sg13g2_tiehi _19155__539 (.L_HI(net539));
 sg13g2_tiehi _19154__540 (.L_HI(net540));
 sg13g2_tiehi _19153__541 (.L_HI(net541));
 sg13g2_tiehi _19152__542 (.L_HI(net542));
 sg13g2_tiehi _19151__543 (.L_HI(net543));
 sg13g2_tiehi _19150__544 (.L_HI(net544));
 sg13g2_tiehi _19149__545 (.L_HI(net545));
 sg13g2_tiehi _19148__546 (.L_HI(net546));
 sg13g2_tiehi _19147__547 (.L_HI(net547));
 sg13g2_tiehi _19146__548 (.L_HI(net548));
 sg13g2_tiehi _19145__549 (.L_HI(net549));
 sg13g2_tiehi _19144__550 (.L_HI(net550));
 sg13g2_tiehi _19143__551 (.L_HI(net551));
 sg13g2_tiehi _19142__552 (.L_HI(net552));
 sg13g2_tiehi _19141__553 (.L_HI(net553));
 sg13g2_tiehi _19140__554 (.L_HI(net554));
 sg13g2_tiehi _19139__555 (.L_HI(net555));
 sg13g2_tiehi _19138__556 (.L_HI(net556));
 sg13g2_tiehi _19137__557 (.L_HI(net557));
 sg13g2_tiehi _19136__558 (.L_HI(net558));
 sg13g2_tiehi _19135__559 (.L_HI(net559));
 sg13g2_tiehi _19134__560 (.L_HI(net560));
 sg13g2_tiehi _19133__561 (.L_HI(net561));
 sg13g2_tiehi _19132__562 (.L_HI(net562));
 sg13g2_tiehi _19131__563 (.L_HI(net563));
 sg13g2_tiehi _19130__564 (.L_HI(net564));
 sg13g2_tiehi _19129__565 (.L_HI(net565));
 sg13g2_tiehi _19128__566 (.L_HI(net566));
 sg13g2_tiehi _19127__567 (.L_HI(net567));
 sg13g2_tiehi _19126__568 (.L_HI(net568));
 sg13g2_tiehi _19125__569 (.L_HI(net569));
 sg13g2_tiehi _19124__570 (.L_HI(net570));
 sg13g2_tiehi _19123__571 (.L_HI(net571));
 sg13g2_tiehi _19122__572 (.L_HI(net572));
 sg13g2_tiehi _19121__573 (.L_HI(net573));
 sg13g2_tiehi _19120__574 (.L_HI(net574));
 sg13g2_tiehi _19119__575 (.L_HI(net575));
 sg13g2_tiehi _19118__576 (.L_HI(net576));
 sg13g2_tiehi _19117__577 (.L_HI(net577));
 sg13g2_tiehi _19116__578 (.L_HI(net578));
 sg13g2_tiehi _19115__579 (.L_HI(net579));
 sg13g2_tiehi _19114__580 (.L_HI(net580));
 sg13g2_tiehi _19113__581 (.L_HI(net581));
 sg13g2_tiehi _19112__582 (.L_HI(net582));
 sg13g2_tiehi _19111__583 (.L_HI(net583));
 sg13g2_tiehi _19110__584 (.L_HI(net584));
 sg13g2_tiehi _19109__585 (.L_HI(net585));
 sg13g2_tiehi _19108__586 (.L_HI(net586));
 sg13g2_tiehi _19107__587 (.L_HI(net587));
 sg13g2_tiehi _19106__588 (.L_HI(net588));
 sg13g2_tiehi _19105__589 (.L_HI(net589));
 sg13g2_tiehi _19104__590 (.L_HI(net590));
 sg13g2_tiehi _19103__591 (.L_HI(net591));
 sg13g2_tiehi _19102__592 (.L_HI(net592));
 sg13g2_tiehi _19101__593 (.L_HI(net593));
 sg13g2_tiehi _19100__594 (.L_HI(net594));
 sg13g2_tiehi _19099__595 (.L_HI(net595));
 sg13g2_tiehi _19098__596 (.L_HI(net596));
 sg13g2_tiehi _19097__597 (.L_HI(net597));
 sg13g2_tiehi _19096__598 (.L_HI(net598));
 sg13g2_tiehi _19095__599 (.L_HI(net599));
 sg13g2_tiehi _19094__600 (.L_HI(net600));
 sg13g2_tiehi _19093__601 (.L_HI(net601));
 sg13g2_tiehi _19092__602 (.L_HI(net602));
 sg13g2_tiehi _19091__603 (.L_HI(net603));
 sg13g2_tiehi _19090__604 (.L_HI(net604));
 sg13g2_tiehi _19089__605 (.L_HI(net605));
 sg13g2_tiehi _19088__606 (.L_HI(net606));
 sg13g2_tiehi _19087__607 (.L_HI(net607));
 sg13g2_tiehi _19086__608 (.L_HI(net608));
 sg13g2_tiehi _19085__609 (.L_HI(net609));
 sg13g2_tiehi _19084__610 (.L_HI(net610));
 sg13g2_tiehi _19083__611 (.L_HI(net611));
 sg13g2_tiehi _19082__612 (.L_HI(net612));
 sg13g2_tiehi _19081__613 (.L_HI(net613));
 sg13g2_tiehi _19080__614 (.L_HI(net614));
 sg13g2_tiehi _19079__615 (.L_HI(net615));
 sg13g2_tiehi _19078__616 (.L_HI(net616));
 sg13g2_tiehi _19077__617 (.L_HI(net617));
 sg13g2_tiehi _19076__618 (.L_HI(net618));
 sg13g2_tiehi _19075__619 (.L_HI(net619));
 sg13g2_tiehi _19074__620 (.L_HI(net620));
 sg13g2_tiehi _19073__621 (.L_HI(net621));
 sg13g2_tiehi _19072__622 (.L_HI(net622));
 sg13g2_tiehi _19071__623 (.L_HI(net623));
 sg13g2_tiehi _19070__624 (.L_HI(net624));
 sg13g2_tiehi _19069__625 (.L_HI(net625));
 sg13g2_tiehi _19068__626 (.L_HI(net626));
 sg13g2_tiehi _19067__627 (.L_HI(net627));
 sg13g2_tiehi _19066__628 (.L_HI(net628));
 sg13g2_tiehi _19065__629 (.L_HI(net629));
 sg13g2_tiehi _19064__630 (.L_HI(net630));
 sg13g2_tiehi _19063__631 (.L_HI(net631));
 sg13g2_tiehi _19062__632 (.L_HI(net632));
 sg13g2_tiehi _19061__633 (.L_HI(net633));
 sg13g2_tiehi _19060__634 (.L_HI(net634));
 sg13g2_tiehi _19059__635 (.L_HI(net635));
 sg13g2_tiehi _19058__636 (.L_HI(net636));
 sg13g2_tiehi _19057__637 (.L_HI(net637));
 sg13g2_tiehi _19056__638 (.L_HI(net638));
 sg13g2_tiehi _19055__639 (.L_HI(net639));
 sg13g2_tiehi _19047__640 (.L_HI(net640));
 sg13g2_tiehi _19046__641 (.L_HI(net641));
 sg13g2_tiehi _19045__642 (.L_HI(net642));
 sg13g2_tiehi _19044__643 (.L_HI(net643));
 sg13g2_tiehi _19043__644 (.L_HI(net644));
 sg13g2_tiehi _19042__645 (.L_HI(net645));
 sg13g2_tiehi _19041__646 (.L_HI(net646));
 sg13g2_tiehi _19040__647 (.L_HI(net647));
 sg13g2_tiehi _19039__648 (.L_HI(net648));
 sg13g2_tiehi _19038__649 (.L_HI(net649));
 sg13g2_tiehi _19037__650 (.L_HI(net650));
 sg13g2_tiehi _19036__651 (.L_HI(net651));
 sg13g2_tiehi _19035__652 (.L_HI(net652));
 sg13g2_tiehi _19034__653 (.L_HI(net653));
 sg13g2_tiehi _19033__654 (.L_HI(net654));
 sg13g2_tiehi _19032__655 (.L_HI(net655));
 sg13g2_tiehi _19031__656 (.L_HI(net656));
 sg13g2_tiehi _19030__657 (.L_HI(net657));
 sg13g2_tiehi _19029__658 (.L_HI(net658));
 sg13g2_tiehi _19028__659 (.L_HI(net659));
 sg13g2_tiehi _19027__660 (.L_HI(net660));
 sg13g2_tiehi _19026__661 (.L_HI(net661));
 sg13g2_tiehi _19025__662 (.L_HI(net662));
 sg13g2_tiehi _19024__663 (.L_HI(net663));
 sg13g2_tiehi _19023__664 (.L_HI(net664));
 sg13g2_tiehi _19022__665 (.L_HI(net665));
 sg13g2_tiehi _19021__666 (.L_HI(net666));
 sg13g2_tiehi _19020__667 (.L_HI(net667));
 sg13g2_tiehi _19019__668 (.L_HI(net668));
 sg13g2_tiehi _19018__669 (.L_HI(net669));
 sg13g2_tiehi _19017__670 (.L_HI(net670));
 sg13g2_tiehi _19016__671 (.L_HI(net671));
 sg13g2_tiehi _19015__672 (.L_HI(net672));
 sg13g2_tiehi _19014__673 (.L_HI(net673));
 sg13g2_tiehi _19013__674 (.L_HI(net674));
 sg13g2_tiehi _19012__675 (.L_HI(net675));
 sg13g2_tiehi _19011__676 (.L_HI(net676));
 sg13g2_tiehi _19010__677 (.L_HI(net677));
 sg13g2_tiehi _19009__678 (.L_HI(net678));
 sg13g2_tiehi _19008__679 (.L_HI(net679));
 sg13g2_tiehi _19007__680 (.L_HI(net680));
 sg13g2_tiehi _19006__681 (.L_HI(net681));
 sg13g2_tiehi _19005__682 (.L_HI(net682));
 sg13g2_tiehi _19004__683 (.L_HI(net683));
 sg13g2_tiehi _19003__684 (.L_HI(net684));
 sg13g2_tiehi _19002__685 (.L_HI(net685));
 sg13g2_tiehi _19001__686 (.L_HI(net686));
 sg13g2_tiehi _19000__687 (.L_HI(net687));
 sg13g2_tiehi _18999__688 (.L_HI(net688));
 sg13g2_tiehi _18384__689 (.L_HI(net689));
 sg13g2_tiehi _19048__690 (.L_HI(net690));
 sg13g2_tiehi _19049__691 (.L_HI(net691));
 sg13g2_tiehi _19050__692 (.L_HI(net692));
 sg13g2_tiehi _19051__693 (.L_HI(net693));
 sg13g2_tiehi _19052__694 (.L_HI(net694));
 sg13g2_tiehi _19053__695 (.L_HI(net695));
 sg13g2_tiehi _18998__696 (.L_HI(net696));
 sg13g2_tiehi _18997__697 (.L_HI(net697));
 sg13g2_tiehi _18996__698 (.L_HI(net698));
 sg13g2_tiehi _18995__699 (.L_HI(net699));
 sg13g2_tiehi _18994__700 (.L_HI(net700));
 sg13g2_tiehi _18993__701 (.L_HI(net701));
 sg13g2_tiehi _18992__702 (.L_HI(net702));
 sg13g2_tiehi _18991__703 (.L_HI(net703));
 sg13g2_tiehi _18990__704 (.L_HI(net704));
 sg13g2_tiehi _18989__705 (.L_HI(net705));
 sg13g2_tiehi _18988__706 (.L_HI(net706));
 sg13g2_tiehi _18987__707 (.L_HI(net707));
 sg13g2_tiehi _18986__708 (.L_HI(net708));
 sg13g2_tiehi _18985__709 (.L_HI(net709));
 sg13g2_tiehi _18984__710 (.L_HI(net710));
 sg13g2_tiehi _18983__711 (.L_HI(net711));
 sg13g2_tiehi _18982__712 (.L_HI(net712));
 sg13g2_tiehi _18981__713 (.L_HI(net713));
 sg13g2_tiehi _18980__714 (.L_HI(net714));
 sg13g2_tiehi _18979__715 (.L_HI(net715));
 sg13g2_tiehi _18978__716 (.L_HI(net716));
 sg13g2_tiehi _18977__717 (.L_HI(net717));
 sg13g2_tiehi _18976__718 (.L_HI(net718));
 sg13g2_tiehi _18975__719 (.L_HI(net719));
 sg13g2_tiehi _18974__720 (.L_HI(net720));
 sg13g2_tiehi _18973__721 (.L_HI(net721));
 sg13g2_tiehi _18972__722 (.L_HI(net722));
 sg13g2_tiehi _18971__723 (.L_HI(net723));
 sg13g2_tiehi _18970__724 (.L_HI(net724));
 sg13g2_tiehi _18969__725 (.L_HI(net725));
 sg13g2_tiehi _20481__726 (.L_HI(net726));
 sg13g2_tiehi _18968__727 (.L_HI(net727));
 sg13g2_tiehi _20480__728 (.L_HI(net728));
 sg13g2_tiehi _18967__729 (.L_HI(net729));
 sg13g2_tiehi _20479__730 (.L_HI(net730));
 sg13g2_tiehi _18966__731 (.L_HI(net731));
 sg13g2_tiehi _20478__732 (.L_HI(net732));
 sg13g2_tiehi _18965__733 (.L_HI(net733));
 sg13g2_tiehi _20477__734 (.L_HI(net734));
 sg13g2_tiehi _18964__735 (.L_HI(net735));
 sg13g2_tiehi _20476__736 (.L_HI(net736));
 sg13g2_tiehi _18963__737 (.L_HI(net737));
 sg13g2_tiehi _20475__738 (.L_HI(net738));
 sg13g2_tiehi _18962__739 (.L_HI(net739));
 sg13g2_tiehi _20474__740 (.L_HI(net740));
 sg13g2_tiehi _18961__741 (.L_HI(net741));
 sg13g2_tiehi _20473__742 (.L_HI(net742));
 sg13g2_tiehi _18960__743 (.L_HI(net743));
 sg13g2_tiehi _20472__744 (.L_HI(net744));
 sg13g2_tiehi _18959__745 (.L_HI(net745));
 sg13g2_tiehi _20471__746 (.L_HI(net746));
 sg13g2_tiehi _18958__747 (.L_HI(net747));
 sg13g2_tiehi _20470__748 (.L_HI(net748));
 sg13g2_tiehi _18957__749 (.L_HI(net749));
 sg13g2_tiehi _20469__750 (.L_HI(net750));
 sg13g2_tiehi _18956__751 (.L_HI(net751));
 sg13g2_tiehi _20468__752 (.L_HI(net752));
 sg13g2_tiehi _18955__753 (.L_HI(net753));
 sg13g2_tiehi _20467__754 (.L_HI(net754));
 sg13g2_tiehi _18954__755 (.L_HI(net755));
 sg13g2_tiehi _20466__756 (.L_HI(net756));
 sg13g2_tiehi _18953__757 (.L_HI(net757));
 sg13g2_tiehi _18952__758 (.L_HI(net758));
 sg13g2_tiehi _18951__759 (.L_HI(net759));
 sg13g2_tiehi _18950__760 (.L_HI(net760));
 sg13g2_tiehi _18949__761 (.L_HI(net761));
 sg13g2_tiehi _18948__762 (.L_HI(net762));
 sg13g2_tiehi _18947__763 (.L_HI(net763));
 sg13g2_tiehi _18946__764 (.L_HI(net764));
 sg13g2_tiehi _18945__765 (.L_HI(net765));
 sg13g2_tiehi _20465__766 (.L_HI(net766));
 sg13g2_tiehi _18944__767 (.L_HI(net767));
 sg13g2_tiehi _20464__768 (.L_HI(net768));
 sg13g2_tiehi _18943__769 (.L_HI(net769));
 sg13g2_tiehi _20463__770 (.L_HI(net770));
 sg13g2_tiehi _18942__771 (.L_HI(net771));
 sg13g2_tiehi _20462__772 (.L_HI(net772));
 sg13g2_tiehi _18941__773 (.L_HI(net773));
 sg13g2_tiehi _20461__774 (.L_HI(net774));
 sg13g2_tiehi _18940__775 (.L_HI(net775));
 sg13g2_tiehi _20460__776 (.L_HI(net776));
 sg13g2_tiehi _18939__777 (.L_HI(net777));
 sg13g2_tiehi _20459__778 (.L_HI(net778));
 sg13g2_tiehi _18938__779 (.L_HI(net779));
 sg13g2_tiehi _20458__780 (.L_HI(net780));
 sg13g2_tiehi _18937__781 (.L_HI(net781));
 sg13g2_tiehi _20457__782 (.L_HI(net782));
 sg13g2_tiehi _18936__783 (.L_HI(net783));
 sg13g2_tiehi _20456__784 (.L_HI(net784));
 sg13g2_tiehi _18935__785 (.L_HI(net785));
 sg13g2_tiehi _20455__786 (.L_HI(net786));
 sg13g2_tiehi _18934__787 (.L_HI(net787));
 sg13g2_tiehi _20454__788 (.L_HI(net788));
 sg13g2_tiehi _18933__789 (.L_HI(net789));
 sg13g2_tiehi _20453__790 (.L_HI(net790));
 sg13g2_tiehi _18932__791 (.L_HI(net791));
 sg13g2_tiehi _20452__792 (.L_HI(net792));
 sg13g2_tiehi _18931__793 (.L_HI(net793));
 sg13g2_tiehi _20451__794 (.L_HI(net794));
 sg13g2_tiehi _18930__795 (.L_HI(net795));
 sg13g2_tiehi _20450__796 (.L_HI(net796));
 sg13g2_tiehi _18929__797 (.L_HI(net797));
 sg13g2_tiehi _20449__798 (.L_HI(net798));
 sg13g2_tiehi _18928__799 (.L_HI(net799));
 sg13g2_tiehi _20448__800 (.L_HI(net800));
 sg13g2_tiehi _18927__801 (.L_HI(net801));
 sg13g2_tiehi _20447__802 (.L_HI(net802));
 sg13g2_tiehi _18926__803 (.L_HI(net803));
 sg13g2_tiehi _20446__804 (.L_HI(net804));
 sg13g2_tiehi _18925__805 (.L_HI(net805));
 sg13g2_tiehi _20445__806 (.L_HI(net806));
 sg13g2_tiehi _18924__807 (.L_HI(net807));
 sg13g2_tiehi _20444__808 (.L_HI(net808));
 sg13g2_tiehi _18923__809 (.L_HI(net809));
 sg13g2_tiehi _20443__810 (.L_HI(net810));
 sg13g2_tiehi _18922__811 (.L_HI(net811));
 sg13g2_tiehi _20442__812 (.L_HI(net812));
 sg13g2_tiehi _18921__813 (.L_HI(net813));
 sg13g2_tiehi _20441__814 (.L_HI(net814));
 sg13g2_tiehi _18920__815 (.L_HI(net815));
 sg13g2_tiehi _20440__816 (.L_HI(net816));
 sg13g2_tiehi _18919__817 (.L_HI(net817));
 sg13g2_tiehi _20439__818 (.L_HI(net818));
 sg13g2_tiehi _18918__819 (.L_HI(net819));
 sg13g2_tiehi _20438__820 (.L_HI(net820));
 sg13g2_tiehi _18917__821 (.L_HI(net821));
 sg13g2_tiehi _20437__822 (.L_HI(net822));
 sg13g2_tiehi _18916__823 (.L_HI(net823));
 sg13g2_tiehi _20436__824 (.L_HI(net824));
 sg13g2_tiehi _18915__825 (.L_HI(net825));
 sg13g2_tiehi _20435__826 (.L_HI(net826));
 sg13g2_tiehi _18914__827 (.L_HI(net827));
 sg13g2_tiehi _20434__828 (.L_HI(net828));
 sg13g2_tiehi _18913__829 (.L_HI(net829));
 sg13g2_tiehi _20433__830 (.L_HI(net830));
 sg13g2_tiehi _18912__831 (.L_HI(net831));
 sg13g2_tiehi _20432__832 (.L_HI(net832));
 sg13g2_tiehi _18911__833 (.L_HI(net833));
 sg13g2_tiehi _20431__834 (.L_HI(net834));
 sg13g2_tiehi _18910__835 (.L_HI(net835));
 sg13g2_tiehi _20430__836 (.L_HI(net836));
 sg13g2_tiehi _18909__837 (.L_HI(net837));
 sg13g2_tiehi _20429__838 (.L_HI(net838));
 sg13g2_tiehi _18908__839 (.L_HI(net839));
 sg13g2_tiehi _20428__840 (.L_HI(net840));
 sg13g2_tiehi _18907__841 (.L_HI(net841));
 sg13g2_tiehi _20427__842 (.L_HI(net842));
 sg13g2_tiehi _18906__843 (.L_HI(net843));
 sg13g2_tiehi _20426__844 (.L_HI(net844));
 sg13g2_tiehi _18905__845 (.L_HI(net845));
 sg13g2_tiehi _18904__846 (.L_HI(net846));
 sg13g2_tiehi _18903__847 (.L_HI(net847));
 sg13g2_tiehi _18902__848 (.L_HI(net848));
 sg13g2_tiehi _18901__849 (.L_HI(net849));
 sg13g2_tiehi _18900__850 (.L_HI(net850));
 sg13g2_tiehi _18899__851 (.L_HI(net851));
 sg13g2_tiehi _18898__852 (.L_HI(net852));
 sg13g2_tiehi _18897__853 (.L_HI(net853));
 sg13g2_tiehi _18896__854 (.L_HI(net854));
 sg13g2_tiehi _18895__855 (.L_HI(net855));
 sg13g2_tiehi _18894__856 (.L_HI(net856));
 sg13g2_tiehi _18893__857 (.L_HI(net857));
 sg13g2_tiehi _18892__858 (.L_HI(net858));
 sg13g2_tiehi _18891__859 (.L_HI(net859));
 sg13g2_tiehi _18890__860 (.L_HI(net860));
 sg13g2_tiehi _18889__861 (.L_HI(net861));
 sg13g2_tiehi _18888__862 (.L_HI(net862));
 sg13g2_tiehi _18887__863 (.L_HI(net863));
 sg13g2_tiehi _18886__864 (.L_HI(net864));
 sg13g2_tiehi _18885__865 (.L_HI(net865));
 sg13g2_tiehi _18884__866 (.L_HI(net866));
 sg13g2_tiehi _18883__867 (.L_HI(net867));
 sg13g2_tiehi _18882__868 (.L_HI(net868));
 sg13g2_tiehi _18881__869 (.L_HI(net869));
 sg13g2_tiehi _18880__870 (.L_HI(net870));
 sg13g2_tiehi _18879__871 (.L_HI(net871));
 sg13g2_tiehi _18878__872 (.L_HI(net872));
 sg13g2_tiehi _18877__873 (.L_HI(net873));
 sg13g2_tiehi _18876__874 (.L_HI(net874));
 sg13g2_tiehi _18875__875 (.L_HI(net875));
 sg13g2_tiehi _18874__876 (.L_HI(net876));
 sg13g2_tiehi _18873__877 (.L_HI(net877));
 sg13g2_tiehi _18872__878 (.L_HI(net878));
 sg13g2_tiehi _18871__879 (.L_HI(net879));
 sg13g2_tiehi _18870__880 (.L_HI(net880));
 sg13g2_tiehi _18869__881 (.L_HI(net881));
 sg13g2_tiehi _18868__882 (.L_HI(net882));
 sg13g2_tiehi _18867__883 (.L_HI(net883));
 sg13g2_tiehi _18866__884 (.L_HI(net884));
 sg13g2_tiehi _18865__885 (.L_HI(net885));
 sg13g2_tiehi _18864__886 (.L_HI(net886));
 sg13g2_tiehi _18863__887 (.L_HI(net887));
 sg13g2_tiehi _18862__888 (.L_HI(net888));
 sg13g2_tiehi _18861__889 (.L_HI(net889));
 sg13g2_tiehi _18860__890 (.L_HI(net890));
 sg13g2_tiehi _18859__891 (.L_HI(net891));
 sg13g2_tiehi _18858__892 (.L_HI(net892));
 sg13g2_tiehi _18857__893 (.L_HI(net893));
 sg13g2_tiehi _18856__894 (.L_HI(net894));
 sg13g2_tiehi _18855__895 (.L_HI(net895));
 sg13g2_tiehi _18854__896 (.L_HI(net896));
 sg13g2_tiehi _18853__897 (.L_HI(net897));
 sg13g2_tiehi _18852__898 (.L_HI(net898));
 sg13g2_tiehi _18851__899 (.L_HI(net899));
 sg13g2_tiehi _18850__900 (.L_HI(net900));
 sg13g2_tiehi _18849__901 (.L_HI(net901));
 sg13g2_tiehi _18848__902 (.L_HI(net902));
 sg13g2_tiehi _18847__903 (.L_HI(net903));
 sg13g2_tiehi _18846__904 (.L_HI(net904));
 sg13g2_tiehi _18845__905 (.L_HI(net905));
 sg13g2_tiehi _18844__906 (.L_HI(net906));
 sg13g2_tiehi _18843__907 (.L_HI(net907));
 sg13g2_tiehi _18842__908 (.L_HI(net908));
 sg13g2_tiehi _18841__909 (.L_HI(net909));
 sg13g2_tiehi _18840__910 (.L_HI(net910));
 sg13g2_tiehi _18839__911 (.L_HI(net911));
 sg13g2_tiehi _18838__912 (.L_HI(net912));
 sg13g2_tiehi _18837__913 (.L_HI(net913));
 sg13g2_tiehi _18836__914 (.L_HI(net914));
 sg13g2_tiehi _18835__915 (.L_HI(net915));
 sg13g2_tiehi _18834__916 (.L_HI(net916));
 sg13g2_tiehi _18833__917 (.L_HI(net917));
 sg13g2_tiehi _18832__918 (.L_HI(net918));
 sg13g2_tiehi _18831__919 (.L_HI(net919));
 sg13g2_tiehi _18830__920 (.L_HI(net920));
 sg13g2_tiehi _18829__921 (.L_HI(net921));
 sg13g2_tiehi _18828__922 (.L_HI(net922));
 sg13g2_tiehi _18827__923 (.L_HI(net923));
 sg13g2_tiehi _18826__924 (.L_HI(net924));
 sg13g2_tiehi _18825__925 (.L_HI(net925));
 sg13g2_tiehi _18824__926 (.L_HI(net926));
 sg13g2_tiehi _18823__927 (.L_HI(net927));
 sg13g2_tiehi _18822__928 (.L_HI(net928));
 sg13g2_tiehi _18821__929 (.L_HI(net929));
 sg13g2_tiehi _18820__930 (.L_HI(net930));
 sg13g2_tiehi _18819__931 (.L_HI(net931));
 sg13g2_tiehi _18818__932 (.L_HI(net932));
 sg13g2_tiehi _18817__933 (.L_HI(net933));
 sg13g2_tiehi _18816__934 (.L_HI(net934));
 sg13g2_tiehi _18815__935 (.L_HI(net935));
 sg13g2_tiehi _18814__936 (.L_HI(net936));
 sg13g2_tiehi _18813__937 (.L_HI(net937));
 sg13g2_tiehi _18812__938 (.L_HI(net938));
 sg13g2_tiehi _18811__939 (.L_HI(net939));
 sg13g2_tiehi _18810__940 (.L_HI(net940));
 sg13g2_tiehi _18809__941 (.L_HI(net941));
 sg13g2_tiehi _18808__942 (.L_HI(net942));
 sg13g2_tiehi _18807__943 (.L_HI(net943));
 sg13g2_tiehi _18806__944 (.L_HI(net944));
 sg13g2_tiehi _18805__945 (.L_HI(net945));
 sg13g2_tiehi _18804__946 (.L_HI(net946));
 sg13g2_tiehi _18803__947 (.L_HI(net947));
 sg13g2_tiehi _18802__948 (.L_HI(net948));
 sg13g2_tiehi _18801__949 (.L_HI(net949));
 sg13g2_tiehi _18800__950 (.L_HI(net950));
 sg13g2_tiehi _18799__951 (.L_HI(net951));
 sg13g2_tiehi _18798__952 (.L_HI(net952));
 sg13g2_tiehi _18797__953 (.L_HI(net953));
 sg13g2_tiehi _18796__954 (.L_HI(net954));
 sg13g2_tiehi _18795__955 (.L_HI(net955));
 sg13g2_tiehi _18794__956 (.L_HI(net956));
 sg13g2_tiehi _18793__957 (.L_HI(net957));
 sg13g2_tiehi _18792__958 (.L_HI(net958));
 sg13g2_tiehi _18791__959 (.L_HI(net959));
 sg13g2_tiehi _18790__960 (.L_HI(net960));
 sg13g2_tiehi _18789__961 (.L_HI(net961));
 sg13g2_tiehi _18788__962 (.L_HI(net962));
 sg13g2_tiehi _18787__963 (.L_HI(net963));
 sg13g2_tiehi _18786__964 (.L_HI(net964));
 sg13g2_tiehi _18785__965 (.L_HI(net965));
 sg13g2_tiehi _18784__966 (.L_HI(net966));
 sg13g2_tiehi _18783__967 (.L_HI(net967));
 sg13g2_tiehi _18782__968 (.L_HI(net968));
 sg13g2_tiehi _18781__969 (.L_HI(net969));
 sg13g2_tiehi _18780__970 (.L_HI(net970));
 sg13g2_tiehi _18779__971 (.L_HI(net971));
 sg13g2_tiehi _18778__972 (.L_HI(net972));
 sg13g2_tiehi _18777__973 (.L_HI(net973));
 sg13g2_tiehi _18776__974 (.L_HI(net974));
 sg13g2_tiehi _18775__975 (.L_HI(net975));
 sg13g2_tiehi _18774__976 (.L_HI(net976));
 sg13g2_tiehi _18773__977 (.L_HI(net977));
 sg13g2_tiehi _18772__978 (.L_HI(net978));
 sg13g2_tiehi _18771__979 (.L_HI(net979));
 sg13g2_tiehi _18770__980 (.L_HI(net980));
 sg13g2_tiehi _18769__981 (.L_HI(net981));
 sg13g2_tiehi _18768__982 (.L_HI(net982));
 sg13g2_tiehi _18767__983 (.L_HI(net983));
 sg13g2_tiehi _18766__984 (.L_HI(net984));
 sg13g2_tiehi _18765__985 (.L_HI(net985));
 sg13g2_tiehi _18764__986 (.L_HI(net986));
 sg13g2_tiehi _18763__987 (.L_HI(net987));
 sg13g2_tiehi _18762__988 (.L_HI(net988));
 sg13g2_tiehi _18761__989 (.L_HI(net989));
 sg13g2_tiehi _18760__990 (.L_HI(net990));
 sg13g2_tiehi _18759__991 (.L_HI(net991));
 sg13g2_tiehi _18758__992 (.L_HI(net992));
 sg13g2_tiehi _18757__993 (.L_HI(net993));
 sg13g2_tiehi _18756__994 (.L_HI(net994));
 sg13g2_tiehi _18755__995 (.L_HI(net995));
 sg13g2_tiehi _18754__996 (.L_HI(net996));
 sg13g2_tiehi _18753__997 (.L_HI(net997));
 sg13g2_tiehi _18752__998 (.L_HI(net998));
 sg13g2_tiehi _18751__999 (.L_HI(net999));
 sg13g2_tiehi _18750__1000 (.L_HI(net1000));
 sg13g2_tiehi _18749__1001 (.L_HI(net1001));
 sg13g2_tiehi _18748__1002 (.L_HI(net1002));
 sg13g2_tiehi _18747__1003 (.L_HI(net1003));
 sg13g2_tiehi _18746__1004 (.L_HI(net1004));
 sg13g2_tiehi _18745__1005 (.L_HI(net1005));
 sg13g2_tiehi _18744__1006 (.L_HI(net1006));
 sg13g2_tiehi _18743__1007 (.L_HI(net1007));
 sg13g2_tiehi _18742__1008 (.L_HI(net1008));
 sg13g2_tiehi _18741__1009 (.L_HI(net1009));
 sg13g2_tiehi _18740__1010 (.L_HI(net1010));
 sg13g2_tiehi _18739__1011 (.L_HI(net1011));
 sg13g2_tiehi _18738__1012 (.L_HI(net1012));
 sg13g2_tiehi _18737__1013 (.L_HI(net1013));
 sg13g2_tiehi _18736__1014 (.L_HI(net1014));
 sg13g2_tiehi _18735__1015 (.L_HI(net1015));
 sg13g2_tiehi _18734__1016 (.L_HI(net1016));
 sg13g2_tiehi _18733__1017 (.L_HI(net1017));
 sg13g2_tiehi _18732__1018 (.L_HI(net1018));
 sg13g2_tiehi _18731__1019 (.L_HI(net1019));
 sg13g2_tiehi _18730__1020 (.L_HI(net1020));
 sg13g2_tiehi _18729__1021 (.L_HI(net1021));
 sg13g2_tiehi _18728__1022 (.L_HI(net1022));
 sg13g2_tiehi _18727__1023 (.L_HI(net1023));
 sg13g2_tiehi _18726__1024 (.L_HI(net1024));
 sg13g2_tiehi _18725__1025 (.L_HI(net1025));
 sg13g2_tiehi _18724__1026 (.L_HI(net1026));
 sg13g2_tiehi _18723__1027 (.L_HI(net1027));
 sg13g2_tiehi _18722__1028 (.L_HI(net1028));
 sg13g2_tiehi _18721__1029 (.L_HI(net1029));
 sg13g2_tiehi _18720__1030 (.L_HI(net1030));
 sg13g2_tiehi _18719__1031 (.L_HI(net1031));
 sg13g2_tiehi _18718__1032 (.L_HI(net1032));
 sg13g2_tiehi _18717__1033 (.L_HI(net1033));
 sg13g2_tiehi _18716__1034 (.L_HI(net1034));
 sg13g2_tiehi _18715__1035 (.L_HI(net1035));
 sg13g2_tiehi _18714__1036 (.L_HI(net1036));
 sg13g2_tiehi _18713__1037 (.L_HI(net1037));
 sg13g2_tiehi _18712__1038 (.L_HI(net1038));
 sg13g2_tiehi _18711__1039 (.L_HI(net1039));
 sg13g2_tiehi _18710__1040 (.L_HI(net1040));
 sg13g2_tiehi _18709__1041 (.L_HI(net1041));
 sg13g2_tiehi _18708__1042 (.L_HI(net1042));
 sg13g2_tiehi _18707__1043 (.L_HI(net1043));
 sg13g2_tiehi _18706__1044 (.L_HI(net1044));
 sg13g2_tiehi _18705__1045 (.L_HI(net1045));
 sg13g2_tiehi _18704__1046 (.L_HI(net1046));
 sg13g2_tiehi _18703__1047 (.L_HI(net1047));
 sg13g2_tiehi _18702__1048 (.L_HI(net1048));
 sg13g2_tiehi _18701__1049 (.L_HI(net1049));
 sg13g2_tiehi _18700__1050 (.L_HI(net1050));
 sg13g2_tiehi _18699__1051 (.L_HI(net1051));
 sg13g2_tiehi _18698__1052 (.L_HI(net1052));
 sg13g2_tiehi _18697__1053 (.L_HI(net1053));
 sg13g2_tiehi _18696__1054 (.L_HI(net1054));
 sg13g2_tiehi _18695__1055 (.L_HI(net1055));
 sg13g2_tiehi _18694__1056 (.L_HI(net1056));
 sg13g2_tiehi _18693__1057 (.L_HI(net1057));
 sg13g2_tiehi _18692__1058 (.L_HI(net1058));
 sg13g2_tiehi _18691__1059 (.L_HI(net1059));
 sg13g2_tiehi _18690__1060 (.L_HI(net1060));
 sg13g2_tiehi _18689__1061 (.L_HI(net1061));
 sg13g2_tiehi _18688__1062 (.L_HI(net1062));
 sg13g2_tiehi _18687__1063 (.L_HI(net1063));
 sg13g2_tiehi _18686__1064 (.L_HI(net1064));
 sg13g2_tiehi _18685__1065 (.L_HI(net1065));
 sg13g2_tiehi _18684__1066 (.L_HI(net1066));
 sg13g2_tiehi _18683__1067 (.L_HI(net1067));
 sg13g2_tiehi _18682__1068 (.L_HI(net1068));
 sg13g2_tiehi _18681__1069 (.L_HI(net1069));
 sg13g2_tiehi _18680__1070 (.L_HI(net1070));
 sg13g2_tiehi _18679__1071 (.L_HI(net1071));
 sg13g2_tiehi _18678__1072 (.L_HI(net1072));
 sg13g2_tiehi _18677__1073 (.L_HI(net1073));
 sg13g2_tiehi _18676__1074 (.L_HI(net1074));
 sg13g2_tiehi _18675__1075 (.L_HI(net1075));
 sg13g2_tiehi _18674__1076 (.L_HI(net1076));
 sg13g2_tiehi _18673__1077 (.L_HI(net1077));
 sg13g2_tiehi _18672__1078 (.L_HI(net1078));
 sg13g2_tiehi _18671__1079 (.L_HI(net1079));
 sg13g2_tiehi _18670__1080 (.L_HI(net1080));
 sg13g2_tiehi _18669__1081 (.L_HI(net1081));
 sg13g2_tiehi _18668__1082 (.L_HI(net1082));
 sg13g2_tiehi _18667__1083 (.L_HI(net1083));
 sg13g2_tiehi _18666__1084 (.L_HI(net1084));
 sg13g2_tiehi _18665__1085 (.L_HI(net1085));
 sg13g2_tiehi _18664__1086 (.L_HI(net1086));
 sg13g2_tiehi _18663__1087 (.L_HI(net1087));
 sg13g2_tiehi _18662__1088 (.L_HI(net1088));
 sg13g2_tiehi _18661__1089 (.L_HI(net1089));
 sg13g2_tiehi _18660__1090 (.L_HI(net1090));
 sg13g2_tiehi _18659__1091 (.L_HI(net1091));
 sg13g2_tiehi _18658__1092 (.L_HI(net1092));
 sg13g2_tiehi _18657__1093 (.L_HI(net1093));
 sg13g2_tiehi _18656__1094 (.L_HI(net1094));
 sg13g2_tiehi _18655__1095 (.L_HI(net1095));
 sg13g2_tiehi _18654__1096 (.L_HI(net1096));
 sg13g2_tiehi _18653__1097 (.L_HI(net1097));
 sg13g2_tiehi _18652__1098 (.L_HI(net1098));
 sg13g2_tiehi _18651__1099 (.L_HI(net1099));
 sg13g2_tiehi _18650__1100 (.L_HI(net1100));
 sg13g2_tiehi _18649__1101 (.L_HI(net1101));
 sg13g2_tiehi _18648__1102 (.L_HI(net1102));
 sg13g2_tiehi _18647__1103 (.L_HI(net1103));
 sg13g2_tiehi _18646__1104 (.L_HI(net1104));
 sg13g2_tiehi _18645__1105 (.L_HI(net1105));
 sg13g2_tiehi _18644__1106 (.L_HI(net1106));
 sg13g2_tiehi _18643__1107 (.L_HI(net1107));
 sg13g2_tiehi _18642__1108 (.L_HI(net1108));
 sg13g2_tiehi _18641__1109 (.L_HI(net1109));
 sg13g2_tiehi _18640__1110 (.L_HI(net1110));
 sg13g2_tiehi _18639__1111 (.L_HI(net1111));
 sg13g2_tiehi _18638__1112 (.L_HI(net1112));
 sg13g2_tiehi _18637__1113 (.L_HI(net1113));
 sg13g2_tiehi _18636__1114 (.L_HI(net1114));
 sg13g2_tiehi _18635__1115 (.L_HI(net1115));
 sg13g2_tiehi _18634__1116 (.L_HI(net1116));
 sg13g2_tiehi _18633__1117 (.L_HI(net1117));
 sg13g2_tiehi _18632__1118 (.L_HI(net1118));
 sg13g2_tiehi _18631__1119 (.L_HI(net1119));
 sg13g2_tiehi _18630__1120 (.L_HI(net1120));
 sg13g2_tiehi _18629__1121 (.L_HI(net1121));
 sg13g2_tiehi _18628__1122 (.L_HI(net1122));
 sg13g2_tiehi _18627__1123 (.L_HI(net1123));
 sg13g2_tiehi _18626__1124 (.L_HI(net1124));
 sg13g2_tiehi _18625__1125 (.L_HI(net1125));
 sg13g2_tiehi _18624__1126 (.L_HI(net1126));
 sg13g2_tiehi _18623__1127 (.L_HI(net1127));
 sg13g2_tiehi _18622__1128 (.L_HI(net1128));
 sg13g2_tiehi _18621__1129 (.L_HI(net1129));
 sg13g2_tiehi _18620__1130 (.L_HI(net1130));
 sg13g2_tiehi _18619__1131 (.L_HI(net1131));
 sg13g2_tiehi _18618__1132 (.L_HI(net1132));
 sg13g2_tiehi _18617__1133 (.L_HI(net1133));
 sg13g2_tiehi _18616__1134 (.L_HI(net1134));
 sg13g2_tiehi _18615__1135 (.L_HI(net1135));
 sg13g2_tiehi _18614__1136 (.L_HI(net1136));
 sg13g2_tiehi _18613__1137 (.L_HI(net1137));
 sg13g2_tiehi _18612__1138 (.L_HI(net1138));
 sg13g2_tiehi _18611__1139 (.L_HI(net1139));
 sg13g2_tiehi _18610__1140 (.L_HI(net1140));
 sg13g2_tiehi _18609__1141 (.L_HI(net1141));
 sg13g2_tiehi _18608__1142 (.L_HI(net1142));
 sg13g2_tiehi _18607__1143 (.L_HI(net1143));
 sg13g2_tiehi _18606__1144 (.L_HI(net1144));
 sg13g2_tiehi _18605__1145 (.L_HI(net1145));
 sg13g2_tiehi _18604__1146 (.L_HI(net1146));
 sg13g2_tiehi _18603__1147 (.L_HI(net1147));
 sg13g2_tiehi _18602__1148 (.L_HI(net1148));
 sg13g2_tiehi _18601__1149 (.L_HI(net1149));
 sg13g2_tiehi _18600__1150 (.L_HI(net1150));
 sg13g2_tiehi _18599__1151 (.L_HI(net1151));
 sg13g2_tiehi _18598__1152 (.L_HI(net1152));
 sg13g2_tiehi _18597__1153 (.L_HI(net1153));
 sg13g2_tiehi _18596__1154 (.L_HI(net1154));
 sg13g2_tiehi _18595__1155 (.L_HI(net1155));
 sg13g2_tiehi _18594__1156 (.L_HI(net1156));
 sg13g2_tiehi _18593__1157 (.L_HI(net1157));
 sg13g2_tiehi _18592__1158 (.L_HI(net1158));
 sg13g2_tiehi _18591__1159 (.L_HI(net1159));
 sg13g2_tiehi _18590__1160 (.L_HI(net1160));
 sg13g2_tiehi _18589__1161 (.L_HI(net1161));
 sg13g2_tiehi _18588__1162 (.L_HI(net1162));
 sg13g2_tiehi _18587__1163 (.L_HI(net1163));
 sg13g2_tiehi _18586__1164 (.L_HI(net1164));
 sg13g2_tiehi _18585__1165 (.L_HI(net1165));
 sg13g2_tiehi _18584__1166 (.L_HI(net1166));
 sg13g2_tiehi _18583__1167 (.L_HI(net1167));
 sg13g2_tiehi _18582__1168 (.L_HI(net1168));
 sg13g2_tiehi _18581__1169 (.L_HI(net1169));
 sg13g2_tiehi _18580__1170 (.L_HI(net1170));
 sg13g2_tiehi _18579__1171 (.L_HI(net1171));
 sg13g2_tiehi _18578__1172 (.L_HI(net1172));
 sg13g2_tiehi _18577__1173 (.L_HI(net1173));
 sg13g2_tiehi _18576__1174 (.L_HI(net1174));
 sg13g2_tiehi _18575__1175 (.L_HI(net1175));
 sg13g2_tiehi _18574__1176 (.L_HI(net1176));
 sg13g2_tiehi _18573__1177 (.L_HI(net1177));
 sg13g2_tiehi _18572__1178 (.L_HI(net1178));
 sg13g2_tiehi _18571__1179 (.L_HI(net1179));
 sg13g2_tiehi _18570__1180 (.L_HI(net1180));
 sg13g2_tiehi _18569__1181 (.L_HI(net1181));
 sg13g2_tiehi _18568__1182 (.L_HI(net1182));
 sg13g2_tiehi _18567__1183 (.L_HI(net1183));
 sg13g2_tiehi _18566__1184 (.L_HI(net1184));
 sg13g2_tiehi _18565__1185 (.L_HI(net1185));
 sg13g2_tiehi _18564__1186 (.L_HI(net1186));
 sg13g2_tiehi _18563__1187 (.L_HI(net1187));
 sg13g2_tiehi _18562__1188 (.L_HI(net1188));
 sg13g2_tiehi _18561__1189 (.L_HI(net1189));
 sg13g2_tiehi _18560__1190 (.L_HI(net1190));
 sg13g2_tiehi _18559__1191 (.L_HI(net1191));
 sg13g2_tiehi _18558__1192 (.L_HI(net1192));
 sg13g2_tiehi _18557__1193 (.L_HI(net1193));
 sg13g2_tiehi _18556__1194 (.L_HI(net1194));
 sg13g2_tiehi _18555__1195 (.L_HI(net1195));
 sg13g2_tiehi _18554__1196 (.L_HI(net1196));
 sg13g2_tiehi _18553__1197 (.L_HI(net1197));
 sg13g2_tiehi _18552__1198 (.L_HI(net1198));
 sg13g2_tiehi _18551__1199 (.L_HI(net1199));
 sg13g2_tiehi _18550__1200 (.L_HI(net1200));
 sg13g2_tiehi _18549__1201 (.L_HI(net1201));
 sg13g2_tiehi _18548__1202 (.L_HI(net1202));
 sg13g2_tiehi _18547__1203 (.L_HI(net1203));
 sg13g2_tiehi _18546__1204 (.L_HI(net1204));
 sg13g2_tiehi _18545__1205 (.L_HI(net1205));
 sg13g2_tiehi _18544__1206 (.L_HI(net1206));
 sg13g2_tiehi _18543__1207 (.L_HI(net1207));
 sg13g2_tiehi _18542__1208 (.L_HI(net1208));
 sg13g2_tiehi _18541__1209 (.L_HI(net1209));
 sg13g2_tiehi _18540__1210 (.L_HI(net1210));
 sg13g2_tiehi _18539__1211 (.L_HI(net1211));
 sg13g2_tiehi _18538__1212 (.L_HI(net1212));
 sg13g2_tiehi _18537__1213 (.L_HI(net1213));
 sg13g2_tiehi _18536__1214 (.L_HI(net1214));
 sg13g2_tiehi _18535__1215 (.L_HI(net1215));
 sg13g2_tiehi _18534__1216 (.L_HI(net1216));
 sg13g2_tiehi _18533__1217 (.L_HI(net1217));
 sg13g2_tiehi _18532__1218 (.L_HI(net1218));
 sg13g2_tiehi _18531__1219 (.L_HI(net1219));
 sg13g2_tiehi _18530__1220 (.L_HI(net1220));
 sg13g2_tiehi _18529__1221 (.L_HI(net1221));
 sg13g2_tiehi _18528__1222 (.L_HI(net1222));
 sg13g2_tiehi _18527__1223 (.L_HI(net1223));
 sg13g2_tiehi _18526__1224 (.L_HI(net1224));
 sg13g2_tiehi _18525__1225 (.L_HI(net1225));
 sg13g2_tiehi _18524__1226 (.L_HI(net1226));
 sg13g2_tiehi _18523__1227 (.L_HI(net1227));
 sg13g2_tiehi _18522__1228 (.L_HI(net1228));
 sg13g2_tiehi _18521__1229 (.L_HI(net1229));
 sg13g2_tiehi _18520__1230 (.L_HI(net1230));
 sg13g2_tiehi _18519__1231 (.L_HI(net1231));
 sg13g2_tiehi _18518__1232 (.L_HI(net1232));
 sg13g2_tiehi _18517__1233 (.L_HI(net1233));
 sg13g2_tiehi _18516__1234 (.L_HI(net1234));
 sg13g2_tiehi _18515__1235 (.L_HI(net1235));
 sg13g2_tiehi _18514__1236 (.L_HI(net1236));
 sg13g2_tiehi _18513__1237 (.L_HI(net1237));
 sg13g2_tiehi _18512__1238 (.L_HI(net1238));
 sg13g2_tiehi _18511__1239 (.L_HI(net1239));
 sg13g2_tiehi _18510__1240 (.L_HI(net1240));
 sg13g2_tiehi _18509__1241 (.L_HI(net1241));
 sg13g2_tiehi _18508__1242 (.L_HI(net1242));
 sg13g2_tiehi _18507__1243 (.L_HI(net1243));
 sg13g2_tiehi _18506__1244 (.L_HI(net1244));
 sg13g2_tiehi _18505__1245 (.L_HI(net1245));
 sg13g2_tiehi _18504__1246 (.L_HI(net1246));
 sg13g2_tiehi _18503__1247 (.L_HI(net1247));
 sg13g2_tiehi _18502__1248 (.L_HI(net1248));
 sg13g2_tiehi _18501__1249 (.L_HI(net1249));
 sg13g2_tiehi _18500__1250 (.L_HI(net1250));
 sg13g2_tiehi _18499__1251 (.L_HI(net1251));
 sg13g2_tiehi _18498__1252 (.L_HI(net1252));
 sg13g2_tiehi _18497__1253 (.L_HI(net1253));
 sg13g2_tiehi _18496__1254 (.L_HI(net1254));
 sg13g2_tiehi _18495__1255 (.L_HI(net1255));
 sg13g2_tiehi _18494__1256 (.L_HI(net1256));
 sg13g2_tiehi _18493__1257 (.L_HI(net1257));
 sg13g2_tiehi _18492__1258 (.L_HI(net1258));
 sg13g2_tiehi _18491__1259 (.L_HI(net1259));
 sg13g2_tiehi _18490__1260 (.L_HI(net1260));
 sg13g2_tiehi _18489__1261 (.L_HI(net1261));
 sg13g2_tiehi _18488__1262 (.L_HI(net1262));
 sg13g2_tiehi _18487__1263 (.L_HI(net1263));
 sg13g2_tiehi _18486__1264 (.L_HI(net1264));
 sg13g2_tiehi _18485__1265 (.L_HI(net1265));
 sg13g2_tiehi _18484__1266 (.L_HI(net1266));
 sg13g2_tiehi _18483__1267 (.L_HI(net1267));
 sg13g2_tiehi _18482__1268 (.L_HI(net1268));
 sg13g2_tiehi _18481__1269 (.L_HI(net1269));
 sg13g2_tiehi _18480__1270 (.L_HI(net1270));
 sg13g2_tiehi _18479__1271 (.L_HI(net1271));
 sg13g2_tiehi _18478__1272 (.L_HI(net1272));
 sg13g2_tiehi _18477__1273 (.L_HI(net1273));
 sg13g2_tiehi _18476__1274 (.L_HI(net1274));
 sg13g2_tiehi _18475__1275 (.L_HI(net1275));
 sg13g2_tiehi _18474__1276 (.L_HI(net1276));
 sg13g2_tiehi _18473__1277 (.L_HI(net1277));
 sg13g2_tiehi _18472__1278 (.L_HI(net1278));
 sg13g2_tiehi _18471__1279 (.L_HI(net1279));
 sg13g2_tiehi _18470__1280 (.L_HI(net1280));
 sg13g2_tiehi _18469__1281 (.L_HI(net1281));
 sg13g2_tiehi _18468__1282 (.L_HI(net1282));
 sg13g2_tiehi _18467__1283 (.L_HI(net1283));
 sg13g2_tiehi _18466__1284 (.L_HI(net1284));
 sg13g2_tiehi _18465__1285 (.L_HI(net1285));
 sg13g2_tiehi _18464__1286 (.L_HI(net1286));
 sg13g2_tiehi _18463__1287 (.L_HI(net1287));
 sg13g2_tiehi _18462__1288 (.L_HI(net1288));
 sg13g2_tiehi _18461__1289 (.L_HI(net1289));
 sg13g2_tiehi _18460__1290 (.L_HI(net1290));
 sg13g2_tiehi _18459__1291 (.L_HI(net1291));
 sg13g2_tiehi _18458__1292 (.L_HI(net1292));
 sg13g2_tiehi _18457__1293 (.L_HI(net1293));
 sg13g2_tiehi _18456__1294 (.L_HI(net1294));
 sg13g2_tiehi _18455__1295 (.L_HI(net1295));
 sg13g2_tiehi _18454__1296 (.L_HI(net1296));
 sg13g2_tiehi _18453__1297 (.L_HI(net1297));
 sg13g2_tiehi _18452__1298 (.L_HI(net1298));
 sg13g2_tiehi _18451__1299 (.L_HI(net1299));
 sg13g2_tiehi _18450__1300 (.L_HI(net1300));
 sg13g2_tiehi _18449__1301 (.L_HI(net1301));
 sg13g2_tiehi _18448__1302 (.L_HI(net1302));
 sg13g2_tiehi _18447__1303 (.L_HI(net1303));
 sg13g2_tiehi _18446__1304 (.L_HI(net1304));
 sg13g2_tiehi _18445__1305 (.L_HI(net1305));
 sg13g2_tiehi _18444__1306 (.L_HI(net1306));
 sg13g2_tiehi _18443__1307 (.L_HI(net1307));
 sg13g2_tiehi _18442__1308 (.L_HI(net1308));
 sg13g2_tiehi _18441__1309 (.L_HI(net1309));
 sg13g2_tiehi _18440__1310 (.L_HI(net1310));
 sg13g2_tiehi _18439__1311 (.L_HI(net1311));
 sg13g2_tiehi _18438__1312 (.L_HI(net1312));
 sg13g2_tiehi _18437__1313 (.L_HI(net1313));
 sg13g2_tiehi _18436__1314 (.L_HI(net1314));
 sg13g2_tiehi _18435__1315 (.L_HI(net1315));
 sg13g2_tiehi _18434__1316 (.L_HI(net1316));
 sg13g2_tiehi _18433__1317 (.L_HI(net1317));
 sg13g2_tiehi _18432__1318 (.L_HI(net1318));
 sg13g2_tiehi _18431__1319 (.L_HI(net1319));
 sg13g2_tiehi _18430__1320 (.L_HI(net1320));
 sg13g2_tiehi _18429__1321 (.L_HI(net1321));
 sg13g2_tiehi _18428__1322 (.L_HI(net1322));
 sg13g2_tiehi _18427__1323 (.L_HI(net1323));
 sg13g2_tiehi _18426__1324 (.L_HI(net1324));
 sg13g2_tiehi _18425__1325 (.L_HI(net1325));
 sg13g2_tiehi _18424__1326 (.L_HI(net1326));
 sg13g2_tiehi _18423__1327 (.L_HI(net1327));
 sg13g2_tiehi _18422__1328 (.L_HI(net1328));
 sg13g2_tiehi _18421__1329 (.L_HI(net1329));
 sg13g2_tiehi _18420__1330 (.L_HI(net1330));
 sg13g2_tiehi _18419__1331 (.L_HI(net1331));
 sg13g2_tiehi _18418__1332 (.L_HI(net1332));
 sg13g2_tiehi _18417__1333 (.L_HI(net1333));
 sg13g2_tiehi _18416__1334 (.L_HI(net1334));
 sg13g2_tiehi _18415__1335 (.L_HI(net1335));
 sg13g2_tiehi _18414__1336 (.L_HI(net1336));
 sg13g2_tiehi _18413__1337 (.L_HI(net1337));
 sg13g2_tiehi _18412__1338 (.L_HI(net1338));
 sg13g2_tiehi _18411__1339 (.L_HI(net1339));
 sg13g2_tiehi _18410__1340 (.L_HI(net1340));
 sg13g2_tiehi _18409__1341 (.L_HI(net1341));
 sg13g2_tiehi _18408__1342 (.L_HI(net1342));
 sg13g2_tiehi _18407__1343 (.L_HI(net1343));
 sg13g2_tiehi _18406__1344 (.L_HI(net1344));
 sg13g2_tiehi _18405__1345 (.L_HI(net1345));
 sg13g2_tiehi _18404__1346 (.L_HI(net1346));
 sg13g2_tiehi _18403__1347 (.L_HI(net1347));
 sg13g2_tiehi _18402__1348 (.L_HI(net1348));
 sg13g2_tiehi _18401__1349 (.L_HI(net1349));
 sg13g2_tiehi _18400__1350 (.L_HI(net1350));
 sg13g2_tiehi _18399__1351 (.L_HI(net1351));
 sg13g2_tiehi _18398__1352 (.L_HI(net1352));
 sg13g2_tiehi _18397__1353 (.L_HI(net1353));
 sg13g2_tiehi _18396__1354 (.L_HI(net1354));
 sg13g2_tiehi _18395__1355 (.L_HI(net1355));
 sg13g2_tiehi _18394__1356 (.L_HI(net1356));
 sg13g2_tiehi _18393__1357 (.L_HI(net1357));
 sg13g2_tiehi _18392__1358 (.L_HI(net1358));
 sg13g2_tiehi _18391__1359 (.L_HI(net1359));
 sg13g2_tiehi _18390__1360 (.L_HI(net1360));
 sg13g2_tiehi _18389__1361 (.L_HI(net1361));
 sg13g2_tiehi _18388__1362 (.L_HI(net1362));
 sg13g2_tiehi _18387__1363 (.L_HI(net1363));
 sg13g2_tiehi _18386__1364 (.L_HI(net1364));
 sg13g2_tiehi _18385__1365 (.L_HI(net1365));
 sg13g2_tiehi _20425__1366 (.L_HI(net1366));
 sg13g2_tiehi _20424__1367 (.L_HI(net1367));
 sg13g2_tiehi _20423__1368 (.L_HI(net1368));
 sg13g2_tiehi _20422__1369 (.L_HI(net1369));
 sg13g2_tiehi _20421__1370 (.L_HI(net1370));
 sg13g2_tiehi _20420__1371 (.L_HI(net1371));
 sg13g2_tiehi _20419__1372 (.L_HI(net1372));
 sg13g2_tiehi _20418__1373 (.L_HI(net1373));
 sg13g2_tiehi _20417__1374 (.L_HI(net1374));
 sg13g2_tiehi _20416__1375 (.L_HI(net1375));
 sg13g2_tiehi _20415__1376 (.L_HI(net1376));
 sg13g2_tiehi _20414__1377 (.L_HI(net1377));
 sg13g2_tiehi _20413__1378 (.L_HI(net1378));
 sg13g2_tiehi _20412__1379 (.L_HI(net1379));
 sg13g2_tiehi _20411__1380 (.L_HI(net1380));
 sg13g2_tiehi _20410__1381 (.L_HI(net1381));
 sg13g2_tiehi _20409__1382 (.L_HI(net1382));
 sg13g2_tiehi _20408__1383 (.L_HI(net1383));
 sg13g2_tiehi _20407__1384 (.L_HI(net1384));
 sg13g2_tiehi _20406__1385 (.L_HI(net1385));
 sg13g2_tiehi _20405__1386 (.L_HI(net1386));
 sg13g2_tiehi _20404__1387 (.L_HI(net1387));
 sg13g2_tiehi _20403__1388 (.L_HI(net1388));
 sg13g2_tiehi _20402__1389 (.L_HI(net1389));
 sg13g2_tiehi _20401__1390 (.L_HI(net1390));
 sg13g2_tiehi _20400__1391 (.L_HI(net1391));
 sg13g2_tiehi _20399__1392 (.L_HI(net1392));
 sg13g2_tiehi _20398__1393 (.L_HI(net1393));
 sg13g2_tiehi _20397__1394 (.L_HI(net1394));
 sg13g2_tiehi _20396__1395 (.L_HI(net1395));
 sg13g2_tiehi _20395__1396 (.L_HI(net1396));
 sg13g2_tiehi _20394__1397 (.L_HI(net1397));
 sg13g2_tiehi _20393__1398 (.L_HI(net1398));
 sg13g2_tiehi _20392__1399 (.L_HI(net1399));
 sg13g2_tiehi _20391__1400 (.L_HI(net1400));
 sg13g2_tiehi _20390__1401 (.L_HI(net1401));
 sg13g2_tiehi _20389__1402 (.L_HI(net1402));
 sg13g2_tiehi _20388__1403 (.L_HI(net1403));
 sg13g2_tiehi _20387__1404 (.L_HI(net1404));
 sg13g2_tiehi _20386__1405 (.L_HI(net1405));
 sg13g2_tiehi _20385__1406 (.L_HI(net1406));
 sg13g2_tiehi _20384__1407 (.L_HI(net1407));
 sg13g2_tiehi _20383__1408 (.L_HI(net1408));
 sg13g2_tiehi _20382__1409 (.L_HI(net1409));
 sg13g2_tiehi _20381__1410 (.L_HI(net1410));
 sg13g2_tiehi _20380__1411 (.L_HI(net1411));
 sg13g2_tiehi _20379__1412 (.L_HI(net1412));
 sg13g2_tiehi _20378__1413 (.L_HI(net1413));
 sg13g2_tiehi _20377__1414 (.L_HI(net1414));
 sg13g2_tiehi _20376__1415 (.L_HI(net1415));
 sg13g2_tiehi _20375__1416 (.L_HI(net1416));
 sg13g2_tiehi _20374__1417 (.L_HI(net1417));
 sg13g2_tiehi _20373__1418 (.L_HI(net1418));
 sg13g2_tiehi _20372__1419 (.L_HI(net1419));
 sg13g2_tiehi _20371__1420 (.L_HI(net1420));
 sg13g2_tiehi _20370__1421 (.L_HI(net1421));
 sg13g2_tiehi _20369__1422 (.L_HI(net1422));
 sg13g2_tiehi _20368__1423 (.L_HI(net1423));
 sg13g2_tiehi _20367__1424 (.L_HI(net1424));
 sg13g2_tiehi _20366__1425 (.L_HI(net1425));
 sg13g2_tiehi _20365__1426 (.L_HI(net1426));
 sg13g2_tiehi _20364__1427 (.L_HI(net1427));
 sg13g2_tiehi _20363__1428 (.L_HI(net1428));
 sg13g2_tiehi _20362__1429 (.L_HI(net1429));
 sg13g2_tiehi _20361__1430 (.L_HI(net1430));
 sg13g2_tiehi _20360__1431 (.L_HI(net1431));
 sg13g2_tiehi _20359__1432 (.L_HI(net1432));
 sg13g2_tiehi _20358__1433 (.L_HI(net1433));
 sg13g2_tiehi _20357__1434 (.L_HI(net1434));
 sg13g2_tiehi _20356__1435 (.L_HI(net1435));
 sg13g2_tiehi _20355__1436 (.L_HI(net1436));
 sg13g2_tiehi _20354__1437 (.L_HI(net1437));
 sg13g2_tiehi _20353__1438 (.L_HI(net1438));
 sg13g2_tiehi _20352__1439 (.L_HI(net1439));
 sg13g2_tiehi _20351__1440 (.L_HI(net1440));
 sg13g2_tiehi _20350__1441 (.L_HI(net1441));
 sg13g2_tiehi _20349__1442 (.L_HI(net1442));
 sg13g2_tiehi _20348__1443 (.L_HI(net1443));
 sg13g2_tiehi _20347__1444 (.L_HI(net1444));
 sg13g2_tiehi _20346__1445 (.L_HI(net1445));
 sg13g2_tiehi _20345__1446 (.L_HI(net1446));
 sg13g2_tiehi _20344__1447 (.L_HI(net1447));
 sg13g2_tiehi _20343__1448 (.L_HI(net1448));
 sg13g2_tiehi _20342__1449 (.L_HI(net1449));
 sg13g2_tiehi _20341__1450 (.L_HI(net1450));
 sg13g2_tiehi _20340__1451 (.L_HI(net1451));
 sg13g2_tiehi _20339__1452 (.L_HI(net1452));
 sg13g2_tiehi _20338__1453 (.L_HI(net1453));
 sg13g2_tiehi _20337__1454 (.L_HI(net1454));
 sg13g2_tiehi _20336__1455 (.L_HI(net1455));
 sg13g2_tiehi _20335__1456 (.L_HI(net1456));
 sg13g2_tiehi _20334__1457 (.L_HI(net1457));
 sg13g2_tiehi _20333__1458 (.L_HI(net1458));
 sg13g2_tiehi _20332__1459 (.L_HI(net1459));
 sg13g2_tiehi _20331__1460 (.L_HI(net1460));
 sg13g2_tiehi _20330__1461 (.L_HI(net1461));
 sg13g2_tiehi _20329__1462 (.L_HI(net1462));
 sg13g2_tiehi _20328__1463 (.L_HI(net1463));
 sg13g2_tiehi _20327__1464 (.L_HI(net1464));
 sg13g2_tiehi _20326__1465 (.L_HI(net1465));
 sg13g2_tiehi _20325__1466 (.L_HI(net1466));
 sg13g2_tiehi _20324__1467 (.L_HI(net1467));
 sg13g2_tiehi _20323__1468 (.L_HI(net1468));
 sg13g2_tiehi _20322__1469 (.L_HI(net1469));
 sg13g2_tiehi _20321__1470 (.L_HI(net1470));
 sg13g2_tiehi _20320__1471 (.L_HI(net1471));
 sg13g2_tiehi _20319__1472 (.L_HI(net1472));
 sg13g2_tiehi _20318__1473 (.L_HI(net1473));
 sg13g2_tiehi _20317__1474 (.L_HI(net1474));
 sg13g2_tiehi _20316__1475 (.L_HI(net1475));
 sg13g2_tiehi _20315__1476 (.L_HI(net1476));
 sg13g2_tiehi _20314__1477 (.L_HI(net1477));
 sg13g2_tiehi _20313__1478 (.L_HI(net1478));
 sg13g2_tiehi _20312__1479 (.L_HI(net1479));
 sg13g2_tiehi _20311__1480 (.L_HI(net1480));
 sg13g2_tiehi _20310__1481 (.L_HI(net1481));
 sg13g2_tiehi _20309__1482 (.L_HI(net1482));
 sg13g2_tiehi _20308__1483 (.L_HI(net1483));
 sg13g2_tiehi _20307__1484 (.L_HI(net1484));
 sg13g2_tiehi _20306__1485 (.L_HI(net1485));
 sg13g2_tiehi _20305__1486 (.L_HI(net1486));
 sg13g2_tiehi _20304__1487 (.L_HI(net1487));
 sg13g2_tiehi _20303__1488 (.L_HI(net1488));
 sg13g2_tiehi _20302__1489 (.L_HI(net1489));
 sg13g2_tiehi _20301__1490 (.L_HI(net1490));
 sg13g2_tiehi _20300__1491 (.L_HI(net1491));
 sg13g2_tiehi _20299__1492 (.L_HI(net1492));
 sg13g2_tiehi _20298__1493 (.L_HI(net1493));
 sg13g2_tiehi _20297__1494 (.L_HI(net1494));
 sg13g2_tiehi _20296__1495 (.L_HI(net1495));
 sg13g2_tiehi _20295__1496 (.L_HI(net1496));
 sg13g2_tiehi _20294__1497 (.L_HI(net1497));
 sg13g2_tiehi _20293__1498 (.L_HI(net1498));
 sg13g2_tiehi _20292__1499 (.L_HI(net1499));
 sg13g2_tiehi _20291__1500 (.L_HI(net1500));
 sg13g2_tiehi _20290__1501 (.L_HI(net1501));
 sg13g2_tiehi _20289__1502 (.L_HI(net1502));
 sg13g2_tiehi _20288__1503 (.L_HI(net1503));
 sg13g2_tiehi _20287__1504 (.L_HI(net1504));
 sg13g2_tiehi _20286__1505 (.L_HI(net1505));
 sg13g2_tiehi _20285__1506 (.L_HI(net1506));
 sg13g2_tiehi _20284__1507 (.L_HI(net1507));
 sg13g2_tiehi _20283__1508 (.L_HI(net1508));
 sg13g2_tiehi _20282__1509 (.L_HI(net1509));
 sg13g2_tiehi _20281__1510 (.L_HI(net1510));
 sg13g2_tiehi _20280__1511 (.L_HI(net1511));
 sg13g2_tiehi _20279__1512 (.L_HI(net1512));
 sg13g2_tiehi _20278__1513 (.L_HI(net1513));
 sg13g2_tiehi _20277__1514 (.L_HI(net1514));
 sg13g2_tiehi _20276__1515 (.L_HI(net1515));
 sg13g2_tiehi _20275__1516 (.L_HI(net1516));
 sg13g2_tiehi _20274__1517 (.L_HI(net1517));
 sg13g2_tiehi _20273__1518 (.L_HI(net1518));
 sg13g2_tiehi _20272__1519 (.L_HI(net1519));
 sg13g2_tiehi _20271__1520 (.L_HI(net1520));
 sg13g2_tiehi _20270__1521 (.L_HI(net1521));
 sg13g2_tiehi _20269__1522 (.L_HI(net1522));
 sg13g2_tiehi _20268__1523 (.L_HI(net1523));
 sg13g2_tiehi _20267__1524 (.L_HI(net1524));
 sg13g2_tiehi _20266__1525 (.L_HI(net1525));
 sg13g2_tiehi _20265__1526 (.L_HI(net1526));
 sg13g2_tiehi _20264__1527 (.L_HI(net1527));
 sg13g2_tiehi _20263__1528 (.L_HI(net1528));
 sg13g2_tiehi _20262__1529 (.L_HI(net1529));
 sg13g2_tiehi _20261__1530 (.L_HI(net1530));
 sg13g2_tiehi _20260__1531 (.L_HI(net1531));
 sg13g2_tiehi _20259__1532 (.L_HI(net1532));
 sg13g2_tiehi _20258__1533 (.L_HI(net1533));
 sg13g2_tiehi _20257__1534 (.L_HI(net1534));
 sg13g2_tiehi _20256__1535 (.L_HI(net1535));
 sg13g2_tiehi _20255__1536 (.L_HI(net1536));
 sg13g2_tiehi _20254__1537 (.L_HI(net1537));
 sg13g2_tiehi _20253__1538 (.L_HI(net1538));
 sg13g2_tiehi _20252__1539 (.L_HI(net1539));
 sg13g2_tiehi _20251__1540 (.L_HI(net1540));
 sg13g2_tiehi _20250__1541 (.L_HI(net1541));
 sg13g2_tiehi _20249__1542 (.L_HI(net1542));
 sg13g2_tiehi _20248__1543 (.L_HI(net1543));
 sg13g2_tiehi _20247__1544 (.L_HI(net1544));
 sg13g2_tiehi _20246__1545 (.L_HI(net1545));
 sg13g2_tiehi _20245__1546 (.L_HI(net1546));
 sg13g2_tiehi _20244__1547 (.L_HI(net1547));
 sg13g2_tiehi _20243__1548 (.L_HI(net1548));
 sg13g2_tiehi _20242__1549 (.L_HI(net1549));
 sg13g2_tiehi _20241__1550 (.L_HI(net1550));
 sg13g2_tiehi _20240__1551 (.L_HI(net1551));
 sg13g2_tiehi _20239__1552 (.L_HI(net1552));
 sg13g2_tiehi _20238__1553 (.L_HI(net1553));
 sg13g2_tiehi _20237__1554 (.L_HI(net1554));
 sg13g2_tiehi _20236__1555 (.L_HI(net1555));
 sg13g2_tiehi _20235__1556 (.L_HI(net1556));
 sg13g2_tiehi _20234__1557 (.L_HI(net1557));
 sg13g2_tiehi _20233__1558 (.L_HI(net1558));
 sg13g2_tiehi _20232__1559 (.L_HI(net1559));
 sg13g2_tiehi _20231__1560 (.L_HI(net1560));
 sg13g2_tiehi _20230__1561 (.L_HI(net1561));
 sg13g2_tiehi _20229__1562 (.L_HI(net1562));
 sg13g2_tiehi _20228__1563 (.L_HI(net1563));
 sg13g2_tiehi _20227__1564 (.L_HI(net1564));
 sg13g2_tiehi _20226__1565 (.L_HI(net1565));
 sg13g2_tiehi _20225__1566 (.L_HI(net1566));
 sg13g2_tiehi _20224__1567 (.L_HI(net1567));
 sg13g2_tiehi _20223__1568 (.L_HI(net1568));
 sg13g2_tiehi _20222__1569 (.L_HI(net1569));
 sg13g2_tiehi _20221__1570 (.L_HI(net1570));
 sg13g2_tiehi _20220__1571 (.L_HI(net1571));
 sg13g2_tiehi _20219__1572 (.L_HI(net1572));
 sg13g2_tiehi _20218__1573 (.L_HI(net1573));
 sg13g2_tiehi _20217__1574 (.L_HI(net1574));
 sg13g2_tiehi _20216__1575 (.L_HI(net1575));
 sg13g2_tiehi _20215__1576 (.L_HI(net1576));
 sg13g2_tiehi _20214__1577 (.L_HI(net1577));
 sg13g2_tiehi _20213__1578 (.L_HI(net1578));
 sg13g2_tiehi _20212__1579 (.L_HI(net1579));
 sg13g2_tiehi _20211__1580 (.L_HI(net1580));
 sg13g2_tiehi _20210__1581 (.L_HI(net1581));
 sg13g2_tiehi _20209__1582 (.L_HI(net1582));
 sg13g2_tiehi _20208__1583 (.L_HI(net1583));
 sg13g2_tiehi _20207__1584 (.L_HI(net1584));
 sg13g2_tiehi _20206__1585 (.L_HI(net1585));
 sg13g2_tiehi _20205__1586 (.L_HI(net1586));
 sg13g2_tiehi _20204__1587 (.L_HI(net1587));
 sg13g2_tiehi _20203__1588 (.L_HI(net1588));
 sg13g2_tiehi _20202__1589 (.L_HI(net1589));
 sg13g2_tiehi _20201__1590 (.L_HI(net1590));
 sg13g2_tiehi _20200__1591 (.L_HI(net1591));
 sg13g2_tiehi _20199__1592 (.L_HI(net1592));
 sg13g2_tiehi _20198__1593 (.L_HI(net1593));
 sg13g2_tiehi _20197__1594 (.L_HI(net1594));
 sg13g2_tiehi _20196__1595 (.L_HI(net1595));
 sg13g2_tiehi _20195__1596 (.L_HI(net1596));
 sg13g2_tiehi _20194__1597 (.L_HI(net1597));
 sg13g2_tiehi _20193__1598 (.L_HI(net1598));
 sg13g2_tiehi _20192__1599 (.L_HI(net1599));
 sg13g2_tiehi _20191__1600 (.L_HI(net1600));
 sg13g2_tiehi _20190__1601 (.L_HI(net1601));
 sg13g2_tiehi _20189__1602 (.L_HI(net1602));
 sg13g2_tiehi _20188__1603 (.L_HI(net1603));
 sg13g2_tiehi _20187__1604 (.L_HI(net1604));
 sg13g2_tiehi _20186__1605 (.L_HI(net1605));
 sg13g2_tiehi _20185__1606 (.L_HI(net1606));
 sg13g2_tiehi _20184__1607 (.L_HI(net1607));
 sg13g2_tiehi _20183__1608 (.L_HI(net1608));
 sg13g2_tiehi _20182__1609 (.L_HI(net1609));
 sg13g2_tiehi _20181__1610 (.L_HI(net1610));
 sg13g2_tiehi _20180__1611 (.L_HI(net1611));
 sg13g2_tiehi _20179__1612 (.L_HI(net1612));
 sg13g2_tiehi _20178__1613 (.L_HI(net1613));
 sg13g2_tiehi _20177__1614 (.L_HI(net1614));
 sg13g2_tiehi _20176__1615 (.L_HI(net1615));
 sg13g2_tiehi _20175__1616 (.L_HI(net1616));
 sg13g2_tiehi _20174__1617 (.L_HI(net1617));
 sg13g2_tiehi _20173__1618 (.L_HI(net1618));
 sg13g2_tiehi _20172__1619 (.L_HI(net1619));
 sg13g2_tiehi _20171__1620 (.L_HI(net1620));
 sg13g2_tiehi _20170__1621 (.L_HI(net1621));
 sg13g2_tiehi _20169__1622 (.L_HI(net1622));
 sg13g2_tiehi _20168__1623 (.L_HI(net1623));
 sg13g2_tiehi _20167__1624 (.L_HI(net1624));
 sg13g2_tiehi _20166__1625 (.L_HI(net1625));
 sg13g2_tiehi _20165__1626 (.L_HI(net1626));
 sg13g2_tiehi _20164__1627 (.L_HI(net1627));
 sg13g2_tiehi _20163__1628 (.L_HI(net1628));
 sg13g2_tiehi _20162__1629 (.L_HI(net1629));
 sg13g2_tiehi _20161__1630 (.L_HI(net1630));
 sg13g2_tiehi _20160__1631 (.L_HI(net1631));
 sg13g2_tiehi _20159__1632 (.L_HI(net1632));
 sg13g2_tiehi _20158__1633 (.L_HI(net1633));
 sg13g2_tiehi _20157__1634 (.L_HI(net1634));
 sg13g2_tiehi _20156__1635 (.L_HI(net1635));
 sg13g2_tiehi _20155__1636 (.L_HI(net1636));
 sg13g2_tiehi _20154__1637 (.L_HI(net1637));
 sg13g2_tiehi _20153__1638 (.L_HI(net1638));
 sg13g2_tiehi _20152__1639 (.L_HI(net1639));
 sg13g2_tiehi _20151__1640 (.L_HI(net1640));
 sg13g2_tiehi _20150__1641 (.L_HI(net1641));
 sg13g2_tiehi _20149__1642 (.L_HI(net1642));
 sg13g2_tiehi _20148__1643 (.L_HI(net1643));
 sg13g2_tiehi _20147__1644 (.L_HI(net1644));
 sg13g2_tiehi _20146__1645 (.L_HI(net1645));
 sg13g2_tiehi _20145__1646 (.L_HI(net1646));
 sg13g2_tiehi _20144__1647 (.L_HI(net1647));
 sg13g2_tiehi _20143__1648 (.L_HI(net1648));
 sg13g2_tiehi _20142__1649 (.L_HI(net1649));
 sg13g2_tiehi _20141__1650 (.L_HI(net1650));
 sg13g2_tiehi _20140__1651 (.L_HI(net1651));
 sg13g2_tiehi _20139__1652 (.L_HI(net1652));
 sg13g2_tiehi _20138__1653 (.L_HI(net1653));
 sg13g2_tiehi _20137__1654 (.L_HI(net1654));
 sg13g2_tiehi _20136__1655 (.L_HI(net1655));
 sg13g2_tiehi _20135__1656 (.L_HI(net1656));
 sg13g2_tiehi _20134__1657 (.L_HI(net1657));
 sg13g2_tiehi _20133__1658 (.L_HI(net1658));
 sg13g2_tiehi _20132__1659 (.L_HI(net1659));
 sg13g2_tiehi _20131__1660 (.L_HI(net1660));
 sg13g2_tiehi _20130__1661 (.L_HI(net1661));
 sg13g2_tiehi _20129__1662 (.L_HI(net1662));
 sg13g2_tiehi _20128__1663 (.L_HI(net1663));
 sg13g2_tiehi _20127__1664 (.L_HI(net1664));
 sg13g2_tiehi _20126__1665 (.L_HI(net1665));
 sg13g2_tiehi _20125__1666 (.L_HI(net1666));
 sg13g2_tiehi _20124__1667 (.L_HI(net1667));
 sg13g2_tiehi _20123__1668 (.L_HI(net1668));
 sg13g2_tiehi _20122__1669 (.L_HI(net1669));
 sg13g2_tiehi _20121__1670 (.L_HI(net1670));
 sg13g2_tiehi _20120__1671 (.L_HI(net1671));
 sg13g2_tiehi _20119__1672 (.L_HI(net1672));
 sg13g2_tiehi _20118__1673 (.L_HI(net1673));
 sg13g2_tiehi _20117__1674 (.L_HI(net1674));
 sg13g2_tiehi _20116__1675 (.L_HI(net1675));
 sg13g2_tiehi _20115__1676 (.L_HI(net1676));
 sg13g2_tiehi _20114__1677 (.L_HI(net1677));
 sg13g2_tiehi _20113__1678 (.L_HI(net1678));
 sg13g2_tiehi _20112__1679 (.L_HI(net1679));
 sg13g2_tiehi _20111__1680 (.L_HI(net1680));
 sg13g2_tiehi _20110__1681 (.L_HI(net1681));
 sg13g2_tiehi _20109__1682 (.L_HI(net1682));
 sg13g2_tiehi _20108__1683 (.L_HI(net1683));
 sg13g2_tiehi _20107__1684 (.L_HI(net1684));
 sg13g2_tiehi _20106__1685 (.L_HI(net1685));
 sg13g2_tiehi _20105__1686 (.L_HI(net1686));
 sg13g2_tiehi _20104__1687 (.L_HI(net1687));
 sg13g2_tiehi _20103__1688 (.L_HI(net1688));
 sg13g2_tiehi _20102__1689 (.L_HI(net1689));
 sg13g2_tiehi _20101__1690 (.L_HI(net1690));
 sg13g2_tiehi _20100__1691 (.L_HI(net1691));
 sg13g2_tiehi _20099__1692 (.L_HI(net1692));
 sg13g2_tiehi _20098__1693 (.L_HI(net1693));
 sg13g2_tiehi _20097__1694 (.L_HI(net1694));
 sg13g2_tiehi _20096__1695 (.L_HI(net1695));
 sg13g2_tiehi _20095__1696 (.L_HI(net1696));
 sg13g2_tiehi _20094__1697 (.L_HI(net1697));
 sg13g2_tiehi _20093__1698 (.L_HI(net1698));
 sg13g2_tiehi _20092__1699 (.L_HI(net1699));
 sg13g2_tiehi _20091__1700 (.L_HI(net1700));
 sg13g2_tiehi _20090__1701 (.L_HI(net1701));
 sg13g2_tiehi _20089__1702 (.L_HI(net1702));
 sg13g2_tiehi _20088__1703 (.L_HI(net1703));
 sg13g2_tiehi _20087__1704 (.L_HI(net1704));
 sg13g2_tiehi _20086__1705 (.L_HI(net1705));
 sg13g2_tiehi _20085__1706 (.L_HI(net1706));
 sg13g2_tiehi _20084__1707 (.L_HI(net1707));
 sg13g2_tiehi _20083__1708 (.L_HI(net1708));
 sg13g2_tiehi _20082__1709 (.L_HI(net1709));
 sg13g2_tiehi _20081__1710 (.L_HI(net1710));
 sg13g2_tiehi _20080__1711 (.L_HI(net1711));
 sg13g2_tiehi _20079__1712 (.L_HI(net1712));
 sg13g2_tiehi _20078__1713 (.L_HI(net1713));
 sg13g2_tiehi _20077__1714 (.L_HI(net1714));
 sg13g2_tiehi _20076__1715 (.L_HI(net1715));
 sg13g2_tiehi _20075__1716 (.L_HI(net1716));
 sg13g2_tiehi _20074__1717 (.L_HI(net1717));
 sg13g2_tiehi _20073__1718 (.L_HI(net1718));
 sg13g2_tiehi _20072__1719 (.L_HI(net1719));
 sg13g2_tiehi _20071__1720 (.L_HI(net1720));
 sg13g2_tiehi _20070__1721 (.L_HI(net1721));
 sg13g2_tiehi _20069__1722 (.L_HI(net1722));
 sg13g2_tiehi _20068__1723 (.L_HI(net1723));
 sg13g2_tiehi _20067__1724 (.L_HI(net1724));
 sg13g2_tiehi _20066__1725 (.L_HI(net1725));
 sg13g2_tiehi _20065__1726 (.L_HI(net1726));
 sg13g2_tiehi _20064__1727 (.L_HI(net1727));
 sg13g2_tiehi _20063__1728 (.L_HI(net1728));
 sg13g2_tiehi _20062__1729 (.L_HI(net1729));
 sg13g2_tiehi _20061__1730 (.L_HI(net1730));
 sg13g2_tiehi _20060__1731 (.L_HI(net1731));
 sg13g2_tiehi _20059__1732 (.L_HI(net1732));
 sg13g2_tiehi _20058__1733 (.L_HI(net1733));
 sg13g2_tiehi _20057__1734 (.L_HI(net1734));
 sg13g2_tiehi _20056__1735 (.L_HI(net1735));
 sg13g2_tiehi _20055__1736 (.L_HI(net1736));
 sg13g2_tiehi _20054__1737 (.L_HI(net1737));
 sg13g2_tiehi _20053__1738 (.L_HI(net1738));
 sg13g2_tiehi _20052__1739 (.L_HI(net1739));
 sg13g2_tiehi _20051__1740 (.L_HI(net1740));
 sg13g2_tiehi _20050__1741 (.L_HI(net1741));
 sg13g2_tiehi _20049__1742 (.L_HI(net1742));
 sg13g2_tiehi _20048__1743 (.L_HI(net1743));
 sg13g2_tiehi _20047__1744 (.L_HI(net1744));
 sg13g2_tiehi _20046__1745 (.L_HI(net1745));
 sg13g2_tiehi _20045__1746 (.L_HI(net1746));
 sg13g2_tiehi _20044__1747 (.L_HI(net1747));
 sg13g2_tiehi _20043__1748 (.L_HI(net1748));
 sg13g2_tiehi _20042__1749 (.L_HI(net1749));
 sg13g2_tiehi _20041__1750 (.L_HI(net1750));
 sg13g2_tiehi _20040__1751 (.L_HI(net1751));
 sg13g2_tiehi _20039__1752 (.L_HI(net1752));
 sg13g2_tiehi _20038__1753 (.L_HI(net1753));
 sg13g2_tiehi _20037__1754 (.L_HI(net1754));
 sg13g2_tiehi _20036__1755 (.L_HI(net1755));
 sg13g2_tiehi _20035__1756 (.L_HI(net1756));
 sg13g2_tiehi _20034__1757 (.L_HI(net1757));
 sg13g2_tiehi _20033__1758 (.L_HI(net1758));
 sg13g2_tiehi _20032__1759 (.L_HI(net1759));
 sg13g2_tiehi _20031__1760 (.L_HI(net1760));
 sg13g2_tiehi _20030__1761 (.L_HI(net1761));
 sg13g2_tiehi _20029__1762 (.L_HI(net1762));
 sg13g2_tiehi _20028__1763 (.L_HI(net1763));
 sg13g2_tiehi _20027__1764 (.L_HI(net1764));
 sg13g2_tiehi _20026__1765 (.L_HI(net1765));
 sg13g2_tiehi _20025__1766 (.L_HI(net1766));
 sg13g2_tiehi _20024__1767 (.L_HI(net1767));
 sg13g2_tiehi _20023__1768 (.L_HI(net1768));
 sg13g2_tiehi _20022__1769 (.L_HI(net1769));
 sg13g2_tiehi _20021__1770 (.L_HI(net1770));
 sg13g2_tiehi _20020__1771 (.L_HI(net1771));
 sg13g2_tiehi _20019__1772 (.L_HI(net1772));
 sg13g2_tiehi _20018__1773 (.L_HI(net1773));
 sg13g2_tiehi _20017__1774 (.L_HI(net1774));
 sg13g2_tiehi _20016__1775 (.L_HI(net1775));
 sg13g2_tiehi _20015__1776 (.L_HI(net1776));
 sg13g2_tiehi _20014__1777 (.L_HI(net1777));
 sg13g2_tiehi _20013__1778 (.L_HI(net1778));
 sg13g2_tiehi _20012__1779 (.L_HI(net1779));
 sg13g2_tiehi _20011__1780 (.L_HI(net1780));
 sg13g2_tiehi _20010__1781 (.L_HI(net1781));
 sg13g2_tiehi _20009__1782 (.L_HI(net1782));
 sg13g2_tiehi _20008__1783 (.L_HI(net1783));
 sg13g2_tiehi _20007__1784 (.L_HI(net1784));
 sg13g2_tiehi _20006__1785 (.L_HI(net1785));
 sg13g2_tiehi _20005__1786 (.L_HI(net1786));
 sg13g2_tiehi _20004__1787 (.L_HI(net1787));
 sg13g2_tiehi _20003__1788 (.L_HI(net1788));
 sg13g2_tiehi _20002__1789 (.L_HI(net1789));
 sg13g2_tiehi _20001__1790 (.L_HI(net1790));
 sg13g2_tiehi _20000__1791 (.L_HI(net1791));
 sg13g2_tiehi _19999__1792 (.L_HI(net1792));
 sg13g2_tiehi _19998__1793 (.L_HI(net1793));
 sg13g2_tiehi _19997__1794 (.L_HI(net1794));
 sg13g2_tiehi _19996__1795 (.L_HI(net1795));
 sg13g2_tiehi _19995__1796 (.L_HI(net1796));
 sg13g2_tiehi _19994__1797 (.L_HI(net1797));
 sg13g2_tiehi _19993__1798 (.L_HI(net1798));
 sg13g2_tiehi _19992__1799 (.L_HI(net1799));
 sg13g2_tiehi _19991__1800 (.L_HI(net1800));
 sg13g2_tiehi _19990__1801 (.L_HI(net1801));
 sg13g2_tiehi _19989__1802 (.L_HI(net1802));
 sg13g2_tiehi _19988__1803 (.L_HI(net1803));
 sg13g2_tiehi _19987__1804 (.L_HI(net1804));
 sg13g2_tiehi _19986__1805 (.L_HI(net1805));
 sg13g2_tiehi _19985__1806 (.L_HI(net1806));
 sg13g2_tiehi _19984__1807 (.L_HI(net1807));
 sg13g2_tiehi _19983__1808 (.L_HI(net1808));
 sg13g2_tiehi _19982__1809 (.L_HI(net1809));
 sg13g2_tiehi _19981__1810 (.L_HI(net1810));
 sg13g2_tiehi _19980__1811 (.L_HI(net1811));
 sg13g2_tiehi _19979__1812 (.L_HI(net1812));
 sg13g2_tiehi _19978__1813 (.L_HI(net1813));
 sg13g2_tiehi _19977__1814 (.L_HI(net1814));
 sg13g2_tiehi _19976__1815 (.L_HI(net1815));
 sg13g2_tiehi _19975__1816 (.L_HI(net1816));
 sg13g2_tiehi _19974__1817 (.L_HI(net1817));
 sg13g2_tiehi _19973__1818 (.L_HI(net1818));
 sg13g2_tiehi _19972__1819 (.L_HI(net1819));
 sg13g2_tiehi _19971__1820 (.L_HI(net1820));
 sg13g2_tiehi _19970__1821 (.L_HI(net1821));
 sg13g2_tiehi _19969__1822 (.L_HI(net1822));
 sg13g2_tiehi _19968__1823 (.L_HI(net1823));
 sg13g2_tiehi _19967__1824 (.L_HI(net1824));
 sg13g2_tiehi _19966__1825 (.L_HI(net1825));
 sg13g2_tiehi _19965__1826 (.L_HI(net1826));
 sg13g2_tiehi _19964__1827 (.L_HI(net1827));
 sg13g2_tiehi _19963__1828 (.L_HI(net1828));
 sg13g2_tiehi _19962__1829 (.L_HI(net1829));
 sg13g2_tiehi _19961__1830 (.L_HI(net1830));
 sg13g2_tiehi _19960__1831 (.L_HI(net1831));
 sg13g2_tiehi _19959__1832 (.L_HI(net1832));
 sg13g2_tiehi _19958__1833 (.L_HI(net1833));
 sg13g2_tiehi _19957__1834 (.L_HI(net1834));
 sg13g2_tiehi _19956__1835 (.L_HI(net1835));
 sg13g2_tiehi _19955__1836 (.L_HI(net1836));
 sg13g2_tiehi _19954__1837 (.L_HI(net1837));
 sg13g2_tiehi _19953__1838 (.L_HI(net1838));
 sg13g2_tiehi _19952__1839 (.L_HI(net1839));
 sg13g2_tiehi _19951__1840 (.L_HI(net1840));
 sg13g2_tiehi _19950__1841 (.L_HI(net1841));
 sg13g2_tiehi _19949__1842 (.L_HI(net1842));
 sg13g2_tiehi _19948__1843 (.L_HI(net1843));
 sg13g2_tiehi _19947__1844 (.L_HI(net1844));
 sg13g2_tiehi _19946__1845 (.L_HI(net1845));
 sg13g2_tiehi _19945__1846 (.L_HI(net1846));
 sg13g2_tiehi _19944__1847 (.L_HI(net1847));
 sg13g2_tiehi _19943__1848 (.L_HI(net1848));
 sg13g2_tiehi _19942__1849 (.L_HI(net1849));
 sg13g2_tiehi _19941__1850 (.L_HI(net1850));
 sg13g2_tiehi _19940__1851 (.L_HI(net1851));
 sg13g2_tiehi _19939__1852 (.L_HI(net1852));
 sg13g2_tiehi _19938__1853 (.L_HI(net1853));
 sg13g2_tiehi _19937__1854 (.L_HI(net1854));
 sg13g2_tiehi _19936__1855 (.L_HI(net1855));
 sg13g2_tiehi _19935__1856 (.L_HI(net1856));
 sg13g2_tiehi _19934__1857 (.L_HI(net1857));
 sg13g2_tiehi _19933__1858 (.L_HI(net1858));
 sg13g2_tiehi _19932__1859 (.L_HI(net1859));
 sg13g2_tiehi _19931__1860 (.L_HI(net1860));
 sg13g2_tiehi _19930__1861 (.L_HI(net1861));
 sg13g2_tiehi _19929__1862 (.L_HI(net1862));
 sg13g2_tiehi _19928__1863 (.L_HI(net1863));
 sg13g2_tiehi _19927__1864 (.L_HI(net1864));
 sg13g2_tiehi _19926__1865 (.L_HI(net1865));
 sg13g2_tiehi _19925__1866 (.L_HI(net1866));
 sg13g2_tiehi _19924__1867 (.L_HI(net1867));
 sg13g2_tiehi _19923__1868 (.L_HI(net1868));
 sg13g2_tiehi _19922__1869 (.L_HI(net1869));
 sg13g2_tiehi _19921__1870 (.L_HI(net1870));
 sg13g2_tiehi _19920__1871 (.L_HI(net1871));
 sg13g2_tiehi _19919__1872 (.L_HI(net1872));
 sg13g2_tiehi _19918__1873 (.L_HI(net1873));
 sg13g2_tiehi _19917__1874 (.L_HI(net1874));
 sg13g2_tiehi _19916__1875 (.L_HI(net1875));
 sg13g2_tiehi _19915__1876 (.L_HI(net1876));
 sg13g2_tiehi _19914__1877 (.L_HI(net1877));
 sg13g2_tiehi _19913__1878 (.L_HI(net1878));
 sg13g2_tiehi _19912__1879 (.L_HI(net1879));
 sg13g2_tiehi _19911__1880 (.L_HI(net1880));
 sg13g2_tiehi _19910__1881 (.L_HI(net1881));
 sg13g2_tiehi _19909__1882 (.L_HI(net1882));
 sg13g2_tiehi _19908__1883 (.L_HI(net1883));
 sg13g2_tiehi _19907__1884 (.L_HI(net1884));
 sg13g2_tiehi _19906__1885 (.L_HI(net1885));
 sg13g2_tiehi _19905__1886 (.L_HI(net1886));
 sg13g2_tiehi _19904__1887 (.L_HI(net1887));
 sg13g2_tiehi _19903__1888 (.L_HI(net1888));
 sg13g2_tiehi _19902__1889 (.L_HI(net1889));
 sg13g2_tiehi _19901__1890 (.L_HI(net1890));
 sg13g2_tiehi _19900__1891 (.L_HI(net1891));
 sg13g2_tiehi _19899__1892 (.L_HI(net1892));
 sg13g2_tiehi _19898__1893 (.L_HI(net1893));
 sg13g2_tiehi _19897__1894 (.L_HI(net1894));
 sg13g2_tiehi _19896__1895 (.L_HI(net1895));
 sg13g2_tiehi _19895__1896 (.L_HI(net1896));
 sg13g2_tiehi _19894__1897 (.L_HI(net1897));
 sg13g2_tiehi _19893__1898 (.L_HI(net1898));
 sg13g2_tiehi _19892__1899 (.L_HI(net1899));
 sg13g2_tiehi _19891__1900 (.L_HI(net1900));
 sg13g2_tiehi _19890__1901 (.L_HI(net1901));
 sg13g2_tiehi _19889__1902 (.L_HI(net1902));
 sg13g2_tiehi _19888__1903 (.L_HI(net1903));
 sg13g2_tiehi _19887__1904 (.L_HI(net1904));
 sg13g2_tiehi _19886__1905 (.L_HI(net1905));
 sg13g2_tiehi _19885__1906 (.L_HI(net1906));
 sg13g2_tiehi _19884__1907 (.L_HI(net1907));
 sg13g2_tiehi _19883__1908 (.L_HI(net1908));
 sg13g2_tiehi _19882__1909 (.L_HI(net1909));
 sg13g2_tiehi _19881__1910 (.L_HI(net1910));
 sg13g2_tiehi _19880__1911 (.L_HI(net1911));
 sg13g2_tiehi _19879__1912 (.L_HI(net1912));
 sg13g2_tiehi _19878__1913 (.L_HI(net1913));
 sg13g2_tiehi _19877__1914 (.L_HI(net1914));
 sg13g2_tiehi _19876__1915 (.L_HI(net1915));
 sg13g2_tiehi _19875__1916 (.L_HI(net1916));
 sg13g2_tiehi _19874__1917 (.L_HI(net1917));
 sg13g2_tiehi _19873__1918 (.L_HI(net1918));
 sg13g2_tiehi _19872__1919 (.L_HI(net1919));
 sg13g2_tiehi _19871__1920 (.L_HI(net1920));
 sg13g2_tiehi _19870__1921 (.L_HI(net1921));
 sg13g2_tiehi _19869__1922 (.L_HI(net1922));
 sg13g2_tiehi _19868__1923 (.L_HI(net1923));
 sg13g2_tiehi _19867__1924 (.L_HI(net1924));
 sg13g2_tiehi _19866__1925 (.L_HI(net1925));
 sg13g2_tiehi _19865__1926 (.L_HI(net1926));
 sg13g2_tiehi _19864__1927 (.L_HI(net1927));
 sg13g2_tiehi _19863__1928 (.L_HI(net1928));
 sg13g2_tiehi _19862__1929 (.L_HI(net1929));
 sg13g2_tiehi _19861__1930 (.L_HI(net1930));
 sg13g2_tiehi _19860__1931 (.L_HI(net1931));
 sg13g2_tiehi _19859__1932 (.L_HI(net1932));
 sg13g2_tiehi _19858__1933 (.L_HI(net1933));
 sg13g2_tiehi _19857__1934 (.L_HI(net1934));
 sg13g2_tiehi _19856__1935 (.L_HI(net1935));
 sg13g2_tiehi _19855__1936 (.L_HI(net1936));
 sg13g2_tiehi _19854__1937 (.L_HI(net1937));
 sg13g2_tiehi _19853__1938 (.L_HI(net1938));
 sg13g2_tiehi _19852__1939 (.L_HI(net1939));
 sg13g2_tiehi _19851__1940 (.L_HI(net1940));
 sg13g2_tiehi _19850__1941 (.L_HI(net1941));
 sg13g2_tiehi _19849__1942 (.L_HI(net1942));
 sg13g2_tiehi _19848__1943 (.L_HI(net1943));
 sg13g2_tiehi _19847__1944 (.L_HI(net1944));
 sg13g2_tiehi _19846__1945 (.L_HI(net1945));
 sg13g2_tiehi _19845__1946 (.L_HI(net1946));
 sg13g2_tiehi _19844__1947 (.L_HI(net1947));
 sg13g2_tiehi _19843__1948 (.L_HI(net1948));
 sg13g2_tiehi _19842__1949 (.L_HI(net1949));
 sg13g2_tiehi _19841__1950 (.L_HI(net1950));
 sg13g2_tiehi _19840__1951 (.L_HI(net1951));
 sg13g2_tiehi _19839__1952 (.L_HI(net1952));
 sg13g2_tiehi _19838__1953 (.L_HI(net1953));
 sg13g2_tiehi _19837__1954 (.L_HI(net1954));
 sg13g2_tiehi _19836__1955 (.L_HI(net1955));
 sg13g2_tiehi _19835__1956 (.L_HI(net1956));
 sg13g2_tiehi _19834__1957 (.L_HI(net1957));
 sg13g2_tiehi _19833__1958 (.L_HI(net1958));
 sg13g2_tiehi _19832__1959 (.L_HI(net1959));
 sg13g2_tiehi _19831__1960 (.L_HI(net1960));
 sg13g2_tiehi _19830__1961 (.L_HI(net1961));
 sg13g2_tiehi _19829__1962 (.L_HI(net1962));
 sg13g2_tiehi _19828__1963 (.L_HI(net1963));
 sg13g2_tiehi _19827__1964 (.L_HI(net1964));
 sg13g2_tiehi _19826__1965 (.L_HI(net1965));
 sg13g2_tiehi _19825__1966 (.L_HI(net1966));
 sg13g2_tiehi _19824__1967 (.L_HI(net1967));
 sg13g2_tiehi _19823__1968 (.L_HI(net1968));
 sg13g2_tiehi _19822__1969 (.L_HI(net1969));
 sg13g2_tiehi _19821__1970 (.L_HI(net1970));
 sg13g2_tiehi _19820__1971 (.L_HI(net1971));
 sg13g2_tiehi _19819__1972 (.L_HI(net1972));
 sg13g2_tiehi _19818__1973 (.L_HI(net1973));
 sg13g2_tiehi _19817__1974 (.L_HI(net1974));
 sg13g2_tiehi _19816__1975 (.L_HI(net1975));
 sg13g2_tiehi _19815__1976 (.L_HI(net1976));
 sg13g2_tiehi _19814__1977 (.L_HI(net1977));
 sg13g2_tiehi _19813__1978 (.L_HI(net1978));
 sg13g2_tiehi _19812__1979 (.L_HI(net1979));
 sg13g2_tiehi _19811__1980 (.L_HI(net1980));
 sg13g2_tiehi _19810__1981 (.L_HI(net1981));
 sg13g2_tiehi _19809__1982 (.L_HI(net1982));
 sg13g2_tiehi _19808__1983 (.L_HI(net1983));
 sg13g2_tiehi _19807__1984 (.L_HI(net1984));
 sg13g2_tiehi _19806__1985 (.L_HI(net1985));
 sg13g2_tiehi _19805__1986 (.L_HI(net1986));
 sg13g2_tiehi _19804__1987 (.L_HI(net1987));
 sg13g2_tiehi _19803__1988 (.L_HI(net1988));
 sg13g2_tiehi _19802__1989 (.L_HI(net1989));
 sg13g2_tiehi _19801__1990 (.L_HI(net1990));
 sg13g2_tiehi _19800__1991 (.L_HI(net1991));
 sg13g2_tiehi _19799__1992 (.L_HI(net1992));
 sg13g2_tiehi _19798__1993 (.L_HI(net1993));
 sg13g2_tiehi _19797__1994 (.L_HI(net1994));
 sg13g2_tiehi _19796__1995 (.L_HI(net1995));
 sg13g2_tiehi _19795__1996 (.L_HI(net1996));
 sg13g2_tiehi _19794__1997 (.L_HI(net1997));
 sg13g2_tiehi _19793__1998 (.L_HI(net1998));
 sg13g2_tiehi _19792__1999 (.L_HI(net1999));
 sg13g2_tiehi _19791__2000 (.L_HI(net2000));
 sg13g2_tiehi _19790__2001 (.L_HI(net2001));
 sg13g2_tiehi _19789__2002 (.L_HI(net2002));
 sg13g2_tiehi _19788__2003 (.L_HI(net2003));
 sg13g2_tiehi _19787__2004 (.L_HI(net2004));
 sg13g2_tiehi _19786__2005 (.L_HI(net2005));
 sg13g2_tiehi _19785__2006 (.L_HI(net2006));
 sg13g2_tiehi _19784__2007 (.L_HI(net2007));
 sg13g2_tiehi _19783__2008 (.L_HI(net2008));
 sg13g2_tiehi _19782__2009 (.L_HI(net2009));
 sg13g2_tiehi _19781__2010 (.L_HI(net2010));
 sg13g2_tiehi _19780__2011 (.L_HI(net2011));
 sg13g2_tiehi _19779__2012 (.L_HI(net2012));
 sg13g2_tiehi _19778__2013 (.L_HI(net2013));
 sg13g2_tiehi _19777__2014 (.L_HI(net2014));
 sg13g2_tiehi _19776__2015 (.L_HI(net2015));
 sg13g2_tiehi _19775__2016 (.L_HI(net2016));
 sg13g2_tiehi _19774__2017 (.L_HI(net2017));
 sg13g2_tiehi _19773__2018 (.L_HI(net2018));
 sg13g2_tiehi _19772__2019 (.L_HI(net2019));
 sg13g2_tiehi _19771__2020 (.L_HI(net2020));
 sg13g2_tiehi _19770__2021 (.L_HI(net2021));
 sg13g2_tiehi _19769__2022 (.L_HI(net2022));
 sg13g2_tiehi _19768__2023 (.L_HI(net2023));
 sg13g2_tiehi _19767__2024 (.L_HI(net2024));
 sg13g2_tiehi _19766__2025 (.L_HI(net2025));
 sg13g2_tiehi _19765__2026 (.L_HI(net2026));
 sg13g2_tiehi _19764__2027 (.L_HI(net2027));
 sg13g2_tiehi _19763__2028 (.L_HI(net2028));
 sg13g2_tiehi _19762__2029 (.L_HI(net2029));
 sg13g2_tiehi _19761__2030 (.L_HI(net2030));
 sg13g2_tiehi _19760__2031 (.L_HI(net2031));
 sg13g2_tiehi _19759__2032 (.L_HI(net2032));
 sg13g2_tiehi _19758__2033 (.L_HI(net2033));
 sg13g2_tiehi _19757__2034 (.L_HI(net2034));
 sg13g2_tiehi _19756__2035 (.L_HI(net2035));
 sg13g2_tiehi _19755__2036 (.L_HI(net2036));
 sg13g2_tiehi _19754__2037 (.L_HI(net2037));
 sg13g2_tiehi _19753__2038 (.L_HI(net2038));
 sg13g2_tiehi _19752__2039 (.L_HI(net2039));
 sg13g2_tiehi _19751__2040 (.L_HI(net2040));
 sg13g2_tiehi _19750__2041 (.L_HI(net2041));
 sg13g2_tiehi _19749__2042 (.L_HI(net2042));
 sg13g2_tiehi _19748__2043 (.L_HI(net2043));
 sg13g2_tiehi _19747__2044 (.L_HI(net2044));
 sg13g2_tiehi _19746__2045 (.L_HI(net2045));
 sg13g2_tiehi _19745__2046 (.L_HI(net2046));
 sg13g2_tiehi _19744__2047 (.L_HI(net2047));
 sg13g2_tiehi _19743__2048 (.L_HI(net2048));
 sg13g2_tiehi _19742__2049 (.L_HI(net2049));
 sg13g2_tiehi _19741__2050 (.L_HI(net2050));
 sg13g2_tiehi _19740__2051 (.L_HI(net2051));
 sg13g2_tiehi _19739__2052 (.L_HI(net2052));
 sg13g2_tiehi _19738__2053 (.L_HI(net2053));
 sg13g2_tiehi _19737__2054 (.L_HI(net2054));
 sg13g2_tiehi _19736__2055 (.L_HI(net2055));
 sg13g2_tiehi _19735__2056 (.L_HI(net2056));
 sg13g2_tiehi _19734__2057 (.L_HI(net2057));
 sg13g2_tiehi _19733__2058 (.L_HI(net2058));
 sg13g2_tiehi _19732__2059 (.L_HI(net2059));
 sg13g2_tiehi _19731__2060 (.L_HI(net2060));
 sg13g2_tiehi _19730__2061 (.L_HI(net2061));
 sg13g2_tiehi _19729__2062 (.L_HI(net2062));
 sg13g2_tiehi _19728__2063 (.L_HI(net2063));
 sg13g2_tiehi _19727__2064 (.L_HI(net2064));
 sg13g2_tiehi _19726__2065 (.L_HI(net2065));
 sg13g2_tiehi _19725__2066 (.L_HI(net2066));
 sg13g2_tiehi _19724__2067 (.L_HI(net2067));
 sg13g2_tiehi _19723__2068 (.L_HI(net2068));
 sg13g2_tiehi _19722__2069 (.L_HI(net2069));
 sg13g2_tiehi _19721__2070 (.L_HI(net2070));
 sg13g2_tiehi _19720__2071 (.L_HI(net2071));
 sg13g2_tiehi _19719__2072 (.L_HI(net2072));
 sg13g2_tiehi _19718__2073 (.L_HI(net2073));
 sg13g2_tiehi _19717__2074 (.L_HI(net2074));
 sg13g2_tiehi _19716__2075 (.L_HI(net2075));
 sg13g2_tiehi _19715__2076 (.L_HI(net2076));
 sg13g2_tiehi _19714__2077 (.L_HI(net2077));
 sg13g2_tiehi _19713__2078 (.L_HI(net2078));
 sg13g2_tiehi _19712__2079 (.L_HI(net2079));
 sg13g2_tiehi _19711__2080 (.L_HI(net2080));
 sg13g2_tiehi _19710__2081 (.L_HI(net2081));
 sg13g2_tiehi _19709__2082 (.L_HI(net2082));
 sg13g2_tiehi _19708__2083 (.L_HI(net2083));
 sg13g2_tiehi _19707__2084 (.L_HI(net2084));
 sg13g2_tiehi _19706__2085 (.L_HI(net2085));
 sg13g2_tiehi _19705__2086 (.L_HI(net2086));
 sg13g2_tiehi _19704__2087 (.L_HI(net2087));
 sg13g2_tiehi _19703__2088 (.L_HI(net2088));
 sg13g2_tiehi _19702__2089 (.L_HI(net2089));
 sg13g2_tiehi _19701__2090 (.L_HI(net2090));
 sg13g2_tiehi _19700__2091 (.L_HI(net2091));
 sg13g2_tiehi _19699__2092 (.L_HI(net2092));
 sg13g2_tiehi _19698__2093 (.L_HI(net2093));
 sg13g2_tiehi _19697__2094 (.L_HI(net2094));
 sg13g2_tiehi _19696__2095 (.L_HI(net2095));
 sg13g2_tiehi _19695__2096 (.L_HI(net2096));
 sg13g2_tiehi _19694__2097 (.L_HI(net2097));
 sg13g2_tiehi _19693__2098 (.L_HI(net2098));
 sg13g2_tiehi _19692__2099 (.L_HI(net2099));
 sg13g2_tiehi _19691__2100 (.L_HI(net2100));
 sg13g2_tiehi _19690__2101 (.L_HI(net2101));
 sg13g2_tiehi _19689__2102 (.L_HI(net2102));
 sg13g2_tiehi _19688__2103 (.L_HI(net2103));
 sg13g2_tiehi _19687__2104 (.L_HI(net2104));
 sg13g2_tiehi _19686__2105 (.L_HI(net2105));
 sg13g2_tiehi _19685__2106 (.L_HI(net2106));
 sg13g2_tiehi _19684__2107 (.L_HI(net2107));
 sg13g2_tiehi _19683__2108 (.L_HI(net2108));
 sg13g2_tiehi _19682__2109 (.L_HI(net2109));
 sg13g2_tiehi _19681__2110 (.L_HI(net2110));
 sg13g2_tiehi _19680__2111 (.L_HI(net2111));
 sg13g2_tiehi _19679__2112 (.L_HI(net2112));
 sg13g2_tiehi _19678__2113 (.L_HI(net2113));
 sg13g2_tiehi _19677__2114 (.L_HI(net2114));
 sg13g2_tiehi _19676__2115 (.L_HI(net2115));
 sg13g2_tiehi _19675__2116 (.L_HI(net2116));
 sg13g2_tiehi _19674__2117 (.L_HI(net2117));
 sg13g2_tiehi _19673__2118 (.L_HI(net2118));
 sg13g2_tiehi _19672__2119 (.L_HI(net2119));
 sg13g2_tiehi _19671__2120 (.L_HI(net2120));
 sg13g2_tiehi _19670__2121 (.L_HI(net2121));
 sg13g2_tiehi _19669__2122 (.L_HI(net2122));
 sg13g2_tiehi _19668__2123 (.L_HI(net2123));
 sg13g2_tiehi _19667__2124 (.L_HI(net2124));
 sg13g2_tiehi _19666__2125 (.L_HI(net2125));
 sg13g2_tiehi _19665__2126 (.L_HI(net2126));
 sg13g2_tiehi _19664__2127 (.L_HI(net2127));
 sg13g2_tiehi _19663__2128 (.L_HI(net2128));
 sg13g2_tiehi _19662__2129 (.L_HI(net2129));
 sg13g2_tiehi tt_um_urish_sic1_2130 (.L_HI(net2130));
 sg13g2_tiehi tt_um_urish_sic1_2131 (.L_HI(net2131));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_urish_sic1_13 (.L_LO(net13));
 sg13g2_tielo tt_um_urish_sic1_14 (.L_LO(net14));
 sg13g2_tielo tt_um_urish_sic1_15 (.L_LO(net15));
 sg13g2_tielo tt_um_urish_sic1_16 (.L_LO(net16));
 sg13g2_tielo tt_um_urish_sic1_17 (.L_LO(net17));
 sg13g2_tielo tt_um_urish_sic1_18 (.L_LO(net18));
 sg13g2_tielo tt_um_urish_sic1_19 (.L_LO(net19));
 sg13g2_tielo tt_um_urish_sic1_20 (.L_LO(net20));
 sg13g2_tielo tt_um_urish_sic1_21 (.L_LO(net21));
 sg13g2_tielo tt_um_urish_sic1_22 (.L_LO(net22));
 sg13g2_tielo tt_um_urish_sic1_23 (.L_LO(net23));
 sg13g2_tiehi _19661__24 (.L_HI(net24));
 sg13g2_buf_4 _22610_ (.X(uio_out[1]),
    .A(halted));
 sg13g2_buf_4 _22611_ (.X(uio_out[4]),
    .A(\mem.out_strobe ));
 sg13g2_buf_2 fanout4673 (.A(_02810_),
    .X(net4673));
 sg13g2_buf_2 fanout4674 (.A(_02810_),
    .X(net4674));
 sg13g2_buf_2 fanout4675 (.A(_02405_),
    .X(net4675));
 sg13g2_buf_2 fanout4676 (.A(_02405_),
    .X(net4676));
 sg13g2_buf_2 fanout4677 (.A(_02396_),
    .X(net4677));
 sg13g2_buf_2 fanout4678 (.A(_02396_),
    .X(net4678));
 sg13g2_buf_2 fanout4679 (.A(net4680),
    .X(net4679));
 sg13g2_buf_2 fanout4680 (.A(_02387_),
    .X(net4680));
 sg13g2_buf_2 fanout4681 (.A(net4682),
    .X(net4681));
 sg13g2_buf_4 fanout4682 (.X(net4682),
    .A(_02378_));
 sg13g2_buf_2 fanout4683 (.A(net4685),
    .X(net4683));
 sg13g2_buf_1 fanout4684 (.A(net4685),
    .X(net4684));
 sg13g2_buf_2 fanout4685 (.A(_02369_),
    .X(net4685));
 sg13g2_buf_2 fanout4686 (.A(net4688),
    .X(net4686));
 sg13g2_buf_1 fanout4687 (.A(net4688),
    .X(net4687));
 sg13g2_buf_2 fanout4688 (.A(_02360_),
    .X(net4688));
 sg13g2_buf_2 fanout4689 (.A(_02351_),
    .X(net4689));
 sg13g2_buf_4 fanout4690 (.X(net4690),
    .A(_02351_));
 sg13g2_buf_2 fanout4691 (.A(net4692),
    .X(net4691));
 sg13g2_buf_2 fanout4692 (.A(_02342_),
    .X(net4692));
 sg13g2_buf_2 fanout4693 (.A(net4694),
    .X(net4693));
 sg13g2_buf_2 fanout4694 (.A(_02333_),
    .X(net4694));
 sg13g2_buf_2 fanout4695 (.A(_02324_),
    .X(net4695));
 sg13g2_buf_2 fanout4696 (.A(_02324_),
    .X(net4696));
 sg13g2_buf_2 fanout4697 (.A(_02315_),
    .X(net4697));
 sg13g2_buf_2 fanout4698 (.A(_02315_),
    .X(net4698));
 sg13g2_buf_2 fanout4699 (.A(_02306_),
    .X(net4699));
 sg13g2_buf_2 fanout4700 (.A(_02306_),
    .X(net4700));
 sg13g2_buf_2 fanout4701 (.A(_02297_),
    .X(net4701));
 sg13g2_buf_2 fanout4702 (.A(_02297_),
    .X(net4702));
 sg13g2_buf_2 fanout4703 (.A(_02288_),
    .X(net4703));
 sg13g2_buf_2 fanout4704 (.A(_02288_),
    .X(net4704));
 sg13g2_buf_2 fanout4705 (.A(net4706),
    .X(net4705));
 sg13g2_buf_2 fanout4706 (.A(_02279_),
    .X(net4706));
 sg13g2_buf_2 fanout4707 (.A(_06949_),
    .X(net4707));
 sg13g2_buf_2 fanout4708 (.A(_06949_),
    .X(net4708));
 sg13g2_buf_2 fanout4709 (.A(_06859_),
    .X(net4709));
 sg13g2_buf_2 fanout4710 (.A(_06859_),
    .X(net4710));
 sg13g2_buf_2 fanout4711 (.A(_06805_),
    .X(net4711));
 sg13g2_buf_2 fanout4712 (.A(_06805_),
    .X(net4712));
 sg13g2_buf_2 fanout4713 (.A(net4714),
    .X(net4713));
 sg13g2_buf_2 fanout4714 (.A(_06796_),
    .X(net4714));
 sg13g2_buf_2 fanout4715 (.A(_06787_),
    .X(net4715));
 sg13g2_buf_2 fanout4716 (.A(_06787_),
    .X(net4716));
 sg13g2_buf_2 fanout4717 (.A(net4718),
    .X(net4717));
 sg13g2_buf_2 fanout4718 (.A(_06778_),
    .X(net4718));
 sg13g2_buf_2 fanout4719 (.A(net4720),
    .X(net4719));
 sg13g2_buf_2 fanout4720 (.A(_06769_),
    .X(net4720));
 sg13g2_buf_2 fanout4721 (.A(_06760_),
    .X(net4721));
 sg13g2_buf_2 fanout4722 (.A(_06760_),
    .X(net4722));
 sg13g2_buf_2 fanout4723 (.A(_06751_),
    .X(net4723));
 sg13g2_buf_2 fanout4724 (.A(_06751_),
    .X(net4724));
 sg13g2_buf_2 fanout4725 (.A(_06742_),
    .X(net4725));
 sg13g2_buf_2 fanout4726 (.A(_06742_),
    .X(net4726));
 sg13g2_buf_2 fanout4727 (.A(_06724_),
    .X(net4727));
 sg13g2_buf_2 fanout4728 (.A(_06724_),
    .X(net4728));
 sg13g2_buf_2 fanout4729 (.A(net4730),
    .X(net4729));
 sg13g2_buf_2 fanout4730 (.A(_06715_),
    .X(net4730));
 sg13g2_buf_2 fanout4731 (.A(_06706_),
    .X(net4731));
 sg13g2_buf_2 fanout4732 (.A(_06706_),
    .X(net4732));
 sg13g2_buf_2 fanout4733 (.A(_06697_),
    .X(net4733));
 sg13g2_buf_2 fanout4734 (.A(_06697_),
    .X(net4734));
 sg13g2_buf_2 fanout4735 (.A(_06688_),
    .X(net4735));
 sg13g2_buf_2 fanout4736 (.A(_06688_),
    .X(net4736));
 sg13g2_buf_2 fanout4737 (.A(_06679_),
    .X(net4737));
 sg13g2_buf_2 fanout4738 (.A(_06679_),
    .X(net4738));
 sg13g2_buf_2 fanout4739 (.A(net4740),
    .X(net4739));
 sg13g2_buf_2 fanout4740 (.A(net4741),
    .X(net4740));
 sg13g2_buf_2 fanout4741 (.A(_06661_),
    .X(net4741));
 sg13g2_buf_2 fanout4742 (.A(net4743),
    .X(net4742));
 sg13g2_buf_2 fanout4743 (.A(_06589_),
    .X(net4743));
 sg13g2_buf_2 fanout4744 (.A(_06499_),
    .X(net4744));
 sg13g2_buf_2 fanout4745 (.A(_06499_),
    .X(net4745));
 sg13g2_buf_2 fanout4746 (.A(_06337_),
    .X(net4746));
 sg13g2_buf_2 fanout4747 (.A(_06337_),
    .X(net4747));
 sg13g2_buf_2 fanout4748 (.A(_06290_),
    .X(net4748));
 sg13g2_buf_2 fanout4749 (.A(_06290_),
    .X(net4749));
 sg13g2_buf_2 fanout4750 (.A(_06094_),
    .X(net4750));
 sg13g2_buf_2 fanout4751 (.A(_06094_),
    .X(net4751));
 sg13g2_buf_2 fanout4752 (.A(_06085_),
    .X(net4752));
 sg13g2_buf_2 fanout4753 (.A(_06085_),
    .X(net4753));
 sg13g2_buf_2 fanout4754 (.A(_06008_),
    .X(net4754));
 sg13g2_buf_2 fanout4755 (.A(_06008_),
    .X(net4755));
 sg13g2_buf_2 fanout4756 (.A(_03621_),
    .X(net4756));
 sg13g2_buf_2 fanout4757 (.A(_03621_),
    .X(net4757));
 sg13g2_buf_2 fanout4758 (.A(_03612_),
    .X(net4758));
 sg13g2_buf_2 fanout4759 (.A(_03612_),
    .X(net4759));
 sg13g2_buf_2 fanout4760 (.A(_03594_),
    .X(net4760));
 sg13g2_buf_2 fanout4761 (.A(_03594_),
    .X(net4761));
 sg13g2_buf_2 fanout4762 (.A(_03477_),
    .X(net4762));
 sg13g2_buf_2 fanout4763 (.A(_03477_),
    .X(net4763));
 sg13g2_buf_2 fanout4764 (.A(net4765),
    .X(net4764));
 sg13g2_buf_4 fanout4765 (.X(net4765),
    .A(_03242_));
 sg13g2_buf_2 fanout4766 (.A(_03171_),
    .X(net4766));
 sg13g2_buf_2 fanout4767 (.A(_03171_),
    .X(net4767));
 sg13g2_buf_2 fanout4768 (.A(net4769),
    .X(net4768));
 sg13g2_buf_2 fanout4769 (.A(_03162_),
    .X(net4769));
 sg13g2_buf_2 fanout4770 (.A(net4771),
    .X(net4770));
 sg13g2_buf_2 fanout4771 (.A(_03141_),
    .X(net4771));
 sg13g2_buf_2 fanout4772 (.A(net4773),
    .X(net4772));
 sg13g2_buf_2 fanout4773 (.A(_03130_),
    .X(net4773));
 sg13g2_buf_2 fanout4774 (.A(net4775),
    .X(net4774));
 sg13g2_buf_2 fanout4775 (.A(_03121_),
    .X(net4775));
 sg13g2_buf_2 fanout4776 (.A(net4777),
    .X(net4776));
 sg13g2_buf_2 fanout4777 (.A(_03110_),
    .X(net4777));
 sg13g2_buf_2 fanout4778 (.A(net4779),
    .X(net4778));
 sg13g2_buf_2 fanout4779 (.A(_03099_),
    .X(net4779));
 sg13g2_buf_2 fanout4780 (.A(net4781),
    .X(net4780));
 sg13g2_buf_2 fanout4781 (.A(_03090_),
    .X(net4781));
 sg13g2_buf_2 fanout4782 (.A(_03081_),
    .X(net4782));
 sg13g2_buf_2 fanout4783 (.A(_03081_),
    .X(net4783));
 sg13g2_buf_2 fanout4784 (.A(_03036_),
    .X(net4784));
 sg13g2_buf_2 fanout4785 (.A(_03036_),
    .X(net4785));
 sg13g2_buf_2 fanout4786 (.A(_03027_),
    .X(net4786));
 sg13g2_buf_2 fanout4787 (.A(_03027_),
    .X(net4787));
 sg13g2_buf_2 fanout4788 (.A(_02993_),
    .X(net4788));
 sg13g2_buf_2 fanout4789 (.A(_02993_),
    .X(net4789));
 sg13g2_buf_2 fanout4790 (.A(_02792_),
    .X(net4790));
 sg13g2_buf_2 fanout4791 (.A(_02792_),
    .X(net4791));
 sg13g2_buf_2 fanout4792 (.A(net4793),
    .X(net4792));
 sg13g2_buf_2 fanout4793 (.A(_02783_),
    .X(net4793));
 sg13g2_buf_2 fanout4794 (.A(_02765_),
    .X(net4794));
 sg13g2_buf_2 fanout4795 (.A(_02765_),
    .X(net4795));
 sg13g2_buf_4 fanout4796 (.X(net4796),
    .A(_02756_));
 sg13g2_buf_2 fanout4797 (.A(_02756_),
    .X(net4797));
 sg13g2_buf_2 fanout4798 (.A(_02747_),
    .X(net4798));
 sg13g2_buf_2 fanout4799 (.A(_02747_),
    .X(net4799));
 sg13g2_buf_2 fanout4800 (.A(_02720_),
    .X(net4800));
 sg13g2_buf_2 fanout4801 (.A(_02720_),
    .X(net4801));
 sg13g2_buf_2 fanout4802 (.A(net4803),
    .X(net4802));
 sg13g2_buf_2 fanout4803 (.A(_02711_),
    .X(net4803));
 sg13g2_buf_2 fanout4804 (.A(_02702_),
    .X(net4804));
 sg13g2_buf_2 fanout4805 (.A(_02702_),
    .X(net4805));
 sg13g2_buf_4 fanout4806 (.X(net4806),
    .A(_02693_));
 sg13g2_buf_2 fanout4807 (.A(_02693_),
    .X(net4807));
 sg13g2_buf_2 fanout4808 (.A(net4809),
    .X(net4808));
 sg13g2_buf_2 fanout4809 (.A(_02684_),
    .X(net4809));
 sg13g2_buf_2 fanout4810 (.A(net4811),
    .X(net4810));
 sg13g2_buf_2 fanout4811 (.A(_02675_),
    .X(net4811));
 sg13g2_buf_2 fanout4812 (.A(_02666_),
    .X(net4812));
 sg13g2_buf_2 fanout4813 (.A(_02666_),
    .X(net4813));
 sg13g2_buf_2 fanout4814 (.A(net4815),
    .X(net4814));
 sg13g2_buf_2 fanout4815 (.A(_02657_),
    .X(net4815));
 sg13g2_buf_2 fanout4816 (.A(net4817),
    .X(net4816));
 sg13g2_buf_2 fanout4817 (.A(_02648_),
    .X(net4817));
 sg13g2_buf_2 fanout4818 (.A(net4820),
    .X(net4818));
 sg13g2_buf_1 fanout4819 (.A(net4820),
    .X(net4819));
 sg13g2_buf_2 fanout4820 (.A(_02639_),
    .X(net4820));
 sg13g2_buf_2 fanout4821 (.A(net4823),
    .X(net4821));
 sg13g2_buf_1 fanout4822 (.A(net4823),
    .X(net4822));
 sg13g2_buf_2 fanout4823 (.A(_02630_),
    .X(net4823));
 sg13g2_buf_2 fanout4824 (.A(_02621_),
    .X(net4824));
 sg13g2_buf_2 fanout4825 (.A(_02621_),
    .X(net4825));
 sg13g2_buf_2 fanout4826 (.A(net4827),
    .X(net4826));
 sg13g2_buf_4 fanout4827 (.X(net4827),
    .A(_02612_));
 sg13g2_buf_2 fanout4828 (.A(_02603_),
    .X(net4828));
 sg13g2_buf_2 fanout4829 (.A(_02603_),
    .X(net4829));
 sg13g2_buf_2 fanout4830 (.A(_02594_),
    .X(net4830));
 sg13g2_buf_2 fanout4831 (.A(_02594_),
    .X(net4831));
 sg13g2_buf_2 fanout4832 (.A(_02585_),
    .X(net4832));
 sg13g2_buf_2 fanout4833 (.A(_02585_),
    .X(net4833));
 sg13g2_buf_2 fanout4834 (.A(net4835),
    .X(net4834));
 sg13g2_buf_2 fanout4835 (.A(_02576_),
    .X(net4835));
 sg13g2_buf_2 fanout4836 (.A(net4837),
    .X(net4836));
 sg13g2_buf_2 fanout4837 (.A(_02567_),
    .X(net4837));
 sg13g2_buf_2 fanout4838 (.A(net4839),
    .X(net4838));
 sg13g2_buf_4 fanout4839 (.X(net4839),
    .A(_02558_));
 sg13g2_buf_2 fanout4840 (.A(net4841),
    .X(net4840));
 sg13g2_buf_2 fanout4841 (.A(_02540_),
    .X(net4841));
 sg13g2_buf_2 fanout4842 (.A(net4843),
    .X(net4842));
 sg13g2_buf_2 fanout4843 (.A(_02531_),
    .X(net4843));
 sg13g2_buf_2 fanout4844 (.A(net4845),
    .X(net4844));
 sg13g2_buf_2 fanout4845 (.A(_02522_),
    .X(net4845));
 sg13g2_buf_2 fanout4846 (.A(net4847),
    .X(net4846));
 sg13g2_buf_2 fanout4847 (.A(_02513_),
    .X(net4847));
 sg13g2_buf_2 fanout4848 (.A(net4849),
    .X(net4848));
 sg13g2_buf_2 fanout4849 (.A(_02504_),
    .X(net4849));
 sg13g2_buf_2 fanout4850 (.A(_02495_),
    .X(net4850));
 sg13g2_buf_2 fanout4851 (.A(_02495_),
    .X(net4851));
 sg13g2_buf_2 fanout4852 (.A(_02486_),
    .X(net4852));
 sg13g2_buf_2 fanout4853 (.A(_02486_),
    .X(net4853));
 sg13g2_buf_2 fanout4854 (.A(net4855),
    .X(net4854));
 sg13g2_buf_2 fanout4855 (.A(_02477_),
    .X(net4855));
 sg13g2_buf_2 fanout4856 (.A(net4857),
    .X(net4856));
 sg13g2_buf_2 fanout4857 (.A(_02468_),
    .X(net4857));
 sg13g2_buf_2 fanout4858 (.A(net4859),
    .X(net4858));
 sg13g2_buf_2 fanout4859 (.A(_02459_),
    .X(net4859));
 sg13g2_buf_2 fanout4860 (.A(net4861),
    .X(net4860));
 sg13g2_buf_2 fanout4861 (.A(_02450_),
    .X(net4861));
 sg13g2_buf_2 fanout4862 (.A(_02441_),
    .X(net4862));
 sg13g2_buf_2 fanout4863 (.A(_02441_),
    .X(net4863));
 sg13g2_buf_2 fanout4864 (.A(_02432_),
    .X(net4864));
 sg13g2_buf_2 fanout4865 (.A(_02432_),
    .X(net4865));
 sg13g2_buf_2 fanout4866 (.A(_02423_),
    .X(net4866));
 sg13g2_buf_2 fanout4867 (.A(_02423_),
    .X(net4867));
 sg13g2_buf_2 fanout4868 (.A(_02414_),
    .X(net4868));
 sg13g2_buf_2 fanout4869 (.A(_02414_),
    .X(net4869));
 sg13g2_buf_2 fanout4870 (.A(net4871),
    .X(net4870));
 sg13g2_buf_2 fanout4871 (.A(_02270_),
    .X(net4871));
 sg13g2_buf_2 fanout4872 (.A(_02252_),
    .X(net4872));
 sg13g2_buf_2 fanout4873 (.A(_02252_),
    .X(net4873));
 sg13g2_buf_2 fanout4874 (.A(_02243_),
    .X(net4874));
 sg13g2_buf_2 fanout4875 (.A(_02243_),
    .X(net4875));
 sg13g2_buf_2 fanout4876 (.A(_02234_),
    .X(net4876));
 sg13g2_buf_2 fanout4877 (.A(_02234_),
    .X(net4877));
 sg13g2_buf_2 fanout4878 (.A(_02225_),
    .X(net4878));
 sg13g2_buf_2 fanout4879 (.A(_02225_),
    .X(net4879));
 sg13g2_buf_2 fanout4880 (.A(_02216_),
    .X(net4880));
 sg13g2_buf_2 fanout4881 (.A(_02216_),
    .X(net4881));
 sg13g2_buf_2 fanout4882 (.A(_02207_),
    .X(net4882));
 sg13g2_buf_2 fanout4883 (.A(_02207_),
    .X(net4883));
 sg13g2_buf_2 fanout4884 (.A(net4885),
    .X(net4884));
 sg13g2_buf_2 fanout4885 (.A(_02198_),
    .X(net4885));
 sg13g2_buf_2 fanout4886 (.A(net4887),
    .X(net4886));
 sg13g2_buf_2 fanout4887 (.A(_02189_),
    .X(net4887));
 sg13g2_buf_2 fanout4888 (.A(_02180_),
    .X(net4888));
 sg13g2_buf_2 fanout4889 (.A(_02180_),
    .X(net4889));
 sg13g2_buf_4 fanout4890 (.X(net4890),
    .A(_02171_));
 sg13g2_buf_2 fanout4891 (.A(_02171_),
    .X(net4891));
 sg13g2_buf_2 fanout4892 (.A(_02162_),
    .X(net4892));
 sg13g2_buf_2 fanout4893 (.A(_02162_),
    .X(net4893));
 sg13g2_buf_4 fanout4894 (.X(net4894),
    .A(_02153_));
 sg13g2_buf_2 fanout4895 (.A(_02153_),
    .X(net4895));
 sg13g2_buf_2 fanout4896 (.A(_02144_),
    .X(net4896));
 sg13g2_buf_2 fanout4897 (.A(_02144_),
    .X(net4897));
 sg13g2_buf_2 fanout4898 (.A(net4899),
    .X(net4898));
 sg13g2_buf_2 fanout4899 (.A(_02135_),
    .X(net4899));
 sg13g2_buf_2 fanout4900 (.A(net4901),
    .X(net4900));
 sg13g2_buf_2 fanout4901 (.A(_02126_),
    .X(net4901));
 sg13g2_buf_2 fanout4902 (.A(net4903),
    .X(net4902));
 sg13g2_buf_2 fanout4903 (.A(_07084_),
    .X(net4903));
 sg13g2_buf_2 fanout4904 (.A(net4905),
    .X(net4904));
 sg13g2_buf_2 fanout4905 (.A(_07075_),
    .X(net4905));
 sg13g2_buf_2 fanout4906 (.A(net4907),
    .X(net4906));
 sg13g2_buf_2 fanout4907 (.A(_07066_),
    .X(net4907));
 sg13g2_buf_4 fanout4908 (.X(net4908),
    .A(_07057_));
 sg13g2_buf_2 fanout4909 (.A(_07057_),
    .X(net4909));
 sg13g2_buf_2 fanout4910 (.A(net4911),
    .X(net4910));
 sg13g2_buf_2 fanout4911 (.A(_07048_),
    .X(net4911));
 sg13g2_buf_4 fanout4912 (.X(net4912),
    .A(_07039_));
 sg13g2_buf_2 fanout4913 (.A(_07039_),
    .X(net4913));
 sg13g2_buf_2 fanout4914 (.A(net4915),
    .X(net4914));
 sg13g2_buf_2 fanout4915 (.A(_07030_),
    .X(net4915));
 sg13g2_buf_2 fanout4916 (.A(_07021_),
    .X(net4916));
 sg13g2_buf_2 fanout4917 (.A(_07021_),
    .X(net4917));
 sg13g2_buf_2 fanout4918 (.A(_07012_),
    .X(net4918));
 sg13g2_buf_2 fanout4919 (.A(_07012_),
    .X(net4919));
 sg13g2_buf_2 fanout4920 (.A(net4921),
    .X(net4920));
 sg13g2_buf_2 fanout4921 (.A(_07003_),
    .X(net4921));
 sg13g2_buf_2 fanout4922 (.A(net4923),
    .X(net4922));
 sg13g2_buf_2 fanout4923 (.A(_06994_),
    .X(net4923));
 sg13g2_buf_2 fanout4924 (.A(net4925),
    .X(net4924));
 sg13g2_buf_2 fanout4925 (.A(_06985_),
    .X(net4925));
 sg13g2_buf_2 fanout4926 (.A(net4927),
    .X(net4926));
 sg13g2_buf_2 fanout4927 (.A(_06958_),
    .X(net4927));
 sg13g2_buf_4 fanout4928 (.X(net4928),
    .A(_06940_));
 sg13g2_buf_2 fanout4929 (.A(_06940_),
    .X(net4929));
 sg13g2_buf_2 fanout4930 (.A(_06931_),
    .X(net4930));
 sg13g2_buf_2 fanout4931 (.A(_06931_),
    .X(net4931));
 sg13g2_buf_4 fanout4932 (.X(net4932),
    .A(net4933));
 sg13g2_buf_2 fanout4933 (.A(_06922_),
    .X(net4933));
 sg13g2_buf_2 fanout4934 (.A(_06913_),
    .X(net4934));
 sg13g2_buf_2 fanout4935 (.A(_06913_),
    .X(net4935));
 sg13g2_buf_2 fanout4936 (.A(_06904_),
    .X(net4936));
 sg13g2_buf_2 fanout4937 (.A(_06904_),
    .X(net4937));
 sg13g2_buf_2 fanout4938 (.A(net4939),
    .X(net4938));
 sg13g2_buf_2 fanout4939 (.A(_06895_),
    .X(net4939));
 sg13g2_buf_2 fanout4940 (.A(_06886_),
    .X(net4940));
 sg13g2_buf_2 fanout4941 (.A(_06886_),
    .X(net4941));
 sg13g2_buf_2 fanout4942 (.A(net4943),
    .X(net4942));
 sg13g2_buf_2 fanout4943 (.A(_06877_),
    .X(net4943));
 sg13g2_buf_2 fanout4944 (.A(net4945),
    .X(net4944));
 sg13g2_buf_2 fanout4945 (.A(_06868_),
    .X(net4945));
 sg13g2_buf_2 fanout4946 (.A(net4947),
    .X(net4946));
 sg13g2_buf_2 fanout4947 (.A(_06850_),
    .X(net4947));
 sg13g2_buf_2 fanout4948 (.A(net4949),
    .X(net4948));
 sg13g2_buf_2 fanout4949 (.A(_06841_),
    .X(net4949));
 sg13g2_buf_2 fanout4950 (.A(net4951),
    .X(net4950));
 sg13g2_buf_2 fanout4951 (.A(_06814_),
    .X(net4951));
 sg13g2_buf_2 fanout4952 (.A(net4953),
    .X(net4952));
 sg13g2_buf_2 fanout4953 (.A(_06733_),
    .X(net4953));
 sg13g2_buf_2 fanout4954 (.A(_06670_),
    .X(net4954));
 sg13g2_buf_2 fanout4955 (.A(_06670_),
    .X(net4955));
 sg13g2_buf_2 fanout4956 (.A(net4957),
    .X(net4956));
 sg13g2_buf_2 fanout4957 (.A(net4958),
    .X(net4957));
 sg13g2_buf_2 fanout4958 (.A(_06652_),
    .X(net4958));
 sg13g2_buf_2 fanout4959 (.A(net4961),
    .X(net4959));
 sg13g2_buf_1 fanout4960 (.A(net4961),
    .X(net4960));
 sg13g2_buf_2 fanout4961 (.A(_06643_),
    .X(net4961));
 sg13g2_buf_2 fanout4962 (.A(net4964),
    .X(net4962));
 sg13g2_buf_1 fanout4963 (.A(net4964),
    .X(net4963));
 sg13g2_buf_2 fanout4964 (.A(_06634_),
    .X(net4964));
 sg13g2_buf_2 fanout4965 (.A(net4966),
    .X(net4965));
 sg13g2_buf_2 fanout4966 (.A(_06625_),
    .X(net4966));
 sg13g2_buf_2 fanout4967 (.A(net4968),
    .X(net4967));
 sg13g2_buf_2 fanout4968 (.A(_06616_),
    .X(net4968));
 sg13g2_buf_2 fanout4969 (.A(net4970),
    .X(net4969));
 sg13g2_buf_2 fanout4970 (.A(_06607_),
    .X(net4970));
 sg13g2_buf_2 fanout4971 (.A(net4972),
    .X(net4971));
 sg13g2_buf_4 fanout4972 (.X(net4972),
    .A(_06598_));
 sg13g2_buf_2 fanout4973 (.A(net4974),
    .X(net4973));
 sg13g2_buf_4 fanout4974 (.X(net4974),
    .A(_06580_));
 sg13g2_buf_2 fanout4975 (.A(net4976),
    .X(net4975));
 sg13g2_buf_4 fanout4976 (.X(net4976),
    .A(_06571_));
 sg13g2_buf_2 fanout4977 (.A(_06562_),
    .X(net4977));
 sg13g2_buf_4 fanout4978 (.X(net4978),
    .A(_06562_));
 sg13g2_buf_2 fanout4979 (.A(_06553_),
    .X(net4979));
 sg13g2_buf_2 fanout4980 (.A(_06553_),
    .X(net4980));
 sg13g2_buf_2 fanout4981 (.A(_06544_),
    .X(net4981));
 sg13g2_buf_2 fanout4982 (.A(_06544_),
    .X(net4982));
 sg13g2_buf_2 fanout4983 (.A(net4984),
    .X(net4983));
 sg13g2_buf_4 fanout4984 (.X(net4984),
    .A(_06535_));
 sg13g2_buf_4 fanout4985 (.X(net4985),
    .A(net4986));
 sg13g2_buf_2 fanout4986 (.A(_06526_),
    .X(net4986));
 sg13g2_buf_2 fanout4987 (.A(net4988),
    .X(net4987));
 sg13g2_buf_2 fanout4988 (.A(_06508_),
    .X(net4988));
 sg13g2_buf_4 fanout4989 (.X(net4989),
    .A(_06490_));
 sg13g2_buf_2 fanout4990 (.A(_06490_),
    .X(net4990));
 sg13g2_buf_2 fanout4991 (.A(_06481_),
    .X(net4991));
 sg13g2_buf_2 fanout4992 (.A(_06481_),
    .X(net4992));
 sg13g2_buf_2 fanout4993 (.A(net4994),
    .X(net4993));
 sg13g2_buf_2 fanout4994 (.A(_06472_),
    .X(net4994));
 sg13g2_buf_2 fanout4995 (.A(_06463_),
    .X(net4995));
 sg13g2_buf_2 fanout4996 (.A(_06463_),
    .X(net4996));
 sg13g2_buf_2 fanout4997 (.A(_06454_),
    .X(net4997));
 sg13g2_buf_2 fanout4998 (.A(_06454_),
    .X(net4998));
 sg13g2_buf_2 fanout4999 (.A(net5001),
    .X(net4999));
 sg13g2_buf_1 fanout5000 (.A(net5001),
    .X(net5000));
 sg13g2_buf_2 fanout5001 (.A(_06445_),
    .X(net5001));
 sg13g2_buf_2 fanout5002 (.A(net5004),
    .X(net5002));
 sg13g2_buf_1 fanout5003 (.A(net5004),
    .X(net5003));
 sg13g2_buf_2 fanout5004 (.A(_06436_),
    .X(net5004));
 sg13g2_buf_2 fanout5005 (.A(net5007),
    .X(net5005));
 sg13g2_buf_1 fanout5006 (.A(net5007),
    .X(net5006));
 sg13g2_buf_2 fanout5007 (.A(_06427_),
    .X(net5007));
 sg13g2_buf_2 fanout5008 (.A(net5010),
    .X(net5008));
 sg13g2_buf_2 fanout5009 (.A(net5010),
    .X(net5009));
 sg13g2_buf_2 fanout5010 (.A(_06418_),
    .X(net5010));
 sg13g2_buf_2 fanout5011 (.A(net5012),
    .X(net5011));
 sg13g2_buf_2 fanout5012 (.A(_06409_),
    .X(net5012));
 sg13g2_buf_4 fanout5013 (.X(net5013),
    .A(_06382_));
 sg13g2_buf_2 fanout5014 (.A(_06382_),
    .X(net5014));
 sg13g2_buf_2 fanout5015 (.A(_06364_),
    .X(net5015));
 sg13g2_buf_2 fanout5016 (.A(_06364_),
    .X(net5016));
 sg13g2_buf_2 fanout5017 (.A(_06355_),
    .X(net5017));
 sg13g2_buf_2 fanout5018 (.A(_06355_),
    .X(net5018));
 sg13g2_buf_2 fanout5019 (.A(_06346_),
    .X(net5019));
 sg13g2_buf_2 fanout5020 (.A(_06346_),
    .X(net5020));
 sg13g2_buf_2 fanout5021 (.A(net5022),
    .X(net5021));
 sg13g2_buf_2 fanout5022 (.A(_06328_),
    .X(net5022));
 sg13g2_buf_4 fanout5023 (.X(net5023),
    .A(_06319_));
 sg13g2_buf_2 fanout5024 (.A(_06319_),
    .X(net5024));
 sg13g2_buf_2 fanout5025 (.A(net5026),
    .X(net5025));
 sg13g2_buf_2 fanout5026 (.A(_06299_),
    .X(net5026));
 sg13g2_buf_2 fanout5027 (.A(net5028),
    .X(net5027));
 sg13g2_buf_2 fanout5028 (.A(_06281_),
    .X(net5028));
 sg13g2_buf_2 fanout5029 (.A(_06272_),
    .X(net5029));
 sg13g2_buf_2 fanout5030 (.A(_06272_),
    .X(net5030));
 sg13g2_buf_2 fanout5031 (.A(net5032),
    .X(net5031));
 sg13g2_buf_2 fanout5032 (.A(_06254_),
    .X(net5032));
 sg13g2_buf_2 fanout5033 (.A(net5034),
    .X(net5033));
 sg13g2_buf_2 fanout5034 (.A(_06244_),
    .X(net5034));
 sg13g2_buf_2 fanout5035 (.A(_06235_),
    .X(net5035));
 sg13g2_buf_2 fanout5036 (.A(_06235_),
    .X(net5036));
 sg13g2_buf_2 fanout5037 (.A(_06226_),
    .X(net5037));
 sg13g2_buf_2 fanout5038 (.A(_06226_),
    .X(net5038));
 sg13g2_buf_2 fanout5039 (.A(net5040),
    .X(net5039));
 sg13g2_buf_2 fanout5040 (.A(_06217_),
    .X(net5040));
 sg13g2_buf_2 fanout5041 (.A(_06208_),
    .X(net5041));
 sg13g2_buf_2 fanout5042 (.A(_06208_),
    .X(net5042));
 sg13g2_buf_2 fanout5043 (.A(net5044),
    .X(net5043));
 sg13g2_buf_2 fanout5044 (.A(_06198_),
    .X(net5044));
 sg13g2_buf_2 fanout5045 (.A(_06197_),
    .X(net5045));
 sg13g2_buf_2 fanout5046 (.A(_06197_),
    .X(net5046));
 sg13g2_buf_2 fanout5047 (.A(_06188_),
    .X(net5047));
 sg13g2_buf_2 fanout5048 (.A(_06188_),
    .X(net5048));
 sg13g2_buf_2 fanout5049 (.A(net5050),
    .X(net5049));
 sg13g2_buf_2 fanout5050 (.A(_06179_),
    .X(net5050));
 sg13g2_buf_4 fanout5051 (.X(net5051),
    .A(_06169_));
 sg13g2_buf_2 fanout5052 (.A(_06169_),
    .X(net5052));
 sg13g2_buf_2 fanout5053 (.A(_06150_),
    .X(net5053));
 sg13g2_buf_2 fanout5054 (.A(_06150_),
    .X(net5054));
 sg13g2_buf_2 fanout5055 (.A(_06130_),
    .X(net5055));
 sg13g2_buf_2 fanout5056 (.A(_06130_),
    .X(net5056));
 sg13g2_buf_2 fanout5057 (.A(_06121_),
    .X(net5057));
 sg13g2_buf_2 fanout5058 (.A(_06121_),
    .X(net5058));
 sg13g2_buf_2 fanout5059 (.A(_06112_),
    .X(net5059));
 sg13g2_buf_2 fanout5060 (.A(_06112_),
    .X(net5060));
 sg13g2_buf_2 fanout5061 (.A(net5062),
    .X(net5061));
 sg13g2_buf_2 fanout5062 (.A(_06103_),
    .X(net5062));
 sg13g2_buf_4 fanout5063 (.X(net5063),
    .A(net5064));
 sg13g2_buf_2 fanout5064 (.A(_03630_),
    .X(net5064));
 sg13g2_buf_2 fanout5065 (.A(net5067),
    .X(net5065));
 sg13g2_buf_1 fanout5066 (.A(net5067),
    .X(net5066));
 sg13g2_buf_2 fanout5067 (.A(_03603_),
    .X(net5067));
 sg13g2_buf_2 fanout5068 (.A(net5069),
    .X(net5068));
 sg13g2_buf_2 fanout5069 (.A(_03585_),
    .X(net5069));
 sg13g2_buf_2 fanout5070 (.A(net5071),
    .X(net5070));
 sg13g2_buf_2 fanout5071 (.A(_03576_),
    .X(net5071));
 sg13g2_buf_2 fanout5072 (.A(net5073),
    .X(net5072));
 sg13g2_buf_2 fanout5073 (.A(_03567_),
    .X(net5073));
 sg13g2_buf_2 fanout5074 (.A(_03558_),
    .X(net5074));
 sg13g2_buf_2 fanout5075 (.A(_03558_),
    .X(net5075));
 sg13g2_buf_2 fanout5076 (.A(_03549_),
    .X(net5076));
 sg13g2_buf_2 fanout5077 (.A(_03549_),
    .X(net5077));
 sg13g2_buf_2 fanout5078 (.A(net5079),
    .X(net5078));
 sg13g2_buf_2 fanout5079 (.A(_03540_),
    .X(net5079));
 sg13g2_buf_2 fanout5080 (.A(_03531_),
    .X(net5080));
 sg13g2_buf_2 fanout5081 (.A(_03531_),
    .X(net5081));
 sg13g2_buf_2 fanout5082 (.A(_03522_),
    .X(net5082));
 sg13g2_buf_2 fanout5083 (.A(_03522_),
    .X(net5083));
 sg13g2_buf_2 fanout5084 (.A(net5085),
    .X(net5084));
 sg13g2_buf_2 fanout5085 (.A(_03504_),
    .X(net5085));
 sg13g2_buf_2 fanout5086 (.A(net5087),
    .X(net5086));
 sg13g2_buf_2 fanout5087 (.A(_03495_),
    .X(net5087));
 sg13g2_buf_2 fanout5088 (.A(_03468_),
    .X(net5088));
 sg13g2_buf_2 fanout5089 (.A(_03468_),
    .X(net5089));
 sg13g2_buf_2 fanout5090 (.A(net5091),
    .X(net5090));
 sg13g2_buf_2 fanout5091 (.A(_03457_),
    .X(net5091));
 sg13g2_buf_4 fanout5092 (.X(net5092),
    .A(_03448_));
 sg13g2_buf_2 fanout5093 (.A(_03448_),
    .X(net5093));
 sg13g2_buf_4 fanout5094 (.X(net5094),
    .A(net5095));
 sg13g2_buf_2 fanout5095 (.A(_03439_),
    .X(net5095));
 sg13g2_buf_2 fanout5096 (.A(_03430_),
    .X(net5096));
 sg13g2_buf_2 fanout5097 (.A(_03430_),
    .X(net5097));
 sg13g2_buf_2 fanout5098 (.A(_03421_),
    .X(net5098));
 sg13g2_buf_2 fanout5099 (.A(_03421_),
    .X(net5099));
 sg13g2_buf_2 fanout5100 (.A(net5101),
    .X(net5100));
 sg13g2_buf_2 fanout5101 (.A(_03412_),
    .X(net5101));
 sg13g2_buf_2 fanout5102 (.A(_03403_),
    .X(net5102));
 sg13g2_buf_2 fanout5103 (.A(_03403_),
    .X(net5103));
 sg13g2_buf_2 fanout5104 (.A(net5105),
    .X(net5104));
 sg13g2_buf_2 fanout5105 (.A(_03394_),
    .X(net5105));
 sg13g2_buf_2 fanout5106 (.A(net5107),
    .X(net5106));
 sg13g2_buf_2 fanout5107 (.A(_03385_),
    .X(net5107));
 sg13g2_buf_2 fanout5108 (.A(_03376_),
    .X(net5108));
 sg13g2_buf_2 fanout5109 (.A(_03376_),
    .X(net5109));
 sg13g2_buf_2 fanout5110 (.A(net5111),
    .X(net5110));
 sg13g2_buf_2 fanout5111 (.A(_03365_),
    .X(net5111));
 sg13g2_buf_2 fanout5112 (.A(_03354_),
    .X(net5112));
 sg13g2_buf_2 fanout5113 (.A(_03354_),
    .X(net5113));
 sg13g2_buf_2 fanout5114 (.A(net5115),
    .X(net5114));
 sg13g2_buf_2 fanout5115 (.A(_03344_),
    .X(net5115));
 sg13g2_buf_2 fanout5116 (.A(_03295_),
    .X(net5116));
 sg13g2_buf_1 fanout5117 (.A(_03295_),
    .X(net5117));
 sg13g2_buf_2 fanout5118 (.A(_03279_),
    .X(net5118));
 sg13g2_buf_2 fanout5119 (.A(_03279_),
    .X(net5119));
 sg13g2_buf_2 fanout5120 (.A(_03269_),
    .X(net5120));
 sg13g2_buf_2 fanout5121 (.A(_03269_),
    .X(net5121));
 sg13g2_buf_2 fanout5122 (.A(_03260_),
    .X(net5122));
 sg13g2_buf_2 fanout5123 (.A(_03260_),
    .X(net5123));
 sg13g2_buf_2 fanout5124 (.A(_03251_),
    .X(net5124));
 sg13g2_buf_2 fanout5125 (.A(_03251_),
    .X(net5125));
 sg13g2_buf_2 fanout5126 (.A(_03233_),
    .X(net5126));
 sg13g2_buf_2 fanout5127 (.A(_03233_),
    .X(net5127));
 sg13g2_buf_2 fanout5128 (.A(net5129),
    .X(net5128));
 sg13g2_buf_4 fanout5129 (.X(net5129),
    .A(_03224_));
 sg13g2_buf_2 fanout5130 (.A(_03214_),
    .X(net5130));
 sg13g2_buf_2 fanout5131 (.A(_03214_),
    .X(net5131));
 sg13g2_buf_2 fanout5132 (.A(net5133),
    .X(net5132));
 sg13g2_buf_2 fanout5133 (.A(_03202_),
    .X(net5133));
 sg13g2_buf_2 fanout5134 (.A(net5135),
    .X(net5134));
 sg13g2_buf_2 fanout5135 (.A(_03191_),
    .X(net5135));
 sg13g2_buf_2 fanout5136 (.A(net5137),
    .X(net5136));
 sg13g2_buf_2 fanout5137 (.A(_03182_),
    .X(net5137));
 sg13g2_buf_4 fanout5138 (.X(net5138),
    .A(_03161_));
 sg13g2_buf_2 fanout5139 (.A(_03161_),
    .X(net5139));
 sg13g2_buf_2 fanout5140 (.A(net5141),
    .X(net5140));
 sg13g2_buf_2 fanout5141 (.A(_03150_),
    .X(net5141));
 sg13g2_buf_4 fanout5142 (.X(net5142),
    .A(net5143));
 sg13g2_buf_2 fanout5143 (.A(_03077_),
    .X(net5143));
 sg13g2_buf_2 fanout5144 (.A(_03068_),
    .X(net5144));
 sg13g2_buf_2 fanout5145 (.A(_03068_),
    .X(net5145));
 sg13g2_buf_2 fanout5146 (.A(net5147),
    .X(net5146));
 sg13g2_buf_2 fanout5147 (.A(_03057_),
    .X(net5147));
 sg13g2_buf_2 fanout5148 (.A(net5149),
    .X(net5148));
 sg13g2_buf_2 fanout5149 (.A(_03048_),
    .X(net5149));
 sg13g2_buf_2 fanout5150 (.A(net5151),
    .X(net5150));
 sg13g2_buf_2 fanout5151 (.A(_03018_),
    .X(net5151));
 sg13g2_buf_2 fanout5152 (.A(net5153),
    .X(net5152));
 sg13g2_buf_2 fanout5153 (.A(_03005_),
    .X(net5153));
 sg13g2_buf_2 fanout5154 (.A(net5155),
    .X(net5154));
 sg13g2_buf_2 fanout5155 (.A(_02992_),
    .X(net5155));
 sg13g2_buf_2 fanout5156 (.A(_02982_),
    .X(net5156));
 sg13g2_buf_4 fanout5157 (.X(net5157),
    .A(_02982_));
 sg13g2_buf_2 fanout5158 (.A(_02969_),
    .X(net5158));
 sg13g2_buf_2 fanout5159 (.A(_02969_),
    .X(net5159));
 sg13g2_buf_2 fanout5160 (.A(net5161),
    .X(net5160));
 sg13g2_buf_2 fanout5161 (.A(_02952_),
    .X(net5161));
 sg13g2_buf_2 fanout5162 (.A(_02801_),
    .X(net5162));
 sg13g2_buf_2 fanout5163 (.A(_02801_),
    .X(net5163));
 sg13g2_buf_2 fanout5164 (.A(_02774_),
    .X(net5164));
 sg13g2_buf_2 fanout5165 (.A(_02774_),
    .X(net5165));
 sg13g2_buf_2 fanout5166 (.A(_02738_),
    .X(net5166));
 sg13g2_buf_2 fanout5167 (.A(_02738_),
    .X(net5167));
 sg13g2_buf_2 fanout5168 (.A(net5169),
    .X(net5168));
 sg13g2_buf_2 fanout5169 (.A(_02729_),
    .X(net5169));
 sg13g2_buf_2 fanout5170 (.A(net5171),
    .X(net5170));
 sg13g2_buf_2 fanout5171 (.A(_02549_),
    .X(net5171));
 sg13g2_buf_2 fanout5172 (.A(_02261_),
    .X(net5172));
 sg13g2_buf_2 fanout5173 (.A(_02261_),
    .X(net5173));
 sg13g2_buf_2 fanout5174 (.A(_07093_),
    .X(net5174));
 sg13g2_buf_2 fanout5175 (.A(_07093_),
    .X(net5175));
 sg13g2_buf_2 fanout5176 (.A(net5177),
    .X(net5176));
 sg13g2_buf_2 fanout5177 (.A(_06976_),
    .X(net5177));
 sg13g2_buf_2 fanout5178 (.A(_06967_),
    .X(net5178));
 sg13g2_buf_2 fanout5179 (.A(_06967_),
    .X(net5179));
 sg13g2_buf_2 fanout5180 (.A(net5181),
    .X(net5180));
 sg13g2_buf_2 fanout5181 (.A(_06832_),
    .X(net5181));
 sg13g2_buf_2 fanout5182 (.A(net5183),
    .X(net5182));
 sg13g2_buf_2 fanout5183 (.A(_06823_),
    .X(net5183));
 sg13g2_buf_2 fanout5184 (.A(net5185),
    .X(net5184));
 sg13g2_buf_2 fanout5185 (.A(_06517_),
    .X(net5185));
 sg13g2_buf_2 fanout5186 (.A(_06400_),
    .X(net5186));
 sg13g2_buf_2 fanout5187 (.A(_06400_),
    .X(net5187));
 sg13g2_buf_2 fanout5188 (.A(_06391_),
    .X(net5188));
 sg13g2_buf_2 fanout5189 (.A(_06391_),
    .X(net5189));
 sg13g2_buf_2 fanout5190 (.A(_06373_),
    .X(net5190));
 sg13g2_buf_2 fanout5191 (.A(_06373_),
    .X(net5191));
 sg13g2_buf_2 fanout5192 (.A(_06263_),
    .X(net5192));
 sg13g2_buf_2 fanout5193 (.A(_06263_),
    .X(net5193));
 sg13g2_buf_4 fanout5194 (.X(net5194),
    .A(_06253_));
 sg13g2_buf_2 fanout5195 (.A(_06253_),
    .X(net5195));
 sg13g2_buf_4 fanout5196 (.X(net5196),
    .A(net5197));
 sg13g2_buf_4 fanout5197 (.X(net5197),
    .A(_06207_));
 sg13g2_buf_2 fanout5198 (.A(net5199),
    .X(net5198));
 sg13g2_buf_4 fanout5199 (.X(net5199),
    .A(_06178_));
 sg13g2_buf_2 fanout5200 (.A(_06160_),
    .X(net5200));
 sg13g2_buf_2 fanout5201 (.A(_06160_),
    .X(net5201));
 sg13g2_buf_4 fanout5202 (.X(net5202),
    .A(net5203));
 sg13g2_buf_4 fanout5203 (.X(net5203),
    .A(_06159_));
 sg13g2_buf_2 fanout5204 (.A(_06141_),
    .X(net5204));
 sg13g2_buf_2 fanout5205 (.A(_06141_),
    .X(net5205));
 sg13g2_buf_2 fanout5206 (.A(net5207),
    .X(net5206));
 sg13g2_buf_2 fanout5207 (.A(_03513_),
    .X(net5207));
 sg13g2_buf_2 fanout5208 (.A(net5209),
    .X(net5208));
 sg13g2_buf_2 fanout5209 (.A(_03486_),
    .X(net5209));
 sg13g2_buf_4 fanout5210 (.X(net5210),
    .A(_03364_));
 sg13g2_buf_2 fanout5211 (.A(net5212),
    .X(net5211));
 sg13g2_buf_2 fanout5212 (.A(_03278_),
    .X(net5212));
 sg13g2_buf_4 fanout5213 (.X(net5213),
    .A(_03223_));
 sg13g2_buf_4 fanout5214 (.X(net5214),
    .A(_03223_));
 sg13g2_buf_4 fanout5215 (.X(net5215),
    .A(net5216));
 sg13g2_buf_2 fanout5216 (.A(_03213_),
    .X(net5216));
 sg13g2_buf_4 fanout5217 (.X(net5217),
    .A(net5219));
 sg13g2_buf_1 fanout5218 (.A(net5219),
    .X(net5218));
 sg13g2_buf_2 fanout5219 (.A(_03181_),
    .X(net5219));
 sg13g2_buf_4 fanout5220 (.X(net5220),
    .A(net5221));
 sg13g2_buf_4 fanout5221 (.X(net5221),
    .A(_02991_));
 sg13g2_buf_4 fanout5222 (.X(net5222),
    .A(_02968_));
 sg13g2_buf_4 fanout5223 (.X(net5223),
    .A(_02951_));
 sg13g2_buf_2 fanout5224 (.A(_02951_),
    .X(net5224));
 sg13g2_buf_2 fanout5225 (.A(net5226),
    .X(net5225));
 sg13g2_buf_2 fanout5226 (.A(_06310_),
    .X(net5226));
 sg13g2_buf_8 fanout5227 (.A(_02965_),
    .X(net5227));
 sg13g2_buf_2 fanout5228 (.A(_02965_),
    .X(net5228));
 sg13g2_buf_8 fanout5229 (.A(_02948_),
    .X(net5229));
 sg13g2_buf_4 fanout5230 (.X(net5230),
    .A(_02948_));
 sg13g2_buf_2 fanout5231 (.A(net5232),
    .X(net5231));
 sg13g2_buf_2 fanout5232 (.A(_06017_),
    .X(net5232));
 sg13g2_buf_2 fanout5233 (.A(_05965_),
    .X(net5233));
 sg13g2_buf_16 fanout5234 (.X(net5234),
    .A(_03200_));
 sg13g2_buf_16 fanout5235 (.X(net5235),
    .A(_03108_));
 sg13g2_buf_8 fanout5236 (.A(_03066_),
    .X(net5236));
 sg13g2_buf_8 fanout5237 (.A(_03047_),
    .X(net5237));
 sg13g2_buf_8 fanout5238 (.A(_03047_),
    .X(net5238));
 sg13g2_buf_16 fanout5239 (.X(net5239),
    .A(_03016_));
 sg13g2_buf_8 fanout5240 (.A(net5241),
    .X(net5240));
 sg13g2_buf_16 fanout5241 (.X(net5241),
    .A(_03003_));
 sg13g2_buf_16 fanout5242 (.X(net5242),
    .A(_02980_));
 sg13g2_buf_16 fanout5243 (.X(net5243),
    .A(_02963_));
 sg13g2_buf_16 fanout5244 (.X(net5244),
    .A(_02938_));
 sg13g2_buf_16 fanout5245 (.X(net5245),
    .A(_03466_));
 sg13g2_buf_8 fanout5246 (.A(_03374_),
    .X(net5246));
 sg13g2_buf_4 fanout5247 (.X(net5247),
    .A(_03374_));
 sg13g2_buf_8 fanout5248 (.A(_03353_),
    .X(net5248));
 sg13g2_buf_8 fanout5249 (.A(_03353_),
    .X(net5249));
 sg13g2_buf_4 fanout5250 (.X(net5250),
    .A(_03291_));
 sg13g2_buf_8 fanout5251 (.A(_03211_),
    .X(net5251));
 sg13g2_buf_16 fanout5252 (.X(net5252),
    .A(_03140_));
 sg13g2_buf_16 fanout5253 (.X(net5253),
    .A(_03119_));
 sg13g2_buf_16 fanout5254 (.X(net5254),
    .A(_03080_));
 sg13g2_buf_2 fanout5255 (.A(_02898_),
    .X(net5255));
 sg13g2_buf_2 fanout5256 (.A(_02898_),
    .X(net5256));
 sg13g2_buf_4 fanout5257 (.X(net5257),
    .A(_03290_));
 sg13g2_buf_4 fanout5258 (.X(net5258),
    .A(_03160_));
 sg13g2_buf_8 fanout5259 (.A(_02950_),
    .X(net5259));
 sg13g2_buf_2 fanout5260 (.A(net5261),
    .X(net5260));
 sg13g2_buf_2 fanout5261 (.A(_02842_),
    .X(net5261));
 sg13g2_buf_8 fanout5262 (.A(_02839_),
    .X(net5262));
 sg13g2_buf_2 fanout5263 (.A(_02839_),
    .X(net5263));
 sg13g2_buf_8 fanout5264 (.A(net5267),
    .X(net5264));
 sg13g2_buf_4 fanout5265 (.X(net5265),
    .A(net5267));
 sg13g2_buf_4 fanout5266 (.X(net5266),
    .A(net5267));
 sg13g2_buf_8 fanout5267 (.A(_02838_),
    .X(net5267));
 sg13g2_buf_4 fanout5268 (.X(net5268),
    .A(net5269));
 sg13g2_buf_8 fanout5269 (.A(net5270),
    .X(net5269));
 sg13g2_buf_8 fanout5270 (.A(_02837_),
    .X(net5270));
 sg13g2_buf_4 fanout5271 (.X(net5271),
    .A(net5272));
 sg13g2_buf_4 fanout5272 (.X(net5272),
    .A(net5275));
 sg13g2_buf_8 fanout5273 (.A(net5275),
    .X(net5273));
 sg13g2_buf_4 fanout5274 (.X(net5274),
    .A(net5275));
 sg13g2_buf_4 fanout5275 (.X(net5275),
    .A(_02837_));
 sg13g2_buf_2 fanout5276 (.A(net5278),
    .X(net5276));
 sg13g2_buf_2 fanout5277 (.A(net5278),
    .X(net5277));
 sg13g2_buf_4 fanout5278 (.X(net5278),
    .A(net5286));
 sg13g2_buf_4 fanout5279 (.X(net5279),
    .A(net5286));
 sg13g2_buf_4 fanout5280 (.X(net5280),
    .A(net5286));
 sg13g2_buf_4 fanout5281 (.X(net5281),
    .A(net5282));
 sg13g2_buf_4 fanout5282 (.X(net5282),
    .A(net5285));
 sg13g2_buf_4 fanout5283 (.X(net5283),
    .A(net5284));
 sg13g2_buf_4 fanout5284 (.X(net5284),
    .A(net5285));
 sg13g2_buf_2 fanout5285 (.A(net5286),
    .X(net5285));
 sg13g2_buf_4 fanout5286 (.X(net5286),
    .A(_02836_));
 sg13g2_buf_4 fanout5287 (.X(net5287),
    .A(net5288));
 sg13g2_buf_4 fanout5288 (.X(net5288),
    .A(net5289));
 sg13g2_buf_4 fanout5289 (.X(net5289),
    .A(net5297));
 sg13g2_buf_4 fanout5290 (.X(net5290),
    .A(net5297));
 sg13g2_buf_4 fanout5291 (.X(net5291),
    .A(net5297));
 sg13g2_buf_4 fanout5292 (.X(net5292),
    .A(net5294));
 sg13g2_buf_4 fanout5293 (.X(net5293),
    .A(net5294));
 sg13g2_buf_2 fanout5294 (.A(net5296),
    .X(net5294));
 sg13g2_buf_8 fanout5295 (.A(net5296),
    .X(net5295));
 sg13g2_buf_4 fanout5296 (.X(net5296),
    .A(net5297));
 sg13g2_buf_4 fanout5297 (.X(net5297),
    .A(_02836_));
 sg13g2_buf_4 fanout5298 (.X(net5298),
    .A(net5301));
 sg13g2_buf_4 fanout5299 (.X(net5299),
    .A(net5301));
 sg13g2_buf_2 fanout5300 (.A(net5301),
    .X(net5300));
 sg13g2_buf_2 fanout5301 (.A(net5309),
    .X(net5301));
 sg13g2_buf_4 fanout5302 (.X(net5302),
    .A(net5303));
 sg13g2_buf_4 fanout5303 (.X(net5303),
    .A(net5309));
 sg13g2_buf_4 fanout5304 (.X(net5304),
    .A(net5305));
 sg13g2_buf_2 fanout5305 (.A(net5309),
    .X(net5305));
 sg13g2_buf_2 fanout5306 (.A(net5308),
    .X(net5306));
 sg13g2_buf_4 fanout5307 (.X(net5307),
    .A(net5308));
 sg13g2_buf_2 fanout5308 (.A(net5309),
    .X(net5308));
 sg13g2_buf_8 fanout5309 (.A(net5322),
    .X(net5309));
 sg13g2_buf_2 fanout5310 (.A(net5311),
    .X(net5310));
 sg13g2_buf_2 fanout5311 (.A(net5322),
    .X(net5311));
 sg13g2_buf_2 fanout5312 (.A(net5314),
    .X(net5312));
 sg13g2_buf_2 fanout5313 (.A(net5314),
    .X(net5313));
 sg13g2_buf_4 fanout5314 (.X(net5314),
    .A(net5322));
 sg13g2_buf_4 fanout5315 (.X(net5315),
    .A(net5317));
 sg13g2_buf_4 fanout5316 (.X(net5316),
    .A(net5317));
 sg13g2_buf_2 fanout5317 (.A(net5321),
    .X(net5317));
 sg13g2_buf_2 fanout5318 (.A(net5321),
    .X(net5318));
 sg13g2_buf_2 fanout5319 (.A(net5321),
    .X(net5319));
 sg13g2_buf_4 fanout5320 (.X(net5320),
    .A(net5321));
 sg13g2_buf_2 fanout5321 (.A(net5322),
    .X(net5321));
 sg13g2_buf_2 fanout5322 (.A(net5347),
    .X(net5322));
 sg13g2_buf_4 fanout5323 (.X(net5323),
    .A(net5324));
 sg13g2_buf_4 fanout5324 (.X(net5324),
    .A(net5327));
 sg13g2_buf_4 fanout5325 (.X(net5325),
    .A(net5326));
 sg13g2_buf_4 fanout5326 (.X(net5326),
    .A(net5327));
 sg13g2_buf_4 fanout5327 (.X(net5327),
    .A(net5347));
 sg13g2_buf_4 fanout5328 (.X(net5328),
    .A(net5329));
 sg13g2_buf_4 fanout5329 (.X(net5329),
    .A(net5333));
 sg13g2_buf_2 fanout5330 (.A(net5333),
    .X(net5330));
 sg13g2_buf_2 fanout5331 (.A(net5332),
    .X(net5331));
 sg13g2_buf_4 fanout5332 (.X(net5332),
    .A(net5333));
 sg13g2_buf_2 fanout5333 (.A(net5347),
    .X(net5333));
 sg13g2_buf_2 fanout5334 (.A(net5335),
    .X(net5334));
 sg13g2_buf_2 fanout5335 (.A(net5346),
    .X(net5335));
 sg13g2_buf_2 fanout5336 (.A(net5346),
    .X(net5336));
 sg13g2_buf_4 fanout5337 (.X(net5337),
    .A(net5338));
 sg13g2_buf_4 fanout5338 (.X(net5338),
    .A(net5339));
 sg13g2_buf_4 fanout5339 (.X(net5339),
    .A(net5346));
 sg13g2_buf_2 fanout5340 (.A(net5343),
    .X(net5340));
 sg13g2_buf_4 fanout5341 (.X(net5341),
    .A(net5343));
 sg13g2_buf_1 fanout5342 (.A(net5343),
    .X(net5342));
 sg13g2_buf_2 fanout5343 (.A(net5346),
    .X(net5343));
 sg13g2_buf_4 fanout5344 (.X(net5344),
    .A(net5346));
 sg13g2_buf_2 fanout5345 (.A(net5346),
    .X(net5345));
 sg13g2_buf_8 fanout5346 (.A(net5347),
    .X(net5346));
 sg13g2_buf_8 fanout5347 (.A(_02835_),
    .X(net5347));
 sg13g2_buf_4 fanout5348 (.X(net5348),
    .A(net5349));
 sg13g2_buf_4 fanout5349 (.X(net5349),
    .A(net5352));
 sg13g2_buf_4 fanout5350 (.X(net5350),
    .A(net5352));
 sg13g2_buf_2 fanout5351 (.A(net5352),
    .X(net5351));
 sg13g2_buf_4 fanout5352 (.X(net5352),
    .A(net5369));
 sg13g2_buf_2 fanout5353 (.A(net5354),
    .X(net5353));
 sg13g2_buf_4 fanout5354 (.X(net5354),
    .A(net5369));
 sg13g2_buf_4 fanout5355 (.X(net5355),
    .A(net5356));
 sg13g2_buf_4 fanout5356 (.X(net5356),
    .A(net5369));
 sg13g2_buf_4 fanout5357 (.X(net5357),
    .A(net5360));
 sg13g2_buf_4 fanout5358 (.X(net5358),
    .A(net5359));
 sg13g2_buf_4 fanout5359 (.X(net5359),
    .A(net5360));
 sg13g2_buf_4 fanout5360 (.X(net5360),
    .A(net5369));
 sg13g2_buf_4 fanout5361 (.X(net5361),
    .A(net5364));
 sg13g2_buf_4 fanout5362 (.X(net5362),
    .A(net5364));
 sg13g2_buf_2 fanout5363 (.A(net5364),
    .X(net5363));
 sg13g2_buf_4 fanout5364 (.X(net5364),
    .A(net5369));
 sg13g2_buf_4 fanout5365 (.X(net5365),
    .A(net5366));
 sg13g2_buf_4 fanout5366 (.X(net5366),
    .A(net5368));
 sg13g2_buf_4 fanout5367 (.X(net5367),
    .A(net5368));
 sg13g2_buf_4 fanout5368 (.X(net5368),
    .A(net5369));
 sg13g2_buf_8 fanout5369 (.A(_02834_),
    .X(net5369));
 sg13g2_buf_4 fanout5370 (.X(net5370),
    .A(net5371));
 sg13g2_buf_4 fanout5371 (.X(net5371),
    .A(net5384));
 sg13g2_buf_2 fanout5372 (.A(net5376),
    .X(net5372));
 sg13g2_buf_2 fanout5373 (.A(net5376),
    .X(net5373));
 sg13g2_buf_4 fanout5374 (.X(net5374),
    .A(net5376));
 sg13g2_buf_2 fanout5375 (.A(net5376),
    .X(net5375));
 sg13g2_buf_2 fanout5376 (.A(net5384),
    .X(net5376));
 sg13g2_buf_4 fanout5377 (.X(net5377),
    .A(net5384));
 sg13g2_buf_2 fanout5378 (.A(net5379),
    .X(net5378));
 sg13g2_buf_2 fanout5379 (.A(net5384),
    .X(net5379));
 sg13g2_buf_2 fanout5380 (.A(net5383),
    .X(net5380));
 sg13g2_buf_4 fanout5381 (.X(net5381),
    .A(net5383));
 sg13g2_buf_2 fanout5382 (.A(net5383),
    .X(net5382));
 sg13g2_buf_2 fanout5383 (.A(net5384),
    .X(net5383));
 sg13g2_buf_8 fanout5384 (.A(net5395),
    .X(net5384));
 sg13g2_buf_4 fanout5385 (.X(net5385),
    .A(net5386));
 sg13g2_buf_4 fanout5386 (.X(net5386),
    .A(net5387));
 sg13g2_buf_4 fanout5387 (.X(net5387),
    .A(net5395));
 sg13g2_buf_2 fanout5388 (.A(net5390),
    .X(net5388));
 sg13g2_buf_4 fanout5389 (.X(net5389),
    .A(net5390));
 sg13g2_buf_2 fanout5390 (.A(net5395),
    .X(net5390));
 sg13g2_buf_2 fanout5391 (.A(net5392),
    .X(net5391));
 sg13g2_buf_4 fanout5392 (.X(net5392),
    .A(net5394));
 sg13g2_buf_4 fanout5393 (.X(net5393),
    .A(net5394));
 sg13g2_buf_2 fanout5394 (.A(net5395),
    .X(net5394));
 sg13g2_buf_4 fanout5395 (.X(net5395),
    .A(_02833_));
 sg13g2_buf_4 fanout5396 (.X(net5396),
    .A(net5398));
 sg13g2_buf_2 fanout5397 (.A(net5398),
    .X(net5397));
 sg13g2_buf_2 fanout5398 (.A(net5408),
    .X(net5398));
 sg13g2_buf_4 fanout5399 (.X(net5399),
    .A(net5401));
 sg13g2_buf_2 fanout5400 (.A(net5401),
    .X(net5400));
 sg13g2_buf_2 fanout5401 (.A(net5408),
    .X(net5401));
 sg13g2_buf_4 fanout5402 (.X(net5402),
    .A(net5404));
 sg13g2_buf_4 fanout5403 (.X(net5403),
    .A(net5404));
 sg13g2_buf_4 fanout5404 (.X(net5404),
    .A(net5408));
 sg13g2_buf_4 fanout5405 (.X(net5405),
    .A(net5407));
 sg13g2_buf_4 fanout5406 (.X(net5406),
    .A(net5407));
 sg13g2_buf_4 fanout5407 (.X(net5407),
    .A(net5408));
 sg13g2_buf_2 fanout5408 (.A(_02833_),
    .X(net5408));
 sg13g2_buf_4 fanout5409 (.X(net5409),
    .A(net5411));
 sg13g2_buf_2 fanout5410 (.A(net5411),
    .X(net5410));
 sg13g2_buf_4 fanout5411 (.X(net5411),
    .A(net5422));
 sg13g2_buf_4 fanout5412 (.X(net5412),
    .A(net5413));
 sg13g2_buf_4 fanout5413 (.X(net5413),
    .A(net5422));
 sg13g2_buf_4 fanout5414 (.X(net5414),
    .A(net5422));
 sg13g2_buf_4 fanout5415 (.X(net5415),
    .A(net5418));
 sg13g2_buf_2 fanout5416 (.A(net5417),
    .X(net5416));
 sg13g2_buf_4 fanout5417 (.X(net5417),
    .A(net5418));
 sg13g2_buf_2 fanout5418 (.A(net5422),
    .X(net5418));
 sg13g2_buf_4 fanout5419 (.X(net5419),
    .A(net5421));
 sg13g2_buf_4 fanout5420 (.X(net5420),
    .A(net5421));
 sg13g2_buf_2 fanout5421 (.A(net5422),
    .X(net5421));
 sg13g2_buf_4 fanout5422 (.X(net5422),
    .A(_02833_));
 sg13g2_buf_2 fanout5423 (.A(net5425),
    .X(net5423));
 sg13g2_buf_2 fanout5424 (.A(net5425),
    .X(net5424));
 sg13g2_buf_2 fanout5425 (.A(net5467),
    .X(net5425));
 sg13g2_buf_2 fanout5426 (.A(net5427),
    .X(net5426));
 sg13g2_buf_4 fanout5427 (.X(net5427),
    .A(net5467));
 sg13g2_buf_2 fanout5428 (.A(net5429),
    .X(net5428));
 sg13g2_buf_2 fanout5429 (.A(net5430),
    .X(net5429));
 sg13g2_buf_2 fanout5430 (.A(net5433),
    .X(net5430));
 sg13g2_buf_4 fanout5431 (.X(net5431),
    .A(net5433));
 sg13g2_buf_4 fanout5432 (.X(net5432),
    .A(net5433));
 sg13g2_buf_4 fanout5433 (.X(net5433),
    .A(net5439));
 sg13g2_buf_4 fanout5434 (.X(net5434),
    .A(net5439));
 sg13g2_buf_4 fanout5435 (.X(net5435),
    .A(net5439));
 sg13g2_buf_4 fanout5436 (.X(net5436),
    .A(net5438));
 sg13g2_buf_2 fanout5437 (.A(net5438),
    .X(net5437));
 sg13g2_buf_4 fanout5438 (.X(net5438),
    .A(net5439));
 sg13g2_buf_4 fanout5439 (.X(net5439),
    .A(net5467));
 sg13g2_buf_4 fanout5440 (.X(net5440),
    .A(net5442));
 sg13g2_buf_4 fanout5441 (.X(net5441),
    .A(net5442));
 sg13g2_buf_2 fanout5442 (.A(net5466),
    .X(net5442));
 sg13g2_buf_4 fanout5443 (.X(net5443),
    .A(net5444));
 sg13g2_buf_2 fanout5444 (.A(net5445),
    .X(net5444));
 sg13g2_buf_4 fanout5445 (.X(net5445),
    .A(net5466));
 sg13g2_buf_4 fanout5446 (.X(net5446),
    .A(net5448));
 sg13g2_buf_2 fanout5447 (.A(net5448),
    .X(net5447));
 sg13g2_buf_4 fanout5448 (.X(net5448),
    .A(net5453));
 sg13g2_buf_4 fanout5449 (.X(net5449),
    .A(net5450));
 sg13g2_buf_1 fanout5450 (.A(net5453),
    .X(net5450));
 sg13g2_buf_2 fanout5451 (.A(net5453),
    .X(net5451));
 sg13g2_buf_2 fanout5452 (.A(net5453),
    .X(net5452));
 sg13g2_buf_4 fanout5453 (.X(net5453),
    .A(net5466));
 sg13g2_buf_4 fanout5454 (.X(net5454),
    .A(net5465));
 sg13g2_buf_2 fanout5455 (.A(net5465),
    .X(net5455));
 sg13g2_buf_4 fanout5456 (.X(net5456),
    .A(net5458));
 sg13g2_buf_4 fanout5457 (.X(net5457),
    .A(net5458));
 sg13g2_buf_4 fanout5458 (.X(net5458),
    .A(net5465));
 sg13g2_buf_4 fanout5459 (.X(net5459),
    .A(net5464));
 sg13g2_buf_4 fanout5460 (.X(net5460),
    .A(net5462));
 sg13g2_buf_1 fanout5461 (.A(net5462),
    .X(net5461));
 sg13g2_buf_2 fanout5462 (.A(net5464),
    .X(net5462));
 sg13g2_buf_4 fanout5463 (.X(net5463),
    .A(net5464));
 sg13g2_buf_4 fanout5464 (.X(net5464),
    .A(net5465));
 sg13g2_buf_4 fanout5465 (.X(net5465),
    .A(net5466));
 sg13g2_buf_4 fanout5466 (.X(net5466),
    .A(net5467));
 sg13g2_buf_8 fanout5467 (.A(_02827_),
    .X(net5467));
 sg13g2_buf_4 fanout5468 (.X(net5468),
    .A(net5469));
 sg13g2_buf_2 fanout5469 (.A(net5470),
    .X(net5469));
 sg13g2_buf_2 fanout5470 (.A(net5512),
    .X(net5470));
 sg13g2_buf_4 fanout5471 (.X(net5471),
    .A(net5472));
 sg13g2_buf_4 fanout5472 (.X(net5472),
    .A(net5512));
 sg13g2_buf_4 fanout5473 (.X(net5473),
    .A(net5476));
 sg13g2_buf_2 fanout5474 (.A(net5476),
    .X(net5474));
 sg13g2_buf_4 fanout5475 (.X(net5475),
    .A(net5476));
 sg13g2_buf_4 fanout5476 (.X(net5476),
    .A(net5484));
 sg13g2_buf_4 fanout5477 (.X(net5477),
    .A(net5484));
 sg13g2_buf_4 fanout5478 (.X(net5478),
    .A(net5479));
 sg13g2_buf_4 fanout5479 (.X(net5479),
    .A(net5484));
 sg13g2_buf_4 fanout5480 (.X(net5480),
    .A(net5484));
 sg13g2_buf_2 fanout5481 (.A(net5484),
    .X(net5481));
 sg13g2_buf_2 fanout5482 (.A(net5483),
    .X(net5482));
 sg13g2_buf_4 fanout5483 (.X(net5483),
    .A(net5484));
 sg13g2_buf_4 fanout5484 (.X(net5484),
    .A(net5512));
 sg13g2_buf_4 fanout5485 (.X(net5485),
    .A(net5488));
 sg13g2_buf_1 fanout5486 (.A(net5488),
    .X(net5486));
 sg13g2_buf_4 fanout5487 (.X(net5487),
    .A(net5488));
 sg13g2_buf_2 fanout5488 (.A(net5511),
    .X(net5488));
 sg13g2_buf_4 fanout5489 (.X(net5489),
    .A(net5490));
 sg13g2_buf_4 fanout5490 (.X(net5490),
    .A(net5491));
 sg13g2_buf_4 fanout5491 (.X(net5491),
    .A(net5511));
 sg13g2_buf_4 fanout5492 (.X(net5492),
    .A(net5499));
 sg13g2_buf_2 fanout5493 (.A(net5499),
    .X(net5493));
 sg13g2_buf_4 fanout5494 (.X(net5494),
    .A(net5499));
 sg13g2_buf_4 fanout5495 (.X(net5495),
    .A(net5496));
 sg13g2_buf_2 fanout5496 (.A(net5498),
    .X(net5496));
 sg13g2_buf_4 fanout5497 (.X(net5497),
    .A(net5498));
 sg13g2_buf_2 fanout5498 (.A(net5499),
    .X(net5498));
 sg13g2_buf_2 fanout5499 (.A(net5511),
    .X(net5499));
 sg13g2_buf_4 fanout5500 (.X(net5500),
    .A(net5501));
 sg13g2_buf_4 fanout5501 (.X(net5501),
    .A(net5506));
 sg13g2_buf_4 fanout5502 (.X(net5502),
    .A(net5506));
 sg13g2_buf_1 fanout5503 (.A(net5506),
    .X(net5503));
 sg13g2_buf_4 fanout5504 (.X(net5504),
    .A(net5506));
 sg13g2_buf_2 fanout5505 (.A(net5506),
    .X(net5505));
 sg13g2_buf_4 fanout5506 (.X(net5506),
    .A(net5511));
 sg13g2_buf_4 fanout5507 (.X(net5507),
    .A(net5509));
 sg13g2_buf_4 fanout5508 (.X(net5508),
    .A(net5509));
 sg13g2_buf_4 fanout5509 (.X(net5509),
    .A(net5510));
 sg13g2_buf_2 fanout5510 (.A(net5511),
    .X(net5510));
 sg13g2_buf_8 fanout5511 (.A(net5512),
    .X(net5511));
 sg13g2_buf_4 fanout5512 (.X(net5512),
    .A(_02826_));
 sg13g2_buf_4 fanout5513 (.X(net5513),
    .A(net5515));
 sg13g2_buf_4 fanout5514 (.X(net5514),
    .A(net5515));
 sg13g2_buf_2 fanout5515 (.A(net5517),
    .X(net5515));
 sg13g2_buf_4 fanout5516 (.X(net5516),
    .A(net5517));
 sg13g2_buf_2 fanout5517 (.A(net5557),
    .X(net5517));
 sg13g2_buf_4 fanout5518 (.X(net5518),
    .A(net5523));
 sg13g2_buf_4 fanout5519 (.X(net5519),
    .A(net5523));
 sg13g2_buf_4 fanout5520 (.X(net5520),
    .A(net5523));
 sg13g2_buf_4 fanout5521 (.X(net5521),
    .A(net5522));
 sg13g2_buf_4 fanout5522 (.X(net5522),
    .A(net5523));
 sg13g2_buf_4 fanout5523 (.X(net5523),
    .A(net5557));
 sg13g2_buf_4 fanout5524 (.X(net5524),
    .A(net5525));
 sg13g2_buf_2 fanout5525 (.A(net5531),
    .X(net5525));
 sg13g2_buf_2 fanout5526 (.A(net5530),
    .X(net5526));
 sg13g2_buf_2 fanout5527 (.A(net5530),
    .X(net5527));
 sg13g2_buf_4 fanout5528 (.X(net5528),
    .A(net5530));
 sg13g2_buf_1 fanout5529 (.A(net5530),
    .X(net5529));
 sg13g2_buf_2 fanout5530 (.A(net5531),
    .X(net5530));
 sg13g2_buf_2 fanout5531 (.A(net5557),
    .X(net5531));
 sg13g2_buf_4 fanout5532 (.X(net5532),
    .A(net5534));
 sg13g2_buf_2 fanout5533 (.A(net5534),
    .X(net5533));
 sg13g2_buf_4 fanout5534 (.X(net5534),
    .A(net5537));
 sg13g2_buf_4 fanout5535 (.X(net5535),
    .A(net5537));
 sg13g2_buf_2 fanout5536 (.A(net5537),
    .X(net5536));
 sg13g2_buf_1 fanout5537 (.A(net5557),
    .X(net5537));
 sg13g2_buf_4 fanout5538 (.X(net5538),
    .A(net5539));
 sg13g2_buf_4 fanout5539 (.X(net5539),
    .A(net5543));
 sg13g2_buf_4 fanout5540 (.X(net5540),
    .A(net5543));
 sg13g2_buf_4 fanout5541 (.X(net5541),
    .A(net5542));
 sg13g2_buf_2 fanout5542 (.A(net5543),
    .X(net5542));
 sg13g2_buf_8 fanout5543 (.A(net5557),
    .X(net5543));
 sg13g2_buf_4 fanout5544 (.X(net5544),
    .A(net5547));
 sg13g2_buf_4 fanout5545 (.X(net5545),
    .A(net5546));
 sg13g2_buf_2 fanout5546 (.A(net5547),
    .X(net5546));
 sg13g2_buf_2 fanout5547 (.A(net5556),
    .X(net5547));
 sg13g2_buf_4 fanout5548 (.X(net5548),
    .A(net5550));
 sg13g2_buf_2 fanout5549 (.A(net5550),
    .X(net5549));
 sg13g2_buf_4 fanout5550 (.X(net5550),
    .A(net5556));
 sg13g2_buf_2 fanout5551 (.A(net5552),
    .X(net5551));
 sg13g2_buf_4 fanout5552 (.X(net5552),
    .A(net5553));
 sg13g2_buf_4 fanout5553 (.X(net5553),
    .A(net5556));
 sg13g2_buf_4 fanout5554 (.X(net5554),
    .A(net5556));
 sg13g2_buf_1 fanout5555 (.A(net5556),
    .X(net5555));
 sg13g2_buf_4 fanout5556 (.X(net5556),
    .A(net5557));
 sg13g2_buf_8 fanout5557 (.A(_02825_),
    .X(net5557));
 sg13g2_buf_4 fanout5558 (.X(net5558),
    .A(net5559));
 sg13g2_buf_4 fanout5559 (.X(net5559),
    .A(net5561));
 sg13g2_buf_4 fanout5560 (.X(net5560),
    .A(net5561));
 sg13g2_buf_2 fanout5561 (.A(net5603),
    .X(net5561));
 sg13g2_buf_4 fanout5562 (.X(net5562),
    .A(net5568));
 sg13g2_buf_2 fanout5563 (.A(net5568),
    .X(net5563));
 sg13g2_buf_4 fanout5564 (.X(net5564),
    .A(net5565));
 sg13g2_buf_2 fanout5565 (.A(net5568),
    .X(net5565));
 sg13g2_buf_4 fanout5566 (.X(net5566),
    .A(net5567));
 sg13g2_buf_4 fanout5567 (.X(net5567),
    .A(net5568));
 sg13g2_buf_4 fanout5568 (.X(net5568),
    .A(net5603));
 sg13g2_buf_4 fanout5569 (.X(net5569),
    .A(net5574));
 sg13g2_buf_4 fanout5570 (.X(net5570),
    .A(net5574));
 sg13g2_buf_4 fanout5571 (.X(net5571),
    .A(net5572));
 sg13g2_buf_4 fanout5572 (.X(net5572),
    .A(net5574));
 sg13g2_buf_1 fanout5573 (.A(net5574),
    .X(net5573));
 sg13g2_buf_2 fanout5574 (.A(net5603),
    .X(net5574));
 sg13g2_buf_2 fanout5575 (.A(net5576),
    .X(net5575));
 sg13g2_buf_2 fanout5576 (.A(net5577),
    .X(net5576));
 sg13g2_buf_4 fanout5577 (.X(net5577),
    .A(net5587));
 sg13g2_buf_4 fanout5578 (.X(net5578),
    .A(net5580));
 sg13g2_buf_1 fanout5579 (.A(net5580),
    .X(net5579));
 sg13g2_buf_4 fanout5580 (.X(net5580),
    .A(net5587));
 sg13g2_buf_4 fanout5581 (.X(net5581),
    .A(net5587));
 sg13g2_buf_2 fanout5582 (.A(net5583),
    .X(net5582));
 sg13g2_buf_4 fanout5583 (.X(net5583),
    .A(net5587));
 sg13g2_buf_2 fanout5584 (.A(net5586),
    .X(net5584));
 sg13g2_buf_1 fanout5585 (.A(net5586),
    .X(net5585));
 sg13g2_buf_2 fanout5586 (.A(net5587),
    .X(net5586));
 sg13g2_buf_4 fanout5587 (.X(net5587),
    .A(net5603));
 sg13g2_buf_4 fanout5588 (.X(net5588),
    .A(net5590));
 sg13g2_buf_4 fanout5589 (.X(net5589),
    .A(net5590));
 sg13g2_buf_2 fanout5590 (.A(net5594),
    .X(net5590));
 sg13g2_buf_4 fanout5591 (.X(net5591),
    .A(net5594));
 sg13g2_buf_2 fanout5592 (.A(net5594),
    .X(net5592));
 sg13g2_buf_4 fanout5593 (.X(net5593),
    .A(net5594));
 sg13g2_buf_2 fanout5594 (.A(net5603),
    .X(net5594));
 sg13g2_buf_4 fanout5595 (.X(net5595),
    .A(net5599));
 sg13g2_buf_1 fanout5596 (.A(net5599),
    .X(net5596));
 sg13g2_buf_4 fanout5597 (.X(net5597),
    .A(net5599));
 sg13g2_buf_1 fanout5598 (.A(net5599),
    .X(net5598));
 sg13g2_buf_2 fanout5599 (.A(net5602),
    .X(net5599));
 sg13g2_buf_4 fanout5600 (.X(net5600),
    .A(net5601));
 sg13g2_buf_4 fanout5601 (.X(net5601),
    .A(net5602));
 sg13g2_buf_4 fanout5602 (.X(net5602),
    .A(net5603));
 sg13g2_buf_8 fanout5603 (.A(_02824_),
    .X(net5603));
 sg13g2_buf_4 fanout5604 (.X(net5604),
    .A(net5608));
 sg13g2_buf_2 fanout5605 (.A(net5608),
    .X(net5605));
 sg13g2_buf_4 fanout5606 (.X(net5606),
    .A(net5608));
 sg13g2_buf_2 fanout5607 (.A(net5608),
    .X(net5607));
 sg13g2_buf_4 fanout5608 (.X(net5608),
    .A(_02823_));
 sg13g2_buf_4 fanout5609 (.X(net5609),
    .A(net5610));
 sg13g2_buf_4 fanout5610 (.X(net5610),
    .A(net5613));
 sg13g2_buf_4 fanout5611 (.X(net5611),
    .A(net5613));
 sg13g2_buf_1 fanout5612 (.A(net5613),
    .X(net5612));
 sg13g2_buf_4 fanout5613 (.X(net5613),
    .A(net5619));
 sg13g2_buf_4 fanout5614 (.X(net5614),
    .A(net5619));
 sg13g2_buf_2 fanout5615 (.A(net5619),
    .X(net5615));
 sg13g2_buf_4 fanout5616 (.X(net5616),
    .A(net5617));
 sg13g2_buf_4 fanout5617 (.X(net5617),
    .A(net5618));
 sg13g2_buf_4 fanout5618 (.X(net5618),
    .A(net5619));
 sg13g2_buf_4 fanout5619 (.X(net5619),
    .A(_02823_));
 sg13g2_buf_2 fanout5620 (.A(net5621),
    .X(net5620));
 sg13g2_buf_2 fanout5621 (.A(net5622),
    .X(net5621));
 sg13g2_buf_2 fanout5622 (.A(net5623),
    .X(net5622));
 sg13g2_buf_4 fanout5623 (.X(net5623),
    .A(net5632));
 sg13g2_buf_4 fanout5624 (.X(net5624),
    .A(net5627));
 sg13g2_buf_2 fanout5625 (.A(net5627),
    .X(net5625));
 sg13g2_buf_4 fanout5626 (.X(net5626),
    .A(net5627));
 sg13g2_buf_2 fanout5627 (.A(net5632),
    .X(net5627));
 sg13g2_buf_2 fanout5628 (.A(net5629),
    .X(net5628));
 sg13g2_buf_4 fanout5629 (.X(net5629),
    .A(net5632));
 sg13g2_buf_4 fanout5630 (.X(net5630),
    .A(net5632));
 sg13g2_buf_2 fanout5631 (.A(net5632),
    .X(net5631));
 sg13g2_buf_4 fanout5632 (.X(net5632),
    .A(net5648));
 sg13g2_buf_4 fanout5633 (.X(net5633),
    .A(net5635));
 sg13g2_buf_4 fanout5634 (.X(net5634),
    .A(net5635));
 sg13g2_buf_4 fanout5635 (.X(net5635),
    .A(net5639));
 sg13g2_buf_4 fanout5636 (.X(net5636),
    .A(net5638));
 sg13g2_buf_1 fanout5637 (.A(net5638),
    .X(net5637));
 sg13g2_buf_4 fanout5638 (.X(net5638),
    .A(net5639));
 sg13g2_buf_2 fanout5639 (.A(net5648),
    .X(net5639));
 sg13g2_buf_4 fanout5640 (.X(net5640),
    .A(net5643));
 sg13g2_buf_4 fanout5641 (.X(net5641),
    .A(net5642));
 sg13g2_buf_4 fanout5642 (.X(net5642),
    .A(net5643));
 sg13g2_buf_2 fanout5643 (.A(net5648),
    .X(net5643));
 sg13g2_buf_4 fanout5644 (.X(net5644),
    .A(net5647));
 sg13g2_buf_1 fanout5645 (.A(net5647),
    .X(net5645));
 sg13g2_buf_4 fanout5646 (.X(net5646),
    .A(net5647));
 sg13g2_buf_2 fanout5647 (.A(net5648),
    .X(net5647));
 sg13g2_buf_8 fanout5648 (.A(_02823_),
    .X(net5648));
 sg13g2_buf_4 fanout5649 (.X(net5649),
    .A(net5653));
 sg13g2_buf_1 fanout5650 (.A(net5653),
    .X(net5650));
 sg13g2_buf_4 fanout5651 (.X(net5651),
    .A(net5653));
 sg13g2_buf_4 fanout5652 (.X(net5652),
    .A(net5653));
 sg13g2_buf_4 fanout5653 (.X(net5653),
    .A(net5693));
 sg13g2_buf_4 fanout5654 (.X(net5654),
    .A(net5664));
 sg13g2_buf_1 fanout5655 (.A(net5664),
    .X(net5655));
 sg13g2_buf_4 fanout5656 (.X(net5656),
    .A(net5660));
 sg13g2_buf_2 fanout5657 (.A(net5659),
    .X(net5657));
 sg13g2_buf_2 fanout5658 (.A(net5659),
    .X(net5658));
 sg13g2_buf_4 fanout5659 (.X(net5659),
    .A(net5660));
 sg13g2_buf_4 fanout5660 (.X(net5660),
    .A(net5664));
 sg13g2_buf_4 fanout5661 (.X(net5661),
    .A(net5664));
 sg13g2_buf_4 fanout5662 (.X(net5662),
    .A(net5663));
 sg13g2_buf_2 fanout5663 (.A(net5664),
    .X(net5663));
 sg13g2_buf_8 fanout5664 (.A(net5693),
    .X(net5664));
 sg13g2_buf_4 fanout5665 (.X(net5665),
    .A(net5669));
 sg13g2_buf_4 fanout5666 (.X(net5666),
    .A(net5669));
 sg13g2_buf_2 fanout5667 (.A(net5668),
    .X(net5667));
 sg13g2_buf_4 fanout5668 (.X(net5668),
    .A(net5669));
 sg13g2_buf_2 fanout5669 (.A(net5677),
    .X(net5669));
 sg13g2_buf_4 fanout5670 (.X(net5670),
    .A(net5673));
 sg13g2_buf_2 fanout5671 (.A(net5673),
    .X(net5671));
 sg13g2_buf_1 fanout5672 (.A(net5673),
    .X(net5672));
 sg13g2_buf_2 fanout5673 (.A(net5677),
    .X(net5673));
 sg13g2_buf_4 fanout5674 (.X(net5674),
    .A(net5675));
 sg13g2_buf_4 fanout5675 (.X(net5675),
    .A(net5677));
 sg13g2_buf_1 fanout5676 (.A(net5677),
    .X(net5676));
 sg13g2_buf_4 fanout5677 (.X(net5677),
    .A(net5693));
 sg13g2_buf_4 fanout5678 (.X(net5678),
    .A(net5680));
 sg13g2_buf_2 fanout5679 (.A(net5680),
    .X(net5679));
 sg13g2_buf_4 fanout5680 (.X(net5680),
    .A(net5685));
 sg13g2_buf_4 fanout5681 (.X(net5681),
    .A(net5685));
 sg13g2_buf_1 fanout5682 (.A(net5685),
    .X(net5682));
 sg13g2_buf_4 fanout5683 (.X(net5683),
    .A(net5684));
 sg13g2_buf_2 fanout5684 (.A(net5685),
    .X(net5684));
 sg13g2_buf_4 fanout5685 (.X(net5685),
    .A(net5693));
 sg13g2_buf_4 fanout5686 (.X(net5686),
    .A(net5687));
 sg13g2_buf_4 fanout5687 (.X(net5687),
    .A(net5692));
 sg13g2_buf_4 fanout5688 (.X(net5688),
    .A(net5689));
 sg13g2_buf_2 fanout5689 (.A(net5692),
    .X(net5689));
 sg13g2_buf_4 fanout5690 (.X(net5690),
    .A(net5692));
 sg13g2_buf_1 fanout5691 (.A(net5692),
    .X(net5691));
 sg13g2_buf_4 fanout5692 (.X(net5692),
    .A(net5693));
 sg13g2_buf_8 fanout5693 (.A(_02822_),
    .X(net5693));
 sg13g2_buf_4 fanout5694 (.X(net5694),
    .A(net5696));
 sg13g2_buf_1 fanout5695 (.A(net5696),
    .X(net5695));
 sg13g2_buf_4 fanout5696 (.X(net5696),
    .A(net5699));
 sg13g2_buf_4 fanout5697 (.X(net5697),
    .A(net5699));
 sg13g2_buf_2 fanout5698 (.A(net5699),
    .X(net5698));
 sg13g2_buf_4 fanout5699 (.X(net5699),
    .A(net5739));
 sg13g2_buf_2 fanout5700 (.A(net5702),
    .X(net5700));
 sg13g2_buf_2 fanout5701 (.A(net5702),
    .X(net5701));
 sg13g2_buf_2 fanout5702 (.A(net5703),
    .X(net5702));
 sg13g2_buf_4 fanout5703 (.X(net5703),
    .A(net5739));
 sg13g2_buf_4 fanout5704 (.X(net5704),
    .A(net5709));
 sg13g2_buf_4 fanout5705 (.X(net5705),
    .A(net5709));
 sg13g2_buf_2 fanout5706 (.A(net5707),
    .X(net5706));
 sg13g2_buf_2 fanout5707 (.A(net5709),
    .X(net5707));
 sg13g2_buf_4 fanout5708 (.X(net5708),
    .A(net5709));
 sg13g2_buf_2 fanout5709 (.A(net5739),
    .X(net5709));
 sg13g2_buf_4 fanout5710 (.X(net5710),
    .A(net5713));
 sg13g2_buf_2 fanout5711 (.A(net5713),
    .X(net5711));
 sg13g2_buf_4 fanout5712 (.X(net5712),
    .A(net5713));
 sg13g2_buf_2 fanout5713 (.A(net5738),
    .X(net5713));
 sg13g2_buf_4 fanout5714 (.X(net5714),
    .A(net5715));
 sg13g2_buf_2 fanout5715 (.A(net5716),
    .X(net5715));
 sg13g2_buf_2 fanout5716 (.A(net5738),
    .X(net5716));
 sg13g2_buf_4 fanout5717 (.X(net5717),
    .A(net5718));
 sg13g2_buf_4 fanout5718 (.X(net5718),
    .A(net5722));
 sg13g2_buf_4 fanout5719 (.X(net5719),
    .A(net5721));
 sg13g2_buf_1 fanout5720 (.A(net5721),
    .X(net5720));
 sg13g2_buf_4 fanout5721 (.X(net5721),
    .A(net5722));
 sg13g2_buf_4 fanout5722 (.X(net5722),
    .A(net5738));
 sg13g2_buf_4 fanout5723 (.X(net5723),
    .A(net5725));
 sg13g2_buf_1 fanout5724 (.A(net5725),
    .X(net5724));
 sg13g2_buf_4 fanout5725 (.X(net5725),
    .A(net5729));
 sg13g2_buf_4 fanout5726 (.X(net5726),
    .A(net5727));
 sg13g2_buf_4 fanout5727 (.X(net5727),
    .A(net5728));
 sg13g2_buf_4 fanout5728 (.X(net5728),
    .A(net5729));
 sg13g2_buf_1 fanout5729 (.A(net5738),
    .X(net5729));
 sg13g2_buf_4 fanout5730 (.X(net5730),
    .A(net5731));
 sg13g2_buf_2 fanout5731 (.A(net5732),
    .X(net5731));
 sg13g2_buf_2 fanout5732 (.A(net5737),
    .X(net5732));
 sg13g2_buf_4 fanout5733 (.X(net5733),
    .A(net5737));
 sg13g2_buf_2 fanout5734 (.A(net5737),
    .X(net5734));
 sg13g2_buf_4 fanout5735 (.X(net5735),
    .A(net5736));
 sg13g2_buf_2 fanout5736 (.A(net5737),
    .X(net5736));
 sg13g2_buf_4 fanout5737 (.X(net5737),
    .A(net5738));
 sg13g2_buf_8 fanout5738 (.A(net5739),
    .X(net5738));
 sg13g2_buf_8 fanout5739 (.A(_02821_),
    .X(net5739));
 sg13g2_buf_2 fanout5740 (.A(net5742),
    .X(net5740));
 sg13g2_buf_4 fanout5741 (.X(net5741),
    .A(net5742));
 sg13g2_buf_4 fanout5742 (.X(net5742),
    .A(net5744));
 sg13g2_buf_4 fanout5743 (.X(net5743),
    .A(net5744));
 sg13g2_buf_4 fanout5744 (.X(net5744),
    .A(net5784));
 sg13g2_buf_4 fanout5745 (.X(net5745),
    .A(net5747));
 sg13g2_buf_4 fanout5746 (.X(net5746),
    .A(net5756));
 sg13g2_buf_2 fanout5747 (.A(net5756),
    .X(net5747));
 sg13g2_buf_2 fanout5748 (.A(net5749),
    .X(net5748));
 sg13g2_buf_4 fanout5749 (.X(net5749),
    .A(net5756));
 sg13g2_buf_4 fanout5750 (.X(net5750),
    .A(net5751));
 sg13g2_buf_4 fanout5751 (.X(net5751),
    .A(net5755));
 sg13g2_buf_2 fanout5752 (.A(net5755),
    .X(net5752));
 sg13g2_buf_1 fanout5753 (.A(net5755),
    .X(net5753));
 sg13g2_buf_4 fanout5754 (.X(net5754),
    .A(net5755));
 sg13g2_buf_4 fanout5755 (.X(net5755),
    .A(net5756));
 sg13g2_buf_2 fanout5756 (.A(net5784),
    .X(net5756));
 sg13g2_buf_4 fanout5757 (.X(net5757),
    .A(net5758));
 sg13g2_buf_4 fanout5758 (.X(net5758),
    .A(net5769));
 sg13g2_buf_2 fanout5759 (.A(net5760),
    .X(net5759));
 sg13g2_buf_2 fanout5760 (.A(net5761),
    .X(net5760));
 sg13g2_buf_4 fanout5761 (.X(net5761),
    .A(net5769));
 sg13g2_buf_4 fanout5762 (.X(net5762),
    .A(net5763));
 sg13g2_buf_4 fanout5763 (.X(net5763),
    .A(net5769));
 sg13g2_buf_1 fanout5764 (.A(net5769),
    .X(net5764));
 sg13g2_buf_4 fanout5765 (.X(net5765),
    .A(net5768));
 sg13g2_buf_4 fanout5766 (.X(net5766),
    .A(net5768));
 sg13g2_buf_2 fanout5767 (.A(net5768),
    .X(net5767));
 sg13g2_buf_2 fanout5768 (.A(net5769),
    .X(net5768));
 sg13g2_buf_4 fanout5769 (.X(net5769),
    .A(net5784));
 sg13g2_buf_4 fanout5770 (.X(net5770),
    .A(net5772));
 sg13g2_buf_2 fanout5771 (.A(net5772),
    .X(net5771));
 sg13g2_buf_4 fanout5772 (.X(net5772),
    .A(net5777));
 sg13g2_buf_4 fanout5773 (.X(net5773),
    .A(net5776));
 sg13g2_buf_1 fanout5774 (.A(net5776),
    .X(net5774));
 sg13g2_buf_4 fanout5775 (.X(net5775),
    .A(net5776));
 sg13g2_buf_4 fanout5776 (.X(net5776),
    .A(net5777));
 sg13g2_buf_2 fanout5777 (.A(net5784),
    .X(net5777));
 sg13g2_buf_2 fanout5778 (.A(net5783),
    .X(net5778));
 sg13g2_buf_4 fanout5779 (.X(net5779),
    .A(net5782));
 sg13g2_buf_2 fanout5780 (.A(net5782),
    .X(net5780));
 sg13g2_buf_2 fanout5781 (.A(net5782),
    .X(net5781));
 sg13g2_buf_2 fanout5782 (.A(net5783),
    .X(net5782));
 sg13g2_buf_2 fanout5783 (.A(net5784),
    .X(net5783));
 sg13g2_buf_8 fanout5784 (.A(_02820_),
    .X(net5784));
 sg13g2_buf_2 fanout5785 (.A(net5786),
    .X(net5785));
 sg13g2_buf_2 fanout5786 (.A(net4244),
    .X(net5786));
 sg13g2_buf_2 fanout5787 (.A(net5789),
    .X(net5787));
 sg13g2_buf_2 fanout5788 (.A(net5789),
    .X(net5788));
 sg13g2_buf_2 fanout5789 (.A(net4254),
    .X(net5789));
 sg13g2_buf_2 fanout5790 (.A(net5791),
    .X(net5790));
 sg13g2_buf_2 fanout5791 (.A(\state[3] ),
    .X(net5791));
 sg13g2_buf_2 fanout5792 (.A(net5793),
    .X(net5792));
 sg13g2_buf_1 fanout5793 (.A(\state[3] ),
    .X(net5793));
 sg13g2_buf_2 fanout5794 (.A(net5796),
    .X(net5794));
 sg13g2_buf_2 fanout5795 (.A(net5796),
    .X(net5795));
 sg13g2_buf_2 fanout5796 (.A(\state[2] ),
    .X(net5796));
 sg13g2_buf_2 fanout5797 (.A(net5800),
    .X(net5797));
 sg13g2_buf_2 fanout5798 (.A(net5800),
    .X(net5798));
 sg13g2_buf_4 fanout5799 (.X(net5799),
    .A(net5800));
 sg13g2_buf_2 fanout5800 (.A(\state[1] ),
    .X(net5800));
 sg13g2_buf_8 fanout5801 (.A(\mem.addr[7] ),
    .X(net5801));
 sg13g2_buf_8 fanout5802 (.A(\mem.addr[6] ),
    .X(net5802));
 sg13g2_buf_2 fanout5803 (.A(\mem.addr[6] ),
    .X(net5803));
 sg13g2_buf_2 fanout5804 (.A(\mem.addr[4] ),
    .X(net5804));
 sg13g2_buf_2 fanout5805 (.A(\mem.addr[1] ),
    .X(net5805));
 sg13g2_buf_4 fanout5806 (.X(net5806),
    .A(\mem.addr[0] ));
 sg13g2_buf_4 fanout5807 (.X(net5807),
    .A(net5808));
 sg13g2_buf_4 fanout5808 (.X(net5808),
    .A(_00006_));
 sg13g2_buf_2 fanout5809 (.A(net5810),
    .X(net5809));
 sg13g2_buf_4 fanout5810 (.X(net5810),
    .A(net5811));
 sg13g2_buf_4 fanout5811 (.X(net5811),
    .A(_00005_));
 sg13g2_buf_2 fanout5812 (.A(net5813),
    .X(net5812));
 sg13g2_buf_2 fanout5813 (.A(net5814),
    .X(net5813));
 sg13g2_buf_2 fanout5814 (.A(net5815),
    .X(net5814));
 sg13g2_buf_4 fanout5815 (.X(net5815),
    .A(_00005_));
 sg13g2_buf_4 fanout5816 (.X(net5816),
    .A(net5819));
 sg13g2_buf_4 fanout5817 (.X(net5817),
    .A(net5819));
 sg13g2_buf_2 fanout5818 (.A(net5819),
    .X(net5818));
 sg13g2_buf_2 fanout5819 (.A(net5826),
    .X(net5819));
 sg13g2_buf_8 fanout5820 (.A(net5826),
    .X(net5820));
 sg13g2_buf_4 fanout5821 (.X(net5821),
    .A(net5822));
 sg13g2_buf_8 fanout5822 (.A(net5825),
    .X(net5822));
 sg13g2_buf_4 fanout5823 (.X(net5823),
    .A(net5824));
 sg13g2_buf_8 fanout5824 (.A(net5825),
    .X(net5824));
 sg13g2_buf_4 fanout5825 (.X(net5825),
    .A(net5826));
 sg13g2_buf_2 fanout5826 (.A(_00004_),
    .X(net5826));
 sg13g2_buf_4 fanout5827 (.X(net5827),
    .A(net5828));
 sg13g2_buf_8 fanout5828 (.A(net5837),
    .X(net5828));
 sg13g2_buf_2 fanout5829 (.A(net5837),
    .X(net5829));
 sg13g2_buf_2 fanout5830 (.A(net5837),
    .X(net5830));
 sg13g2_buf_4 fanout5831 (.X(net5831),
    .A(net5836));
 sg13g2_buf_2 fanout5832 (.A(net5836),
    .X(net5832));
 sg13g2_buf_4 fanout5833 (.X(net5833),
    .A(net5835));
 sg13g2_buf_2 fanout5834 (.A(net5835),
    .X(net5834));
 sg13g2_buf_4 fanout5835 (.X(net5835),
    .A(net5836));
 sg13g2_buf_4 fanout5836 (.X(net5836),
    .A(net5837));
 sg13g2_buf_4 fanout5837 (.X(net5837),
    .A(net5849));
 sg13g2_buf_8 fanout5838 (.A(net5842),
    .X(net5838));
 sg13g2_buf_2 fanout5839 (.A(net5842),
    .X(net5839));
 sg13g2_buf_4 fanout5840 (.X(net5840),
    .A(net5841));
 sg13g2_buf_4 fanout5841 (.X(net5841),
    .A(net5842));
 sg13g2_buf_4 fanout5842 (.X(net5842),
    .A(net5849));
 sg13g2_buf_4 fanout5843 (.X(net5843),
    .A(net5845));
 sg13g2_buf_2 fanout5844 (.A(net5845),
    .X(net5844));
 sg13g2_buf_4 fanout5845 (.X(net5845),
    .A(net5849));
 sg13g2_buf_4 fanout5846 (.X(net5846),
    .A(net5848));
 sg13g2_buf_4 fanout5847 (.X(net5847),
    .A(net5848));
 sg13g2_buf_4 fanout5848 (.X(net5848),
    .A(net5849));
 sg13g2_buf_8 fanout5849 (.A(_00003_),
    .X(net5849));
 sg13g2_buf_4 fanout5850 (.X(net5850),
    .A(net5856));
 sg13g2_buf_2 fanout5851 (.A(net5856),
    .X(net5851));
 sg13g2_buf_4 fanout5852 (.X(net5852),
    .A(net5853));
 sg13g2_buf_4 fanout5853 (.X(net5853),
    .A(net5856));
 sg13g2_buf_4 fanout5854 (.X(net5854),
    .A(net5855));
 sg13g2_buf_4 fanout5855 (.X(net5855),
    .A(net5856));
 sg13g2_buf_4 fanout5856 (.X(net5856),
    .A(net5884));
 sg13g2_buf_4 fanout5857 (.X(net5857),
    .A(net5860));
 sg13g2_buf_2 fanout5858 (.A(net5859),
    .X(net5858));
 sg13g2_buf_2 fanout5859 (.A(net5860),
    .X(net5859));
 sg13g2_buf_2 fanout5860 (.A(net5884),
    .X(net5860));
 sg13g2_buf_4 fanout5861 (.X(net5861),
    .A(net5864));
 sg13g2_buf_4 fanout5862 (.X(net5862),
    .A(net5863));
 sg13g2_buf_4 fanout5863 (.X(net5863),
    .A(net5864));
 sg13g2_buf_2 fanout5864 (.A(net5884),
    .X(net5864));
 sg13g2_buf_4 fanout5865 (.X(net5865),
    .A(net5874));
 sg13g2_buf_2 fanout5866 (.A(net5874),
    .X(net5866));
 sg13g2_buf_4 fanout5867 (.X(net5867),
    .A(net5868));
 sg13g2_buf_4 fanout5868 (.X(net5868),
    .A(net5874));
 sg13g2_buf_4 fanout5869 (.X(net5869),
    .A(net5873));
 sg13g2_buf_4 fanout5870 (.X(net5870),
    .A(net5873));
 sg13g2_buf_2 fanout5871 (.A(net5872),
    .X(net5871));
 sg13g2_buf_4 fanout5872 (.X(net5872),
    .A(net5873));
 sg13g2_buf_4 fanout5873 (.X(net5873),
    .A(net5874));
 sg13g2_buf_2 fanout5874 (.A(net5884),
    .X(net5874));
 sg13g2_buf_4 fanout5875 (.X(net5875),
    .A(net5883));
 sg13g2_buf_4 fanout5876 (.X(net5876),
    .A(net5883));
 sg13g2_buf_4 fanout5877 (.X(net5877),
    .A(net5879));
 sg13g2_buf_2 fanout5878 (.A(net5879),
    .X(net5878));
 sg13g2_buf_2 fanout5879 (.A(net5883),
    .X(net5879));
 sg13g2_buf_4 fanout5880 (.X(net5880),
    .A(net5883));
 sg13g2_buf_4 fanout5881 (.X(net5881),
    .A(net5882));
 sg13g2_buf_4 fanout5882 (.X(net5882),
    .A(net5883));
 sg13g2_buf_8 fanout5883 (.A(net5884),
    .X(net5883));
 sg13g2_buf_8 fanout5884 (.A(_00002_),
    .X(net5884));
 sg13g2_buf_4 fanout5885 (.X(net5885),
    .A(net5887));
 sg13g2_buf_4 fanout5886 (.X(net5886),
    .A(net5887));
 sg13g2_buf_2 fanout5887 (.A(net5914),
    .X(net5887));
 sg13g2_buf_2 fanout5888 (.A(net5891),
    .X(net5888));
 sg13g2_buf_2 fanout5889 (.A(net5891),
    .X(net5889));
 sg13g2_buf_4 fanout5890 (.X(net5890),
    .A(net5891));
 sg13g2_buf_2 fanout5891 (.A(net5914),
    .X(net5891));
 sg13g2_buf_2 fanout5892 (.A(net5894),
    .X(net5892));
 sg13g2_buf_1 fanout5893 (.A(net5894),
    .X(net5893));
 sg13g2_buf_2 fanout5894 (.A(net5896),
    .X(net5894));
 sg13g2_buf_4 fanout5895 (.X(net5895),
    .A(net5896));
 sg13g2_buf_2 fanout5896 (.A(net5900),
    .X(net5896));
 sg13g2_buf_4 fanout5897 (.X(net5897),
    .A(net5900));
 sg13g2_buf_2 fanout5898 (.A(net5899),
    .X(net5898));
 sg13g2_buf_2 fanout5899 (.A(net5900),
    .X(net5899));
 sg13g2_buf_2 fanout5900 (.A(net5914),
    .X(net5900));
 sg13g2_buf_4 fanout5901 (.X(net5901),
    .A(net5907));
 sg13g2_buf_2 fanout5902 (.A(net5907),
    .X(net5902));
 sg13g2_buf_2 fanout5903 (.A(net5907),
    .X(net5903));
 sg13g2_buf_2 fanout5904 (.A(net5907),
    .X(net5904));
 sg13g2_buf_2 fanout5905 (.A(net5906),
    .X(net5905));
 sg13g2_buf_2 fanout5906 (.A(net5907),
    .X(net5906));
 sg13g2_buf_2 fanout5907 (.A(net5914),
    .X(net5907));
 sg13g2_buf_2 fanout5908 (.A(net5913),
    .X(net5908));
 sg13g2_buf_2 fanout5909 (.A(net5913),
    .X(net5909));
 sg13g2_buf_2 fanout5910 (.A(net5913),
    .X(net5910));
 sg13g2_buf_2 fanout5911 (.A(net5913),
    .X(net5911));
 sg13g2_buf_2 fanout5912 (.A(net5913),
    .X(net5912));
 sg13g2_buf_2 fanout5913 (.A(net5914),
    .X(net5913));
 sg13g2_buf_4 fanout5914 (.X(net5914),
    .A(net6004));
 sg13g2_buf_4 fanout5915 (.X(net5915),
    .A(net5916));
 sg13g2_buf_4 fanout5916 (.X(net5916),
    .A(net5942));
 sg13g2_buf_4 fanout5917 (.X(net5917),
    .A(net5919));
 sg13g2_buf_4 fanout5918 (.X(net5918),
    .A(net5919));
 sg13g2_buf_2 fanout5919 (.A(net5942),
    .X(net5919));
 sg13g2_buf_4 fanout5920 (.X(net5920),
    .A(net5924));
 sg13g2_buf_4 fanout5921 (.X(net5921),
    .A(net5924));
 sg13g2_buf_4 fanout5922 (.X(net5922),
    .A(net5924));
 sg13g2_buf_2 fanout5923 (.A(net5924),
    .X(net5923));
 sg13g2_buf_2 fanout5924 (.A(net5942),
    .X(net5924));
 sg13g2_buf_2 fanout5925 (.A(net5932),
    .X(net5925));
 sg13g2_buf_2 fanout5926 (.A(net5932),
    .X(net5926));
 sg13g2_buf_4 fanout5927 (.X(net5927),
    .A(net5932));
 sg13g2_buf_4 fanout5928 (.X(net5928),
    .A(net5931));
 sg13g2_buf_1 fanout5929 (.A(net5931),
    .X(net5929));
 sg13g2_buf_2 fanout5930 (.A(net5931),
    .X(net5930));
 sg13g2_buf_2 fanout5931 (.A(net5932),
    .X(net5931));
 sg13g2_buf_2 fanout5932 (.A(net5941),
    .X(net5932));
 sg13g2_buf_4 fanout5933 (.X(net5933),
    .A(net5935));
 sg13g2_buf_2 fanout5934 (.A(net5941),
    .X(net5934));
 sg13g2_buf_2 fanout5935 (.A(net5941),
    .X(net5935));
 sg13g2_buf_4 fanout5936 (.X(net5936),
    .A(net5937));
 sg13g2_buf_4 fanout5937 (.X(net5937),
    .A(net5940));
 sg13g2_buf_2 fanout5938 (.A(net5940),
    .X(net5938));
 sg13g2_buf_2 fanout5939 (.A(net5940),
    .X(net5939));
 sg13g2_buf_2 fanout5940 (.A(net5941),
    .X(net5940));
 sg13g2_buf_2 fanout5941 (.A(net5942),
    .X(net5941));
 sg13g2_buf_2 fanout5942 (.A(net6004),
    .X(net5942));
 sg13g2_buf_4 fanout5943 (.X(net5943),
    .A(net5945));
 sg13g2_buf_4 fanout5944 (.X(net5944),
    .A(net5945));
 sg13g2_buf_4 fanout5945 (.X(net5945),
    .A(net5971));
 sg13g2_buf_2 fanout5946 (.A(net5949),
    .X(net5946));
 sg13g2_buf_4 fanout5947 (.X(net5947),
    .A(net5949));
 sg13g2_buf_2 fanout5948 (.A(net5949),
    .X(net5948));
 sg13g2_buf_2 fanout5949 (.A(net5971),
    .X(net5949));
 sg13g2_buf_4 fanout5950 (.X(net5950),
    .A(net5954));
 sg13g2_buf_4 fanout5951 (.X(net5951),
    .A(net5954));
 sg13g2_buf_4 fanout5952 (.X(net5952),
    .A(net5953));
 sg13g2_buf_4 fanout5953 (.X(net5953),
    .A(net5954));
 sg13g2_buf_2 fanout5954 (.A(net5971),
    .X(net5954));
 sg13g2_buf_4 fanout5955 (.X(net5955),
    .A(net5957));
 sg13g2_buf_1 fanout5956 (.A(net5957),
    .X(net5956));
 sg13g2_buf_4 fanout5957 (.X(net5957),
    .A(net5962));
 sg13g2_buf_2 fanout5958 (.A(net5961),
    .X(net5958));
 sg13g2_buf_4 fanout5959 (.X(net5959),
    .A(net5961));
 sg13g2_buf_2 fanout5960 (.A(net5961),
    .X(net5960));
 sg13g2_buf_2 fanout5961 (.A(net5962),
    .X(net5961));
 sg13g2_buf_2 fanout5962 (.A(net5971),
    .X(net5962));
 sg13g2_buf_4 fanout5963 (.X(net5963),
    .A(net5965));
 sg13g2_buf_4 fanout5964 (.X(net5964),
    .A(net5965));
 sg13g2_buf_2 fanout5965 (.A(net5971),
    .X(net5965));
 sg13g2_buf_4 fanout5966 (.X(net5966),
    .A(net5970));
 sg13g2_buf_1 fanout5967 (.A(net5970),
    .X(net5967));
 sg13g2_buf_4 fanout5968 (.X(net5968),
    .A(net5970));
 sg13g2_buf_2 fanout5969 (.A(net5970),
    .X(net5969));
 sg13g2_buf_2 fanout5970 (.A(net5971),
    .X(net5970));
 sg13g2_buf_4 fanout5971 (.X(net5971),
    .A(net6004));
 sg13g2_buf_4 fanout5972 (.X(net5972),
    .A(net5974));
 sg13g2_buf_4 fanout5973 (.X(net5973),
    .A(net5974));
 sg13g2_buf_2 fanout5974 (.A(net5986),
    .X(net5974));
 sg13g2_buf_4 fanout5975 (.X(net5975),
    .A(net5977));
 sg13g2_buf_4 fanout5976 (.X(net5976),
    .A(net5977));
 sg13g2_buf_2 fanout5977 (.A(net5986),
    .X(net5977));
 sg13g2_buf_4 fanout5978 (.X(net5978),
    .A(net5980));
 sg13g2_buf_2 fanout5979 (.A(net5980),
    .X(net5979));
 sg13g2_buf_2 fanout5980 (.A(net5986),
    .X(net5980));
 sg13g2_buf_4 fanout5981 (.X(net5981),
    .A(net5985));
 sg13g2_buf_1 fanout5982 (.A(net5985),
    .X(net5982));
 sg13g2_buf_4 fanout5983 (.X(net5983),
    .A(net5985));
 sg13g2_buf_2 fanout5984 (.A(net5985),
    .X(net5984));
 sg13g2_buf_2 fanout5985 (.A(net5986),
    .X(net5985));
 sg13g2_buf_4 fanout5986 (.X(net5986),
    .A(net6004));
 sg13g2_buf_2 fanout5987 (.A(net5988),
    .X(net5987));
 sg13g2_buf_2 fanout5988 (.A(net5989),
    .X(net5988));
 sg13g2_buf_4 fanout5989 (.X(net5989),
    .A(net6003));
 sg13g2_buf_2 fanout5990 (.A(net5994),
    .X(net5990));
 sg13g2_buf_2 fanout5991 (.A(net5994),
    .X(net5991));
 sg13g2_buf_2 fanout5992 (.A(net5993),
    .X(net5992));
 sg13g2_buf_4 fanout5993 (.X(net5993),
    .A(net5994));
 sg13g2_buf_2 fanout5994 (.A(net6003),
    .X(net5994));
 sg13g2_buf_4 fanout5995 (.X(net5995),
    .A(net5998));
 sg13g2_buf_4 fanout5996 (.X(net5996),
    .A(net5998));
 sg13g2_buf_1 fanout5997 (.A(net5998),
    .X(net5997));
 sg13g2_buf_2 fanout5998 (.A(net6003),
    .X(net5998));
 sg13g2_buf_4 fanout5999 (.X(net5999),
    .A(net6000));
 sg13g2_buf_4 fanout6000 (.X(net6000),
    .A(net6002));
 sg13g2_buf_4 fanout6001 (.X(net6001),
    .A(net6002));
 sg13g2_buf_2 fanout6002 (.A(net6003),
    .X(net6002));
 sg13g2_buf_4 fanout6003 (.X(net6003),
    .A(net6004));
 sg13g2_buf_8 fanout6004 (.A(_00001_),
    .X(net6004));
 sg13g2_buf_8 fanout6005 (.A(net6007),
    .X(net6005));
 sg13g2_buf_8 fanout6006 (.A(net6007),
    .X(net6006));
 sg13g2_buf_4 fanout6007 (.X(net6007),
    .A(net6014));
 sg13g2_buf_2 fanout6008 (.A(net6011),
    .X(net6008));
 sg13g2_buf_1 fanout6009 (.A(net6011),
    .X(net6009));
 sg13g2_buf_4 fanout6010 (.X(net6010),
    .A(net6011));
 sg13g2_buf_2 fanout6011 (.A(net6014),
    .X(net6011));
 sg13g2_buf_4 fanout6012 (.X(net6012),
    .A(net6014));
 sg13g2_buf_2 fanout6013 (.A(net6014),
    .X(net6013));
 sg13g2_buf_2 fanout6014 (.A(net6045),
    .X(net6014));
 sg13g2_buf_2 fanout6015 (.A(net6017),
    .X(net6015));
 sg13g2_buf_2 fanout6016 (.A(net6017),
    .X(net6016));
 sg13g2_buf_4 fanout6017 (.X(net6017),
    .A(net6020));
 sg13g2_buf_8 fanout6018 (.A(net6020),
    .X(net6018));
 sg13g2_buf_4 fanout6019 (.X(net6019),
    .A(net6020));
 sg13g2_buf_2 fanout6020 (.A(net6045),
    .X(net6020));
 sg13g2_buf_4 fanout6021 (.X(net6021),
    .A(net6025));
 sg13g2_buf_4 fanout6022 (.X(net6022),
    .A(net6025));
 sg13g2_buf_4 fanout6023 (.X(net6023),
    .A(net6024));
 sg13g2_buf_2 fanout6024 (.A(net6025),
    .X(net6024));
 sg13g2_buf_2 fanout6025 (.A(net6045),
    .X(net6025));
 sg13g2_buf_2 fanout6026 (.A(net6027),
    .X(net6026));
 sg13g2_buf_2 fanout6027 (.A(net6044),
    .X(net6027));
 sg13g2_buf_4 fanout6028 (.X(net6028),
    .A(net6044));
 sg13g2_buf_2 fanout6029 (.A(net6034),
    .X(net6029));
 sg13g2_buf_4 fanout6030 (.X(net6030),
    .A(net6034));
 sg13g2_buf_2 fanout6031 (.A(net6032),
    .X(net6031));
 sg13g2_buf_2 fanout6032 (.A(net6033),
    .X(net6032));
 sg13g2_buf_2 fanout6033 (.A(net6034),
    .X(net6033));
 sg13g2_buf_2 fanout6034 (.A(net6044),
    .X(net6034));
 sg13g2_buf_2 fanout6035 (.A(net6037),
    .X(net6035));
 sg13g2_buf_2 fanout6036 (.A(net6037),
    .X(net6036));
 sg13g2_buf_2 fanout6037 (.A(net6044),
    .X(net6037));
 sg13g2_buf_2 fanout6038 (.A(net6039),
    .X(net6038));
 sg13g2_buf_2 fanout6039 (.A(net6044),
    .X(net6039));
 sg13g2_buf_4 fanout6040 (.X(net6040),
    .A(net6043));
 sg13g2_buf_4 fanout6041 (.X(net6041),
    .A(net6043));
 sg13g2_buf_2 fanout6042 (.A(net6043),
    .X(net6042));
 sg13g2_buf_2 fanout6043 (.A(net6044),
    .X(net6043));
 sg13g2_buf_4 fanout6044 (.X(net6044),
    .A(net6045));
 sg13g2_buf_4 fanout6045 (.X(net6045),
    .A(net6174));
 sg13g2_buf_4 fanout6046 (.X(net6046),
    .A(net6049));
 sg13g2_buf_1 fanout6047 (.A(net6049),
    .X(net6047));
 sg13g2_buf_8 fanout6048 (.A(net6049),
    .X(net6048));
 sg13g2_buf_2 fanout6049 (.A(net6062),
    .X(net6049));
 sg13g2_buf_2 fanout6050 (.A(net6054),
    .X(net6050));
 sg13g2_buf_2 fanout6051 (.A(net6054),
    .X(net6051));
 sg13g2_buf_4 fanout6052 (.X(net6052),
    .A(net6053));
 sg13g2_buf_8 fanout6053 (.A(net6054),
    .X(net6053));
 sg13g2_buf_2 fanout6054 (.A(net6062),
    .X(net6054));
 sg13g2_buf_4 fanout6055 (.X(net6055),
    .A(net6057));
 sg13g2_buf_8 fanout6056 (.A(net6057),
    .X(net6056));
 sg13g2_buf_4 fanout6057 (.X(net6057),
    .A(net6062));
 sg13g2_buf_4 fanout6058 (.X(net6058),
    .A(net6061));
 sg13g2_buf_1 fanout6059 (.A(net6061),
    .X(net6059));
 sg13g2_buf_4 fanout6060 (.X(net6060),
    .A(net6061));
 sg13g2_buf_4 fanout6061 (.X(net6061),
    .A(net6062));
 sg13g2_buf_4 fanout6062 (.X(net6062),
    .A(net6174));
 sg13g2_buf_4 fanout6063 (.X(net6063),
    .A(net6073));
 sg13g2_buf_2 fanout6064 (.A(net6073),
    .X(net6064));
 sg13g2_buf_4 fanout6065 (.X(net6065),
    .A(net6067));
 sg13g2_buf_2 fanout6066 (.A(net6067),
    .X(net6066));
 sg13g2_buf_2 fanout6067 (.A(net6073),
    .X(net6067));
 sg13g2_buf_4 fanout6068 (.X(net6068),
    .A(net6070));
 sg13g2_buf_4 fanout6069 (.X(net6069),
    .A(net6073));
 sg13g2_buf_2 fanout6070 (.A(net6073),
    .X(net6070));
 sg13g2_buf_2 fanout6071 (.A(net6072),
    .X(net6071));
 sg13g2_buf_4 fanout6072 (.X(net6072),
    .A(net6073));
 sg13g2_buf_4 fanout6073 (.X(net6073),
    .A(net6084));
 sg13g2_buf_2 fanout6074 (.A(net6075),
    .X(net6074));
 sg13g2_buf_4 fanout6075 (.X(net6075),
    .A(net6078));
 sg13g2_buf_4 fanout6076 (.X(net6076),
    .A(net6077));
 sg13g2_buf_4 fanout6077 (.X(net6077),
    .A(net6078));
 sg13g2_buf_2 fanout6078 (.A(net6084),
    .X(net6078));
 sg13g2_buf_4 fanout6079 (.X(net6079),
    .A(net6080));
 sg13g2_buf_4 fanout6080 (.X(net6080),
    .A(net6084));
 sg13g2_buf_4 fanout6081 (.X(net6081),
    .A(net6083));
 sg13g2_buf_2 fanout6082 (.A(net6083),
    .X(net6082));
 sg13g2_buf_4 fanout6083 (.X(net6083),
    .A(net6084));
 sg13g2_buf_2 fanout6084 (.A(net6174),
    .X(net6084));
 sg13g2_buf_4 fanout6085 (.X(net6085),
    .A(net6089));
 sg13g2_buf_4 fanout6086 (.X(net6086),
    .A(net6089));
 sg13g2_buf_4 fanout6087 (.X(net6087),
    .A(net6089));
 sg13g2_buf_2 fanout6088 (.A(net6089),
    .X(net6088));
 sg13g2_buf_2 fanout6089 (.A(net6094),
    .X(net6089));
 sg13g2_buf_4 fanout6090 (.X(net6090),
    .A(net6091));
 sg13g2_buf_4 fanout6091 (.X(net6091),
    .A(net6094));
 sg13g2_buf_4 fanout6092 (.X(net6092),
    .A(net6093));
 sg13g2_buf_4 fanout6093 (.X(net6093),
    .A(net6094));
 sg13g2_buf_2 fanout6094 (.A(net6104),
    .X(net6094));
 sg13g2_buf_8 fanout6095 (.A(net6098),
    .X(net6095));
 sg13g2_buf_4 fanout6096 (.X(net6096),
    .A(net6097));
 sg13g2_buf_4 fanout6097 (.X(net6097),
    .A(net6098));
 sg13g2_buf_4 fanout6098 (.X(net6098),
    .A(net6104));
 sg13g2_buf_2 fanout6099 (.A(net6100),
    .X(net6099));
 sg13g2_buf_4 fanout6100 (.X(net6100),
    .A(net6104));
 sg13g2_buf_4 fanout6101 (.X(net6101),
    .A(net6103));
 sg13g2_buf_2 fanout6102 (.A(net6103),
    .X(net6102));
 sg13g2_buf_2 fanout6103 (.A(net6104),
    .X(net6103));
 sg13g2_buf_2 fanout6104 (.A(net6174),
    .X(net6104));
 sg13g2_buf_2 fanout6105 (.A(net6106),
    .X(net6105));
 sg13g2_buf_4 fanout6106 (.X(net6106),
    .A(net6115));
 sg13g2_buf_4 fanout6107 (.X(net6107),
    .A(net6115));
 sg13g2_buf_2 fanout6108 (.A(net6115),
    .X(net6108));
 sg13g2_buf_2 fanout6109 (.A(net6112),
    .X(net6109));
 sg13g2_buf_4 fanout6110 (.X(net6110),
    .A(net6112));
 sg13g2_buf_2 fanout6111 (.A(net6112),
    .X(net6111));
 sg13g2_buf_2 fanout6112 (.A(net6115),
    .X(net6112));
 sg13g2_buf_4 fanout6113 (.X(net6113),
    .A(net6114));
 sg13g2_buf_4 fanout6114 (.X(net6114),
    .A(net6115));
 sg13g2_buf_4 fanout6115 (.X(net6115),
    .A(net6129));
 sg13g2_buf_4 fanout6116 (.X(net6116),
    .A(net6120));
 sg13g2_buf_4 fanout6117 (.X(net6117),
    .A(net6120));
 sg13g2_buf_2 fanout6118 (.A(net6119),
    .X(net6118));
 sg13g2_buf_4 fanout6119 (.X(net6119),
    .A(net6120));
 sg13g2_buf_2 fanout6120 (.A(net6129),
    .X(net6120));
 sg13g2_buf_4 fanout6121 (.X(net6121),
    .A(net6124));
 sg13g2_buf_4 fanout6122 (.X(net6122),
    .A(net6124));
 sg13g2_buf_1 fanout6123 (.A(net6124),
    .X(net6123));
 sg13g2_buf_2 fanout6124 (.A(net6129),
    .X(net6124));
 sg13g2_buf_4 fanout6125 (.X(net6125),
    .A(net6128));
 sg13g2_buf_2 fanout6126 (.A(net6127),
    .X(net6126));
 sg13g2_buf_4 fanout6127 (.X(net6127),
    .A(net6128));
 sg13g2_buf_2 fanout6128 (.A(net6129),
    .X(net6128));
 sg13g2_buf_2 fanout6129 (.A(net6174),
    .X(net6129));
 sg13g2_buf_8 fanout6130 (.A(net6133),
    .X(net6130));
 sg13g2_buf_2 fanout6131 (.A(net6133),
    .X(net6131));
 sg13g2_buf_4 fanout6132 (.X(net6132),
    .A(net6133));
 sg13g2_buf_4 fanout6133 (.X(net6133),
    .A(net6173));
 sg13g2_buf_4 fanout6134 (.X(net6134),
    .A(net6137));
 sg13g2_buf_4 fanout6135 (.X(net6135),
    .A(net6137));
 sg13g2_buf_2 fanout6136 (.A(net6137),
    .X(net6136));
 sg13g2_buf_4 fanout6137 (.X(net6137),
    .A(net6173));
 sg13g2_buf_8 fanout6138 (.A(net6148),
    .X(net6138));
 sg13g2_buf_4 fanout6139 (.X(net6139),
    .A(net6148));
 sg13g2_buf_4 fanout6140 (.X(net6140),
    .A(net6141));
 sg13g2_buf_4 fanout6141 (.X(net6141),
    .A(net6148));
 sg13g2_buf_2 fanout6142 (.A(net6144),
    .X(net6142));
 sg13g2_buf_2 fanout6143 (.A(net6144),
    .X(net6143));
 sg13g2_buf_2 fanout6144 (.A(net6148),
    .X(net6144));
 sg13g2_buf_4 fanout6145 (.X(net6145),
    .A(net6147));
 sg13g2_buf_4 fanout6146 (.X(net6146),
    .A(net6147));
 sg13g2_buf_2 fanout6147 (.A(net6148),
    .X(net6147));
 sg13g2_buf_4 fanout6148 (.X(net6148),
    .A(net6173));
 sg13g2_buf_2 fanout6149 (.A(net6151),
    .X(net6149));
 sg13g2_buf_1 fanout6150 (.A(net6151),
    .X(net6150));
 sg13g2_buf_2 fanout6151 (.A(net6154),
    .X(net6151));
 sg13g2_buf_4 fanout6152 (.X(net6152),
    .A(net6153));
 sg13g2_buf_4 fanout6153 (.X(net6153),
    .A(net6154));
 sg13g2_buf_2 fanout6154 (.A(net6172),
    .X(net6154));
 sg13g2_buf_2 fanout6155 (.A(net6157),
    .X(net6155));
 sg13g2_buf_4 fanout6156 (.X(net6156),
    .A(net6157));
 sg13g2_buf_2 fanout6157 (.A(net6172),
    .X(net6157));
 sg13g2_buf_2 fanout6158 (.A(net6160),
    .X(net6158));
 sg13g2_buf_4 fanout6159 (.X(net6159),
    .A(net6160));
 sg13g2_buf_2 fanout6160 (.A(net6172),
    .X(net6160));
 sg13g2_buf_4 fanout6161 (.X(net6161),
    .A(net6162));
 sg13g2_buf_4 fanout6162 (.X(net6162),
    .A(net6165));
 sg13g2_buf_4 fanout6163 (.X(net6163),
    .A(net6164));
 sg13g2_buf_4 fanout6164 (.X(net6164),
    .A(net6165));
 sg13g2_buf_2 fanout6165 (.A(net6172),
    .X(net6165));
 sg13g2_buf_4 fanout6166 (.X(net6166),
    .A(net6169));
 sg13g2_buf_4 fanout6167 (.X(net6167),
    .A(net6169));
 sg13g2_buf_1 fanout6168 (.A(net6169),
    .X(net6168));
 sg13g2_buf_2 fanout6169 (.A(net6172),
    .X(net6169));
 sg13g2_buf_2 fanout6170 (.A(net6171),
    .X(net6170));
 sg13g2_buf_4 fanout6171 (.X(net6171),
    .A(net6172));
 sg13g2_buf_4 fanout6172 (.X(net6172),
    .A(net6173));
 sg13g2_buf_4 fanout6173 (.X(net6173),
    .A(net6174));
 sg13g2_buf_8 fanout6174 (.A(_00000_),
    .X(net6174));
 sg13g2_buf_2 fanout6175 (.A(net6178),
    .X(net6175));
 sg13g2_buf_2 fanout6176 (.A(net6178),
    .X(net6176));
 sg13g2_buf_2 fanout6177 (.A(net6178),
    .X(net6177));
 sg13g2_buf_2 fanout6178 (.A(_02883_),
    .X(net6178));
 sg13g2_buf_2 fanout6179 (.A(net6180),
    .X(net6179));
 sg13g2_buf_2 fanout6180 (.A(uio_in[2]),
    .X(net6180));
 sg13g2_buf_2 fanout6181 (.A(net1),
    .X(net6181));
 sg13g2_buf_2 fanout6182 (.A(net6189),
    .X(net6182));
 sg13g2_buf_2 fanout6183 (.A(net6186),
    .X(net6183));
 sg13g2_buf_2 fanout6184 (.A(net6186),
    .X(net6184));
 sg13g2_buf_2 fanout6185 (.A(net6186),
    .X(net6185));
 sg13g2_buf_1 fanout6186 (.A(net6189),
    .X(net6186));
 sg13g2_buf_2 fanout6187 (.A(net6188),
    .X(net6187));
 sg13g2_buf_2 fanout6188 (.A(net6189),
    .X(net6188));
 sg13g2_buf_2 fanout6189 (.A(net6190),
    .X(net6189));
 sg13g2_buf_2 fanout6190 (.A(net1),
    .X(net6190));
 sg13g2_buf_4 input1 (.X(net1),
    .A(rst_n));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[0]));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[1]));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[2]));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[3]));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[4]));
 sg13g2_buf_4 input7 (.X(net7),
    .A(ui_in[5]));
 sg13g2_buf_4 input8 (.X(net8),
    .A(ui_in[6]));
 sg13g2_buf_4 input9 (.X(net9),
    .A(ui_in[7]));
 sg13g2_buf_4 input10 (.X(net10),
    .A(uio_in[0]));
 sg13g2_buf_4 input11 (.X(net11),
    .A(uio_in[3]));
 sg13g2_tielo tt_um_urish_sic1_12 (.L_LO(net12));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_6_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_6_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_6_3_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_6_3_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_6_6_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_6_6_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_6_6_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_6_4_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_6_1_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_6_1_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_6_4_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_6_4_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_6_4_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_6_5_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_6_5_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_6_5_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_6_5_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_6_7_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_6_7_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_6_7_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_6_6_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_6_7_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_6_12_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_6_12_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_6_12_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_6_24_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_6_24_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_6_13_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_6_13_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_6_26_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_6_26_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_6_24_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_6_24_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_6_24_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_6_25_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_6_25_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_6_19_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_6_19_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_6_18_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_6_18_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_6_18_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_6_18_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_6_17_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_6_17_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_6_17_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_6_19_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_6_19_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_6_22_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_6_20_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_6_20_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_6_17_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_6_20_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_6_20_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_6_21_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_6_21_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_6_21_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_6_21_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_6_23_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_6_23_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_6_23_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_6_23_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_6_22_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_6_22_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_6_22_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_6_28_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_6_28_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_6_29_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_6_29_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_6_29_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_6_29_0_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_6_31_0_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_6_31_0_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_6_31_0_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_6_31_0_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_leaf_82_clk (.A(clknet_6_30_0_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_2 clkbuf_leaf_83_clk (.A(clknet_6_30_0_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_2 clkbuf_leaf_84_clk (.A(clknet_6_30_0_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_2 clkbuf_leaf_85_clk (.A(clknet_6_30_0_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_2 clkbuf_leaf_86_clk (.A(clknet_6_28_0_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_2 clkbuf_leaf_87_clk (.A(clknet_6_28_0_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_2 clkbuf_leaf_88_clk (.A(clknet_6_25_0_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_2 clkbuf_leaf_89_clk (.A(clknet_6_25_0_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_2 clkbuf_leaf_90_clk (.A(clknet_6_27_0_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_2 clkbuf_leaf_91_clk (.A(clknet_6_27_0_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_2 clkbuf_leaf_92_clk (.A(clknet_6_27_0_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_2 clkbuf_leaf_93_clk (.A(clknet_6_27_0_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_2 clkbuf_leaf_94_clk (.A(clknet_6_26_0_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_2 clkbuf_leaf_95_clk (.A(clknet_6_26_0_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_2 clkbuf_leaf_96_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_2 clkbuf_leaf_97_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_2 clkbuf_leaf_98_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_2 clkbuf_leaf_99_clk (.A(clknet_6_49_0_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_2 clkbuf_leaf_100_clk (.A(clknet_6_49_0_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_2 clkbuf_leaf_101_clk (.A(clknet_6_49_0_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_2 clkbuf_leaf_102_clk (.A(clknet_6_51_0_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_2 clkbuf_leaf_103_clk (.A(clknet_6_51_0_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_2 clkbuf_leaf_104_clk (.A(clknet_6_54_0_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_2 clkbuf_leaf_105_clk (.A(clknet_6_54_0_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_2 clkbuf_leaf_106_clk (.A(clknet_6_49_0_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_2 clkbuf_leaf_107_clk (.A(clknet_6_52_0_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_2 clkbuf_leaf_108_clk (.A(clknet_6_52_0_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_2 clkbuf_leaf_109_clk (.A(clknet_6_52_0_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_2 clkbuf_leaf_110_clk (.A(clknet_6_52_0_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_2 clkbuf_leaf_111_clk (.A(clknet_6_53_0_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_2 clkbuf_leaf_112_clk (.A(clknet_6_53_0_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_2 clkbuf_leaf_113_clk (.A(clknet_6_53_0_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_2 clkbuf_leaf_114_clk (.A(clknet_6_53_0_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_2 clkbuf_leaf_115_clk (.A(clknet_6_55_0_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_2 clkbuf_leaf_116_clk (.A(clknet_6_55_0_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_2 clkbuf_leaf_117_clk (.A(clknet_6_55_0_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_2 clkbuf_leaf_118_clk (.A(clknet_6_55_0_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_2 clkbuf_leaf_119_clk (.A(clknet_6_54_0_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_2 clkbuf_leaf_120_clk (.A(clknet_6_54_0_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_2 clkbuf_leaf_121_clk (.A(clknet_6_60_0_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_2 clkbuf_leaf_122_clk (.A(clknet_6_60_0_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_2 clkbuf_leaf_123_clk (.A(clknet_6_61_0_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_2 clkbuf_leaf_124_clk (.A(clknet_6_61_0_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_2 clkbuf_leaf_125_clk (.A(clknet_6_61_0_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_2 clkbuf_leaf_126_clk (.A(clknet_6_61_0_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_2 clkbuf_leaf_127_clk (.A(clknet_6_63_0_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_2 clkbuf_leaf_128_clk (.A(clknet_6_63_0_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_2 clkbuf_leaf_129_clk (.A(clknet_6_63_0_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_2 clkbuf_leaf_130_clk (.A(clknet_6_63_0_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_2 clkbuf_leaf_131_clk (.A(clknet_6_62_0_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_2 clkbuf_leaf_132_clk (.A(clknet_6_62_0_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_2 clkbuf_leaf_133_clk (.A(clknet_6_62_0_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_2 clkbuf_leaf_134_clk (.A(clknet_6_62_0_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_2 clkbuf_leaf_135_clk (.A(clknet_6_60_0_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_2 clkbuf_leaf_136_clk (.A(clknet_6_60_0_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_2 clkbuf_leaf_137_clk (.A(clknet_6_57_0_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_2 clkbuf_leaf_138_clk (.A(clknet_6_59_0_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_2 clkbuf_leaf_139_clk (.A(clknet_6_59_0_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_2 clkbuf_leaf_140_clk (.A(clknet_6_59_0_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_2 clkbuf_leaf_141_clk (.A(clknet_6_59_0_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_2 clkbuf_leaf_142_clk (.A(clknet_6_58_0_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_2 clkbuf_leaf_143_clk (.A(clknet_6_58_0_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_2 clkbuf_leaf_144_clk (.A(clknet_6_58_0_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_2 clkbuf_leaf_145_clk (.A(clknet_6_58_0_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_2 clkbuf_leaf_146_clk (.A(clknet_6_56_0_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_2 clkbuf_leaf_147_clk (.A(clknet_6_56_0_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_2 clkbuf_leaf_148_clk (.A(clknet_6_56_0_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_2 clkbuf_leaf_149_clk (.A(clknet_6_56_0_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_2 clkbuf_leaf_150_clk (.A(clknet_6_57_0_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_2 clkbuf_leaf_151_clk (.A(clknet_6_57_0_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_2 clkbuf_leaf_152_clk (.A(clknet_6_57_0_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_2 clkbuf_leaf_153_clk (.A(clknet_6_51_0_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_2 clkbuf_leaf_154_clk (.A(clknet_6_51_0_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_2 clkbuf_leaf_155_clk (.A(clknet_6_56_0_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_2 clkbuf_leaf_156_clk (.A(clknet_6_50_0_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_2 clkbuf_leaf_157_clk (.A(clknet_6_50_0_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_2 clkbuf_leaf_158_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_2 clkbuf_leaf_159_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_2 clkbuf_leaf_160_clk (.A(clknet_6_37_0_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_2 clkbuf_leaf_161_clk (.A(clknet_6_37_0_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_2 clkbuf_leaf_162_clk (.A(clknet_6_50_0_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_2 clkbuf_leaf_163_clk (.A(clknet_6_50_0_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_2 clkbuf_leaf_164_clk (.A(clknet_6_39_0_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_2 clkbuf_leaf_165_clk (.A(clknet_6_39_0_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_2 clkbuf_leaf_166_clk (.A(clknet_6_39_0_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_2 clkbuf_leaf_167_clk (.A(clknet_6_39_0_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_2 clkbuf_leaf_168_clk (.A(clknet_6_44_0_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_2 clkbuf_leaf_169_clk (.A(clknet_6_44_0_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_2 clkbuf_leaf_170_clk (.A(clknet_6_44_0_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_2 clkbuf_leaf_171_clk (.A(clknet_6_45_0_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_2 clkbuf_leaf_172_clk (.A(clknet_6_45_0_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_2 clkbuf_leaf_173_clk (.A(clknet_6_45_0_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_2 clkbuf_leaf_174_clk (.A(clknet_6_45_0_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_2 clkbuf_leaf_175_clk (.A(clknet_6_47_0_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_2 clkbuf_leaf_176_clk (.A(clknet_6_47_0_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_2 clkbuf_leaf_177_clk (.A(clknet_6_47_0_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_2 clkbuf_leaf_178_clk (.A(clknet_6_47_0_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_2 clkbuf_leaf_179_clk (.A(clknet_6_46_0_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_2 clkbuf_leaf_180_clk (.A(clknet_6_46_0_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_2 clkbuf_leaf_181_clk (.A(clknet_6_46_0_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_2 clkbuf_leaf_182_clk (.A(clknet_6_46_0_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_2 clkbuf_leaf_183_clk (.A(clknet_6_44_0_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_2 clkbuf_leaf_184_clk (.A(clknet_6_41_0_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_2 clkbuf_leaf_185_clk (.A(clknet_6_41_0_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_2 clkbuf_leaf_186_clk (.A(clknet_6_43_0_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_2 clkbuf_leaf_187_clk (.A(clknet_6_43_0_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_2 clkbuf_leaf_188_clk (.A(clknet_6_43_0_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_2 clkbuf_leaf_189_clk (.A(clknet_6_43_0_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_2 clkbuf_leaf_190_clk (.A(clknet_6_42_0_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_2 clkbuf_leaf_191_clk (.A(clknet_6_42_0_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_2 clkbuf_leaf_192_clk (.A(clknet_6_42_0_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_2 clkbuf_leaf_193_clk (.A(clknet_6_42_0_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_2 clkbuf_leaf_194_clk (.A(clknet_6_40_0_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_2 clkbuf_leaf_195_clk (.A(clknet_6_40_0_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_2 clkbuf_leaf_196_clk (.A(clknet_6_40_0_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_2 clkbuf_leaf_197_clk (.A(clknet_6_40_0_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_2 clkbuf_leaf_198_clk (.A(clknet_6_40_0_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_2 clkbuf_leaf_199_clk (.A(clknet_6_41_0_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_2 clkbuf_leaf_200_clk (.A(clknet_6_41_0_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_2 clkbuf_leaf_201_clk (.A(clknet_6_35_0_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_2 clkbuf_leaf_202_clk (.A(clknet_6_35_0_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_2 clkbuf_leaf_203_clk (.A(clknet_6_35_0_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_2 clkbuf_leaf_204_clk (.A(clknet_6_35_0_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_2 clkbuf_leaf_205_clk (.A(clknet_6_34_0_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_2 clkbuf_leaf_206_clk (.A(clknet_6_34_0_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_2 clkbuf_leaf_207_clk (.A(clknet_6_34_0_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_2 clkbuf_leaf_208_clk (.A(clknet_6_34_0_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_2 clkbuf_leaf_209_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_2 clkbuf_leaf_210_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_2 clkbuf_leaf_211_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_2 clkbuf_leaf_212_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_2 clkbuf_leaf_213_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_2 clkbuf_leaf_214_clk (.A(clknet_6_33_0_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_2 clkbuf_leaf_215_clk (.A(clknet_6_33_0_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_2 clkbuf_leaf_216_clk (.A(clknet_6_33_0_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_2 clkbuf_leaf_217_clk (.A(clknet_6_33_0_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_2 clkbuf_leaf_218_clk (.A(clknet_6_38_0_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_2 clkbuf_leaf_219_clk (.A(clknet_6_38_0_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_2 clkbuf_leaf_220_clk (.A(clknet_6_38_0_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_2 clkbuf_leaf_221_clk (.A(clknet_6_38_0_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_2 clkbuf_leaf_222_clk (.A(clknet_6_36_0_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_2 clkbuf_leaf_223_clk (.A(clknet_6_36_0_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_2 clkbuf_leaf_224_clk (.A(clknet_6_36_0_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_2 clkbuf_leaf_225_clk (.A(clknet_6_36_0_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_2 clkbuf_leaf_226_clk (.A(clknet_6_37_0_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_2 clkbuf_leaf_227_clk (.A(clknet_6_37_0_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_2 clkbuf_leaf_228_clk (.A(clknet_6_15_0_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_2 clkbuf_leaf_229_clk (.A(clknet_6_15_0_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_2 clkbuf_leaf_230_clk (.A(clknet_6_15_0_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_2 clkbuf_leaf_231_clk (.A(clknet_6_14_0_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_2 clkbuf_leaf_232_clk (.A(clknet_6_15_0_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_2 clkbuf_leaf_233_clk (.A(clknet_6_14_0_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_2 clkbuf_leaf_234_clk (.A(clknet_6_13_0_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_2 clkbuf_leaf_235_clk (.A(clknet_6_13_0_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_2 clkbuf_leaf_236_clk (.A(clknet_6_12_0_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_2 clkbuf_leaf_237_clk (.A(clknet_6_9_0_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_2 clkbuf_leaf_238_clk (.A(clknet_6_9_0_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_2 clkbuf_leaf_239_clk (.A(clknet_6_11_0_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_2 clkbuf_leaf_240_clk (.A(clknet_6_14_0_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_2 clkbuf_leaf_241_clk (.A(clknet_6_14_0_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_2 clkbuf_leaf_242_clk (.A(clknet_6_11_0_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_2 clkbuf_leaf_243_clk (.A(clknet_6_11_0_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_2 clkbuf_leaf_244_clk (.A(clknet_6_11_0_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_2 clkbuf_leaf_245_clk (.A(clknet_6_10_0_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_2 clkbuf_leaf_246_clk (.A(clknet_6_10_0_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_2 clkbuf_leaf_247_clk (.A(clknet_6_10_0_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_2 clkbuf_leaf_248_clk (.A(clknet_6_10_0_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_2 clkbuf_leaf_249_clk (.A(clknet_6_8_0_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_2 clkbuf_leaf_250_clk (.A(clknet_6_8_0_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_2 clkbuf_leaf_251_clk (.A(clknet_6_8_0_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_2 clkbuf_leaf_252_clk (.A(clknet_6_8_0_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_2 clkbuf_leaf_253_clk (.A(clknet_6_9_0_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_2 clkbuf_leaf_254_clk (.A(clknet_6_9_0_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_2 clkbuf_leaf_255_clk (.A(clknet_6_3_0_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_2 clkbuf_leaf_256_clk (.A(clknet_6_3_0_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_2 clkbuf_leaf_257_clk (.A(clknet_6_8_0_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_2 clkbuf_leaf_258_clk (.A(clknet_6_2_0_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_2 clkbuf_leaf_259_clk (.A(clknet_6_2_0_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_2 clkbuf_leaf_260_clk (.A(clknet_6_2_0_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_2 clkbuf_leaf_261_clk (.A(clknet_6_2_0_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_2 clkbuf_leaf_262_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_2 clkbuf_leaf_263_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_2 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_2 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_2 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_2 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_2 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_2 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_2 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_2 clkbuf_6_0_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_0_0_clk));
 sg13g2_buf_2 clkbuf_6_1_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_1_0_clk));
 sg13g2_buf_2 clkbuf_6_2_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_2_0_clk));
 sg13g2_buf_2 clkbuf_6_3_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_3_0_clk));
 sg13g2_buf_2 clkbuf_6_4_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_4_0_clk));
 sg13g2_buf_2 clkbuf_6_5_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_5_0_clk));
 sg13g2_buf_2 clkbuf_6_6_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_6_0_clk));
 sg13g2_buf_2 clkbuf_6_7_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_7_0_clk));
 sg13g2_buf_2 clkbuf_6_8_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_8_0_clk));
 sg13g2_buf_2 clkbuf_6_9_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_9_0_clk));
 sg13g2_buf_2 clkbuf_6_10_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_10_0_clk));
 sg13g2_buf_2 clkbuf_6_11_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_11_0_clk));
 sg13g2_buf_2 clkbuf_6_12_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_12_0_clk));
 sg13g2_buf_2 clkbuf_6_13_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_13_0_clk));
 sg13g2_buf_2 clkbuf_6_14_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_14_0_clk));
 sg13g2_buf_2 clkbuf_6_15_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_15_0_clk));
 sg13g2_buf_2 clkbuf_6_16_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_16_0_clk));
 sg13g2_buf_2 clkbuf_6_17_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_17_0_clk));
 sg13g2_buf_2 clkbuf_6_18_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_18_0_clk));
 sg13g2_buf_2 clkbuf_6_19_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_19_0_clk));
 sg13g2_buf_2 clkbuf_6_20_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_20_0_clk));
 sg13g2_buf_2 clkbuf_6_21_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_21_0_clk));
 sg13g2_buf_2 clkbuf_6_22_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_22_0_clk));
 sg13g2_buf_2 clkbuf_6_23_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_23_0_clk));
 sg13g2_buf_2 clkbuf_6_24_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_24_0_clk));
 sg13g2_buf_2 clkbuf_6_25_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_25_0_clk));
 sg13g2_buf_2 clkbuf_6_26_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_26_0_clk));
 sg13g2_buf_2 clkbuf_6_27_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_27_0_clk));
 sg13g2_buf_2 clkbuf_6_28_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_28_0_clk));
 sg13g2_buf_2 clkbuf_6_29_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_29_0_clk));
 sg13g2_buf_2 clkbuf_6_30_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_30_0_clk));
 sg13g2_buf_2 clkbuf_6_31_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_31_0_clk));
 sg13g2_buf_2 clkbuf_6_32_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_32_0_clk));
 sg13g2_buf_2 clkbuf_6_33_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_33_0_clk));
 sg13g2_buf_2 clkbuf_6_34_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_34_0_clk));
 sg13g2_buf_2 clkbuf_6_35_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_35_0_clk));
 sg13g2_buf_2 clkbuf_6_36_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_36_0_clk));
 sg13g2_buf_2 clkbuf_6_37_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_37_0_clk));
 sg13g2_buf_2 clkbuf_6_38_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_38_0_clk));
 sg13g2_buf_2 clkbuf_6_39_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_39_0_clk));
 sg13g2_buf_2 clkbuf_6_40_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_40_0_clk));
 sg13g2_buf_2 clkbuf_6_41_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_41_0_clk));
 sg13g2_buf_2 clkbuf_6_42_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_42_0_clk));
 sg13g2_buf_2 clkbuf_6_43_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_43_0_clk));
 sg13g2_buf_2 clkbuf_6_44_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_44_0_clk));
 sg13g2_buf_2 clkbuf_6_45_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_45_0_clk));
 sg13g2_buf_2 clkbuf_6_46_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_46_0_clk));
 sg13g2_buf_2 clkbuf_6_47_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_47_0_clk));
 sg13g2_buf_2 clkbuf_6_48_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_48_0_clk));
 sg13g2_buf_2 clkbuf_6_49_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_49_0_clk));
 sg13g2_buf_2 clkbuf_6_50_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_50_0_clk));
 sg13g2_buf_2 clkbuf_6_51_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_51_0_clk));
 sg13g2_buf_2 clkbuf_6_52_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_52_0_clk));
 sg13g2_buf_2 clkbuf_6_53_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_53_0_clk));
 sg13g2_buf_2 clkbuf_6_54_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_54_0_clk));
 sg13g2_buf_2 clkbuf_6_55_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_55_0_clk));
 sg13g2_buf_2 clkbuf_6_56_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_56_0_clk));
 sg13g2_buf_2 clkbuf_6_57_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_57_0_clk));
 sg13g2_buf_2 clkbuf_6_58_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_58_0_clk));
 sg13g2_buf_2 clkbuf_6_59_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_59_0_clk));
 sg13g2_buf_2 clkbuf_6_60_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_60_0_clk));
 sg13g2_buf_2 clkbuf_6_61_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_61_0_clk));
 sg13g2_buf_2 clkbuf_6_62_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_62_0_clk));
 sg13g2_buf_2 clkbuf_6_63_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_63_0_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_6_1_0_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_6_2_0_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_6_3_0_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_6_4_0_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_6_5_0_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_6_6_0_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_6_7_0_clk));
 sg13g2_buf_2 clkload7 (.A(clknet_6_9_0_clk));
 sg13g2_buf_2 clkload8 (.A(clknet_6_10_0_clk));
 sg13g2_buf_2 clkload9 (.A(clknet_6_11_0_clk));
 sg13g2_buf_2 clkload10 (.A(clknet_6_12_0_clk));
 sg13g2_buf_2 clkload11 (.A(clknet_6_13_0_clk));
 sg13g2_buf_2 clkload12 (.A(clknet_6_14_0_clk));
 sg13g2_buf_2 clkload13 (.A(clknet_6_15_0_clk));
 sg13g2_buf_2 clkload14 (.A(clknet_6_17_0_clk));
 sg13g2_buf_2 clkload15 (.A(clknet_6_18_0_clk));
 sg13g2_buf_2 clkload16 (.A(clknet_6_19_0_clk));
 sg13g2_buf_2 clkload17 (.A(clknet_6_20_0_clk));
 sg13g2_buf_2 clkload18 (.A(clknet_6_21_0_clk));
 sg13g2_buf_2 clkload19 (.A(clknet_6_22_0_clk));
 sg13g2_buf_2 clkload20 (.A(clknet_6_23_0_clk));
 sg13g2_buf_2 clkload21 (.A(clknet_6_25_0_clk));
 sg13g2_buf_2 clkload22 (.A(clknet_6_26_0_clk));
 sg13g2_buf_2 clkload23 (.A(clknet_6_27_0_clk));
 sg13g2_buf_2 clkload24 (.A(clknet_6_28_0_clk));
 sg13g2_buf_2 clkload25 (.A(clknet_6_29_0_clk));
 sg13g2_buf_2 clkload26 (.A(clknet_6_30_0_clk));
 sg13g2_buf_2 clkload27 (.A(clknet_6_31_0_clk));
 sg13g2_buf_2 clkload28 (.A(clknet_6_33_0_clk));
 sg13g2_buf_2 clkload29 (.A(clknet_6_34_0_clk));
 sg13g2_buf_2 clkload30 (.A(clknet_6_35_0_clk));
 sg13g2_buf_2 clkload31 (.A(clknet_6_36_0_clk));
 sg13g2_buf_2 clkload32 (.A(clknet_6_37_0_clk));
 sg13g2_buf_2 clkload33 (.A(clknet_6_38_0_clk));
 sg13g2_buf_2 clkload34 (.A(clknet_6_39_0_clk));
 sg13g2_buf_2 clkload35 (.A(clknet_6_41_0_clk));
 sg13g2_buf_2 clkload36 (.A(clknet_6_42_0_clk));
 sg13g2_buf_2 clkload37 (.A(clknet_6_43_0_clk));
 sg13g2_buf_2 clkload38 (.A(clknet_6_44_0_clk));
 sg13g2_buf_2 clkload39 (.A(clknet_6_45_0_clk));
 sg13g2_buf_2 clkload40 (.A(clknet_6_46_0_clk));
 sg13g2_buf_2 clkload41 (.A(clknet_6_47_0_clk));
 sg13g2_buf_2 clkload42 (.A(clknet_6_49_0_clk));
 sg13g2_buf_2 clkload43 (.A(clknet_6_50_0_clk));
 sg13g2_buf_2 clkload44 (.A(clknet_6_51_0_clk));
 sg13g2_buf_2 clkload45 (.A(clknet_6_52_0_clk));
 sg13g2_buf_2 clkload46 (.A(clknet_6_53_0_clk));
 sg13g2_buf_2 clkload47 (.A(clknet_6_54_0_clk));
 sg13g2_buf_2 clkload48 (.A(clknet_6_55_0_clk));
 sg13g2_buf_2 clkload49 (.A(clknet_6_57_0_clk));
 sg13g2_buf_2 clkload50 (.A(clknet_6_58_0_clk));
 sg13g2_buf_2 clkload51 (.A(clknet_6_59_0_clk));
 sg13g2_buf_2 clkload52 (.A(clknet_6_60_0_clk));
 sg13g2_buf_2 clkload53 (.A(clknet_6_61_0_clk));
 sg13g2_buf_2 clkload54 (.A(clknet_6_62_0_clk));
 sg13g2_buf_2 clkload55 (.A(clknet_6_63_0_clk));
 sg13g2_inv_4 clkload56 (.A(clknet_leaf_263_clk));
 sg13g2_inv_1 clkload57 (.A(clknet_leaf_160_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mem.mem[220][5] ),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mem.mem[100][0] ),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mem.mem[180][3] ),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold4 (.A(\mem.mem[172][3] ),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mem.mem[154][7] ),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mem.mem[226][3] ),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold7 (.A(\mem.wr_en ),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold8 (.A(_00804_),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mem.mem[236][6] ),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold10 (.A(\mem.mem[110][0] ),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold11 (.A(\mem.mem[52][0] ),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mem.mem[170][3] ),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mem.mem[148][4] ),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold14 (.A(\mem.mem[188][3] ),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold15 (.A(\mem.mem[148][3] ),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold16 (.A(\mem.mem[128][6] ),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold17 (.A(\mem.mem[96][0] ),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold18 (.A(\mem.mem[148][7] ),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold19 (.A(\mem.mem[188][7] ),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold20 (.A(\mem.mem[180][7] ),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold21 (.A(\mem.mem[84][0] ),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold22 (.A(\mem.mem[168][3] ),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold23 (.A(\mem.mem[192][4] ),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold24 (.A(\mem.mem[224][3] ),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold25 (.A(\mem.mem[222][1] ),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold26 (.A(\mem.mem[56][0] ),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold27 (.A(\mem.mem[158][1] ),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold28 (.A(\mem.mem[156][7] ),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold29 (.A(\mem.mem[86][0] ),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold30 (.A(\mem.mem[208][5] ),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold31 (.A(\mem.mem[54][0] ),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold32 (.A(\mem.mem[164][3] ),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold33 (.A(\mem.mem[30][0] ),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold34 (.A(\mem.mem[126][1] ),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold35 (.A(\mem.mem[164][7] ),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mem.mem[86][7] ),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mem.mem[236][7] ),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold38 (.A(\mem.mem[58][0] ),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold39 (.A(\mem.mem[166][3] ),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold40 (.A(\mem.mem[232][4] ),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold41 (.A(\mem.mem[184][4] ),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold42 (.A(\mem.mem[46][3] ),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold43 (.A(\mem.mem[92][0] ),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold44 (.A(\mem.mem[46][0] ),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold45 (.A(\mem.mem[114][0] ),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold46 (.A(\mem.mem[228][3] ),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold47 (.A(\mem.mem[110][3] ),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold48 (.A(\mem.mem[228][6] ),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold49 (.A(\mem.mem[160][7] ),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold50 (.A(\mem.mem[184][3] ),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold51 (.A(\mem.mem[46][2] ),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold52 (.A(\mem.mem[52][1] ),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold53 (.A(\mem.mem[186][0] ),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold54 (.A(\mem.mem[60][1] ),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold55 (.A(\mem.mem[88][1] ),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold56 (.A(\mem.mem[64][0] ),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold57 (.A(\mem.mem[186][4] ),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold58 (.A(\mem.mem[233][1] ),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mem.mem[126][6] ),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold60 (.A(\mem.mem[188][5] ),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mem.mem[60][0] ),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold62 (.A(\mem.mem[85][7] ),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mem.mem[210][6] ),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold64 (.A(\mem.mem[55][1] ),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mem.mem[231][0] ),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold66 (.A(\mem.mem[192][5] ),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mem.mem[179][7] ),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold68 (.A(\mem.mem[80][3] ),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold69 (.A(\mem.mem[116][0] ),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold70 (.A(\mem.mem[186][3] ),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold71 (.A(\mem.mem[231][3] ),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold72 (.A(\mem.mem[122][7] ),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold73 (.A(\mem.mem[90][2] ),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold74 (.A(\mem.mem[177][1] ),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold75 (.A(\mem.mem[220][1] ),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold76 (.A(\mem.mem[50][3] ),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold77 (.A(\mem.mem[150][1] ),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold78 (.A(\mem.mem[108][6] ),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold79 (.A(\mem.mem[114][3] ),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold80 (.A(\mem.mem[71][0] ),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold81 (.A(\mem.mem[39][2] ),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold82 (.A(\mem.mem[215][4] ),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold83 (.A(\mem.mem[192][0] ),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold84 (.A(\mem.mem[235][2] ),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold85 (.A(\mem.mem[158][7] ),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold86 (.A(\mem.mem[122][4] ),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold87 (.A(\mem.mem[234][1] ),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold88 (.A(\mem.mem[71][2] ),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold89 (.A(\mem.mem[246][5] ),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold90 (.A(\mem.mem[119][5] ),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold91 (.A(\mem.mem[93][3] ),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold92 (.A(\mem.mem[246][1] ),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold93 (.A(\mem.mem[89][6] ),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold94 (.A(\mem.mem[88][7] ),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mem.mem[154][0] ),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold96 (.A(\mem.mem[108][7] ),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold97 (.A(\mem.mem[183][4] ),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold98 (.A(\mem.mem[212][4] ),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold99 (.A(\mem.mem[214][2] ),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold100 (.A(\mem.mem[108][1] ),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold101 (.A(\mem.mem[182][3] ),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mem.mem[128][0] ),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold103 (.A(\mem.mem[210][4] ),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold104 (.A(\mem.mem[32][0] ),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold105 (.A(\mem.mem[54][4] ),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold106 (.A(\mem.mem[124][6] ),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold107 (.A(\mem.mem[45][0] ),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold108 (.A(\mem.mem[122][5] ),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold109 (.A(\mem.mem[104][1] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold110 (.A(\mem.mem[212][0] ),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold111 (.A(\mem.mem[58][5] ),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold112 (.A(\mem.mem[80][6] ),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold113 (.A(\mem.mem[62][6] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold114 (.A(\mem.mem[50][6] ),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold115 (.A(\mem.mem[124][3] ),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold116 (.A(\mem.mem[211][3] ),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold117 (.A(\mem.mem[189][4] ),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold118 (.A(\mem.mem[238][1] ),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold119 (.A(\mem.mem[224][6] ),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold120 (.A(\mem.mem[235][6] ),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold121 (.A(\mem.mem[233][2] ),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold122 (.A(\mem.mem[32][5] ),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold123 (.A(\mem.mem[7][5] ),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold124 (.A(\mem.mem[59][4] ),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold125 (.A(\mem.mem[152][7] ),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold126 (.A(\mem.mem[112][7] ),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold127 (.A(\mem.mem[226][7] ),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold128 (.A(\mem.mem[51][0] ),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold129 (.A(\mem.mem[43][1] ),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold130 (.A(\mem.mem[108][0] ),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold131 (.A(\mem.mem[55][6] ),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold132 (.A(\mem.mem[238][3] ),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold133 (.A(\mem.mem[29][7] ),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold134 (.A(\mem.mem[156][0] ),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold135 (.A(\mem.mem[147][2] ),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold136 (.A(\mem.mem[192][2] ),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold137 (.A(\mem.mem[217][7] ),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold138 (.A(\mem.mem[7][3] ),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold139 (.A(\mem.mem[96][6] ),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold140 (.A(\mem.mem[32][1] ),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold141 (.A(\mem.mem[210][5] ),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold142 (.A(\mem.mem[0][5] ),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold143 (.A(\mem.mem[120][6] ),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold144 (.A(\mem.mem[125][6] ),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold145 (.A(\mem.mem[228][5] ),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold146 (.A(\mem.mem[109][3] ),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold147 (.A(\mem.mem[16][5] ),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold148 (.A(\mem.mem[123][3] ),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold149 (.A(\mem.mem[60][5] ),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold150 (.A(\mem.mem[232][0] ),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mem.mem[214][3] ),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold152 (.A(\mem.mem[90][4] ),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold153 (.A(\mem.mem[58][3] ),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold154 (.A(\mem.mem[172][7] ),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold155 (.A(\mem.mem[237][1] ),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold156 (.A(\mem.mem[89][7] ),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold157 (.A(\mem.mem[58][1] ),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold158 (.A(\mem.mem[158][6] ),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold159 (.A(\mem.mem[222][4] ),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold160 (.A(\mem.mem[125][1] ),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold161 (.A(\mem.mem[64][5] ),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold162 (.A(\mem.mem[94][3] ),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold163 (.A(\mem.mem[229][7] ),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold164 (.A(\mem.mem[121][3] ),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold165 (.A(\mem.mem[16][4] ),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold166 (.A(\mem.mem[23][0] ),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold167 (.A(\mem.mem[246][7] ),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold168 (.A(\mem.mem[45][1] ),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold169 (.A(\mem.mem[118][2] ),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold170 (.A(\mem.mem[166][1] ),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold171 (.A(\mem.mem[103][0] ),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold172 (.A(\mem.mem[94][1] ),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold173 (.A(\mem.mem[221][7] ),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold174 (.A(\mem.mem[229][0] ),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold175 (.A(\mem.mem[225][0] ),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold176 (.A(\mem.mem[91][5] ),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold177 (.A(\mem.mem[229][4] ),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold178 (.A(\mem.mem[86][1] ),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold179 (.A(\mem.mem[221][3] ),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold180 (.A(\mem.mem[156][4] ),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold181 (.A(\mem.mem[92][6] ),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold182 (.A(\mem.mem[166][0] ),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold183 (.A(\mem.mem[86][4] ),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold184 (.A(\mem.mem[220][7] ),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold185 (.A(\mem.mem[238][6] ),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold186 (.A(\mem.mem[103][6] ),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold187 (.A(\mem.mem[55][5] ),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold188 (.A(\mem.mem[102][6] ),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold189 (.A(\mem.mem[237][2] ),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold190 (.A(\mem.mem[149][2] ),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold191 (.A(\mem.mem[50][2] ),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold192 (.A(\mem.mem[100][6] ),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold193 (.A(\mem.mem[55][2] ),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold194 (.A(\mem.mem[94][4] ),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold195 (.A(\mem.mem[92][7] ),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold196 (.A(\mem.mem[216][7] ),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold197 (.A(\mem.mem[90][5] ),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold198 (.A(\mem.mem[221][2] ),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold199 (.A(\mem.mem[54][5] ),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold200 (.A(\mem.mem[16][7] ),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold201 (.A(\mem.mem[104][0] ),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold202 (.A(\mem.mem[157][0] ),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold203 (.A(\mem.mem[212][1] ),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold204 (.A(\mem.mem[126][7] ),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold205 (.A(\mem.mem[57][1] ),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold206 (.A(\mem.mem[30][1] ),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold207 (.A(\mem.mem[241][3] ),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold208 (.A(\mem.mem[53][7] ),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold209 (.A(\mem.mem[192][6] ),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold210 (.A(\mem.mem[32][4] ),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold211 (.A(\mem.mem[233][6] ),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold212 (.A(\mem.mem[104][3] ),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold213 (.A(\mem.mem[172][2] ),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold214 (.A(\mem.mem[7][1] ),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold215 (.A(\mem.mem[213][5] ),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold216 (.A(\mem.mem[225][5] ),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold217 (.A(\mem.mem[114][2] ),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold218 (.A(\mem.mem[208][6] ),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold219 (.A(\mem.mem[57][5] ),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold220 (.A(\mem.mem[48][3] ),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold221 (.A(\mem.mem[215][6] ),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold222 (.A(\mem.mem[32][2] ),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold223 (.A(\mem.mem[100][2] ),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold224 (.A(\mem.mem[236][0] ),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold225 (.A(\mem.mem[225][1] ),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold226 (.A(\mem.mem[46][6] ),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold227 (.A(\mem.mem[85][4] ),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold228 (.A(\mem.mem[125][7] ),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold229 (.A(\mem.mem[228][0] ),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold230 (.A(\mem.mem[61][3] ),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold231 (.A(\mem.mem[86][5] ),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold232 (.A(\mem.mem[174][0] ),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold233 (.A(\mem.mem[187][4] ),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold234 (.A(\mem.mem[100][1] ),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold235 (.A(\mem.mem[241][2] ),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold236 (.A(\mem.mem[163][1] ),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold237 (.A(\mem.mem[100][5] ),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold238 (.A(\mem.mem[245][2] ),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold239 (.A(\mem.mem[55][4] ),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold240 (.A(\mem.mem[199][7] ),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold241 (.A(\mem.mem[51][2] ),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold242 (.A(\mem.mem[109][2] ),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold243 (.A(\mem.mem[215][3] ),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold244 (.A(\mem.mem[163][3] ),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold245 (.A(\mem.mem[91][0] ),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold246 (.A(\mem.mem[48][2] ),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold247 (.A(\mem.mem[7][4] ),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold248 (.A(\mem.mem[224][5] ),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold249 (.A(\mem.mem[91][1] ),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold250 (.A(\mem.mem[178][1] ),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold251 (.A(\mem.mem[59][3] ),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold252 (.A(\mem.mem[112][1] ),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold253 (.A(\mem.mem[103][3] ),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold254 (.A(\mem.mem[180][4] ),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold255 (.A(\mem.mem[178][2] ),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold256 (.A(\mem.mem[48][4] ),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold257 (.A(\mem.mem[165][4] ),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold258 (.A(\mem.mem[246][2] ),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold259 (.A(\mem.mem[125][4] ),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold260 (.A(\mem.mem[120][0] ),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold261 (.A(\mem.mem[231][6] ),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold262 (.A(\mem.mem[221][4] ),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold263 (.A(\mem.mem[23][2] ),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold264 (.A(\mem.mem[184][1] ),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold265 (.A(\mem.mem[236][4] ),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold266 (.A(\mem.mem[242][1] ),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold267 (.A(\mem.mem[230][7] ),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold268 (.A(\mem.mem[71][5] ),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold269 (.A(\mem.mem[219][4] ),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold270 (.A(\mem.mem[83][7] ),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold271 (.A(\mem.mem[215][2] ),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold272 (.A(\mem.mem[245][5] ),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold273 (.A(\mem.mem[53][3] ),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold274 (.A(\mem.mem[229][5] ),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold275 (.A(\mem.mem[112][3] ),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold276 (.A(\mem.mem[186][1] ),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold277 (.A(\mem.mem[157][2] ),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold278 (.A(\mem.mem[221][0] ),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold279 (.A(\mem.mem[173][2] ),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold280 (.A(\mem.mem[116][3] ),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold281 (.A(\mem.mem[168][2] ),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold282 (.A(\mem.mem[188][4] ),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold283 (.A(\mem.mem[113][3] ),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold284 (.A(\mem.mem[39][5] ),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold285 (.A(\mem.mem[237][0] ),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold286 (.A(\mem.mem[249][1] ),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold287 (.A(\mem.mem[187][6] ),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold288 (.A(\mem.mem[190][1] ),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold289 (.A(\mem.mem[48][1] ),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold290 (.A(\mem.mem[119][0] ),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold291 (.A(\mem.mem[242][2] ),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold292 (.A(\mem.mem[43][5] ),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold293 (.A(\mem.mem[90][1] ),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold294 (.A(\mem.mem[107][3] ),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold295 (.A(\mem.mem[51][3] ),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold296 (.A(\mem.mem[182][0] ),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold297 (.A(\mem.mem[216][5] ),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold298 (.A(\mem.mem[165][3] ),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold299 (.A(\mem.mem[241][5] ),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold300 (.A(\mem.mem[113][5] ),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold301 (.A(\mem.mem[225][2] ),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold302 (.A(\mem.mem[230][6] ),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold303 (.A(\mem.mem[231][4] ),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold304 (.A(\mem.mem[119][3] ),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold305 (.A(\mem.mem[153][1] ),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold306 (.A(\mem.mem[56][3] ),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold307 (.A(\mem.mem[209][7] ),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold308 (.A(\mem.mem[218][6] ),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold309 (.A(\mem.mem[108][2] ),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold310 (.A(\mem.mem[217][5] ),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold311 (.A(\mem.mem[249][6] ),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold312 (.A(\mem.mem[117][6] ),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold313 (.A(\mem.mem[220][0] ),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold314 (.A(\mem.mem[169][2] ),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold315 (.A(\mem.mem[84][4] ),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold316 (.A(\mem.mem[114][4] ),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold317 (.A(\mem.mem[184][7] ),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold318 (.A(\mem.mem[49][1] ),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold319 (.A(\mem.mem[101][5] ),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold320 (.A(\mem.mem[188][6] ),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold321 (.A(\mem.mem[58][6] ),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold322 (.A(\mem.mem[227][1] ),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold323 (.A(\mem.mem[91][3] ),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold324 (.A(\mem.mem[50][1] ),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold325 (.A(\mem.mem[99][5] ),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold326 (.A(\mem.mem[169][3] ),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold327 (.A(\mem.mem[103][5] ),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold328 (.A(\mem.mem[232][2] ),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold329 (.A(\mem.mem[39][7] ),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold330 (.A(\mem.mem[32][6] ),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold331 (.A(\mem.mem[30][6] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold332 (.A(\mem.mem[148][2] ),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold333 (.A(\mem.mem[209][0] ),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold334 (.A(\mem.mem[23][3] ),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold335 (.A(\mem.mem[150][5] ),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold336 (.A(\mem.mem[86][3] ),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold337 (.A(\mem.mem[84][6] ),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold338 (.A(\mem.mem[208][3] ),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold339 (.A(\mem.mem[158][0] ),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold340 (.A(\mem.mem[103][1] ),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold341 (.A(\mem.mem[180][6] ),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold342 (.A(\mem.mem[112][0] ),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold343 (.A(\mem.mem[29][1] ),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold344 (.A(\mem.mem[234][4] ),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold345 (.A(\mem.mem[217][2] ),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold346 (.A(\mem.mem[247][5] ),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold347 (.A(\mem.mem[215][1] ),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold348 (.A(\mem.mem[213][6] ),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold349 (.A(\mem.mem[51][7] ),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold350 (.A(\mem.mem[222][7] ),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold351 (.A(\mem.mem[118][3] ),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold352 (.A(\mem.mem[221][5] ),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold353 (.A(\mem.mem[177][3] ),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold354 (.A(\mem.mem[166][5] ),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold355 (.A(\mem.mem[185][2] ),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold356 (.A(\mem.mem[236][1] ),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold357 (.A(\mem.mem[168][0] ),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold358 (.A(\mem.mem[99][0] ),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold359 (.A(\mem.mem[213][3] ),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold360 (.A(\mem.mem[39][1] ),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold361 (.A(\mem.mem[167][2] ),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold362 (.A(\mem.mem[152][0] ),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold363 (.A(\mem.mem[27][4] ),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold364 (.A(\mem.mem[114][6] ),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold365 (.A(\mem.mem[90][7] ),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold366 (.A(\mem.mem[116][2] ),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold367 (.A(\mem.mem[232][6] ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold368 (.A(\mem.mem[123][0] ),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold369 (.A(\mem.mem[190][4] ),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold370 (.A(\mem.mem[226][0] ),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold371 (.A(\mem.mem[236][5] ),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold372 (.A(\mem.mem[182][5] ),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold373 (.A(\mem.mem[124][5] ),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold374 (.A(\mem.mem[228][2] ),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold375 (.A(\mem.mem[84][5] ),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold376 (.A(\mem.mem[171][1] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold377 (.A(\mem.mem[220][4] ),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold378 (.A(\mem.mem[213][7] ),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold379 (.A(\mem.mem[222][5] ),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold380 (.A(\mem.mem[128][7] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold381 (.A(\mem.mem[151][0] ),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold382 (.A(\mem.mem[80][4] ),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold383 (.A(\mem.mem[151][2] ),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold384 (.A(\mem.mem[71][3] ),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold385 (.A(\mem.mem[61][5] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold386 (.A(\mem.mem[238][5] ),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold387 (.A(\mem.mem[185][4] ),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold388 (.A(\mem.mem[7][2] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold389 (.A(\mem.mem[51][5] ),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold390 (.A(\mem.mem[179][5] ),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold391 (.A(\mem.mem[108][4] ),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold392 (.A(\mem.mem[119][6] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold393 (.A(\mem.mem[157][6] ),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold394 (.A(\mem.mem[245][4] ),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold395 (.A(\mem.mem[170][6] ),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold396 (.A(\mem.mem[176][6] ),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold397 (.A(\mem.mem[231][7] ),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold398 (.A(\mem.mem[154][2] ),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold399 (.A(\mem.mem[241][6] ),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold400 (.A(\mem.mem[234][7] ),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold401 (.A(\mem.mem[112][4] ),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold402 (.A(\mem.mem[115][0] ),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold403 (.A(\mem.mem[48][7] ),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold404 (.A(\mem.mem[171][7] ),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold405 (.A(\mem.mem[123][1] ),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold406 (.A(\mem.mem[106][3] ),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold407 (.A(\mem.mem[212][6] ),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold408 (.A(\mem.mem[124][2] ),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold409 (.A(\mem.mem[104][4] ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold410 (.A(\mem.mem[208][2] ),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold411 (.A(\mem.mem[181][1] ),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold412 (.A(\mem.mem[105][1] ),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold413 (.A(\mem.mem[213][2] ),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold414 (.A(\mem.mem[29][2] ),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold415 (.A(\mem.mem[92][1] ),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold416 (.A(\mem.mem[90][0] ),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold417 (.A(\mem.mem[163][6] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold418 (.A(\mem.mem[219][2] ),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold419 (.A(\mem.mem[85][2] ),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold420 (.A(\mem.mem[160][5] ),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold421 (.A(\mem.mem[171][0] ),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold422 (.A(\mem.mem[167][5] ),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold423 (.A(\mem.mem[183][0] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold424 (.A(\mem.mem[247][2] ),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold425 (.A(\mem.mem[50][5] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold426 (.A(\mem.mem[245][6] ),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold427 (.A(\mem.mem[23][5] ),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold428 (.A(\mem.mem[199][6] ),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold429 (.A(\mem.mem[123][6] ),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold430 (.A(\mem.mem[247][4] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold431 (.A(\mem.mem[105][7] ),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold432 (.A(\mem.mem[220][3] ),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold433 (.A(\mem.mem[247][3] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold434 (.A(\mem.mem[144][1] ),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold435 (.A(\mem.mem[49][7] ),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold436 (.A(\mem.mem[151][4] ),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold437 (.A(\mem.mem[230][5] ),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold438 (.A(\mem.mem[190][6] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold439 (.A(\mem.mem[250][6] ),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold440 (.A(\mem.mem[233][3] ),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold441 (.A(\mem.mem[149][1] ),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold442 (.A(\mem.mem[89][3] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold443 (.A(\mem.mem[229][2] ),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold444 (.A(\mem.mem[180][0] ),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold445 (.A(\mem.mem[209][1] ),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold446 (.A(\mem.mem[119][4] ),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold447 (.A(\mem.mem[226][1] ),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold448 (.A(\mem.mem[164][0] ),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold449 (.A(\mem.mem[242][0] ),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold450 (.A(\mem.mem[178][3] ),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold451 (.A(\mem.mem[147][6] ),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold452 (.A(\mem.mem[71][6] ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold453 (.A(\mem.mem[115][1] ),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold454 (.A(\mem.mem[187][2] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold455 (.A(\mem.mem[183][6] ),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold456 (.A(\mem.mem[228][4] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold457 (.A(\mem.mem[154][4] ),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold458 (.A(\mem.mem[216][1] ),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold459 (.A(\mem.mem[49][6] ),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold460 (.A(\mem.mem[119][1] ),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold461 (.A(\mem.mem[182][2] ),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold462 (.A(\mem.mem[212][3] ),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold463 (.A(\mem.mem[118][4] ),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold464 (.A(\mem.mem[180][5] ),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold465 (.A(\mem.mem[216][6] ),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold466 (.A(\mem.mem[71][4] ),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold467 (.A(\mem.mem[224][7] ),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold468 (.A(\mem.mem[94][7] ),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold469 (.A(\mem.mem[55][7] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold470 (.A(\mem.mem[233][0] ),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold471 (.A(\mem.mem[113][7] ),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold472 (.A(\mem.mem[160][3] ),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold473 (.A(\mem.mem[144][4] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold474 (.A(\mem.mem[147][7] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold475 (.A(\mem.mem[96][1] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold476 (.A(\mem.mem[102][5] ),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold477 (.A(\mem.mem[158][5] ),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold478 (.A(\mem.mem[238][4] ),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold479 (.A(\mem.mem[176][7] ),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold480 (.A(\mem.mem[54][2] ),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold481 (.A(\mem.mem[29][3] ),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold482 (.A(\mem.mem[249][2] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold483 (.A(\mem.mem[163][4] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold484 (.A(\mem.mem[177][5] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold485 (.A(\mem.mem[105][6] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold486 (.A(\mem.mem[168][4] ),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold487 (.A(\mem.mem[249][4] ),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold488 (.A(\mem.mem[96][3] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold489 (.A(\mem.mem[114][5] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold490 (.A(\mem.mem[106][1] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold491 (.A(\mem.mem[155][2] ),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold492 (.A(\mem.mem[54][7] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold493 (.A(\mem.mem[174][1] ),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold494 (.A(\mem.mem[61][2] ),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold495 (.A(\mem.mem[153][4] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold496 (.A(\mem.mem[209][6] ),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold497 (.A(\mem.mem[155][5] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold498 (.A(\mem.mem[176][2] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold499 (.A(\mem.mem[227][4] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold500 (.A(\mem.mem[123][5] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold501 (.A(\mem.mem[93][5] ),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold502 (.A(\mem.mem[64][6] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold503 (.A(\mem.mem[246][4] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold504 (.A(\mem.mem[117][4] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold505 (.A(\mem.mem[121][0] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold506 (.A(\mem.mem[124][7] ),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold507 (.A(\mem.mem[121][7] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold508 (.A(\mem.mem[186][5] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold509 (.A(\mem.mem[185][0] ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold510 (.A(\mem.mem[85][5] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold511 (.A(\mem.mem[90][6] ),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold512 (.A(\mem.mem[177][2] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold513 (.A(\mem.mem[182][1] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold514 (.A(\mem.mem[179][1] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold515 (.A(\mem.mem[23][7] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold516 (.A(\mem.mem[238][7] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold517 (.A(\mem.mem[92][5] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold518 (.A(\mem.mem[237][7] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold519 (.A(\mem.mem[210][3] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold520 (.A(\mem.mem[89][4] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold521 (.A(\mem.mem[144][2] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold522 (.A(\mem.mem[107][5] ),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold523 (.A(\mem.mem[135][5] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold524 (.A(\mem.mem[160][2] ),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold525 (.A(\mem.mem[211][0] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold526 (.A(\mem.mem[53][6] ),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold527 (.A(\mem.mem[225][4] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold528 (.A(\mem.mem[105][3] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold529 (.A(\mem.mem[45][3] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold530 (.A(\mem.mem[179][0] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold531 (.A(\mem.mem[188][2] ),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold532 (.A(\mem.mem[46][4] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold533 (.A(\mem.mem[222][3] ),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold534 (.A(\mem.mem[183][7] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold535 (.A(\mem.mem[242][4] ),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold536 (.A(\mem.mem[238][0] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold537 (.A(\mem.mem[99][7] ),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold538 (.A(\mem.mem[187][5] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold539 (.A(\mem.mem[178][6] ),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold540 (.A(\mem.mem[172][0] ),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold541 (.A(\mem.mem[56][2] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold542 (.A(\mem.mem[236][2] ),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold543 (.A(\mem.mem[91][6] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold544 (.A(\mem.mem[88][2] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold545 (.A(\mem.mem[128][3] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold546 (.A(\mem.mem[59][6] ),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold547 (.A(\mem.mem[121][2] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold548 (.A(\mem.mem[221][6] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold549 (.A(\mem.mem[173][4] ),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold550 (.A(\mem.mem[0][0] ),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold551 (.A(\mem.mem[118][6] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold552 (.A(\mem.mem[178][0] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold553 (.A(\mem.mem[165][0] ),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold554 (.A(\mem.mem[250][4] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold555 (.A(\mem.mem[212][7] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold556 (.A(\mem.mem[176][5] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold557 (.A(\mem.mem[177][0] ),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold558 (.A(\mem.mem[30][3] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold559 (.A(\mem.mem[117][7] ),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold560 (.A(\mem.mem[222][2] ),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold561 (.A(\mem.mem[100][7] ),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold562 (.A(\mem.mem[208][0] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold563 (.A(\mem.mem[173][1] ),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold564 (.A(\mem.mem[115][4] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold565 (.A(\mem.mem[210][1] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold566 (.A(\mem.mem[169][6] ),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold567 (.A(\mem.mem[58][7] ),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold568 (.A(\mem.mem[186][2] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold569 (.A(\mem.mem[160][4] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold570 (.A(\mem.mem[148][1] ),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold571 (.A(\mem.mem[213][0] ),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold572 (.A(\mem.mem[181][0] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold573 (.A(\mem.mem[227][5] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold574 (.A(\mem.mem[182][6] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold575 (.A(\mem.mem[224][0] ),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold576 (.A(\mem.mem[235][3] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold577 (.A(\mem.mem[112][5] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold578 (.A(\mem.mem[153][3] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold579 (.A(\mem.mem[96][4] ),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold580 (.A(\mem.mem[215][0] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold581 (.A(\mem.mem[44][6] ),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold582 (.A(\mem.mem[54][3] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold583 (.A(\mem.mem[119][2] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold584 (.A(\mem.mem[184][0] ),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold585 (.A(\mem.mem[165][2] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold586 (.A(\mem.mem[122][2] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold587 (.A(\mem.mem[23][1] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold588 (.A(\mem.mem[128][5] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold589 (.A(\mem.mem[170][5] ),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold590 (.A(\mem.mem[181][2] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold591 (.A(\mem.mem[199][1] ),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold592 (.A(\mem.mem[115][2] ),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold593 (.A(\mem.mem[184][2] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold594 (.A(\mem.mem[154][6] ),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold595 (.A(\mem.mem[164][1] ),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold596 (.A(\mem.mem[110][6] ),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold597 (.A(\mem.mem[184][6] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold598 (.A(\mem.mem[246][3] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold599 (.A(\mem.mem[120][7] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold600 (.A(\mem.mem[176][0] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold601 (.A(\mem.mem[59][1] ),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold602 (.A(\mem.mem[103][4] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold603 (.A(\mem.mem[186][6] ),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold604 (.A(\mem.mem[110][5] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold605 (.A(\mem.mem[237][3] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold606 (.A(\mem.mem[59][5] ),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold607 (.A(\mem.mem[57][7] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold608 (.A(\mem.mem[169][1] ),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold609 (.A(\mem.mem[106][5] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold610 (.A(\mem.mem[45][5] ),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold611 (.A(\mem.mem[247][7] ),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold612 (.A(\mem.mem[140][3] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold613 (.A(\mem.mem[176][4] ),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold614 (.A(\mem.mem[170][4] ),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold615 (.A(\mem.mem[93][6] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold616 (.A(\mem.mem[124][1] ),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold617 (.A(\mem.mem[211][2] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold618 (.A(\mem.mem[181][3] ),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold619 (.A(\mem.mem[103][2] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold620 (.A(\mem.mem[165][1] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold621 (.A(\mem.mem[174][4] ),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold622 (.A(\mem.mem[230][4] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold623 (.A(\mem.mem[218][4] ),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold624 (.A(\mem.mem[0][3] ),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold625 (.A(\mem.mem[189][7] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold626 (.A(\mem.mem[99][2] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold627 (.A(\mem.mem[249][0] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold628 (.A(\mem.mem[107][2] ),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold629 (.A(\mem.mem[115][7] ),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold630 (.A(\mem.mem[102][4] ),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold631 (.A(\mem.mem[164][4] ),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold632 (.A(\mem.mem[209][2] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold633 (.A(\mem.mem[91][4] ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold634 (.A(\mem.mem[157][1] ),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold635 (.A(\mem.mem[241][4] ),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold636 (.A(\mem.mem[23][6] ),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold637 (.A(\mem.mem[85][1] ),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold638 (.A(\mem.mem[218][0] ),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold639 (.A(\mem.mem[46][7] ),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold640 (.A(\mem.mem[4][0] ),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold641 (.A(\mem.mem[158][2] ),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold642 (.A(\mem.mem[114][7] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold643 (.A(\mem.mem[192][1] ),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold644 (.A(\mem.mem[169][7] ),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold645 (.A(\mem.mem[178][4] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold646 (.A(\mem.mem[98][0] ),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold647 (.A(\mem.mem[157][4] ),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold648 (.A(\mem.mem[155][7] ),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold649 (.A(\mem.mem[211][7] ),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold650 (.A(\mem.mem[217][1] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold651 (.A(\mem.mem[186][7] ),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold652 (.A(\mem.mem[155][1] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold653 (.A(\mem.mem[199][2] ),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold654 (.A(\mem.mem[247][6] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold655 (.A(\mem.mem[50][0] ),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold656 (.A(\mem.mem[171][5] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold657 (.A(\mem.mem[48][5] ),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold658 (.A(\mem.mem[126][2] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold659 (.A(\mem.mem[105][0] ),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold660 (.A(\mem.mem[61][1] ),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold661 (.A(\mem.mem[187][1] ),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold662 (.A(\mem.mem[52][7] ),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold663 (.A(\mem.mem[22][1] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold664 (.A(\mem.mem[219][3] ),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold665 (.A(\mem.mem[116][6] ),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold666 (.A(\mem.mem[165][5] ),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold667 (.A(\mem.mem[209][3] ),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold668 (.A(\mem.mem[227][7] ),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold669 (.A(\mem.mem[105][4] ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold670 (.A(\mem.mem[62][4] ),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold671 (.A(\mem.mem[230][0] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold672 (.A(\mem.mem[150][2] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold673 (.A(\mem.mem[120][5] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold674 (.A(\mem.mem[166][4] ),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold675 (.A(\mem.mem[27][3] ),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold676 (.A(\mem.mem[227][3] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold677 (.A(\mem.mem[216][3] ),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold678 (.A(\mem.mem[174][7] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold679 (.A(\mem.mem[94][0] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold680 (.A(\mem.mem[222][6] ),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold681 (.A(\mem.mem[7][7] ),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold682 (.A(\mem.mem[149][5] ),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold683 (.A(\mem.mem[214][4] ),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold684 (.A(\mem.mem[245][0] ),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold685 (.A(\mem.mem[168][1] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold686 (.A(\mem.mem[183][5] ),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold687 (.A(\mem.mem[247][0] ),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold688 (.A(\mem.mem[101][7] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold689 (.A(\mem.mem[250][5] ),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold690 (.A(\mem.mem[177][6] ),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold691 (.A(\mem.mem[110][1] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold692 (.A(\mem.mem[109][7] ),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold693 (.A(\mem.mem[99][4] ),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold694 (.A(\mem.mem[102][2] ),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold695 (.A(\mem.mem[228][1] ),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold696 (.A(\mem.mem[174][5] ),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold697 (.A(\mem.mem[113][1] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold698 (.A(\mem.mem[78][7] ),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold699 (.A(\mem.mem[227][0] ),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold700 (.A(\mem.mem[188][1] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold701 (.A(\mem.mem[23][4] ),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold702 (.A(\mem.mem[231][5] ),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold703 (.A(\mem.mem[169][5] ),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold704 (.A(\mem.mem[83][1] ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold705 (.A(\mem.mem[250][1] ),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold706 (.A(\mem.mem[220][6] ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold707 (.A(\mem.mem[46][1] ),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold708 (.A(\mem.mem[87][5] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold709 (.A(\mem.mem[64][7] ),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold710 (.A(\mem.mem[241][1] ),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold711 (.A(\mem.mem[217][6] ),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold712 (.A(\mem.mem[211][6] ),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold713 (.A(\mem.mem[85][0] ),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold714 (.A(\mem.mem[27][2] ),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold715 (.A(\mem.mem[181][7] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold716 (.A(\mem.mem[83][5] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold717 (.A(\mem.mem[50][7] ),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold718 (.A(\mem.mem[55][0] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold719 (.A(\mem.mem[83][2] ),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold720 (.A(\mem.mem[144][7] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold721 (.A(\mem.mem[171][6] ),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold722 (.A(\mem.mem[227][6] ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold723 (.A(\mem.mem[16][1] ),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold724 (.A(\mem.mem[150][0] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold725 (.A(\mem.mem[171][3] ),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold726 (.A(\mem.mem[80][5] ),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold727 (.A(\mem.mem[27][6] ),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold728 (.A(\mem.mem[91][7] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold729 (.A(\mem.mem[100][4] ),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold730 (.A(\mem.mem[149][0] ),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold731 (.A(\mem.mem[190][3] ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold732 (.A(\mem.mem[115][5] ),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold733 (.A(\mem.mem[194][5] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold734 (.A(\mem.mem[80][2] ),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold735 (.A(\mem.mem[182][4] ),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold736 (.A(\mem.mem[44][7] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold737 (.A(\mem.mem[125][0] ),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold738 (.A(\mem.mem[214][7] ),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold739 (.A(\mem.mem[245][1] ),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold740 (.A(\mem.mem[22][6] ),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold741 (.A(\mem.mem[87][2] ),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold742 (.A(\mem.mem[151][3] ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold743 (.A(\mem.mem[166][2] ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold744 (.A(\mem.mem[177][7] ),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold745 (.A(\mem.mem[102][7] ),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold746 (.A(\mem.mem[164][5] ),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold747 (.A(\mem.mem[179][3] ),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold748 (.A(\mem.mem[83][4] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold749 (.A(\mem.mem[225][6] ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold750 (.A(\mem.mem[52][2] ),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold751 (.A(\mem.mem[71][1] ),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold752 (.A(\mem.mem[32][3] ),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold753 (.A(\mem.mem[214][6] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold754 (.A(\mem.mem[101][4] ),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold755 (.A(\mem.mem[96][7] ),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold756 (.A(\mem.mem[92][4] ),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold757 (.A(\mem.mem[103][7] ),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold758 (.A(\mem.mem[216][2] ),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold759 (.A(\mem.mem[152][6] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold760 (.A(\mem.mem[190][5] ),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold761 (.A(\mem.mem[87][1] ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold762 (.A(\mem.mem[83][3] ),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold763 (.A(\mem.mem[235][5] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold764 (.A(\mem.mem[119][7] ),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold765 (.A(\mem.mem[64][1] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold766 (.A(\mem.mem[230][3] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold767 (.A(\mem.mem[190][2] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold768 (.A(\mem.mem[61][7] ),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold769 (.A(\mem.mem[158][3] ),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold770 (.A(\mem.mem[152][5] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold771 (.A(\mem.mem[120][4] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold772 (.A(\mem.mem[170][1] ),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold773 (.A(\mem.mem[116][5] ),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold774 (.A(\mem.mem[53][5] ),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold775 (.A(\mem.mem[149][6] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold776 (.A(\mem.mem[113][2] ),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold777 (.A(\mem.mem[154][5] ),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold778 (.A(\mem.mem[104][6] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold779 (.A(\mem.mem[74][0] ),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold780 (.A(\mem.mem[117][1] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold781 (.A(\mem.mem[78][5] ),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold782 (.A(\mem.mem[61][4] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold783 (.A(\mem.mem[85][3] ),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold784 (.A(\mem.mem[30][4] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold785 (.A(\mem.mem[185][3] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold786 (.A(\mem.mem[61][0] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold787 (.A(\mem.mem[179][4] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold788 (.A(\mem.mem[122][3] ),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold789 (.A(\mem.mem[233][7] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold790 (.A(\mem.mem[163][5] ),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold791 (.A(\mem.mem[199][5] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold792 (.A(\mem.mem[155][3] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold793 (.A(\mem.mem[60][2] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold794 (.A(\mem.mem[170][7] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold795 (.A(\mem.mem[233][5] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold796 (.A(\mem.mem[214][1] ),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold797 (.A(\mem.mem[179][6] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold798 (.A(\mem.mem[16][3] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold799 (.A(\mem.mem[209][5] ),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold800 (.A(\mem.mem[228][7] ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold801 (.A(\mem.mem[224][1] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold802 (.A(\mem.mem[234][6] ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold803 (.A(\mem.mem[178][5] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold804 (.A(\mem.mem[45][4] ),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold805 (.A(\mem.mem[174][2] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold806 (.A(\mem.mem[244][1] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold807 (.A(\mem.mem[173][0] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold808 (.A(\mem.mem[122][6] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold809 (.A(\mem.mem[118][7] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold810 (.A(\mem.mem[154][1] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold811 (.A(\mem.mem[29][4] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold812 (.A(\mem.mem[123][4] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold813 (.A(\mem.mem[59][2] ),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold814 (.A(\mem.mem[101][3] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold815 (.A(\mem.mem[27][1] ),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold816 (.A(\mem.mem[86][2] ),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold817 (.A(\mem.mem[121][4] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold818 (.A(\mem.mem[170][0] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold819 (.A(\mem.mem[116][4] ),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold820 (.A(\mem.mem[62][0] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold821 (.A(\mem.mem[211][4] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold822 (.A(\mem.mem[49][0] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold823 (.A(\mem.mem[135][0] ),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold824 (.A(\mem.mem[210][7] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold825 (.A(\mem.mem[30][2] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold826 (.A(\mem.mem[117][2] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold827 (.A(\mem.mem[106][2] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold828 (.A(\mem.mem[216][0] ),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold829 (.A(\mem.mem[99][3] ),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold830 (.A(\mem.mem[93][0] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold831 (.A(\mem.mem[124][0] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold832 (.A(\mem.mem[164][2] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold833 (.A(\mem.mem[105][2] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold834 (.A(\mem.mem[92][2] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold835 (.A(\mem.mem[46][5] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold836 (.A(\mem.mem[232][1] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold837 (.A(\mem.mem[214][5] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold838 (.A(\mem.mem[185][1] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold839 (.A(\mem.mem[39][4] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold840 (.A(\mem.mem[234][0] ),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold841 (.A(\mem.mem[0][2] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold842 (.A(\mem.mem[89][0] ),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold843 (.A(\mem.mem[234][3] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold844 (.A(\mem.mem[213][4] ),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold845 (.A(\mem.mem[189][5] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold846 (.A(\mem.mem[80][1] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold847 (.A(\mem.mem[96][2] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold848 (.A(\mem.mem[125][2] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold849 (.A(\mem.mem[176][3] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold850 (.A(\mem.mem[210][0] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold851 (.A(\mem.mem[32][7] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold852 (.A(\mem.mem[208][7] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold853 (.A(\mem.mem[196][6] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold854 (.A(\mem.mem[155][0] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold855 (.A(\mem.mem[85][6] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold856 (.A(\mem.mem[231][2] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold857 (.A(\mem.mem[135][1] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold858 (.A(\mem.mem[45][2] ),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold859 (.A(\mem.mem[242][3] ),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold860 (.A(\mem.mem[156][6] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold861 (.A(\mem.mem[91][2] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold862 (.A(\mem.mem[0][6] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold863 (.A(\mem.mem[118][5] ),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold864 (.A(\mem.mem[109][1] ),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold865 (.A(\mem.mem[93][1] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold866 (.A(\mem.mem[49][4] ),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold867 (.A(\mem.mem[185][6] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold868 (.A(\mem.mem[144][0] ),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold869 (.A(\mem.mem[27][0] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold870 (.A(\mem.mem[198][4] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold871 (.A(\mem.mem[92][3] ),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold872 (.A(\mem.mem[225][7] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold873 (.A(\mem.mem[104][2] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold874 (.A(\mem.mem[189][2] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold875 (.A(\mem.mem[176][1] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold876 (.A(\mem.mem[64][2] ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold877 (.A(\mem.mem[151][1] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold878 (.A(\mem.mem[49][2] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold879 (.A(\mem.mem[245][3] ),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold880 (.A(\mem.mem[110][2] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold881 (.A(\mem.mem[209][4] ),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold882 (.A(\mem.mem[149][3] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold883 (.A(\mem.mem[189][3] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold884 (.A(\mem.mem[60][4] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold885 (.A(\mem.mem[84][3] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold886 (.A(\mem.mem[30][5] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold887 (.A(\mem.mem[163][2] ),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold888 (.A(\mem.mem[114][1] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold889 (.A(\mem.mem[121][1] ),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold890 (.A(\mem.mem[172][6] ),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold891 (.A(\mem.mem[242][5] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold892 (.A(\mem.mem[169][4] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold893 (.A(\mem.mem[94][5] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold894 (.A(\mem.mem[198][6] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold895 (.A(\mem.mem[215][7] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold896 (.A(\mem.mem[150][7] ),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold897 (.A(\mem.mem[219][0] ),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold898 (.A(\mem.mem[60][7] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold899 (.A(\mem.mem[218][1] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold900 (.A(\mem.mem[124][4] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold901 (.A(\mem.mem[181][5] ),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold902 (.A(\mem.mem[39][6] ),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold903 (.A(\mem.mem[43][4] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold904 (.A(\mem.mem[153][0] ),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold905 (.A(\mem.mem[170][2] ),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold906 (.A(\mem.mem[135][6] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold907 (.A(\mem.mem[151][7] ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold908 (.A(\mem.mem[171][2] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold909 (.A(\mem.mem[187][0] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold910 (.A(\mem.mem[155][6] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold911 (.A(\mem.mem[58][2] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold912 (.A(\mem.mem[178][7] ),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold913 (.A(\mem.mem[115][6] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold914 (.A(\mem.mem[89][2] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold915 (.A(\mem.mem[250][0] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold916 (.A(\mem.mem[218][3] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold917 (.A(\mem.mem[101][1] ),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold918 (.A(\mem.mem[128][1] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold919 (.A(\mem.mem[149][4] ),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold920 (.A(\mem.mem[208][1] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold921 (.A(\mem.mem[60][3] ),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold922 (.A(\mem.mem[20][0] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold923 (.A(\mem.mem[56][6] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold924 (.A(\mem.mem[123][7] ),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold925 (.A(\mem.mem[48][6] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold926 (.A(\mem.mem[87][4] ),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold927 (.A(\mem.mem[20][7] ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold928 (.A(\mem.mem[150][4] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold929 (.A(\mem.mem[107][1] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold930 (.A(\mem.mem[108][5] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold931 (.A(\mem.mem[43][6] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold932 (.A(\mem.mem[172][4] ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold933 (.A(\mem.mem[0][1] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold934 (.A(\mem.mem[235][0] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold935 (.A(\mem.mem[50][4] ),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold936 (.A(\mem.mem[177][4] ),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold937 (.A(\mem.mem[88][4] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold938 (.A(\mem.mem[214][0] ),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold939 (.A(\mem.mem[247][1] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold940 (.A(\mem.mem[235][7] ),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold941 (.A(\mem.mem[156][3] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold942 (.A(\mem.mem[117][3] ),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold943 (.A(\mem.mem[219][1] ),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold944 (.A(\mem.mem[134][3] ),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold945 (.A(\mem.mem[61][6] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold946 (.A(\mem.mem[102][3] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold947 (.A(\mem.mem[225][3] ),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold948 (.A(\mem.mem[30][7] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold949 (.A(\mem.mem[184][5] ),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold950 (.A(\mem.mem[76][0] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold951 (.A(\mem.mem[241][0] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold952 (.A(\mem.mem[58][4] ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold953 (.A(\mem.mem[144][5] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold954 (.A(\mem.mem[190][7] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold955 (.A(\mem.mem[126][0] ),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold956 (.A(\mem.mem[43][7] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold957 (.A(\mem.mem[232][5] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold958 (.A(\mem.mem[250][3] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold959 (.A(\mem.mem[192][3] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold960 (.A(\mem.mem[118][0] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold961 (.A(_01045_),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold962 (.A(\mem.mem[88][3] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold963 (.A(\mem.mem[152][4] ),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold964 (.A(\mem.mem[39][3] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold965 (.A(\mem.mem[93][7] ),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold966 (.A(\mem.mem[229][1] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold967 (.A(\mem.mem[49][3] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold968 (.A(\mem.mem[122][0] ),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold969 (.A(\mem.mem[120][1] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold970 (.A(\mem.mem[153][7] ),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold971 (.A(\mem.mem[238][2] ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold972 (.A(\mem.mem[226][6] ),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold973 (.A(\mem.mem[206][3] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold974 (.A(\mem.mem[148][0] ),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold975 (.A(\mem.mem[16][6] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold976 (.A(\mem.mem[28][6] ),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold977 (.A(\mem.mem[173][5] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold978 (.A(\mem.mem[39][0] ),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold979 (.A(\mem.mem[53][4] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold980 (.A(\mem.mem[115][3] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold981 (.A(\mem.mem[150][3] ),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold982 (.A(\mem.mem[93][4] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold983 (.A(\mem.mem[210][2] ),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold984 (.A(\mem.mem[135][2] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold985 (.A(\mem.mem[56][5] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold986 (.A(\mem.mem[163][7] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold987 (.A(\mem.mem[218][5] ),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold988 (.A(\mem.mem[106][0] ),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold989 (.A(\mem.mem[241][7] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold990 (.A(\mem.mem[183][2] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold991 (.A(\mem.mem[99][1] ),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold992 (.A(\mem.mem[121][5] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold993 (.A(\mem.mem[232][3] ),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold994 (.A(\mem.mem[51][6] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold995 (.A(\mem.mem[110][7] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold996 (.A(\mem.mem[224][2] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold997 (.A(\mem.mem[54][1] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold998 (.A(\mem.mem[185][7] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold999 (.A(\mem.mem[224][4] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\mem.mem[217][0] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\mem.mem[169][0] ),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\mem.mem[222][0] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\mem.mem[217][4] ),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\mem.mem[94][6] ),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\mem.mem[53][1] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\mem.mem[104][5] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\mem.mem[167][0] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\mem.mem[229][6] ),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\mem.mem[87][0] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\mem.mem[59][0] ),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\mem.mem[160][6] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\mem.mem[43][3] ),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\mem.mem[125][3] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\mem.mem[118][1] ),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\mem.mem[179][2] ),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\mem.mem[199][3] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\mem.mem[167][3] ),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\mem.mem[56][4] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\mem.mem[160][1] ),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\mem.mem[231][1] ),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\mem.mem[199][0] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\mem.mem[226][4] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\mem.mem[234][5] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\mem.mem[62][2] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\mem.mem[43][2] ),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\mem.mem[113][0] ),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\mem.mem[249][5] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\mem.mem[215][5] ),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\mem.mem[233][4] ),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\mem.mem[219][7] ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\mem.mem[164][6] ),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\mem.mem[99][6] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\mem.mem[94][2] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\mem.mem[162][7] ),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\mem.mem[7][0] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\mem.mem[42][6] ),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\mem.mem[156][5] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\mem.mem[167][1] ),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\mem.mem[192][7] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\mem.mem[232][7] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\mem.mem[83][6] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\mem.mem[237][6] ),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\mem.mem[16][2] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\mem.mem[123][2] ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\mem.mem[174][6] ),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\mem.mem[113][4] ),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\mem.mem[105][5] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\mem.mem[212][2] ),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\mem.mem[29][0] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\mem.mem[148][5] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\mem.mem[106][7] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\mem.mem[90][3] ),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\mem.mem[152][1] ),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\mem.mem[52][5] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\mem.mem[101][6] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\mem.mem[117][5] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\mem.mem[172][5] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\mem.mem[245][7] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\mem.mem[88][0] ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\mem.mem[125][5] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\mem.mem[167][6] ),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\mem.mem[153][5] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\mem.mem[216][4] ),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\mem.mem[135][7] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\mem.mem[126][5] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\mem.mem[29][5] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\mem.mem[132][3] ),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\mem.mem[80][0] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\mem.mem[156][2] ),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\mem.mem[87][3] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\mem.mem[165][6] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\mem.mem[107][6] ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\mem.mem[106][4] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\mem.mem[235][1] ),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\mem.mem[135][3] ),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\mem.mem[27][5] ),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\mem.mem[168][7] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\mem.mem[230][2] ),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\mem.mem[62][1] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\mem.mem[236][3] ),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\mem.mem[96][5] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\mem.mem[250][2] ),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\mem.mem[183][1] ),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\mem.mem[190][0] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\mem.mem[109][5] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\mem.mem[218][2] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\mem.mem[45][6] ),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\mem.mem[153][6] ),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\mem.mem[202][4] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\mem.mem[55][3] ),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\mem.mem[62][3] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\mem.mem[26][4] ),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\mem.mem[51][1] ),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\mem.mem[180][2] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\mem.mem[72][6] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\mem.mem[22][5] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\mem.mem[57][0] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\mem.mem[213][1] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\mem.mem[53][0] ),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\mem.mem[120][2] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\mem.mem[155][4] ),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\mem.mem[211][1] ),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\mem.mem[43][0] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\mem.mem[204][6] ),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\mem.mem[27][7] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\mem.mem[83][0] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\mem.mem[56][7] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\mem.mem[165][7] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\mem.mem[242][7] ),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\mem.mem[45][7] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\mem.mem[180][1] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\mem.mem[121][6] ),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\mem.mem[74][5] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\mem.mem[120][3] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\mem.mem[229][3] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\mem.mem[147][0] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\mem.mem[88][5] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\mem.mem[149][7] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\mem.mem[80][7] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\mem.mem[135][4] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\mem.mem[206][4] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\mem.mem[182][7] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\mem.mem[0][7] ),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\mem.mem[158][4] ),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\mem.mem[107][7] ),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\mem.mem[196][5] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\mem.mem[166][6] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\mem.mem[189][6] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\mem.mem[167][4] ),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\mem.mem[7][6] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\mem.mem[42][3] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\mem.mem[108][3] ),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\mem.mem[250][7] ),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\mem.mem[128][4] ),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\mem.mem[163][0] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\mem.mem[199][4] ),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\mem.mem[188][0] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\mem.mem[128][2] ),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\mem.mem[87][6] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\mem.mem[173][7] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\mem.mem[183][3] ),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\mem.mem[204][3] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\mem.mem[109][4] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\mem.mem[235][4] ),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\mem.mem[110][4] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\mem.mem[218][7] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\mem.mem[57][4] ),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\mem.mem[219][6] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\mem.mem[53][2] ),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\mem.mem[189][0] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\mem.mem[109][6] ),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\mem.mem[71][7] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\mem.mem[217][3] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\mem.mem[181][4] ),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\mem.mem[246][0] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\mem.mem[66][0] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\mem.mem[102][1] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\mem.mem[41][6] ),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\mem.mem[101][2] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\mem.mem[147][5] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\mem.mem[227][2] ),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\mem.mem[191][7] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\mem.mem[193][7] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\mem.mem[212][5] ),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\mem.mem[87][7] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\mem.mem[187][7] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\mem.mem[174][3] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\mem.mem[194][4] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\mem.mem[84][1] ),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\mem.mem[147][1] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\mem.mem[187][3] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\mem.mem[148][6] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\mem.mem[220][2] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\mem.mem[191][6] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\mem.mem[198][7] ),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\mem.mem[57][2] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\mem.mem[226][5] ),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\mem.mem[76][7] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\mem.mem[151][5] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\mem.mem[150][6] ),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\mem.mem[171][4] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\mem.mem[191][5] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\mem.mem[131][1] ),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\mem.mem[116][7] ),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\mem.mem[248][2] ),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\mem.mem[109][0] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\mem.mem[93][2] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\mem.mem[57][6] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\mem.mem[181][6] ),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\mem.mem[134][1] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\mem.mem[126][3] ),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\mem.mem[237][4] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\mem.mem[239][7] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\mem.mem[8][4] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\mem.mem[137][5] ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\mem.mem[239][0] ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\mem.mem[77][3] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\mem.mem[81][5] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\mem.mem[204][0] ),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\mem.mem[12][0] ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\mem.mem[197][2] ),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\mem.mem[134][5] ),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\mem.mem[157][5] ),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\mem.mem[16][0] ),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\mem.mem[113][6] ),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\mem.mem[12][3] ),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\mem.mem[249][3] ),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\mem.mem[3][2] ),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\mem.mem[106][6] ),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\mem.mem[146][5] ),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\mem.mem[74][4] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\mem.mem[29][6] ),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\mem.mem[57][3] ),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\mem.mem[239][6] ),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\mem.mem[66][6] ),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\mem.mem[234][2] ),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\mem.mem[157][7] ),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\mem.mem[24][6] ),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\mem.mem[138][4] ),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\mem.mem[167][7] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\mem.mem[52][3] ),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\mem.mem[17][6] ),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\mem.mem[100][3] ),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\mem.mem[101][0] ),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\mem.mem[36][0] ),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\mem.mem[242][6] ),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\mem.mem[207][6] ),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\mem.mem[140][5] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\mem.mem[185][5] ),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\mem.mem[142][3] ),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\mem.mem[147][3] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\mem.mem[82][4] ),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\mem.mem[13][2] ),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\mem.mem[194][1] ),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\mem.mem[243][5] ),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\mem.mem[162][3] ),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\mem.mem[84][7] ),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\mem.mem[54][6] ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\mem.mem[97][5] ),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\mem.mem[249][7] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\mem.mem[219][5] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\mem.mem[138][2] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\mem.mem[226][2] ),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\mem.mem[168][5] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\mem.mem[211][5] ),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\mem.mem[122][1] ),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\mem.mem[21][6] ),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\mem.mem[89][1] ),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\mem.mem[243][2] ),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\mem.mem[172][1] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\mem.mem[196][3] ),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\mem.mem[60][6] ),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\mem.mem[197][1] ),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\mem.mem[166][7] ),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold1255 (.A(_01436_),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\mem.mem[26][3] ),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\mem.mem[202][1] ),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\mem.mem[37][7] ),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\mem.mem[33][3] ),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\mem.mem[17][3] ),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\mem.mem[194][0] ),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\mem.mem[77][2] ),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\mem.mem[157][3] ),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\mem.mem[1][4] ),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\mem.mem[161][0] ),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\mem.mem[112][2] ),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\mem.mem[5][5] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\mem.mem[73][3] ),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\mem.mem[152][3] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\mem.mem[102][0] ),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\mem.mem[207][5] ),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\mem.mem[28][7] ),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\mem.mem[237][5] ),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\mem.mem[68][0] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\mem.mem[117][0] ),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\mem.mem[18][3] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\mem.mem[252][6] ),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\mem.mem[142][6] ),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\mem.mem[127][7] ),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\mem.mem[76][5] ),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\mem.mem[14][7] ),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\mem.mem[142][0] ),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\mem.mem[141][6] ),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\mem.mem[31][2] ),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\mem.mem[193][2] ),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\mem.mem[139][1] ),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\mem.mem[152][2] ),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\mem.mem[194][7] ),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\mem.mem[137][0] ),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\mem.mem[89][5] ),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\mem.mem[79][6] ),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\mem.mem[244][3] ),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\mem.mem[136][0] ),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\mem.mem[40][4] ),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\mem.mem[144][6] ),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\mem.mem[133][4] ),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\mem.mem[82][5] ),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\mem.mem[33][1] ),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\mem.mem[47][4] ),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\mem.mem[21][1] ),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\mem.mem[252][3] ),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\mem.mem[37][1] ),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\mem.mem[76][2] ),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\mem.mem[133][1] ),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\mem.mem[208][4] ),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold1306 (.A(\mem.mem[221][1] ),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\mem.mem[173][3] ),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\mem.mem[193][3] ),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\mem.mem[6][0] ),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\mem.mem[65][7] ),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\mem.mem[18][5] ),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\mem.mem[8][2] ),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\mem.mem[20][4] ),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\mem.mem[141][4] ),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\mem.mem[72][3] ),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\mem.mem[146][3] ),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\mem.mem[239][2] ),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\mem.mem[12][2] ),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\mem.mem[204][5] ),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\mem.mem[38][0] ),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\mem.mem[70][3] ),
    .X(net3452));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\mem.mem[146][6] ),
    .X(net3453));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\mem.mem[59][7] ),
    .X(net3454));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\mem.mem[72][7] ),
    .X(net3455));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\mem.mem[75][0] ),
    .X(net3456));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\mem.mem[153][2] ),
    .X(net3457));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\mem.mem[15][3] ),
    .X(net3458));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\mem.mem[132][1] ),
    .X(net3459));
 sg13g2_dlygate4sd3_1 hold1329 (.A(\mem.mem[35][1] ),
    .X(net3460));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\mem.mem[33][5] ),
    .X(net3461));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\mem.mem[111][3] ),
    .X(net3462));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\mem.mem[40][6] ),
    .X(net3463));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\mem.mem[137][4] ),
    .X(net3464));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\mem.mem[35][2] ),
    .X(net3465));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\mem.mem[134][7] ),
    .X(net3466));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\mem.mem[243][4] ),
    .X(net3467));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\mem.mem[173][6] ),
    .X(net3468));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\mem.mem[205][5] ),
    .X(net3469));
 sg13g2_dlygate4sd3_1 hold1339 (.A(\mem.mem[37][4] ),
    .X(net3470));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\mem.mem[145][2] ),
    .X(net3471));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\mem.mem[131][6] ),
    .X(net3472));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\mem.mem[111][1] ),
    .X(net3473));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\mem.mem[36][3] ),
    .X(net3474));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\mem.mem[162][2] ),
    .X(net3475));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\mem.mem[162][1] ),
    .X(net3476));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\mem.mem[4][7] ),
    .X(net3477));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\mem.mem[111][7] ),
    .X(net3478));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\mem.mem[207][4] ),
    .X(net3479));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\mem.mem[112][6] ),
    .X(net3480));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\mem.mem[86][6] ),
    .X(net3481));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\mem.mem[44][4] ),
    .X(net3482));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\mem.mem[251][6] ),
    .X(net3483));
 sg13g2_dlygate4sd3_1 hold1353 (.A(\mem.mem[6][5] ),
    .X(net3484));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\mem.mem[127][0] ),
    .X(net3485));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\mem.mem[142][1] ),
    .X(net3486));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\mem.mem[147][4] ),
    .X(net3487));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\mem.mem[168][6] ),
    .X(net3488));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\mem.mem[25][1] ),
    .X(net3489));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\mem.mem[1][5] ),
    .X(net3490));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\mem.mem[67][5] ),
    .X(net3491));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\mem.mem[140][4] ),
    .X(net3492));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\mem.mem[51][4] ),
    .X(net3493));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\mem.mem[34][4] ),
    .X(net3494));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\mem.mem[175][0] ),
    .X(net3495));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\mem.mem[198][3] ),
    .X(net3496));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\mem.mem[28][4] ),
    .X(net3497));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\mem.mem[8][1] ),
    .X(net3498));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\mem.mem[200][5] ),
    .X(net3499));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\mem.mem[19][4] ),
    .X(net3500));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\mem.mem[69][0] ),
    .X(net3501));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\mem.mem[206][5] ),
    .X(net3502));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\mem.mem[197][0] ),
    .X(net3503));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\mem.mem[5][3] ),
    .X(net3504));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\mem.mem[56][1] ),
    .X(net3505));
 sg13g2_dlygate4sd3_1 hold1375 (.A(_00445_),
    .X(net3506));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\mem.mem[66][5] ),
    .X(net3507));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\mem.mem[240][4] ),
    .X(net3508));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\mem.mem[47][5] ),
    .X(net3509));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\mem.mem[14][2] ),
    .X(net3510));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\mem.mem[68][4] ),
    .X(net3511));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\mem.mem[248][1] ),
    .X(net3512));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\mem.mem[203][0] ),
    .X(net3513));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\mem.mem[145][7] ),
    .X(net3514));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\mem.mem[31][1] ),
    .X(net3515));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\mem.mem[14][6] ),
    .X(net3516));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\mem.mem[201][6] ),
    .X(net3517));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\mem.mem[132][7] ),
    .X(net3518));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\mem.mem[161][4] ),
    .X(net3519));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\mem.mem[240][3] ),
    .X(net3520));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\mem.mem[195][3] ),
    .X(net3521));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\mem.mem[14][4] ),
    .X(net3522));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\mem.mem[116][1] ),
    .X(net3523));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\mem.mem[230][1] ),
    .X(net3524));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\mem.mem[143][6] ),
    .X(net3525));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\mem.mem[78][1] ),
    .X(net3526));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\mem.mem[129][5] ),
    .X(net3527));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\mem.mem[67][7] ),
    .X(net3528));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\mem.mem[97][3] ),
    .X(net3529));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\mem.mem[49][5] ),
    .X(net3530));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\mem.mem[14][3] ),
    .X(net3531));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\mem.mem[24][7] ),
    .X(net3532));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\mem.mem[28][0] ),
    .X(net3533));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\mem.mem[66][3] ),
    .X(net3534));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\mem.mem[206][2] ),
    .X(net3535));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\mem.mem[200][6] ),
    .X(net3536));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\mem.mem[204][4] ),
    .X(net3537));
 sg13g2_dlygate4sd3_1 hold1407 (.A(\mem.mem[130][0] ),
    .X(net3538));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\mem.mem[70][1] ),
    .X(net3539));
 sg13g2_dlygate4sd3_1 hold1409 (.A(\mem.mem[9][4] ),
    .X(net3540));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\mem.mem[70][7] ),
    .X(net3541));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\mem.mem[97][6] ),
    .X(net3542));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\mem.mem[0][4] ),
    .X(net3543));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\mem.mem[201][0] ),
    .X(net3544));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\mem.mem[252][4] ),
    .X(net3545));
 sg13g2_dlygate4sd3_1 hold1415 (.A(\mem.mem[98][4] ),
    .X(net3546));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\mem.mem[9][2] ),
    .X(net3547));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\mem.mem[205][3] ),
    .X(net3548));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\mem.mem[42][7] ),
    .X(net3549));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\mem.mem[21][2] ),
    .X(net3550));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\mem.mem[137][7] ),
    .X(net3551));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\mem.mem[142][2] ),
    .X(net3552));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\mem.mem[223][5] ),
    .X(net3553));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\mem.mem[251][7] ),
    .X(net3554));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\mem.mem[246][6] ),
    .X(net3555));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\mem.mem[74][3] ),
    .X(net3556));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\mem.mem[191][0] ),
    .X(net3557));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\mem.mem[143][0] ),
    .X(net3558));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\mem.mem[11][3] ),
    .X(net3559));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\mem.mem[42][2] ),
    .X(net3560));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\mem.mem[131][3] ),
    .X(net3561));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\mem.mem[18][6] ),
    .X(net3562));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\mem.mem[203][1] ),
    .X(net3563));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\mem.mem[223][0] ),
    .X(net3564));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\mem.mem[37][5] ),
    .X(net3565));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\mem.mem[36][6] ),
    .X(net3566));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\mem.mem[132][6] ),
    .X(net3567));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\mem.mem[34][6] ),
    .X(net3568));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\mem.mem[36][2] ),
    .X(net3569));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\mem.mem[12][1] ),
    .X(net3570));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\mem.mem[74][2] ),
    .X(net3571));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\mem.mem[95][3] ),
    .X(net3572));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\mem.mem[18][7] ),
    .X(net3573));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\mem.mem[17][2] ),
    .X(net3574));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\mem.mem[22][4] ),
    .X(net3575));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\mem.mem[47][7] ),
    .X(net3576));
 sg13g2_dlygate4sd3_1 hold1446 (.A(\mem.mem[142][5] ),
    .X(net3577));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\mem.mem[244][0] ),
    .X(net3578));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\mem.mem[197][5] ),
    .X(net3579));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\mem.mem[33][6] ),
    .X(net3580));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\mem.mem[194][3] ),
    .X(net3581));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\mem.mem[156][1] ),
    .X(net3582));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\mem.mem[48][0] ),
    .X(net3583));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\mem.mem[14][0] ),
    .X(net3584));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\mem.mem[17][7] ),
    .X(net3585));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\mem.mem[63][0] ),
    .X(net3586));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\mem.mem[44][0] ),
    .X(net3587));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\mem.mem[136][3] ),
    .X(net3588));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\mem.mem[97][2] ),
    .X(net3589));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\mem.mem[143][7] ),
    .X(net3590));
 sg13g2_dlygate4sd3_1 hold1460 (.A(\mem.mem[248][4] ),
    .X(net3591));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\mem.mem[13][7] ),
    .X(net3592));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\mem.mem[44][5] ),
    .X(net3593));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\mem.mem[77][4] ),
    .X(net3594));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\mem.mem[64][4] ),
    .X(net3595));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\mem.mem[136][6] ),
    .X(net3596));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\mem.mem[130][4] ),
    .X(net3597));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\mem.mem[14][1] ),
    .X(net3598));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\mem.mem[107][4] ),
    .X(net3599));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\mem.mem[4][6] ),
    .X(net3600));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\mem.mem[142][4] ),
    .X(net3601));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\mem.mem[10][6] ),
    .X(net3602));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\mem.mem[44][3] ),
    .X(net3603));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\mem.mem[138][7] ),
    .X(net3604));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\mem.mem[69][7] ),
    .X(net3605));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\mem.mem[72][0] ),
    .X(net3606));
 sg13g2_dlygate4sd3_1 hold1476 (.A(\mem.mem[73][6] ),
    .X(net3607));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\mem.mem[204][2] ),
    .X(net3608));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\mem.mem[64][3] ),
    .X(net3609));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\mem.mem[79][1] ),
    .X(net3610));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\mem.mem[74][1] ),
    .X(net3611));
 sg13g2_dlygate4sd3_1 hold1481 (.A(\mem.mem[22][2] ),
    .X(net3612));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\mem.mem[3][6] ),
    .X(net3613));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\mem.mem[98][7] ),
    .X(net3614));
 sg13g2_dlygate4sd3_1 hold1484 (.A(\mem.mem[196][7] ),
    .X(net3615));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\mem.mem[78][0] ),
    .X(net3616));
 sg13g2_dlygate4sd3_1 hold1486 (.A(\mem.mem[200][3] ),
    .X(net3617));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\mem.mem[203][4] ),
    .X(net3618));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\mem.mem[204][7] ),
    .X(net3619));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\mem.mem[81][3] ),
    .X(net3620));
 sg13g2_dlygate4sd3_1 hold1490 (.A(\mem.mem[248][6] ),
    .X(net3621));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\mem.mem[42][4] ),
    .X(net3622));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\mem.mem[200][0] ),
    .X(net3623));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\mem.mem[240][7] ),
    .X(net3624));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\mem.mem[251][2] ),
    .X(net3625));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\mem.mem[145][0] ),
    .X(net3626));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\mem.mem[65][1] ),
    .X(net3627));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\mem.mem[203][6] ),
    .X(net3628));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\mem.mem[63][1] ),
    .X(net3629));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\mem.mem[197][3] ),
    .X(net3630));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\mem.mem[2][0] ),
    .X(net3631));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\mem.mem[11][0] ),
    .X(net3632));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\mem.mem[111][6] ),
    .X(net3633));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\mem.mem[11][1] ),
    .X(net3634));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\mem.mem[98][3] ),
    .X(net3635));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\mem.mem[98][1] ),
    .X(net3636));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\mem.mem[201][5] ),
    .X(net3637));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\mem.mem[205][6] ),
    .X(net3638));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\mem.mem[38][5] ),
    .X(net3639));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\mem.mem[143][1] ),
    .X(net3640));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\mem.mem[14][5] ),
    .X(net3641));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\mem.mem[200][4] ),
    .X(net3642));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\mem.mem[17][4] ),
    .X(net3643));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\mem.mem[34][1] ),
    .X(net3644));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\mem.mem[13][4] ),
    .X(net3645));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\mem.mem[244][5] ),
    .X(net3646));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\mem.mem[88][6] ),
    .X(net3647));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\mem.mem[44][1] ),
    .X(net3648));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\mem.mem[133][2] ),
    .X(net3649));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\mem.mem[95][1] ),
    .X(net3650));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\mem.mem[136][2] ),
    .X(net3651));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\mem.mem[162][0] ),
    .X(net3652));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\mem.mem[104][7] ),
    .X(net3653));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\mem.mem[21][4] ),
    .X(net3654));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\mem.mem[5][7] ),
    .X(net3655));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\mem.mem[97][1] ),
    .X(net3656));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\mem.mem[17][0] ),
    .X(net3657));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\mem.mem[159][3] ),
    .X(net3658));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\mem.mem[130][1] ),
    .X(net3659));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\mem.mem[65][6] ),
    .X(net3660));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\mem.mem[141][1] ),
    .X(net3661));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\mem.mem[81][6] ),
    .X(net3662));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\mem.mem[193][1] ),
    .X(net3663));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\mem.mem[82][6] ),
    .X(net3664));
 sg13g2_dlygate4sd3_1 hold1534 (.A(\mem.mem[73][5] ),
    .X(net3665));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\mem.mem[25][3] ),
    .X(net3666));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\mem.mem[244][2] ),
    .X(net3667));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\mem.mem[1][1] ),
    .X(net3668));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\mem.mem[205][0] ),
    .X(net3669));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\mem.mem[12][7] ),
    .X(net3670));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\mem.mem[11][7] ),
    .X(net3671));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\mem.mem[141][2] ),
    .X(net3672));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\mem.mem[75][3] ),
    .X(net3673));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\mem.mem[143][3] ),
    .X(net3674));
 sg13g2_dlygate4sd3_1 hold1544 (.A(\mem.mem[252][0] ),
    .X(net3675));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\mem.mem[78][4] ),
    .X(net3676));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\mem.mem[240][6] ),
    .X(net3677));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\mem.mem[201][3] ),
    .X(net3678));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\mem.mem[35][4] ),
    .X(net3679));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\mem.mem[69][1] ),
    .X(net3680));
 sg13g2_dlygate4sd3_1 hold1550 (.A(\mem.mem[143][5] ),
    .X(net3681));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\mem.mem[196][4] ),
    .X(net3682));
 sg13g2_dlygate4sd3_1 hold1552 (.A(\mem.mem[26][7] ),
    .X(net3683));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\mem.mem[79][5] ),
    .X(net3684));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\mem.mem[146][4] ),
    .X(net3685));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\mem.mem[159][1] ),
    .X(net3686));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\mem.mem[205][1] ),
    .X(net3687));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\mem.mem[31][5] ),
    .X(net3688));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\mem.mem[68][5] ),
    .X(net3689));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\mem.mem[127][6] ),
    .X(net3690));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\mem.mem[175][1] ),
    .X(net3691));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\mem.mem[191][2] ),
    .X(net3692));
 sg13g2_dlygate4sd3_1 hold1562 (.A(\mem.mem[15][2] ),
    .X(net3693));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\mem.mem[223][7] ),
    .X(net3694));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\mem.mem[74][6] ),
    .X(net3695));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\mem.mem[138][1] ),
    .X(net3696));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\mem.mem[201][2] ),
    .X(net3697));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\mem.mem[95][6] ),
    .X(net3698));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\mem.mem[252][5] ),
    .X(net3699));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\mem.mem[69][3] ),
    .X(net3700));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\mem.mem[17][5] ),
    .X(net3701));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\mem.mem[203][7] ),
    .X(net3702));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\mem.mem[243][6] ),
    .X(net3703));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\mem.mem[131][0] ),
    .X(net3704));
 sg13g2_dlygate4sd3_1 hold1574 (.A(\mem.mem[206][7] ),
    .X(net3705));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\mem.mem[243][3] ),
    .X(net3706));
 sg13g2_dlygate4sd3_1 hold1576 (.A(\mem.mem[207][3] ),
    .X(net3707));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\mem.mem[159][5] ),
    .X(net3708));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\mem.mem[203][3] ),
    .X(net3709));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\mem.mem[240][5] ),
    .X(net3710));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\mem.mem[98][5] ),
    .X(net3711));
 sg13g2_dlygate4sd3_1 hold1581 (.A(\mem.mem[84][2] ),
    .X(net3712));
 sg13g2_dlygate4sd3_1 hold1582 (.A(_00366_),
    .X(net3713));
 sg13g2_dlygate4sd3_1 hold1583 (.A(\mem.mem[78][2] ),
    .X(net3714));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\mem.mem[63][6] ),
    .X(net3715));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\mem.mem[63][2] ),
    .X(net3716));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\mem.mem[41][4] ),
    .X(net3717));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\mem.mem[75][7] ),
    .X(net3718));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\mem.mem[248][3] ),
    .X(net3719));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\mem.mem[11][4] ),
    .X(net3720));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\mem.mem[111][5] ),
    .X(net3721));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\mem.mem[136][4] ),
    .X(net3722));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\mem.mem[22][3] ),
    .X(net3723));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\mem.mem[77][5] ),
    .X(net3724));
 sg13g2_dlygate4sd3_1 hold1594 (.A(\mem.mem[70][4] ),
    .X(net3725));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\mem.mem[28][1] ),
    .X(net3726));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\mem.mem[146][0] ),
    .X(net3727));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\mem.mem[21][5] ),
    .X(net3728));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\mem.mem[132][0] ),
    .X(net3729));
 sg13g2_dlygate4sd3_1 hold1599 (.A(\mem.mem[77][0] ),
    .X(net3730));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\mem.mem[79][7] ),
    .X(net3731));
 sg13g2_dlygate4sd3_1 hold1601 (.A(\mem.mem[139][2] ),
    .X(net3732));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\mem.mem[67][2] ),
    .X(net3733));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\mem.mem[72][5] ),
    .X(net3734));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\mem.mem[44][2] ),
    .X(net3735));
 sg13g2_dlygate4sd3_1 hold1605 (.A(\mem.mem[161][6] ),
    .X(net3736));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\mem.mem[136][7] ),
    .X(net3737));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\mem.mem[159][2] ),
    .X(net3738));
 sg13g2_dlygate4sd3_1 hold1608 (.A(\mem.mem[107][0] ),
    .X(net3739));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\mem.mem[145][5] ),
    .X(net3740));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\mem.mem[28][2] ),
    .X(net3741));
 sg13g2_dlygate4sd3_1 hold1611 (.A(\mem.mem[244][6] ),
    .X(net3742));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\mem.mem[140][7] ),
    .X(net3743));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\mem.mem[141][0] ),
    .X(net3744));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\mem.mem[69][2] ),
    .X(net3745));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\mem.mem[75][1] ),
    .X(net3746));
 sg13g2_dlygate4sd3_1 hold1616 (.A(\mem.mem[38][3] ),
    .X(net3747));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\mem.mem[73][0] ),
    .X(net3748));
 sg13g2_dlygate4sd3_1 hold1618 (.A(\mem.mem[200][2] ),
    .X(net3749));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\mem.mem[10][2] ),
    .X(net3750));
 sg13g2_dlygate4sd3_1 hold1620 (.A(\mem.mem[191][4] ),
    .X(net3751));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\mem.mem[73][4] ),
    .X(net3752));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\mem.mem[5][0] ),
    .X(net3753));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\mem.mem[131][7] ),
    .X(net3754));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\mem.mem[201][4] ),
    .X(net3755));
 sg13g2_dlygate4sd3_1 hold1625 (.A(\mem.mem[6][4] ),
    .X(net3756));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\mem.mem[138][5] ),
    .X(net3757));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\mem.mem[9][5] ),
    .X(net3758));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\mem.mem[160][0] ),
    .X(net3759));
 sg13g2_dlygate4sd3_1 hold1629 (.A(\mem.mem[2][4] ),
    .X(net3760));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\mem.mem[127][2] ),
    .X(net3761));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\mem.mem[77][7] ),
    .X(net3762));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\mem.mem[98][6] ),
    .X(net3763));
 sg13g2_dlygate4sd3_1 hold1633 (.A(\mem.mem[15][6] ),
    .X(net3764));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\mem.mem[73][2] ),
    .X(net3765));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\mem.mem[10][1] ),
    .X(net3766));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\mem.mem[137][3] ),
    .X(net3767));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\mem.mem[129][0] ),
    .X(net3768));
 sg13g2_dlygate4sd3_1 hold1638 (.A(\mem.mem[70][5] ),
    .X(net3769));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\mem.mem[38][1] ),
    .X(net3770));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\mem.mem[79][4] ),
    .X(net3771));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\mem.mem[22][7] ),
    .X(net3772));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\mem.mem[31][3] ),
    .X(net3773));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\mem.mem[130][5] ),
    .X(net3774));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\mem.mem[139][4] ),
    .X(net3775));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\mem.mem[207][1] ),
    .X(net3776));
 sg13g2_dlygate4sd3_1 hold1646 (.A(\mem.mem[40][5] ),
    .X(net3777));
 sg13g2_dlygate4sd3_1 hold1647 (.A(\mem.mem[81][1] ),
    .X(net3778));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\mem.mem[36][1] ),
    .X(net3779));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\mem.mem[72][2] ),
    .X(net3780));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\mem.mem[73][1] ),
    .X(net3781));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\mem.mem[82][3] ),
    .X(net3782));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\mem.mem[26][5] ),
    .X(net3783));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\mem.mem[151][6] ),
    .X(net3784));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\mem.mem[78][6] ),
    .X(net3785));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\mem.mem[41][7] ),
    .X(net3786));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\mem.mem[127][4] ),
    .X(net3787));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\mem.mem[129][1] ),
    .X(net3788));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\mem.mem[240][2] ),
    .X(net3789));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\mem.mem[197][4] ),
    .X(net3790));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\mem.mem[223][3] ),
    .X(net3791));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\mem.mem[1][0] ),
    .X(net3792));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\mem.mem[11][5] ),
    .X(net3793));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\mem.mem[130][7] ),
    .X(net3794));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\mem.mem[31][4] ),
    .X(net3795));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\mem.mem[73][7] ),
    .X(net3796));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\mem.mem[189][1] ),
    .X(net3797));
 sg13g2_dlygate4sd3_1 hold1667 (.A(\mem.mem[134][2] ),
    .X(net3798));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\mem.mem[25][7] ),
    .X(net3799));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\mem.mem[251][0] ),
    .X(net3800));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\mem.mem[70][2] ),
    .X(net3801));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\mem.mem[47][1] ),
    .X(net3802));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\mem.mem[3][1] ),
    .X(net3803));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\mem.mem[72][4] ),
    .X(net3804));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\mem.mem[159][7] ),
    .X(net3805));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\mem.mem[252][2] ),
    .X(net3806));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\mem.mem[191][1] ),
    .X(net3807));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\mem.mem[18][4] ),
    .X(net3808));
 sg13g2_dlygate4sd3_1 hold1678 (.A(\mem.mem[63][3] ),
    .X(net3809));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\mem.mem[66][7] ),
    .X(net3810));
 sg13g2_dlygate4sd3_1 hold1680 (.A(\mem.mem[24][1] ),
    .X(net3811));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\mem.mem[65][4] ),
    .X(net3812));
 sg13g2_dlygate4sd3_1 hold1682 (.A(\mem.mem[38][6] ),
    .X(net3813));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\mem.mem[251][5] ),
    .X(net3814));
 sg13g2_dlygate4sd3_1 hold1684 (.A(\mem.mem[81][2] ),
    .X(net3815));
 sg13g2_dlygate4sd3_1 hold1685 (.A(\mem.mem[202][3] ),
    .X(net3816));
 sg13g2_dlygate4sd3_1 hold1686 (.A(\mem.mem[35][3] ),
    .X(net3817));
 sg13g2_dlygate4sd3_1 hold1687 (.A(\mem.mem[1][3] ),
    .X(net3818));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\mem.mem[20][3] ),
    .X(net3819));
 sg13g2_dlygate4sd3_1 hold1689 (.A(\mem.mem[67][6] ),
    .X(net3820));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\mem.mem[12][6] ),
    .X(net3821));
 sg13g2_dlygate4sd3_1 hold1691 (.A(\mem.mem[195][7] ),
    .X(net3822));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\mem.mem[6][3] ),
    .X(net3823));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\mem.mem[137][2] ),
    .X(net3824));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\mem.mem[10][4] ),
    .X(net3825));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\mem.mem[204][1] ),
    .X(net3826));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\mem.mem[193][4] ),
    .X(net3827));
 sg13g2_dlygate4sd3_1 hold1697 (.A(\mem.mem[223][6] ),
    .X(net3828));
 sg13g2_dlygate4sd3_1 hold1698 (.A(\mem.mem[15][5] ),
    .X(net3829));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\mem.mem[129][2] ),
    .X(net3830));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\mem.mem[2][1] ),
    .X(net3831));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\mem.mem[34][5] ),
    .X(net3832));
 sg13g2_dlygate4sd3_1 hold1702 (.A(\mem.mem[26][6] ),
    .X(net3833));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\mem.mem[146][7] ),
    .X(net3834));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\mem.mem[6][7] ),
    .X(net3835));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\mem.mem[67][1] ),
    .X(net3836));
 sg13g2_dlygate4sd3_1 hold1706 (.A(\mem.mem[9][1] ),
    .X(net3837));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\mem.mem[200][1] ),
    .X(net3838));
 sg13g2_dlygate4sd3_1 hold1708 (.A(\mem.mem[25][0] ),
    .X(net3839));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\mem.mem[111][2] ),
    .X(net3840));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\mem.mem[243][7] ),
    .X(net3841));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\mem.mem[25][4] ),
    .X(net3842));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\mem.mem[75][4] ),
    .X(net3843));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\mem.mem[63][5] ),
    .X(net3844));
 sg13g2_dlygate4sd3_1 hold1714 (.A(\mem.mem[138][0] ),
    .X(net3845));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\mem.mem[2][5] ),
    .X(net3846));
 sg13g2_dlygate4sd3_1 hold1716 (.A(\mem.mem[13][1] ),
    .X(net3847));
 sg13g2_dlygate4sd3_1 hold1717 (.A(\mem.mem[76][6] ),
    .X(net3848));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\mem.mem[175][6] ),
    .X(net3849));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\mem.mem[195][5] ),
    .X(net3850));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\mem.mem[162][4] ),
    .X(net3851));
 sg13g2_dlygate4sd3_1 hold1721 (.A(\mem.mem[161][7] ),
    .X(net3852));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\mem.mem[202][5] ),
    .X(net3853));
 sg13g2_dlygate4sd3_1 hold1723 (.A(\mem.mem[161][5] ),
    .X(net3854));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\mem.mem[81][0] ),
    .X(net3855));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\mem.mem[207][7] ),
    .X(net3856));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\mem.mem[175][7] ),
    .X(net3857));
 sg13g2_dlygate4sd3_1 hold1727 (.A(\mem.mem[3][5] ),
    .X(net3858));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\mem.mem[24][5] ),
    .X(net3859));
 sg13g2_dlygate4sd3_1 hold1729 (.A(\mem.mem[240][0] ),
    .X(net3860));
 sg13g2_dlygate4sd3_1 hold1730 (.A(\mem.mem[202][2] ),
    .X(net3861));
 sg13g2_dlygate4sd3_1 hold1731 (.A(\mem.mem[36][7] ),
    .X(net3862));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\mem.mem[198][5] ),
    .X(net3863));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\mem.mem[191][3] ),
    .X(net3864));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\mem.mem[82][2] ),
    .X(net3865));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\mem.mem[35][6] ),
    .X(net3866));
 sg13g2_dlygate4sd3_1 hold1736 (.A(\mem.mem[72][1] ),
    .X(net3867));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\mem.mem[126][4] ),
    .X(net3868));
 sg13g2_dlygate4sd3_1 hold1738 (.A(\mem.mem[139][7] ),
    .X(net3869));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\mem.mem[140][2] ),
    .X(net3870));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\mem.mem[19][5] ),
    .X(net3871));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\mem.mem[251][1] ),
    .X(net3872));
 sg13g2_dlygate4sd3_1 hold1742 (.A(\mem.mem[13][6] ),
    .X(net3873));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\mem.mem[131][5] ),
    .X(net3874));
 sg13g2_dlygate4sd3_1 hold1744 (.A(\mem.mem[24][4] ),
    .X(net3875));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\mem.mem[223][4] ),
    .X(net3876));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\mem.mem[20][6] ),
    .X(net3877));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\mem.mem[47][0] ),
    .X(net3878));
 sg13g2_dlygate4sd3_1 hold1748 (.A(\mem.mem[4][5] ),
    .X(net3879));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\mem.mem[41][3] ),
    .X(net3880));
 sg13g2_dlygate4sd3_1 hold1750 (.A(\mem.mem[129][6] ),
    .X(net3881));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\mem.mem[130][3] ),
    .X(net3882));
 sg13g2_dlygate4sd3_1 hold1752 (.A(\mem.mem[18][2] ),
    .X(net3883));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\mem.mem[20][5] ),
    .X(net3884));
 sg13g2_dlygate4sd3_1 hold1754 (.A(\mem.mem[33][0] ),
    .X(net3885));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\mem.mem[95][5] ),
    .X(net3886));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\mem.mem[69][5] ),
    .X(net3887));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\mem.mem[4][4] ),
    .X(net3888));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\mem.mem[41][5] ),
    .X(net3889));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\mem.mem[205][2] ),
    .X(net3890));
 sg13g2_dlygate4sd3_1 hold1760 (.A(\mem.mem[9][3] ),
    .X(net3891));
 sg13g2_dlygate4sd3_1 hold1761 (.A(\mem.mem[15][1] ),
    .X(net3892));
 sg13g2_dlygate4sd3_1 hold1762 (.A(\mem.mem[62][7] ),
    .X(net3893));
 sg13g2_dlygate4sd3_1 hold1763 (.A(_00379_),
    .X(net3894));
 sg13g2_dlygate4sd3_1 hold1764 (.A(\mem.mem[31][0] ),
    .X(net3895));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\mem.mem[25][6] ),
    .X(net3896));
 sg13g2_dlygate4sd3_1 hold1766 (.A(\mem.mem[26][0] ),
    .X(net3897));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\mem.mem[68][2] ),
    .X(net3898));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\mem.mem[18][0] ),
    .X(net3899));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\mem.mem[2][2] ),
    .X(net3900));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\mem.mem[38][4] ),
    .X(net3901));
 sg13g2_dlygate4sd3_1 hold1771 (.A(\C[3] ),
    .X(net3902));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\mem.mem[194][2] ),
    .X(net3903));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\mem.mem[144][3] ),
    .X(net3904));
 sg13g2_dlygate4sd3_1 hold1774 (.A(_01256_),
    .X(net3905));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\mem.mem[244][7] ),
    .X(net3906));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\mem.mem[69][6] ),
    .X(net3907));
 sg13g2_dlygate4sd3_1 hold1777 (.A(\mem.mem[5][6] ),
    .X(net3908));
 sg13g2_dlygate4sd3_1 hold1778 (.A(\mem.mem[240][1] ),
    .X(net3909));
 sg13g2_dlygate4sd3_1 hold1779 (.A(\mem.mem[5][4] ),
    .X(net3910));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\mem.mem[34][2] ),
    .X(net3911));
 sg13g2_dlygate4sd3_1 hold1781 (.A(\mem.mem[37][6] ),
    .X(net3912));
 sg13g2_dlygate4sd3_1 hold1782 (.A(\mem.mem[26][2] ),
    .X(net3913));
 sg13g2_dlygate4sd3_1 hold1783 (.A(\mem.mem[195][1] ),
    .X(net3914));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\mem.mem[10][3] ),
    .X(net3915));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\mem.mem[4][3] ),
    .X(net3916));
 sg13g2_dlygate4sd3_1 hold1786 (.A(\mem.mem[145][4] ),
    .X(net3917));
 sg13g2_dlygate4sd3_1 hold1787 (.A(\mem.mem[35][0] ),
    .X(net3918));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\C[5] ),
    .X(net3919));
 sg13g2_dlygate4sd3_1 hold1789 (.A(_00569_),
    .X(net3920));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\mem.mem[143][4] ),
    .X(net3921));
 sg13g2_dlygate4sd3_1 hold1791 (.A(\mem.mem[223][1] ),
    .X(net3922));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\mem.mem[65][0] ),
    .X(net3923));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\mem.mem[134][0] ),
    .X(net3924));
 sg13g2_dlygate4sd3_1 hold1794 (.A(\mem.mem[239][5] ),
    .X(net3925));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\mem.mem[95][7] ),
    .X(net3926));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\mem.mem[138][6] ),
    .X(net3927));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\mem.mem[77][1] ),
    .X(net3928));
 sg13g2_dlygate4sd3_1 hold1798 (.A(\mem.mem[198][0] ),
    .X(net3929));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\mem.mem[62][5] ),
    .X(net3930));
 sg13g2_dlygate4sd3_1 hold1800 (.A(\mem.mem[132][5] ),
    .X(net3931));
 sg13g2_dlygate4sd3_1 hold1801 (.A(\mem.mem[127][3] ),
    .X(net3932));
 sg13g2_dlygate4sd3_1 hold1802 (.A(\mem.mem[28][5] ),
    .X(net3933));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\mem.mem[37][3] ),
    .X(net3934));
 sg13g2_dlygate4sd3_1 hold1804 (.A(\mem.mem[130][6] ),
    .X(net3935));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\mem.mem[159][0] ),
    .X(net3936));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\mem.mem[161][2] ),
    .X(net3937));
 sg13g2_dlygate4sd3_1 hold1807 (.A(\mem.mem[79][2] ),
    .X(net3938));
 sg13g2_dlygate4sd3_1 hold1808 (.A(\mem.mem[139][0] ),
    .X(net3939));
 sg13g2_dlygate4sd3_1 hold1809 (.A(\mem.mem[67][4] ),
    .X(net3940));
 sg13g2_dlygate4sd3_1 hold1810 (.A(\mem.mem[206][0] ),
    .X(net3941));
 sg13g2_dlygate4sd3_1 hold1811 (.A(\mem.mem[127][1] ),
    .X(net3942));
 sg13g2_dlygate4sd3_1 hold1812 (.A(\mem.mem[66][2] ),
    .X(net3943));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\mem.mem[196][0] ),
    .X(net3944));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\mem.mem[81][7] ),
    .X(net3945));
 sg13g2_dlygate4sd3_1 hold1815 (.A(\mem.mem[34][7] ),
    .X(net3946));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\mem.mem[70][6] ),
    .X(net3947));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\mem.mem[2][6] ),
    .X(net3948));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\mem.mem[95][2] ),
    .X(net3949));
 sg13g2_dlygate4sd3_1 hold1819 (.A(\mem.mem[38][2] ),
    .X(net3950));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\mem.mem[202][7] ),
    .X(net3951));
 sg13g2_dlygate4sd3_1 hold1821 (.A(\mem.mem[13][3] ),
    .X(net3952));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\mem.mem[154][3] ),
    .X(net3953));
 sg13g2_dlygate4sd3_1 hold1823 (.A(\mem.mem[19][3] ),
    .X(net3954));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\mem.mem[25][2] ),
    .X(net3955));
 sg13g2_dlygate4sd3_1 hold1825 (.A(\mem.mem[138][3] ),
    .X(net3956));
 sg13g2_dlygate4sd3_1 hold1826 (.A(\mem.mem[67][3] ),
    .X(net3957));
 sg13g2_dlygate4sd3_1 hold1827 (.A(\mem.mem[41][1] ),
    .X(net3958));
 sg13g2_dlygate4sd3_1 hold1828 (.A(\mem.mem[95][4] ),
    .X(net3959));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\mem.mem[38][7] ),
    .X(net3960));
 sg13g2_dlygate4sd3_1 hold1830 (.A(\mem.mem[34][0] ),
    .X(net3961));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\mem.mem[12][5] ),
    .X(net3962));
 sg13g2_dlygate4sd3_1 hold1832 (.A(\mem.mem[244][4] ),
    .X(net3963));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\mem.mem[130][2] ),
    .X(net3964));
 sg13g2_dlygate4sd3_1 hold1834 (.A(\mem.mem[251][4] ),
    .X(net3965));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\mem.mem[145][3] ),
    .X(net3966));
 sg13g2_dlygate4sd3_1 hold1836 (.A(\mem.mem[196][2] ),
    .X(net3967));
 sg13g2_dlygate4sd3_1 hold1837 (.A(\mem.mem[8][5] ),
    .X(net3968));
 sg13g2_dlygate4sd3_1 hold1838 (.A(\mem.mem[52][4] ),
    .X(net3969));
 sg13g2_dlygate4sd3_1 hold1839 (.A(_00496_),
    .X(net3970));
 sg13g2_dlygate4sd3_1 hold1840 (.A(\mem.mem[19][1] ),
    .X(net3971));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\mem.mem[82][7] ),
    .X(net3972));
 sg13g2_dlygate4sd3_1 hold1842 (.A(\mem.mem[40][2] ),
    .X(net3973));
 sg13g2_dlygate4sd3_1 hold1843 (.A(\mem.mem[67][0] ),
    .X(net3974));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\mem.mem[15][7] ),
    .X(net3975));
 sg13g2_dlygate4sd3_1 hold1845 (.A(\mem.mem[75][5] ),
    .X(net3976));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\mem.mem[2][3] ),
    .X(net3977));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\mem.mem[65][5] ),
    .X(net3978));
 sg13g2_dlygate4sd3_1 hold1848 (.A(\mem.mem[79][3] ),
    .X(net3979));
 sg13g2_dlygate4sd3_1 hold1849 (.A(\mem.mem[1][7] ),
    .X(net3980));
 sg13g2_dlygate4sd3_1 hold1850 (.A(\mem.mem[197][7] ),
    .X(net3981));
 sg13g2_dlygate4sd3_1 hold1851 (.A(\mem.mem[47][2] ),
    .X(net3982));
 sg13g2_dlygate4sd3_1 hold1852 (.A(\mem.mem[5][1] ),
    .X(net3983));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\mem.mem[243][0] ),
    .X(net3984));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\mem.mem[68][1] ),
    .X(net3985));
 sg13g2_dlygate4sd3_1 hold1855 (.A(\mem.mem[97][7] ),
    .X(net3986));
 sg13g2_dlygate4sd3_1 hold1856 (.A(\mem.mem[162][6] ),
    .X(net3987));
 sg13g2_dlygate4sd3_1 hold1857 (.A(\mem.mem[252][1] ),
    .X(net3988));
 sg13g2_dlygate4sd3_1 hold1858 (.A(\mem.mem[12][4] ),
    .X(net3989));
 sg13g2_dlygate4sd3_1 hold1859 (.A(\mem.mem[70][0] ),
    .X(net3990));
 sg13g2_dlygate4sd3_1 hold1860 (.A(\mem.mem[251][3] ),
    .X(net3991));
 sg13g2_dlygate4sd3_1 hold1861 (.A(\mem.mem[40][1] ),
    .X(net3992));
 sg13g2_dlygate4sd3_1 hold1862 (.A(\mem.mem[5][2] ),
    .X(net3993));
 sg13g2_dlygate4sd3_1 hold1863 (.A(\mem.mem[129][4] ),
    .X(net3994));
 sg13g2_dlygate4sd3_1 hold1864 (.A(\mem.mem[74][7] ),
    .X(net3995));
 sg13g2_dlygate4sd3_1 hold1865 (.A(\mem.mem[81][4] ),
    .X(net3996));
 sg13g2_dlygate4sd3_1 hold1866 (.A(\mem.mem[207][0] ),
    .X(net3997));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\mem.mem[1][2] ),
    .X(net3998));
 sg13g2_dlygate4sd3_1 hold1868 (.A(\mem.mem[133][0] ),
    .X(net3999));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\mem.mem[9][6] ),
    .X(net4000));
 sg13g2_dlygate4sd3_1 hold1870 (.A(\mem.mem[203][2] ),
    .X(net4001));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\mem.mem[205][7] ),
    .X(net4002));
 sg13g2_dlygate4sd3_1 hold1872 (.A(\mem.mem[243][1] ),
    .X(net4003));
 sg13g2_dlygate4sd3_1 hold1873 (.A(\mem.mem[134][4] ),
    .X(net4004));
 sg13g2_dlygate4sd3_1 hold1874 (.A(\mem.mem[201][7] ),
    .X(net4005));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\mem.mem[65][3] ),
    .X(net4006));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\mem.mem[47][3] ),
    .X(net4007));
 sg13g2_dlygate4sd3_1 hold1877 (.A(\mem.mem[21][3] ),
    .X(net4008));
 sg13g2_dlygate4sd3_1 hold1878 (.A(\mem.mem[202][6] ),
    .X(net4009));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\mem.mem[76][4] ),
    .X(net4010));
 sg13g2_dlygate4sd3_1 hold1880 (.A(\mem.mem[136][5] ),
    .X(net4011));
 sg13g2_dlygate4sd3_1 hold1881 (.A(\mem.mem[142][7] ),
    .X(net4012));
 sg13g2_dlygate4sd3_1 hold1882 (.A(\mem.mem[78][3] ),
    .X(net4013));
 sg13g2_dlygate4sd3_1 hold1883 (.A(\mem.mem[8][7] ),
    .X(net4014));
 sg13g2_dlygate4sd3_1 hold1884 (.A(\mem.mem[40][0] ),
    .X(net4015));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\mem.mem[76][3] ),
    .X(net4016));
 sg13g2_dlygate4sd3_1 hold1886 (.A(\mem.mem[13][5] ),
    .X(net4017));
 sg13g2_dlygate4sd3_1 hold1887 (.A(\mem.mem[47][6] ),
    .X(net4018));
 sg13g2_dlygate4sd3_1 hold1888 (.A(\mem.mem[131][2] ),
    .X(net4019));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\mem.mem[248][5] ),
    .X(net4020));
 sg13g2_dlygate4sd3_1 hold1890 (.A(\mem.mem[31][7] ),
    .X(net4021));
 sg13g2_dlygate4sd3_1 hold1891 (.A(\mem.mem[141][7] ),
    .X(net4022));
 sg13g2_dlygate4sd3_1 hold1892 (.A(\mem.mem[9][0] ),
    .X(net4023));
 sg13g2_dlygate4sd3_1 hold1893 (.A(\mem.mem[31][6] ),
    .X(net4024));
 sg13g2_dlygate4sd3_1 hold1894 (.A(\mem.mem[129][3] ),
    .X(net4025));
 sg13g2_dlygate4sd3_1 hold1895 (.A(\mem.mem[139][5] ),
    .X(net4026));
 sg13g2_dlygate4sd3_1 hold1896 (.A(\mem.mem[68][7] ),
    .X(net4027));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\mem.mem[137][1] ),
    .X(net4028));
 sg13g2_dlygate4sd3_1 hold1898 (.A(\mem.mem[97][4] ),
    .X(net4029));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\mem.mem[19][2] ),
    .X(net4030));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\mem.mem[139][3] ),
    .X(net4031));
 sg13g2_dlygate4sd3_1 hold1901 (.A(\mem.mem[197][6] ),
    .X(net4032));
 sg13g2_dlygate4sd3_1 hold1902 (.A(\mem.mem[161][1] ),
    .X(net4033));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\mem.mem[20][2] ),
    .X(net4034));
 sg13g2_dlygate4sd3_1 hold1904 (.A(\mem.mem[22][0] ),
    .X(net4035));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\mem.mem[127][5] ),
    .X(net4036));
 sg13g2_dlygate4sd3_1 hold1906 (.A(\mem.mem[24][0] ),
    .X(net4037));
 sg13g2_dlygate4sd3_1 hold1907 (.A(\mem.mem[205][4] ),
    .X(net4038));
 sg13g2_dlygate4sd3_1 hold1908 (.A(\mem.mem[198][2] ),
    .X(net4039));
 sg13g2_dlygate4sd3_1 hold1909 (.A(\mem.mem[95][0] ),
    .X(net4040));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\mem.mem[131][4] ),
    .X(net4041));
 sg13g2_dlygate4sd3_1 hold1911 (.A(\mem.mem[200][7] ),
    .X(net4042));
 sg13g2_dlygate4sd3_1 hold1912 (.A(\mem.mem[159][6] ),
    .X(net4043));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\mem.mem[66][1] ),
    .X(net4044));
 sg13g2_dlygate4sd3_1 hold1914 (.A(\mem.mem[76][1] ),
    .X(net4045));
 sg13g2_dlygate4sd3_1 hold1915 (.A(\mem.mem[68][6] ),
    .X(net4046));
 sg13g2_dlygate4sd3_1 hold1916 (.A(\mem.mem[161][3] ),
    .X(net4047));
 sg13g2_dlygate4sd3_1 hold1917 (.A(\mem.mem[252][7] ),
    .X(net4048));
 sg13g2_dlygate4sd3_1 hold1918 (.A(\mem.mem[4][1] ),
    .X(net4049));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\mem.mem[133][5] ),
    .X(net4050));
 sg13g2_dlygate4sd3_1 hold1920 (.A(\mem.mem[21][0] ),
    .X(net4051));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\mem.mem[68][3] ),
    .X(net4052));
 sg13g2_dlygate4sd3_1 hold1922 (.A(\mem.mem[201][1] ),
    .X(net4053));
 sg13g2_dlygate4sd3_1 hold1923 (.A(\mem.mem[21][7] ),
    .X(net4054));
 sg13g2_dlygate4sd3_1 hold1924 (.A(\mem.mem[140][1] ),
    .X(net4055));
 sg13g2_dlygate4sd3_1 hold1925 (.A(\mem.mem[202][0] ),
    .X(net4056));
 sg13g2_dlygate4sd3_1 hold1926 (.A(\mem.mem[195][6] ),
    .X(net4057));
 sg13g2_dlygate4sd3_1 hold1927 (.A(\mem.mem[79][0] ),
    .X(net4058));
 sg13g2_dlygate4sd3_1 hold1928 (.A(\mem.mem[146][1] ),
    .X(net4059));
 sg13g2_dlygate4sd3_1 hold1929 (.A(\mem.mem[24][3] ),
    .X(net4060));
 sg13g2_dlygate4sd3_1 hold1930 (.A(\mem.mem[145][1] ),
    .X(net4061));
 sg13g2_dlygate4sd3_1 hold1931 (.A(\mem.mem[248][7] ),
    .X(net4062));
 sg13g2_dlygate4sd3_1 hold1932 (.A(\mem.mem[203][5] ),
    .X(net4063));
 sg13g2_dlygate4sd3_1 hold1933 (.A(\mem.mem[77][6] ),
    .X(net4064));
 sg13g2_dlygate4sd3_1 hold1934 (.A(\mem.mem[239][1] ),
    .X(net4065));
 sg13g2_dlygate4sd3_1 hold1935 (.A(\mem.mem[35][5] ),
    .X(net4066));
 sg13g2_dlygate4sd3_1 hold1936 (.A(\mem.mem[41][2] ),
    .X(net4067));
 sg13g2_dlygate4sd3_1 hold1937 (.A(\mem.mem[134][6] ),
    .X(net4068));
 sg13g2_dlygate4sd3_1 hold1938 (.A(\mem.mem[195][4] ),
    .X(net4069));
 sg13g2_dlygate4sd3_1 hold1939 (.A(\mem.mem[10][0] ),
    .X(net4070));
 sg13g2_dlygate4sd3_1 hold1940 (.A(\mem.mem[145][6] ),
    .X(net4071));
 sg13g2_dlygate4sd3_1 hold1941 (.A(\mem.mem[34][3] ),
    .X(net4072));
 sg13g2_dlygate4sd3_1 hold1942 (.A(\mem.mem[195][2] ),
    .X(net4073));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\mem.mem[137][6] ),
    .X(net4074));
 sg13g2_dlygate4sd3_1 hold1944 (.A(\mem.mem[17][1] ),
    .X(net4075));
 sg13g2_dlygate4sd3_1 hold1945 (.A(\mem.mem[41][0] ),
    .X(net4076));
 sg13g2_dlygate4sd3_1 hold1946 (.A(\mem.mem[136][1] ),
    .X(net4077));
 sg13g2_dlygate4sd3_1 hold1947 (.A(\mem.mem[40][3] ),
    .X(net4078));
 sg13g2_dlygate4sd3_1 hold1948 (.A(\mem.mem[15][4] ),
    .X(net4079));
 sg13g2_dlygate4sd3_1 hold1949 (.A(\mem.mem[132][2] ),
    .X(net4080));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\mem.mem[10][7] ),
    .X(net4081));
 sg13g2_dlygate4sd3_1 hold1951 (.A(\mem.mem[33][7] ),
    .X(net4082));
 sg13g2_dlygate4sd3_1 hold1952 (.A(\mem.mem[28][3] ),
    .X(net4083));
 sg13g2_dlygate4sd3_1 hold1953 (.A(\mem.mem[141][5] ),
    .X(net4084));
 sg13g2_dlygate4sd3_1 hold1954 (.A(\mem.mem[207][2] ),
    .X(net4085));
 sg13g2_dlygate4sd3_1 hold1955 (.A(\mem.mem[111][4] ),
    .X(net4086));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\mem.mem[63][7] ),
    .X(net4087));
 sg13g2_dlygate4sd3_1 hold1957 (.A(\mem.mem[42][0] ),
    .X(net4088));
 sg13g2_dlygate4sd3_1 hold1958 (.A(\mem.mem[133][7] ),
    .X(net4089));
 sg13g2_dlygate4sd3_1 hold1959 (.A(\mem.mem[19][7] ),
    .X(net4090));
 sg13g2_dlygate4sd3_1 hold1960 (.A(\mem.mem[175][4] ),
    .X(net4091));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\mem.mem[20][1] ),
    .X(net4092));
 sg13g2_dlygate4sd3_1 hold1962 (.A(\mem.mem[239][4] ),
    .X(net4093));
 sg13g2_dlygate4sd3_1 hold1963 (.A(\mem.mem[18][1] ),
    .X(net4094));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\mem.mem[162][5] ),
    .X(net4095));
 sg13g2_dlygate4sd3_1 hold1965 (.A(\mem.mem[196][1] ),
    .X(net4096));
 sg13g2_dlygate4sd3_1 hold1966 (.A(\mem.mem[8][3] ),
    .X(net4097));
 sg13g2_dlygate4sd3_1 hold1967 (.A(\mem.mem[239][3] ),
    .X(net4098));
 sg13g2_dlygate4sd3_1 hold1968 (.A(\mem.mem[8][0] ),
    .X(net4099));
 sg13g2_dlygate4sd3_1 hold1969 (.A(\mem.mem[159][4] ),
    .X(net4100));
 sg13g2_dlygate4sd3_1 hold1970 (.A(\mem.mem[198][1] ),
    .X(net4101));
 sg13g2_dlygate4sd3_1 hold1971 (.A(\mem.mem[248][0] ),
    .X(net4102));
 sg13g2_dlygate4sd3_1 hold1972 (.A(\mem.mem[223][2] ),
    .X(net4103));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\mem.mem[37][0] ),
    .X(net4104));
 sg13g2_dlygate4sd3_1 hold1974 (.A(\mem.mem[193][0] ),
    .X(net4105));
 sg13g2_dlygate4sd3_1 hold1975 (.A(\mem.mem[24][2] ),
    .X(net4106));
 sg13g2_dlygate4sd3_1 hold1976 (.A(\mem.mem[10][5] ),
    .X(net4107));
 sg13g2_dlygate4sd3_1 hold1977 (.A(\mem.mem[97][0] ),
    .X(net4108));
 sg13g2_dlygate4sd3_1 hold1978 (.A(\mem.mem[15][0] ),
    .X(net4109));
 sg13g2_dlygate4sd3_1 hold1979 (.A(\mem.mem[26][1] ),
    .X(net4110));
 sg13g2_dlygate4sd3_1 hold1980 (.A(\mem.mem[98][2] ),
    .X(net4111));
 sg13g2_dlygate4sd3_1 hold1981 (.A(\mem.mem[75][6] ),
    .X(net4112));
 sg13g2_dlygate4sd3_1 hold1982 (.A(\mem.mem[194][6] ),
    .X(net4113));
 sg13g2_dlygate4sd3_1 hold1983 (.A(\mem.mem[133][3] ),
    .X(net4114));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\mem.mem[4][2] ),
    .X(net4115));
 sg13g2_dlygate4sd3_1 hold1985 (.A(\mem.mem[9][7] ),
    .X(net4116));
 sg13g2_dlygate4sd3_1 hold1986 (.A(\mem.mem[42][1] ),
    .X(net4117));
 sg13g2_dlygate4sd3_1 hold1987 (.A(\mem.mem[146][2] ),
    .X(net4118));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\mem.mem[42][5] ),
    .X(net4119));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\mem.mem[25][5] ),
    .X(net4120));
 sg13g2_dlygate4sd3_1 hold1990 (.A(\mem.mem[36][5] ),
    .X(net4121));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\mem.mem[36][4] ),
    .X(net4122));
 sg13g2_dlygate4sd3_1 hold1992 (.A(\mem.mem[13][0] ),
    .X(net4123));
 sg13g2_dlygate4sd3_1 hold1993 (.A(\mem.mem[6][1] ),
    .X(net4124));
 sg13g2_dlygate4sd3_1 hold1994 (.A(\mem.mem[140][6] ),
    .X(net4125));
 sg13g2_dlygate4sd3_1 hold1995 (.A(\mem.mem[63][4] ),
    .X(net4126));
 sg13g2_dlygate4sd3_1 hold1996 (.A(\mem.mem[3][4] ),
    .X(net4127));
 sg13g2_dlygate4sd3_1 hold1997 (.A(\mem.mem[82][1] ),
    .X(net4128));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\mem.mem[19][6] ),
    .X(net4129));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\mem.mem[2][7] ),
    .X(net4130));
 sg13g2_dlygate4sd3_1 hold2000 (.A(\mem.mem[132][4] ),
    .X(net4131));
 sg13g2_dlygate4sd3_1 hold2001 (.A(\mem.mem[69][4] ),
    .X(net4132));
 sg13g2_dlygate4sd3_1 hold2002 (.A(\mem.mem[19][0] ),
    .X(net4133));
 sg13g2_dlygate4sd3_1 hold2003 (.A(\mem.mem[139][6] ),
    .X(net4134));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\mem.mem[195][0] ),
    .X(net4135));
 sg13g2_dlygate4sd3_1 hold2005 (.A(\mem.mem[75][2] ),
    .X(net4136));
 sg13g2_dlygate4sd3_1 hold2006 (.A(\mem.mem[33][4] ),
    .X(net4137));
 sg13g2_dlygate4sd3_1 hold2007 (.A(\mem.mem[206][6] ),
    .X(net4138));
 sg13g2_dlygate4sd3_1 hold2008 (.A(\mem.mem[35][7] ),
    .X(net4139));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\mem.mem[1][6] ),
    .X(net4140));
 sg13g2_dlygate4sd3_1 hold2010 (.A(\mem.mem[193][5] ),
    .X(net4141));
 sg13g2_dlygate4sd3_1 hold2011 (.A(\mem.mem[111][0] ),
    .X(net4142));
 sg13g2_dlygate4sd3_1 hold2012 (.A(\mem.mem[3][7] ),
    .X(net4143));
 sg13g2_dlygate4sd3_1 hold2013 (.A(\mem.mem[11][6] ),
    .X(net4144));
 sg13g2_dlygate4sd3_1 hold2014 (.A(\mem.mem[129][7] ),
    .X(net4145));
 sg13g2_dlygate4sd3_1 hold2015 (.A(\mem.mem[52][6] ),
    .X(net4146));
 sg13g2_dlygate4sd3_1 hold2016 (.A(_00498_),
    .X(net4147));
 sg13g2_dlygate4sd3_1 hold2017 (.A(\mem.mem[141][3] ),
    .X(net4148));
 sg13g2_dlygate4sd3_1 hold2018 (.A(\mem.mem[175][3] ),
    .X(net4149));
 sg13g2_dlygate4sd3_1 hold2019 (.A(\mem.mem[133][6] ),
    .X(net4150));
 sg13g2_dlygate4sd3_1 hold2020 (.A(\mem.mem[206][1] ),
    .X(net4151));
 sg13g2_dlygate4sd3_1 hold2021 (.A(\mem_A[1] ),
    .X(net4152));
 sg13g2_dlygate4sd3_1 hold2022 (.A(\mem.mem[175][2] ),
    .X(net4153));
 sg13g2_dlygate4sd3_1 hold2023 (.A(\mem.mem[143][2] ),
    .X(net4154));
 sg13g2_dlygate4sd3_1 hold2024 (.A(\mem.mem[33][2] ),
    .X(net4155));
 sg13g2_dlygate4sd3_1 hold2025 (.A(\mem.mem[37][2] ),
    .X(net4156));
 sg13g2_dlygate4sd3_1 hold2026 (.A(\mem.mem[8][6] ),
    .X(net4157));
 sg13g2_dlygate4sd3_1 hold2027 (.A(\mem.mem[3][0] ),
    .X(net4158));
 sg13g2_dlygate4sd3_1 hold2028 (.A(\mem.mem[65][2] ),
    .X(net4159));
 sg13g2_dlygate4sd3_1 hold2029 (.A(\mem.mem[82][0] ),
    .X(net4160));
 sg13g2_dlygate4sd3_1 hold2030 (.A(\mem.mem[6][6] ),
    .X(net4161));
 sg13g2_dlygate4sd3_1 hold2031 (.A(\mem.mem[6][2] ),
    .X(net4162));
 sg13g2_dlygate4sd3_1 hold2032 (.A(\mem.mem[66][4] ),
    .X(net4163));
 sg13g2_dlygate4sd3_1 hold2033 (.A(\mem.mem[140][0] ),
    .X(net4164));
 sg13g2_dlygate4sd3_1 hold2034 (.A(\mem.data_in[5] ),
    .X(net4165));
 sg13g2_dlygate4sd3_1 hold2035 (.A(\mem.mem[193][6] ),
    .X(net4166));
 sg13g2_dlygate4sd3_1 hold2036 (.A(\mem.mem[40][7] ),
    .X(net4167));
 sg13g2_dlygate4sd3_1 hold2037 (.A(\mem.mem[175][5] ),
    .X(net4168));
 sg13g2_dlygate4sd3_1 hold2038 (.A(\C[2] ),
    .X(net4169));
 sg13g2_dlygate4sd3_1 hold2039 (.A(_00566_),
    .X(net4170));
 sg13g2_dlygate4sd3_1 hold2040 (.A(\C[1] ),
    .X(net4171));
 sg13g2_dlygate4sd3_1 hold2041 (.A(_00565_),
    .X(net4172));
 sg13g2_dlygate4sd3_1 hold2042 (.A(\mem.mem[3][3] ),
    .X(net4173));
 sg13g2_dlygate4sd3_1 hold2043 (.A(\C[4] ),
    .X(net4174));
 sg13g2_dlygate4sd3_1 hold2044 (.A(\C[7] ),
    .X(net4175));
 sg13g2_dlygate4sd3_1 hold2045 (.A(_00571_),
    .X(net4176));
 sg13g2_dlygate4sd3_1 hold2046 (.A(\C[6] ),
    .X(net4177));
 sg13g2_dlygate4sd3_1 hold2047 (.A(\A[5] ),
    .X(net4178));
 sg13g2_dlygate4sd3_1 hold2048 (.A(_00553_),
    .X(net4179));
 sg13g2_dlygate4sd3_1 hold2049 (.A(\mem.mem[11][2] ),
    .X(net4180));
 sg13g2_dlygate4sd3_1 hold2050 (.A(\A[3] ),
    .X(net4181));
 sg13g2_dlygate4sd3_1 hold2051 (.A(_00551_),
    .X(net4182));
 sg13g2_dlygate4sd3_1 hold2052 (.A(\A[0] ),
    .X(net4183));
 sg13g2_dlygate4sd3_1 hold2053 (.A(_00548_),
    .X(net4184));
 sg13g2_dlygate4sd3_1 hold2054 (.A(\C[0] ),
    .X(net4185));
 sg13g2_dlygate4sd3_1 hold2055 (.A(_00564_),
    .X(net4186));
 sg13g2_dlygate4sd3_1 hold2056 (.A(\A[4] ),
    .X(net4187));
 sg13g2_dlygate4sd3_1 hold2057 (.A(\A[6] ),
    .X(net4188));
 sg13g2_dlygate4sd3_1 hold2058 (.A(\B[6] ),
    .X(net4189));
 sg13g2_dlygate4sd3_1 hold2059 (.A(_05952_),
    .X(net4190));
 sg13g2_dlygate4sd3_1 hold2060 (.A(_00562_),
    .X(net4191));
 sg13g2_dlygate4sd3_1 hold2061 (.A(\B[5] ),
    .X(net4192));
 sg13g2_dlygate4sd3_1 hold2062 (.A(\B[0] ),
    .X(net4193));
 sg13g2_dlygate4sd3_1 hold2063 (.A(\B[3] ),
    .X(net4194));
 sg13g2_dlygate4sd3_1 hold2064 (.A(\A[1] ),
    .X(net4195));
 sg13g2_dlygate4sd3_1 hold2065 (.A(_00549_),
    .X(net4196));
 sg13g2_dlygate4sd3_1 hold2066 (.A(\A[2] ),
    .X(net4197));
 sg13g2_dlygate4sd3_1 hold2067 (.A(_00550_),
    .X(net4198));
 sg13g2_dlygate4sd3_1 hold2068 (.A(\B[4] ),
    .X(net4199));
 sg13g2_dlygate4sd3_1 hold2069 (.A(\A[7] ),
    .X(net4200));
 sg13g2_dlygate4sd3_1 hold2070 (.A(_05945_),
    .X(net4201));
 sg13g2_dlygate4sd3_1 hold2071 (.A(\B[2] ),
    .X(net4202));
 sg13g2_dlygate4sd3_1 hold2072 (.A(_05948_),
    .X(net4203));
 sg13g2_dlygate4sd3_1 hold2073 (.A(\B[7] ),
    .X(net4204));
 sg13g2_dlygate4sd3_1 hold2074 (.A(\mem_A[0] ),
    .X(net4205));
 sg13g2_dlygate4sd3_1 hold2075 (.A(\B[1] ),
    .X(net4206));
 sg13g2_dlygate4sd3_1 hold2076 (.A(\mem_A[2] ),
    .X(net4207));
 sg13g2_dlygate4sd3_1 hold2077 (.A(\mem_A[4] ),
    .X(net4208));
 sg13g2_dlygate4sd3_1 hold2078 (.A(\mem_A[7] ),
    .X(net4209));
 sg13g2_dlygate4sd3_1 hold2079 (.A(\mem_A[6] ),
    .X(net4210));
 sg13g2_dlygate4sd3_1 hold2080 (.A(\mem.data_in[6] ),
    .X(net4211));
 sg13g2_dlygate4sd3_1 hold2081 (.A(_06070_),
    .X(net4212));
 sg13g2_dlygate4sd3_1 hold2082 (.A(\mem_A[5] ),
    .X(net4213));
 sg13g2_dlygate4sd3_1 hold2083 (.A(_06082_),
    .X(net4214));
 sg13g2_dlygate4sd3_1 hold2084 (.A(\mem_A[3] ),
    .X(net4215));
 sg13g2_dlygate4sd3_1 hold2085 (.A(halted),
    .X(net4216));
 sg13g2_dlygate4sd3_1 hold2086 (.A(_02932_),
    .X(net4217));
 sg13g2_dlygate4sd3_1 hold2087 (.A(\mem.data_in[2] ),
    .X(net4218));
 sg13g2_dlygate4sd3_1 hold2088 (.A(\PC[5] ),
    .X(net4219));
 sg13g2_dlygate4sd3_1 hold2089 (.A(_00577_),
    .X(net4220));
 sg13g2_dlygate4sd3_1 hold2090 (.A(\PC[6] ),
    .X(net4221));
 sg13g2_dlygate4sd3_1 hold2091 (.A(_00578_),
    .X(net4222));
 sg13g2_dlygate4sd3_1 hold2092 (.A(\PC[0] ),
    .X(net4223));
 sg13g2_dlygate4sd3_1 hold2093 (.A(_00572_),
    .X(net4224));
 sg13g2_dlygate4sd3_1 hold2094 (.A(\mem.data_in[1] ),
    .X(net4225));
 sg13g2_dlygate4sd3_1 hold2095 (.A(_06029_),
    .X(net4226));
 sg13g2_dlygate4sd3_1 hold2096 (.A(prev_run),
    .X(net4227));
 sg13g2_dlygate4sd3_1 hold2097 (.A(\mem.data_in[4] ),
    .X(net4228));
 sg13g2_dlygate4sd3_1 hold2098 (.A(_06054_),
    .X(net4229));
 sg13g2_dlygate4sd3_1 hold2099 (.A(\PC[1] ),
    .X(net4230));
 sg13g2_dlygate4sd3_1 hold2100 (.A(\PC[3] ),
    .X(net4231));
 sg13g2_dlygate4sd3_1 hold2101 (.A(\PC[4] ),
    .X(net4232));
 sg13g2_dlygate4sd3_1 hold2102 (.A(_05991_),
    .X(net4233));
 sg13g2_dlygate4sd3_1 hold2103 (.A(\PC[7] ),
    .X(net4234));
 sg13g2_dlygate4sd3_1 hold2104 (.A(_00579_),
    .X(net4235));
 sg13g2_dlygate4sd3_1 hold2105 (.A(_00025_),
    .X(net4236));
 sg13g2_dlygate4sd3_1 hold2106 (.A(_03306_),
    .X(net4237));
 sg13g2_dlygate4sd3_1 hold2107 (.A(\mem.data_in[3] ),
    .X(net4238));
 sg13g2_dlygate4sd3_1 hold2108 (.A(\state[5] ),
    .X(net4239));
 sg13g2_dlygate4sd3_1 hold2109 (.A(\PC[2] ),
    .X(net4240));
 sg13g2_dlygate4sd3_1 hold2110 (.A(uo_out[5]),
    .X(net4241));
 sg13g2_dlygate4sd3_1 hold2111 (.A(uo_out[2]),
    .X(net4242));
 sg13g2_dlygate4sd3_1 hold2112 (.A(uo_out[4]),
    .X(net4243));
 sg13g2_dlygate4sd3_1 hold2113 (.A(\state[6] ),
    .X(net4244));
 sg13g2_dlygate4sd3_1 hold2114 (.A(uo_out[3]),
    .X(net4245));
 sg13g2_dlygate4sd3_1 hold2115 (.A(uo_out[1]),
    .X(net4246));
 sg13g2_dlygate4sd3_1 hold2116 (.A(uo_out[6]),
    .X(net4247));
 sg13g2_dlygate4sd3_1 hold2117 (.A(uo_out[0]),
    .X(net4248));
 sg13g2_dlygate4sd3_1 hold2118 (.A(_00805_),
    .X(net4249));
 sg13g2_dlygate4sd3_1 hold2119 (.A(uo_out[7]),
    .X(net4250));
 sg13g2_dlygate4sd3_1 hold2120 (.A(\mem.data_in[7] ),
    .X(net4251));
 sg13g2_dlygate4sd3_1 hold2121 (.A(\mem.addr[5] ),
    .X(net4252));
 sg13g2_dlygate4sd3_1 hold2122 (.A(\mem.addr[3] ),
    .X(net4253));
 sg13g2_dlygate4sd3_1 hold2123 (.A(\state[4] ),
    .X(net4254));
 sg13g2_dlygate4sd3_1 hold2124 (.A(\A[0] ),
    .X(net4255));
 sg13g2_dlygate4sd3_1 hold2125 (.A(_00580_),
    .X(net4256));
 sg13g2_dlygate4sd3_1 hold2126 (.A(\A[7] ),
    .X(net4257));
 sg13g2_antennanp ANTENNA_1 (.A(_03375_));
 sg13g2_antennanp ANTENNA_2 (.A(_03375_));
 sg13g2_antennanp ANTENNA_3 (.A(_03375_));
 sg13g2_antennanp ANTENNA_4 (.A(_03375_));
 sg13g2_antennanp ANTENNA_5 (.A(_03467_));
 sg13g2_antennanp ANTENNA_6 (.A(_03467_));
 sg13g2_antennanp ANTENNA_7 (.A(_03467_));
 sg13g2_antennanp ANTENNA_8 (.A(_03467_));
 sg13g2_antennanp ANTENNA_9 (.A(_03467_));
 sg13g2_antennanp ANTENNA_10 (.A(_03467_));
 sg13g2_antennanp ANTENNA_11 (.A(_03467_));
 sg13g2_antennanp ANTENNA_12 (.A(_03690_));
 sg13g2_antennanp ANTENNA_13 (.A(_03708_));
 sg13g2_antennanp ANTENNA_14 (.A(_03934_));
 sg13g2_antennanp ANTENNA_15 (.A(_04048_));
 sg13g2_antennanp ANTENNA_16 (.A(_04198_));
 sg13g2_antennanp ANTENNA_17 (.A(_04317_));
 sg13g2_antennanp ANTENNA_18 (.A(_04549_));
 sg13g2_antennanp ANTENNA_19 (.A(_04560_));
 sg13g2_antennanp ANTENNA_20 (.A(_04684_));
 sg13g2_antennanp ANTENNA_21 (.A(_04950_));
 sg13g2_antennanp ANTENNA_22 (.A(_05139_));
 sg13g2_antennanp ANTENNA_23 (.A(_05263_));
 sg13g2_antennanp ANTENNA_24 (.A(_05355_));
 sg13g2_antennanp ANTENNA_25 (.A(_05488_));
 sg13g2_antennanp ANTENNA_26 (.A(_05663_));
 sg13g2_antennanp ANTENNA_27 (.A(_05723_));
 sg13g2_antennanp ANTENNA_28 (.A(clk));
 sg13g2_antennanp ANTENNA_29 (.A(clk));
 sg13g2_antennanp ANTENNA_30 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_31 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_32 (.A(uo_out[5]));
 sg13g2_antennanp ANTENNA_33 (.A(uo_out[5]));
 sg13g2_antennanp ANTENNA_34 (.A(net5244));
 sg13g2_antennanp ANTENNA_35 (.A(net5244));
 sg13g2_antennanp ANTENNA_36 (.A(net5244));
 sg13g2_antennanp ANTENNA_37 (.A(net5244));
 sg13g2_antennanp ANTENNA_38 (.A(net5244));
 sg13g2_antennanp ANTENNA_39 (.A(net5244));
 sg13g2_antennanp ANTENNA_40 (.A(net5244));
 sg13g2_antennanp ANTENNA_41 (.A(net5244));
 sg13g2_antennanp ANTENNA_42 (.A(net5244));
 sg13g2_antennanp ANTENNA_43 (.A(net5244));
 sg13g2_antennanp ANTENNA_44 (.A(net5244));
 sg13g2_antennanp ANTENNA_45 (.A(net5244));
 sg13g2_antennanp ANTENNA_46 (.A(net5244));
 sg13g2_antennanp ANTENNA_47 (.A(net5244));
 sg13g2_antennanp ANTENNA_48 (.A(net5244));
 sg13g2_antennanp ANTENNA_49 (.A(net5244));
 sg13g2_antennanp ANTENNA_50 (.A(net5244));
 sg13g2_antennanp ANTENNA_51 (.A(net5244));
 sg13g2_antennanp ANTENNA_52 (.A(net5244));
 sg13g2_antennanp ANTENNA_53 (.A(net5244));
 sg13g2_antennanp ANTENNA_54 (.A(net5244));
 sg13g2_antennanp ANTENNA_55 (.A(net5244));
 sg13g2_antennanp ANTENNA_56 (.A(net5244));
 sg13g2_antennanp ANTENNA_57 (.A(net5244));
 sg13g2_antennanp ANTENNA_58 (.A(net5244));
 sg13g2_antennanp ANTENNA_59 (.A(net5244));
 sg13g2_antennanp ANTENNA_60 (.A(net5244));
 sg13g2_antennanp ANTENNA_61 (.A(net5244));
 sg13g2_antennanp ANTENNA_62 (.A(net5244));
 sg13g2_antennanp ANTENNA_63 (.A(net5244));
 sg13g2_antennanp ANTENNA_64 (.A(net5244));
 sg13g2_antennanp ANTENNA_65 (.A(net5244));
 sg13g2_antennanp ANTENNA_66 (.A(net5252));
 sg13g2_antennanp ANTENNA_67 (.A(net5252));
 sg13g2_antennanp ANTENNA_68 (.A(net5252));
 sg13g2_antennanp ANTENNA_69 (.A(net5252));
 sg13g2_antennanp ANTENNA_70 (.A(net5252));
 sg13g2_antennanp ANTENNA_71 (.A(net5252));
 sg13g2_antennanp ANTENNA_72 (.A(net5252));
 sg13g2_antennanp ANTENNA_73 (.A(net5252));
 sg13g2_antennanp ANTENNA_74 (.A(net5252));
 sg13g2_antennanp ANTENNA_75 (.A(net5252));
 sg13g2_antennanp ANTENNA_76 (.A(net5252));
 sg13g2_antennanp ANTENNA_77 (.A(net5252));
 sg13g2_antennanp ANTENNA_78 (.A(net5252));
 sg13g2_antennanp ANTENNA_79 (.A(net5252));
 sg13g2_antennanp ANTENNA_80 (.A(net5347));
 sg13g2_antennanp ANTENNA_81 (.A(net5347));
 sg13g2_antennanp ANTENNA_82 (.A(net5347));
 sg13g2_antennanp ANTENNA_83 (.A(net5347));
 sg13g2_antennanp ANTENNA_84 (.A(net5648));
 sg13g2_antennanp ANTENNA_85 (.A(net5648));
 sg13g2_antennanp ANTENNA_86 (.A(net5648));
 sg13g2_antennanp ANTENNA_87 (.A(net5648));
 sg13g2_antennanp ANTENNA_88 (.A(net5648));
 sg13g2_antennanp ANTENNA_89 (.A(net5648));
 sg13g2_antennanp ANTENNA_90 (.A(net5648));
 sg13g2_antennanp ANTENNA_91 (.A(net5648));
 sg13g2_antennanp ANTENNA_92 (.A(net5648));
 sg13g2_antennanp ANTENNA_93 (.A(net5648));
 sg13g2_antennanp ANTENNA_94 (.A(net5648));
 sg13g2_antennanp ANTENNA_95 (.A(net5884));
 sg13g2_antennanp ANTENNA_96 (.A(net5884));
 sg13g2_antennanp ANTENNA_97 (.A(net5884));
 sg13g2_antennanp ANTENNA_98 (.A(net5884));
 sg13g2_antennanp ANTENNA_99 (.A(net5884));
 sg13g2_antennanp ANTENNA_100 (.A(net5884));
 sg13g2_antennanp ANTENNA_101 (.A(net5884));
 sg13g2_antennanp ANTENNA_102 (.A(net5884));
 sg13g2_antennanp ANTENNA_103 (.A(net5884));
 sg13g2_antennanp ANTENNA_104 (.A(_02964_));
 sg13g2_antennanp ANTENNA_105 (.A(_02964_));
 sg13g2_antennanp ANTENNA_106 (.A(_02964_));
 sg13g2_antennanp ANTENNA_107 (.A(_02964_));
 sg13g2_antennanp ANTENNA_108 (.A(_02964_));
 sg13g2_antennanp ANTENNA_109 (.A(_02964_));
 sg13g2_antennanp ANTENNA_110 (.A(_02964_));
 sg13g2_antennanp ANTENNA_111 (.A(_02964_));
 sg13g2_antennanp ANTENNA_112 (.A(_02964_));
 sg13g2_antennanp ANTENNA_113 (.A(_02981_));
 sg13g2_antennanp ANTENNA_114 (.A(_02981_));
 sg13g2_antennanp ANTENNA_115 (.A(_02981_));
 sg13g2_antennanp ANTENNA_116 (.A(_02981_));
 sg13g2_antennanp ANTENNA_117 (.A(_02981_));
 sg13g2_antennanp ANTENNA_118 (.A(_02981_));
 sg13g2_antennanp ANTENNA_119 (.A(_02981_));
 sg13g2_antennanp ANTENNA_120 (.A(_03375_));
 sg13g2_antennanp ANTENNA_121 (.A(_03375_));
 sg13g2_antennanp ANTENNA_122 (.A(_03375_));
 sg13g2_antennanp ANTENNA_123 (.A(_03375_));
 sg13g2_antennanp ANTENNA_124 (.A(_03467_));
 sg13g2_antennanp ANTENNA_125 (.A(_03467_));
 sg13g2_antennanp ANTENNA_126 (.A(_03467_));
 sg13g2_antennanp ANTENNA_127 (.A(_03467_));
 sg13g2_antennanp ANTENNA_128 (.A(_03467_));
 sg13g2_antennanp ANTENNA_129 (.A(_03467_));
 sg13g2_antennanp ANTENNA_130 (.A(_03467_));
 sg13g2_antennanp ANTENNA_131 (.A(_03467_));
 sg13g2_antennanp ANTENNA_132 (.A(_03467_));
 sg13g2_antennanp ANTENNA_133 (.A(_03467_));
 sg13g2_antennanp ANTENNA_134 (.A(_03467_));
 sg13g2_antennanp ANTENNA_135 (.A(_03467_));
 sg13g2_antennanp ANTENNA_136 (.A(_03467_));
 sg13g2_antennanp ANTENNA_137 (.A(_03690_));
 sg13g2_antennanp ANTENNA_138 (.A(_03708_));
 sg13g2_antennanp ANTENNA_139 (.A(_03934_));
 sg13g2_antennanp ANTENNA_140 (.A(_04048_));
 sg13g2_antennanp ANTENNA_141 (.A(_04317_));
 sg13g2_antennanp ANTENNA_142 (.A(_04549_));
 sg13g2_antennanp ANTENNA_143 (.A(_04560_));
 sg13g2_antennanp ANTENNA_144 (.A(_04684_));
 sg13g2_antennanp ANTENNA_145 (.A(_04950_));
 sg13g2_antennanp ANTENNA_146 (.A(_05139_));
 sg13g2_antennanp ANTENNA_147 (.A(_05263_));
 sg13g2_antennanp ANTENNA_148 (.A(_05355_));
 sg13g2_antennanp ANTENNA_149 (.A(_05488_));
 sg13g2_antennanp ANTENNA_150 (.A(_05663_));
 sg13g2_antennanp ANTENNA_151 (.A(_05723_));
 sg13g2_antennanp ANTENNA_152 (.A(clk));
 sg13g2_antennanp ANTENNA_153 (.A(clk));
 sg13g2_antennanp ANTENNA_154 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_155 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_156 (.A(uo_out[5]));
 sg13g2_antennanp ANTENNA_157 (.A(net5230));
 sg13g2_antennanp ANTENNA_158 (.A(net5230));
 sg13g2_antennanp ANTENNA_159 (.A(net5230));
 sg13g2_antennanp ANTENNA_160 (.A(net5230));
 sg13g2_antennanp ANTENNA_161 (.A(net5230));
 sg13g2_antennanp ANTENNA_162 (.A(net5230));
 sg13g2_antennanp ANTENNA_163 (.A(net5230));
 sg13g2_antennanp ANTENNA_164 (.A(net5230));
 sg13g2_antennanp ANTENNA_165 (.A(net5236));
 sg13g2_antennanp ANTENNA_166 (.A(net5236));
 sg13g2_antennanp ANTENNA_167 (.A(net5236));
 sg13g2_antennanp ANTENNA_168 (.A(net5236));
 sg13g2_antennanp ANTENNA_169 (.A(net5236));
 sg13g2_antennanp ANTENNA_170 (.A(net5236));
 sg13g2_antennanp ANTENNA_171 (.A(net5236));
 sg13g2_antennanp ANTENNA_172 (.A(net5236));
 sg13g2_antennanp ANTENNA_173 (.A(net5236));
 sg13g2_antennanp ANTENNA_174 (.A(net5236));
 sg13g2_antennanp ANTENNA_175 (.A(net5236));
 sg13g2_antennanp ANTENNA_176 (.A(net5236));
 sg13g2_antennanp ANTENNA_177 (.A(net5236));
 sg13g2_antennanp ANTENNA_178 (.A(net5236));
 sg13g2_antennanp ANTENNA_179 (.A(net5236));
 sg13g2_antennanp ANTENNA_180 (.A(net5236));
 sg13g2_antennanp ANTENNA_181 (.A(net5236));
 sg13g2_antennanp ANTENNA_182 (.A(net5236));
 sg13g2_antennanp ANTENNA_183 (.A(net5236));
 sg13g2_antennanp ANTENNA_184 (.A(net5236));
 sg13g2_antennanp ANTENNA_185 (.A(net5236));
 sg13g2_antennanp ANTENNA_186 (.A(net5236));
 sg13g2_antennanp ANTENNA_187 (.A(net5236));
 sg13g2_antennanp ANTENNA_188 (.A(net5236));
 sg13g2_antennanp ANTENNA_189 (.A(net5236));
 sg13g2_antennanp ANTENNA_190 (.A(net5236));
 sg13g2_antennanp ANTENNA_191 (.A(net5236));
 sg13g2_antennanp ANTENNA_192 (.A(net5236));
 sg13g2_antennanp ANTENNA_193 (.A(net5236));
 sg13g2_antennanp ANTENNA_194 (.A(net5236));
 sg13g2_antennanp ANTENNA_195 (.A(net5239));
 sg13g2_antennanp ANTENNA_196 (.A(net5239));
 sg13g2_antennanp ANTENNA_197 (.A(net5239));
 sg13g2_antennanp ANTENNA_198 (.A(net5239));
 sg13g2_antennanp ANTENNA_199 (.A(net5239));
 sg13g2_antennanp ANTENNA_200 (.A(net5239));
 sg13g2_antennanp ANTENNA_201 (.A(net5239));
 sg13g2_antennanp ANTENNA_202 (.A(net5239));
 sg13g2_antennanp ANTENNA_203 (.A(net5242));
 sg13g2_antennanp ANTENNA_204 (.A(net5242));
 sg13g2_antennanp ANTENNA_205 (.A(net5242));
 sg13g2_antennanp ANTENNA_206 (.A(net5242));
 sg13g2_antennanp ANTENNA_207 (.A(net5242));
 sg13g2_antennanp ANTENNA_208 (.A(net5242));
 sg13g2_antennanp ANTENNA_209 (.A(net5242));
 sg13g2_antennanp ANTENNA_210 (.A(net5242));
 sg13g2_antennanp ANTENNA_211 (.A(net5244));
 sg13g2_antennanp ANTENNA_212 (.A(net5244));
 sg13g2_antennanp ANTENNA_213 (.A(net5244));
 sg13g2_antennanp ANTENNA_214 (.A(net5244));
 sg13g2_antennanp ANTENNA_215 (.A(net5244));
 sg13g2_antennanp ANTENNA_216 (.A(net5244));
 sg13g2_antennanp ANTENNA_217 (.A(net5244));
 sg13g2_antennanp ANTENNA_218 (.A(net5244));
 sg13g2_antennanp ANTENNA_219 (.A(net5244));
 sg13g2_antennanp ANTENNA_220 (.A(net5244));
 sg13g2_antennanp ANTENNA_221 (.A(net5244));
 sg13g2_antennanp ANTENNA_222 (.A(net5244));
 sg13g2_antennanp ANTENNA_223 (.A(net5244));
 sg13g2_antennanp ANTENNA_224 (.A(net5244));
 sg13g2_antennanp ANTENNA_225 (.A(net5244));
 sg13g2_antennanp ANTENNA_226 (.A(net5244));
 sg13g2_antennanp ANTENNA_227 (.A(net5244));
 sg13g2_antennanp ANTENNA_228 (.A(net5251));
 sg13g2_antennanp ANTENNA_229 (.A(net5251));
 sg13g2_antennanp ANTENNA_230 (.A(net5251));
 sg13g2_antennanp ANTENNA_231 (.A(net5251));
 sg13g2_antennanp ANTENNA_232 (.A(net5251));
 sg13g2_antennanp ANTENNA_233 (.A(net5251));
 sg13g2_antennanp ANTENNA_234 (.A(net5251));
 sg13g2_antennanp ANTENNA_235 (.A(net5251));
 sg13g2_antennanp ANTENNA_236 (.A(net5251));
 sg13g2_antennanp ANTENNA_237 (.A(net5251));
 sg13g2_antennanp ANTENNA_238 (.A(net5251));
 sg13g2_antennanp ANTENNA_239 (.A(net5251));
 sg13g2_antennanp ANTENNA_240 (.A(net5251));
 sg13g2_antennanp ANTENNA_241 (.A(net5286));
 sg13g2_antennanp ANTENNA_242 (.A(net5286));
 sg13g2_antennanp ANTENNA_243 (.A(net5286));
 sg13g2_antennanp ANTENNA_244 (.A(net5286));
 sg13g2_antennanp ANTENNA_245 (.A(net5286));
 sg13g2_antennanp ANTENNA_246 (.A(net5286));
 sg13g2_antennanp ANTENNA_247 (.A(net5286));
 sg13g2_antennanp ANTENNA_248 (.A(net5286));
 sg13g2_antennanp ANTENNA_249 (.A(net5347));
 sg13g2_antennanp ANTENNA_250 (.A(net5347));
 sg13g2_antennanp ANTENNA_251 (.A(net5347));
 sg13g2_antennanp ANTENNA_252 (.A(net5347));
 sg13g2_antennanp ANTENNA_253 (.A(_03375_));
 sg13g2_antennanp ANTENNA_254 (.A(_03375_));
 sg13g2_antennanp ANTENNA_255 (.A(_03375_));
 sg13g2_antennanp ANTENNA_256 (.A(_03375_));
 sg13g2_antennanp ANTENNA_257 (.A(_03467_));
 sg13g2_antennanp ANTENNA_258 (.A(_03467_));
 sg13g2_antennanp ANTENNA_259 (.A(_03467_));
 sg13g2_antennanp ANTENNA_260 (.A(_03467_));
 sg13g2_antennanp ANTENNA_261 (.A(_03467_));
 sg13g2_antennanp ANTENNA_262 (.A(_03467_));
 sg13g2_antennanp ANTENNA_263 (.A(_03467_));
 sg13g2_antennanp ANTENNA_264 (.A(_03467_));
 sg13g2_antennanp ANTENNA_265 (.A(_03467_));
 sg13g2_antennanp ANTENNA_266 (.A(_03467_));
 sg13g2_antennanp ANTENNA_267 (.A(_03467_));
 sg13g2_antennanp ANTENNA_268 (.A(_03467_));
 sg13g2_antennanp ANTENNA_269 (.A(_03467_));
 sg13g2_antennanp ANTENNA_270 (.A(_03467_));
 sg13g2_antennanp ANTENNA_271 (.A(_03467_));
 sg13g2_antennanp ANTENNA_272 (.A(_03467_));
 sg13g2_antennanp ANTENNA_273 (.A(_03690_));
 sg13g2_antennanp ANTENNA_274 (.A(_03708_));
 sg13g2_antennanp ANTENNA_275 (.A(_03934_));
 sg13g2_antennanp ANTENNA_276 (.A(_04048_));
 sg13g2_antennanp ANTENNA_277 (.A(_04317_));
 sg13g2_antennanp ANTENNA_278 (.A(_04560_));
 sg13g2_antennanp ANTENNA_279 (.A(_04684_));
 sg13g2_antennanp ANTENNA_280 (.A(_04950_));
 sg13g2_antennanp ANTENNA_281 (.A(_05012_));
 sg13g2_antennanp ANTENNA_282 (.A(_05139_));
 sg13g2_antennanp ANTENNA_283 (.A(_05263_));
 sg13g2_antennanp ANTENNA_284 (.A(_05355_));
 sg13g2_antennanp ANTENNA_285 (.A(_05488_));
 sg13g2_antennanp ANTENNA_286 (.A(_05723_));
 sg13g2_antennanp ANTENNA_287 (.A(clk));
 sg13g2_antennanp ANTENNA_288 (.A(clk));
 sg13g2_antennanp ANTENNA_289 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_290 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_291 (.A(uo_out[5]));
 sg13g2_antennanp ANTENNA_292 (.A(net5230));
 sg13g2_antennanp ANTENNA_293 (.A(net5230));
 sg13g2_antennanp ANTENNA_294 (.A(net5230));
 sg13g2_antennanp ANTENNA_295 (.A(net5230));
 sg13g2_antennanp ANTENNA_296 (.A(net5230));
 sg13g2_antennanp ANTENNA_297 (.A(net5230));
 sg13g2_antennanp ANTENNA_298 (.A(net5230));
 sg13g2_antennanp ANTENNA_299 (.A(net5230));
 sg13g2_antennanp ANTENNA_300 (.A(net5230));
 sg13g2_antennanp ANTENNA_301 (.A(net5239));
 sg13g2_antennanp ANTENNA_302 (.A(net5239));
 sg13g2_antennanp ANTENNA_303 (.A(net5239));
 sg13g2_antennanp ANTENNA_304 (.A(net5239));
 sg13g2_antennanp ANTENNA_305 (.A(net5239));
 sg13g2_antennanp ANTENNA_306 (.A(net5239));
 sg13g2_antennanp ANTENNA_307 (.A(net5239));
 sg13g2_antennanp ANTENNA_308 (.A(net5239));
 sg13g2_antennanp ANTENNA_309 (.A(net5239));
 sg13g2_antennanp ANTENNA_310 (.A(net5239));
 sg13g2_antennanp ANTENNA_311 (.A(net5239));
 sg13g2_antennanp ANTENNA_312 (.A(net5239));
 sg13g2_antennanp ANTENNA_313 (.A(net5239));
 sg13g2_antennanp ANTENNA_314 (.A(net5239));
 sg13g2_antennanp ANTENNA_315 (.A(net5242));
 sg13g2_antennanp ANTENNA_316 (.A(net5242));
 sg13g2_antennanp ANTENNA_317 (.A(net5242));
 sg13g2_antennanp ANTENNA_318 (.A(net5242));
 sg13g2_antennanp ANTENNA_319 (.A(net5242));
 sg13g2_antennanp ANTENNA_320 (.A(net5242));
 sg13g2_antennanp ANTENNA_321 (.A(net5242));
 sg13g2_antennanp ANTENNA_322 (.A(net5242));
 sg13g2_antennanp ANTENNA_323 (.A(net5242));
 sg13g2_antennanp ANTENNA_324 (.A(net5242));
 sg13g2_antennanp ANTENNA_325 (.A(net5242));
 sg13g2_antennanp ANTENNA_326 (.A(net5242));
 sg13g2_antennanp ANTENNA_327 (.A(net5242));
 sg13g2_antennanp ANTENNA_328 (.A(net5242));
 sg13g2_antennanp ANTENNA_329 (.A(net5242));
 sg13g2_antennanp ANTENNA_330 (.A(net5242));
 sg13g2_antennanp ANTENNA_331 (.A(net5347));
 sg13g2_antennanp ANTENNA_332 (.A(net5347));
 sg13g2_antennanp ANTENNA_333 (.A(net5347));
 sg13g2_antennanp ANTENNA_334 (.A(net5347));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_fill_2 FILLER_0_518 ();
 sg13g2_fill_1 FILLER_0_520 ();
 sg13g2_fill_2 FILLER_0_551 ();
 sg13g2_fill_1 FILLER_0_558 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_fill_1 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_587 ();
 sg13g2_decap_8 FILLER_0_594 ();
 sg13g2_fill_1 FILLER_0_601 ();
 sg13g2_fill_1 FILLER_0_619 ();
 sg13g2_decap_8 FILLER_0_628 ();
 sg13g2_decap_8 FILLER_0_635 ();
 sg13g2_decap_8 FILLER_0_642 ();
 sg13g2_decap_8 FILLER_0_649 ();
 sg13g2_decap_8 FILLER_0_656 ();
 sg13g2_decap_8 FILLER_0_663 ();
 sg13g2_decap_8 FILLER_0_670 ();
 sg13g2_decap_8 FILLER_0_677 ();
 sg13g2_decap_8 FILLER_0_684 ();
 sg13g2_decap_8 FILLER_0_691 ();
 sg13g2_decap_8 FILLER_0_698 ();
 sg13g2_decap_8 FILLER_0_705 ();
 sg13g2_decap_8 FILLER_0_712 ();
 sg13g2_decap_4 FILLER_0_719 ();
 sg13g2_fill_2 FILLER_0_723 ();
 sg13g2_decap_8 FILLER_0_729 ();
 sg13g2_decap_8 FILLER_0_736 ();
 sg13g2_decap_8 FILLER_0_743 ();
 sg13g2_decap_8 FILLER_0_750 ();
 sg13g2_decap_8 FILLER_0_757 ();
 sg13g2_decap_8 FILLER_0_764 ();
 sg13g2_decap_8 FILLER_0_775 ();
 sg13g2_decap_8 FILLER_0_782 ();
 sg13g2_decap_8 FILLER_0_789 ();
 sg13g2_decap_8 FILLER_0_796 ();
 sg13g2_decap_8 FILLER_0_803 ();
 sg13g2_decap_8 FILLER_0_810 ();
 sg13g2_decap_8 FILLER_0_817 ();
 sg13g2_decap_8 FILLER_0_824 ();
 sg13g2_decap_8 FILLER_0_831 ();
 sg13g2_decap_8 FILLER_0_838 ();
 sg13g2_decap_8 FILLER_0_845 ();
 sg13g2_decap_8 FILLER_0_852 ();
 sg13g2_decap_8 FILLER_0_859 ();
 sg13g2_decap_8 FILLER_0_866 ();
 sg13g2_decap_8 FILLER_0_873 ();
 sg13g2_decap_8 FILLER_0_880 ();
 sg13g2_decap_8 FILLER_0_887 ();
 sg13g2_decap_8 FILLER_0_894 ();
 sg13g2_decap_8 FILLER_0_901 ();
 sg13g2_decap_8 FILLER_0_908 ();
 sg13g2_decap_8 FILLER_0_915 ();
 sg13g2_decap_8 FILLER_0_922 ();
 sg13g2_decap_8 FILLER_0_929 ();
 sg13g2_decap_8 FILLER_0_936 ();
 sg13g2_decap_8 FILLER_0_943 ();
 sg13g2_decap_8 FILLER_0_950 ();
 sg13g2_decap_8 FILLER_0_957 ();
 sg13g2_decap_8 FILLER_0_964 ();
 sg13g2_decap_8 FILLER_0_971 ();
 sg13g2_decap_8 FILLER_0_978 ();
 sg13g2_decap_8 FILLER_0_985 ();
 sg13g2_decap_8 FILLER_0_992 ();
 sg13g2_decap_8 FILLER_0_999 ();
 sg13g2_decap_8 FILLER_0_1006 ();
 sg13g2_decap_8 FILLER_0_1013 ();
 sg13g2_decap_8 FILLER_0_1020 ();
 sg13g2_decap_8 FILLER_0_1027 ();
 sg13g2_decap_8 FILLER_0_1034 ();
 sg13g2_decap_8 FILLER_0_1041 ();
 sg13g2_decap_8 FILLER_0_1048 ();
 sg13g2_decap_8 FILLER_0_1055 ();
 sg13g2_decap_8 FILLER_0_1062 ();
 sg13g2_decap_8 FILLER_0_1069 ();
 sg13g2_decap_8 FILLER_0_1076 ();
 sg13g2_decap_8 FILLER_0_1083 ();
 sg13g2_decap_8 FILLER_0_1090 ();
 sg13g2_decap_8 FILLER_0_1097 ();
 sg13g2_decap_8 FILLER_0_1104 ();
 sg13g2_decap_8 FILLER_0_1111 ();
 sg13g2_decap_8 FILLER_0_1118 ();
 sg13g2_decap_8 FILLER_0_1125 ();
 sg13g2_decap_8 FILLER_0_1132 ();
 sg13g2_fill_1 FILLER_0_1139 ();
 sg13g2_fill_2 FILLER_0_1144 ();
 sg13g2_fill_2 FILLER_0_1150 ();
 sg13g2_decap_8 FILLER_0_1161 ();
 sg13g2_decap_8 FILLER_0_1168 ();
 sg13g2_decap_8 FILLER_0_1175 ();
 sg13g2_decap_8 FILLER_0_1182 ();
 sg13g2_fill_2 FILLER_0_1189 ();
 sg13g2_fill_1 FILLER_0_1191 ();
 sg13g2_decap_8 FILLER_0_1196 ();
 sg13g2_decap_8 FILLER_0_1203 ();
 sg13g2_decap_8 FILLER_0_1210 ();
 sg13g2_decap_8 FILLER_0_1217 ();
 sg13g2_decap_8 FILLER_0_1224 ();
 sg13g2_decap_8 FILLER_0_1231 ();
 sg13g2_decap_8 FILLER_0_1238 ();
 sg13g2_decap_8 FILLER_0_1245 ();
 sg13g2_decap_8 FILLER_0_1252 ();
 sg13g2_fill_2 FILLER_0_1316 ();
 sg13g2_fill_1 FILLER_0_1318 ();
 sg13g2_fill_1 FILLER_0_1332 ();
 sg13g2_fill_1 FILLER_0_1355 ();
 sg13g2_fill_2 FILLER_0_1370 ();
 sg13g2_decap_4 FILLER_0_1376 ();
 sg13g2_fill_1 FILLER_0_1380 ();
 sg13g2_decap_4 FILLER_0_1415 ();
 sg13g2_fill_1 FILLER_0_1419 ();
 sg13g2_decap_8 FILLER_0_1425 ();
 sg13g2_decap_8 FILLER_0_1440 ();
 sg13g2_decap_8 FILLER_0_1447 ();
 sg13g2_decap_8 FILLER_0_1454 ();
 sg13g2_decap_8 FILLER_0_1461 ();
 sg13g2_decap_8 FILLER_0_1468 ();
 sg13g2_decap_8 FILLER_0_1475 ();
 sg13g2_decap_8 FILLER_0_1482 ();
 sg13g2_decap_8 FILLER_0_1489 ();
 sg13g2_decap_8 FILLER_0_1496 ();
 sg13g2_decap_8 FILLER_0_1503 ();
 sg13g2_decap_8 FILLER_0_1510 ();
 sg13g2_decap_8 FILLER_0_1517 ();
 sg13g2_fill_2 FILLER_0_1524 ();
 sg13g2_fill_1 FILLER_0_1526 ();
 sg13g2_fill_2 FILLER_0_1563 ();
 sg13g2_fill_1 FILLER_0_1565 ();
 sg13g2_fill_2 FILLER_0_1570 ();
 sg13g2_fill_1 FILLER_0_1572 ();
 sg13g2_fill_2 FILLER_0_1591 ();
 sg13g2_fill_2 FILLER_0_1616 ();
 sg13g2_decap_8 FILLER_0_1682 ();
 sg13g2_decap_8 FILLER_0_1689 ();
 sg13g2_fill_2 FILLER_0_1696 ();
 sg13g2_decap_8 FILLER_0_1702 ();
 sg13g2_fill_1 FILLER_0_1709 ();
 sg13g2_fill_2 FILLER_0_1719 ();
 sg13g2_fill_1 FILLER_0_1721 ();
 sg13g2_decap_8 FILLER_0_1787 ();
 sg13g2_fill_2 FILLER_0_1794 ();
 sg13g2_fill_1 FILLER_0_1796 ();
 sg13g2_decap_8 FILLER_0_1802 ();
 sg13g2_decap_8 FILLER_0_1809 ();
 sg13g2_decap_8 FILLER_0_1816 ();
 sg13g2_decap_8 FILLER_0_1823 ();
 sg13g2_decap_8 FILLER_0_1830 ();
 sg13g2_fill_2 FILLER_0_1837 ();
 sg13g2_fill_1 FILLER_0_1839 ();
 sg13g2_fill_2 FILLER_0_1853 ();
 sg13g2_fill_2 FILLER_0_1881 ();
 sg13g2_fill_1 FILLER_0_1896 ();
 sg13g2_decap_8 FILLER_0_1928 ();
 sg13g2_fill_1 FILLER_0_1935 ();
 sg13g2_fill_2 FILLER_0_1966 ();
 sg13g2_fill_1 FILLER_0_1968 ();
 sg13g2_fill_1 FILLER_0_2008 ();
 sg13g2_decap_8 FILLER_0_2044 ();
 sg13g2_decap_8 FILLER_0_2051 ();
 sg13g2_decap_4 FILLER_0_2058 ();
 sg13g2_fill_2 FILLER_0_2062 ();
 sg13g2_fill_2 FILLER_0_2103 ();
 sg13g2_fill_1 FILLER_0_2105 ();
 sg13g2_fill_2 FILLER_0_2119 ();
 sg13g2_fill_1 FILLER_0_2125 ();
 sg13g2_decap_4 FILLER_0_2165 ();
 sg13g2_fill_2 FILLER_0_2169 ();
 sg13g2_decap_8 FILLER_0_2175 ();
 sg13g2_decap_8 FILLER_0_2208 ();
 sg13g2_decap_8 FILLER_0_2215 ();
 sg13g2_decap_8 FILLER_0_2222 ();
 sg13g2_fill_1 FILLER_0_2229 ();
 sg13g2_decap_8 FILLER_0_2234 ();
 sg13g2_fill_2 FILLER_0_2241 ();
 sg13g2_decap_8 FILLER_0_2247 ();
 sg13g2_decap_8 FILLER_0_2254 ();
 sg13g2_decap_8 FILLER_0_2261 ();
 sg13g2_decap_8 FILLER_0_2268 ();
 sg13g2_decap_8 FILLER_0_2275 ();
 sg13g2_decap_8 FILLER_0_2282 ();
 sg13g2_decap_8 FILLER_0_2289 ();
 sg13g2_decap_8 FILLER_0_2296 ();
 sg13g2_decap_8 FILLER_0_2303 ();
 sg13g2_decap_8 FILLER_0_2310 ();
 sg13g2_decap_8 FILLER_0_2317 ();
 sg13g2_decap_8 FILLER_0_2324 ();
 sg13g2_decap_8 FILLER_0_2331 ();
 sg13g2_decap_8 FILLER_0_2338 ();
 sg13g2_decap_8 FILLER_0_2345 ();
 sg13g2_decap_8 FILLER_0_2352 ();
 sg13g2_decap_8 FILLER_0_2359 ();
 sg13g2_decap_8 FILLER_0_2366 ();
 sg13g2_decap_8 FILLER_0_2373 ();
 sg13g2_decap_8 FILLER_0_2380 ();
 sg13g2_decap_8 FILLER_0_2387 ();
 sg13g2_decap_8 FILLER_0_2394 ();
 sg13g2_decap_8 FILLER_0_2401 ();
 sg13g2_decap_8 FILLER_0_2408 ();
 sg13g2_decap_8 FILLER_0_2415 ();
 sg13g2_decap_8 FILLER_0_2422 ();
 sg13g2_decap_8 FILLER_0_2429 ();
 sg13g2_decap_8 FILLER_0_2436 ();
 sg13g2_decap_8 FILLER_0_2443 ();
 sg13g2_decap_8 FILLER_0_2450 ();
 sg13g2_decap_8 FILLER_0_2457 ();
 sg13g2_decap_8 FILLER_0_2464 ();
 sg13g2_decap_8 FILLER_0_2471 ();
 sg13g2_decap_8 FILLER_0_2478 ();
 sg13g2_decap_8 FILLER_0_2485 ();
 sg13g2_decap_8 FILLER_0_2492 ();
 sg13g2_decap_8 FILLER_0_2499 ();
 sg13g2_decap_8 FILLER_0_2506 ();
 sg13g2_decap_8 FILLER_0_2513 ();
 sg13g2_decap_8 FILLER_0_2520 ();
 sg13g2_decap_8 FILLER_0_2527 ();
 sg13g2_decap_8 FILLER_0_2534 ();
 sg13g2_decap_8 FILLER_0_2541 ();
 sg13g2_decap_8 FILLER_0_2548 ();
 sg13g2_decap_8 FILLER_0_2555 ();
 sg13g2_decap_8 FILLER_0_2562 ();
 sg13g2_decap_8 FILLER_0_2569 ();
 sg13g2_decap_8 FILLER_0_2576 ();
 sg13g2_decap_8 FILLER_0_2583 ();
 sg13g2_decap_8 FILLER_0_2590 ();
 sg13g2_decap_8 FILLER_0_2597 ();
 sg13g2_decap_8 FILLER_0_2604 ();
 sg13g2_decap_8 FILLER_0_2611 ();
 sg13g2_decap_8 FILLER_0_2618 ();
 sg13g2_decap_8 FILLER_0_2625 ();
 sg13g2_decap_8 FILLER_0_2632 ();
 sg13g2_decap_8 FILLER_0_2639 ();
 sg13g2_decap_8 FILLER_0_2646 ();
 sg13g2_decap_8 FILLER_0_2653 ();
 sg13g2_decap_8 FILLER_0_2660 ();
 sg13g2_decap_8 FILLER_0_2667 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_fill_1 FILLER_1_518 ();
 sg13g2_fill_2 FILLER_1_523 ();
 sg13g2_fill_1 FILLER_1_525 ();
 sg13g2_decap_4 FILLER_1_583 ();
 sg13g2_decap_4 FILLER_1_653 ();
 sg13g2_fill_1 FILLER_1_657 ();
 sg13g2_decap_8 FILLER_1_662 ();
 sg13g2_decap_8 FILLER_1_669 ();
 sg13g2_decap_8 FILLER_1_676 ();
 sg13g2_fill_2 FILLER_1_683 ();
 sg13g2_decap_8 FILLER_1_737 ();
 sg13g2_decap_8 FILLER_1_744 ();
 sg13g2_decap_8 FILLER_1_751 ();
 sg13g2_fill_2 FILLER_1_758 ();
 sg13g2_fill_1 FILLER_1_786 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_decap_8 FILLER_1_875 ();
 sg13g2_decap_8 FILLER_1_882 ();
 sg13g2_decap_8 FILLER_1_889 ();
 sg13g2_decap_8 FILLER_1_896 ();
 sg13g2_decap_8 FILLER_1_903 ();
 sg13g2_decap_8 FILLER_1_910 ();
 sg13g2_decap_8 FILLER_1_917 ();
 sg13g2_decap_8 FILLER_1_924 ();
 sg13g2_decap_8 FILLER_1_931 ();
 sg13g2_decap_8 FILLER_1_938 ();
 sg13g2_decap_8 FILLER_1_945 ();
 sg13g2_decap_8 FILLER_1_952 ();
 sg13g2_decap_8 FILLER_1_959 ();
 sg13g2_decap_8 FILLER_1_966 ();
 sg13g2_decap_8 FILLER_1_973 ();
 sg13g2_decap_8 FILLER_1_980 ();
 sg13g2_decap_8 FILLER_1_987 ();
 sg13g2_decap_8 FILLER_1_994 ();
 sg13g2_decap_8 FILLER_1_1001 ();
 sg13g2_decap_8 FILLER_1_1008 ();
 sg13g2_decap_8 FILLER_1_1015 ();
 sg13g2_decap_8 FILLER_1_1022 ();
 sg13g2_fill_1 FILLER_1_1029 ();
 sg13g2_fill_1 FILLER_1_1035 ();
 sg13g2_fill_2 FILLER_1_1040 ();
 sg13g2_fill_2 FILLER_1_1051 ();
 sg13g2_decap_8 FILLER_1_1062 ();
 sg13g2_decap_8 FILLER_1_1069 ();
 sg13g2_decap_4 FILLER_1_1076 ();
 sg13g2_fill_1 FILLER_1_1080 ();
 sg13g2_decap_8 FILLER_1_1089 ();
 sg13g2_decap_4 FILLER_1_1096 ();
 sg13g2_fill_1 FILLER_1_1100 ();
 sg13g2_decap_8 FILLER_1_1105 ();
 sg13g2_decap_8 FILLER_1_1112 ();
 sg13g2_decap_8 FILLER_1_1119 ();
 sg13g2_fill_1 FILLER_1_1126 ();
 sg13g2_decap_8 FILLER_1_1162 ();
 sg13g2_decap_8 FILLER_1_1169 ();
 sg13g2_decap_4 FILLER_1_1176 ();
 sg13g2_fill_1 FILLER_1_1180 ();
 sg13g2_decap_8 FILLER_1_1207 ();
 sg13g2_decap_8 FILLER_1_1214 ();
 sg13g2_decap_8 FILLER_1_1221 ();
 sg13g2_decap_8 FILLER_1_1228 ();
 sg13g2_decap_8 FILLER_1_1235 ();
 sg13g2_decap_8 FILLER_1_1242 ();
 sg13g2_decap_4 FILLER_1_1249 ();
 sg13g2_fill_1 FILLER_1_1253 ();
 sg13g2_fill_2 FILLER_1_1280 ();
 sg13g2_fill_1 FILLER_1_1282 ();
 sg13g2_decap_8 FILLER_1_1448 ();
 sg13g2_decap_8 FILLER_1_1455 ();
 sg13g2_decap_8 FILLER_1_1462 ();
 sg13g2_decap_8 FILLER_1_1469 ();
 sg13g2_decap_8 FILLER_1_1476 ();
 sg13g2_decap_8 FILLER_1_1483 ();
 sg13g2_decap_8 FILLER_1_1490 ();
 sg13g2_decap_8 FILLER_1_1497 ();
 sg13g2_decap_4 FILLER_1_1504 ();
 sg13g2_fill_1 FILLER_1_1508 ();
 sg13g2_fill_2 FILLER_1_1565 ();
 sg13g2_fill_2 FILLER_1_1593 ();
 sg13g2_fill_1 FILLER_1_1647 ();
 sg13g2_decap_8 FILLER_1_1683 ();
 sg13g2_decap_4 FILLER_1_1690 ();
 sg13g2_decap_4 FILLER_1_1720 ();
 sg13g2_fill_1 FILLER_1_1724 ();
 sg13g2_fill_1 FILLER_1_1730 ();
 sg13g2_decap_4 FILLER_1_1783 ();
 sg13g2_decap_4 FILLER_1_1874 ();
 sg13g2_decap_8 FILLER_1_1930 ();
 sg13g2_decap_8 FILLER_1_1937 ();
 sg13g2_fill_1 FILLER_1_1974 ();
 sg13g2_fill_2 FILLER_1_1993 ();
 sg13g2_decap_8 FILLER_1_2047 ();
 sg13g2_decap_4 FILLER_1_2054 ();
 sg13g2_fill_2 FILLER_1_2058 ();
 sg13g2_fill_2 FILLER_1_2077 ();
 sg13g2_fill_1 FILLER_1_2079 ();
 sg13g2_fill_2 FILLER_1_2141 ();
 sg13g2_fill_1 FILLER_1_2143 ();
 sg13g2_fill_2 FILLER_1_2214 ();
 sg13g2_fill_1 FILLER_1_2216 ();
 sg13g2_fill_2 FILLER_1_2247 ();
 sg13g2_fill_1 FILLER_1_2249 ();
 sg13g2_decap_8 FILLER_1_2259 ();
 sg13g2_decap_8 FILLER_1_2266 ();
 sg13g2_decap_8 FILLER_1_2273 ();
 sg13g2_decap_8 FILLER_1_2280 ();
 sg13g2_decap_8 FILLER_1_2287 ();
 sg13g2_decap_8 FILLER_1_2294 ();
 sg13g2_decap_8 FILLER_1_2301 ();
 sg13g2_decap_8 FILLER_1_2308 ();
 sg13g2_decap_8 FILLER_1_2315 ();
 sg13g2_decap_8 FILLER_1_2322 ();
 sg13g2_decap_8 FILLER_1_2329 ();
 sg13g2_decap_8 FILLER_1_2336 ();
 sg13g2_decap_8 FILLER_1_2343 ();
 sg13g2_decap_8 FILLER_1_2350 ();
 sg13g2_decap_8 FILLER_1_2357 ();
 sg13g2_decap_8 FILLER_1_2364 ();
 sg13g2_decap_8 FILLER_1_2371 ();
 sg13g2_decap_8 FILLER_1_2378 ();
 sg13g2_decap_8 FILLER_1_2385 ();
 sg13g2_decap_8 FILLER_1_2392 ();
 sg13g2_decap_8 FILLER_1_2399 ();
 sg13g2_decap_8 FILLER_1_2406 ();
 sg13g2_decap_8 FILLER_1_2413 ();
 sg13g2_decap_8 FILLER_1_2420 ();
 sg13g2_decap_8 FILLER_1_2427 ();
 sg13g2_decap_8 FILLER_1_2434 ();
 sg13g2_decap_8 FILLER_1_2441 ();
 sg13g2_decap_8 FILLER_1_2448 ();
 sg13g2_decap_8 FILLER_1_2455 ();
 sg13g2_decap_8 FILLER_1_2462 ();
 sg13g2_decap_8 FILLER_1_2469 ();
 sg13g2_decap_8 FILLER_1_2476 ();
 sg13g2_decap_8 FILLER_1_2483 ();
 sg13g2_decap_8 FILLER_1_2490 ();
 sg13g2_decap_8 FILLER_1_2497 ();
 sg13g2_decap_8 FILLER_1_2504 ();
 sg13g2_decap_8 FILLER_1_2511 ();
 sg13g2_decap_8 FILLER_1_2518 ();
 sg13g2_decap_8 FILLER_1_2525 ();
 sg13g2_decap_8 FILLER_1_2532 ();
 sg13g2_decap_8 FILLER_1_2539 ();
 sg13g2_decap_8 FILLER_1_2546 ();
 sg13g2_decap_8 FILLER_1_2553 ();
 sg13g2_decap_8 FILLER_1_2560 ();
 sg13g2_decap_8 FILLER_1_2567 ();
 sg13g2_decap_8 FILLER_1_2574 ();
 sg13g2_decap_8 FILLER_1_2581 ();
 sg13g2_decap_8 FILLER_1_2588 ();
 sg13g2_decap_8 FILLER_1_2595 ();
 sg13g2_decap_8 FILLER_1_2602 ();
 sg13g2_decap_8 FILLER_1_2609 ();
 sg13g2_decap_8 FILLER_1_2616 ();
 sg13g2_decap_8 FILLER_1_2623 ();
 sg13g2_decap_8 FILLER_1_2630 ();
 sg13g2_decap_8 FILLER_1_2637 ();
 sg13g2_decap_8 FILLER_1_2644 ();
 sg13g2_decap_8 FILLER_1_2651 ();
 sg13g2_decap_8 FILLER_1_2658 ();
 sg13g2_decap_8 FILLER_1_2665 ();
 sg13g2_fill_2 FILLER_1_2672 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_fill_2 FILLER_2_462 ();
 sg13g2_fill_1 FILLER_2_464 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_501 ();
 sg13g2_fill_2 FILLER_2_552 ();
 sg13g2_fill_2 FILLER_2_614 ();
 sg13g2_fill_1 FILLER_2_616 ();
 sg13g2_fill_2 FILLER_2_664 ();
 sg13g2_decap_4 FILLER_2_679 ();
 sg13g2_fill_1 FILLER_2_683 ();
 sg13g2_fill_1 FILLER_2_697 ();
 sg13g2_fill_1 FILLER_2_774 ();
 sg13g2_fill_2 FILLER_2_788 ();
 sg13g2_fill_2 FILLER_2_799 ();
 sg13g2_fill_1 FILLER_2_801 ();
 sg13g2_decap_8 FILLER_2_806 ();
 sg13g2_decap_4 FILLER_2_813 ();
 sg13g2_fill_2 FILLER_2_817 ();
 sg13g2_decap_4 FILLER_2_845 ();
 sg13g2_fill_1 FILLER_2_849 ();
 sg13g2_decap_4 FILLER_2_858 ();
 sg13g2_fill_2 FILLER_2_867 ();
 sg13g2_decap_8 FILLER_2_873 ();
 sg13g2_decap_8 FILLER_2_880 ();
 sg13g2_decap_8 FILLER_2_887 ();
 sg13g2_decap_8 FILLER_2_894 ();
 sg13g2_decap_8 FILLER_2_901 ();
 sg13g2_decap_8 FILLER_2_908 ();
 sg13g2_decap_8 FILLER_2_915 ();
 sg13g2_decap_8 FILLER_2_922 ();
 sg13g2_decap_8 FILLER_2_929 ();
 sg13g2_decap_8 FILLER_2_936 ();
 sg13g2_decap_8 FILLER_2_943 ();
 sg13g2_decap_8 FILLER_2_950 ();
 sg13g2_decap_8 FILLER_2_957 ();
 sg13g2_decap_8 FILLER_2_964 ();
 sg13g2_decap_8 FILLER_2_971 ();
 sg13g2_decap_8 FILLER_2_978 ();
 sg13g2_decap_8 FILLER_2_985 ();
 sg13g2_decap_8 FILLER_2_992 ();
 sg13g2_decap_8 FILLER_2_999 ();
 sg13g2_decap_8 FILLER_2_1006 ();
 sg13g2_decap_8 FILLER_2_1013 ();
 sg13g2_fill_1 FILLER_2_1020 ();
 sg13g2_fill_2 FILLER_2_1081 ();
 sg13g2_fill_1 FILLER_2_1087 ();
 sg13g2_fill_2 FILLER_2_1102 ();
 sg13g2_fill_1 FILLER_2_1104 ();
 sg13g2_fill_1 FILLER_2_1109 ();
 sg13g2_fill_1 FILLER_2_1136 ();
 sg13g2_fill_2 FILLER_2_1142 ();
 sg13g2_decap_4 FILLER_2_1148 ();
 sg13g2_fill_1 FILLER_2_1152 ();
 sg13g2_fill_1 FILLER_2_1170 ();
 sg13g2_fill_1 FILLER_2_1185 ();
 sg13g2_fill_2 FILLER_2_1221 ();
 sg13g2_fill_1 FILLER_2_1223 ();
 sg13g2_decap_4 FILLER_2_1234 ();
 sg13g2_fill_1 FILLER_2_1238 ();
 sg13g2_fill_2 FILLER_2_1274 ();
 sg13g2_fill_1 FILLER_2_1276 ();
 sg13g2_fill_1 FILLER_2_1286 ();
 sg13g2_fill_1 FILLER_2_1321 ();
 sg13g2_fill_2 FILLER_2_1331 ();
 sg13g2_fill_1 FILLER_2_1333 ();
 sg13g2_decap_4 FILLER_2_1360 ();
 sg13g2_fill_1 FILLER_2_1368 ();
 sg13g2_decap_4 FILLER_2_1373 ();
 sg13g2_fill_1 FILLER_2_1377 ();
 sg13g2_fill_2 FILLER_2_1392 ();
 sg13g2_fill_1 FILLER_2_1394 ();
 sg13g2_fill_2 FILLER_2_1413 ();
 sg13g2_fill_1 FILLER_2_1424 ();
 sg13g2_decap_8 FILLER_2_1460 ();
 sg13g2_decap_8 FILLER_2_1467 ();
 sg13g2_decap_8 FILLER_2_1474 ();
 sg13g2_decap_8 FILLER_2_1481 ();
 sg13g2_fill_1 FILLER_2_1488 ();
 sg13g2_decap_4 FILLER_2_1498 ();
 sg13g2_fill_2 FILLER_2_1502 ();
 sg13g2_decap_8 FILLER_2_1513 ();
 sg13g2_fill_2 FILLER_2_1524 ();
 sg13g2_fill_1 FILLER_2_1526 ();
 sg13g2_fill_2 FILLER_2_1552 ();
 sg13g2_fill_1 FILLER_2_1554 ();
 sg13g2_fill_1 FILLER_2_1581 ();
 sg13g2_decap_4 FILLER_2_1626 ();
 sg13g2_fill_1 FILLER_2_1630 ();
 sg13g2_fill_2 FILLER_2_1649 ();
 sg13g2_fill_1 FILLER_2_1651 ();
 sg13g2_fill_2 FILLER_2_1657 ();
 sg13g2_fill_1 FILLER_2_1659 ();
 sg13g2_fill_2 FILLER_2_1701 ();
 sg13g2_decap_8 FILLER_2_1712 ();
 sg13g2_decap_8 FILLER_2_1719 ();
 sg13g2_decap_4 FILLER_2_1726 ();
 sg13g2_fill_2 FILLER_2_1734 ();
 sg13g2_fill_1 FILLER_2_1788 ();
 sg13g2_fill_2 FILLER_2_1802 ();
 sg13g2_fill_1 FILLER_2_1804 ();
 sg13g2_fill_1 FILLER_2_1827 ();
 sg13g2_fill_2 FILLER_2_1841 ();
 sg13g2_fill_1 FILLER_2_1843 ();
 sg13g2_fill_2 FILLER_2_1853 ();
 sg13g2_fill_1 FILLER_2_1855 ();
 sg13g2_fill_1 FILLER_2_1865 ();
 sg13g2_fill_1 FILLER_2_1870 ();
 sg13g2_fill_2 FILLER_2_1880 ();
 sg13g2_fill_1 FILLER_2_1882 ();
 sg13g2_fill_2 FILLER_2_1888 ();
 sg13g2_decap_4 FILLER_2_1894 ();
 sg13g2_fill_2 FILLER_2_1898 ();
 sg13g2_decap_4 FILLER_2_1925 ();
 sg13g2_fill_1 FILLER_2_1960 ();
 sg13g2_fill_1 FILLER_2_1970 ();
 sg13g2_fill_2 FILLER_2_2011 ();
 sg13g2_fill_1 FILLER_2_2013 ();
 sg13g2_fill_2 FILLER_2_2089 ();
 sg13g2_fill_2 FILLER_2_2165 ();
 sg13g2_fill_1 FILLER_2_2172 ();
 sg13g2_fill_2 FILLER_2_2177 ();
 sg13g2_fill_1 FILLER_2_2179 ();
 sg13g2_fill_1 FILLER_2_2214 ();
 sg13g2_decap_8 FILLER_2_2278 ();
 sg13g2_decap_8 FILLER_2_2285 ();
 sg13g2_decap_8 FILLER_2_2292 ();
 sg13g2_decap_8 FILLER_2_2299 ();
 sg13g2_decap_8 FILLER_2_2306 ();
 sg13g2_decap_8 FILLER_2_2313 ();
 sg13g2_decap_8 FILLER_2_2320 ();
 sg13g2_decap_8 FILLER_2_2327 ();
 sg13g2_decap_8 FILLER_2_2334 ();
 sg13g2_decap_8 FILLER_2_2341 ();
 sg13g2_decap_8 FILLER_2_2348 ();
 sg13g2_decap_8 FILLER_2_2355 ();
 sg13g2_decap_8 FILLER_2_2362 ();
 sg13g2_decap_8 FILLER_2_2369 ();
 sg13g2_decap_8 FILLER_2_2376 ();
 sg13g2_decap_8 FILLER_2_2383 ();
 sg13g2_decap_8 FILLER_2_2390 ();
 sg13g2_decap_8 FILLER_2_2397 ();
 sg13g2_decap_8 FILLER_2_2404 ();
 sg13g2_decap_8 FILLER_2_2411 ();
 sg13g2_decap_8 FILLER_2_2418 ();
 sg13g2_decap_8 FILLER_2_2425 ();
 sg13g2_decap_8 FILLER_2_2432 ();
 sg13g2_decap_8 FILLER_2_2439 ();
 sg13g2_decap_8 FILLER_2_2446 ();
 sg13g2_decap_8 FILLER_2_2453 ();
 sg13g2_decap_8 FILLER_2_2460 ();
 sg13g2_decap_8 FILLER_2_2467 ();
 sg13g2_decap_8 FILLER_2_2474 ();
 sg13g2_decap_8 FILLER_2_2481 ();
 sg13g2_decap_8 FILLER_2_2488 ();
 sg13g2_decap_8 FILLER_2_2495 ();
 sg13g2_decap_8 FILLER_2_2502 ();
 sg13g2_decap_8 FILLER_2_2509 ();
 sg13g2_decap_8 FILLER_2_2516 ();
 sg13g2_decap_8 FILLER_2_2523 ();
 sg13g2_decap_8 FILLER_2_2530 ();
 sg13g2_decap_8 FILLER_2_2537 ();
 sg13g2_decap_8 FILLER_2_2544 ();
 sg13g2_decap_8 FILLER_2_2551 ();
 sg13g2_decap_8 FILLER_2_2558 ();
 sg13g2_decap_8 FILLER_2_2565 ();
 sg13g2_decap_8 FILLER_2_2572 ();
 sg13g2_decap_8 FILLER_2_2579 ();
 sg13g2_decap_8 FILLER_2_2586 ();
 sg13g2_decap_8 FILLER_2_2593 ();
 sg13g2_decap_8 FILLER_2_2600 ();
 sg13g2_decap_8 FILLER_2_2607 ();
 sg13g2_decap_8 FILLER_2_2614 ();
 sg13g2_decap_8 FILLER_2_2621 ();
 sg13g2_decap_8 FILLER_2_2628 ();
 sg13g2_decap_8 FILLER_2_2635 ();
 sg13g2_decap_8 FILLER_2_2642 ();
 sg13g2_decap_8 FILLER_2_2649 ();
 sg13g2_decap_8 FILLER_2_2656 ();
 sg13g2_decap_8 FILLER_2_2663 ();
 sg13g2_decap_4 FILLER_2_2670 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_fill_2 FILLER_3_455 ();
 sg13g2_fill_1 FILLER_3_457 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_4 FILLER_3_483 ();
 sg13g2_fill_1 FILLER_3_487 ();
 sg13g2_decap_4 FILLER_3_519 ();
 sg13g2_fill_2 FILLER_3_523 ();
 sg13g2_fill_2 FILLER_3_534 ();
 sg13g2_fill_1 FILLER_3_536 ();
 sg13g2_fill_1 FILLER_3_567 ();
 sg13g2_fill_1 FILLER_3_600 ();
 sg13g2_fill_1 FILLER_3_630 ();
 sg13g2_fill_1 FILLER_3_640 ();
 sg13g2_fill_2 FILLER_3_650 ();
 sg13g2_fill_1 FILLER_3_652 ();
 sg13g2_decap_4 FILLER_3_688 ();
 sg13g2_fill_1 FILLER_3_692 ();
 sg13g2_fill_2 FILLER_3_738 ();
 sg13g2_fill_1 FILLER_3_770 ();
 sg13g2_fill_1 FILLER_3_802 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_fill_2 FILLER_3_826 ();
 sg13g2_fill_1 FILLER_3_828 ();
 sg13g2_fill_2 FILLER_3_833 ();
 sg13g2_fill_1 FILLER_3_835 ();
 sg13g2_decap_8 FILLER_3_888 ();
 sg13g2_fill_1 FILLER_3_895 ();
 sg13g2_decap_8 FILLER_3_900 ();
 sg13g2_decap_8 FILLER_3_907 ();
 sg13g2_decap_8 FILLER_3_914 ();
 sg13g2_decap_8 FILLER_3_921 ();
 sg13g2_decap_8 FILLER_3_928 ();
 sg13g2_decap_8 FILLER_3_935 ();
 sg13g2_decap_8 FILLER_3_942 ();
 sg13g2_decap_8 FILLER_3_949 ();
 sg13g2_decap_8 FILLER_3_956 ();
 sg13g2_decap_8 FILLER_3_963 ();
 sg13g2_decap_8 FILLER_3_970 ();
 sg13g2_decap_8 FILLER_3_977 ();
 sg13g2_decap_8 FILLER_3_984 ();
 sg13g2_decap_8 FILLER_3_991 ();
 sg13g2_decap_8 FILLER_3_998 ();
 sg13g2_decap_8 FILLER_3_1005 ();
 sg13g2_fill_2 FILLER_3_1017 ();
 sg13g2_fill_1 FILLER_3_1019 ();
 sg13g2_decap_8 FILLER_3_1024 ();
 sg13g2_fill_2 FILLER_3_1031 ();
 sg13g2_fill_2 FILLER_3_1037 ();
 sg13g2_fill_1 FILLER_3_1039 ();
 sg13g2_decap_4 FILLER_3_1045 ();
 sg13g2_fill_2 FILLER_3_1049 ();
 sg13g2_fill_2 FILLER_3_1130 ();
 sg13g2_fill_1 FILLER_3_1141 ();
 sg13g2_fill_2 FILLER_3_1194 ();
 sg13g2_decap_8 FILLER_3_1243 ();
 sg13g2_fill_2 FILLER_3_1272 ();
 sg13g2_fill_1 FILLER_3_1274 ();
 sg13g2_decap_4 FILLER_3_1340 ();
 sg13g2_decap_8 FILLER_3_1348 ();
 sg13g2_decap_4 FILLER_3_1355 ();
 sg13g2_fill_1 FILLER_3_1359 ();
 sg13g2_fill_1 FILLER_3_1391 ();
 sg13g2_fill_2 FILLER_3_1396 ();
 sg13g2_fill_1 FILLER_3_1398 ();
 sg13g2_fill_2 FILLER_3_1433 ();
 sg13g2_fill_1 FILLER_3_1435 ();
 sg13g2_fill_2 FILLER_3_1466 ();
 sg13g2_decap_8 FILLER_3_1542 ();
 sg13g2_decap_4 FILLER_3_1549 ();
 sg13g2_fill_2 FILLER_3_1563 ();
 sg13g2_decap_8 FILLER_3_1600 ();
 sg13g2_fill_2 FILLER_3_1633 ();
 sg13g2_fill_2 FILLER_3_1686 ();
 sg13g2_fill_2 FILLER_3_1723 ();
 sg13g2_fill_2 FILLER_3_1751 ();
 sg13g2_decap_8 FILLER_3_1771 ();
 sg13g2_fill_1 FILLER_3_1936 ();
 sg13g2_fill_2 FILLER_3_1954 ();
 sg13g2_fill_2 FILLER_3_1964 ();
 sg13g2_fill_1 FILLER_3_1980 ();
 sg13g2_fill_1 FILLER_3_1993 ();
 sg13g2_decap_8 FILLER_3_2054 ();
 sg13g2_fill_2 FILLER_3_2061 ();
 sg13g2_fill_1 FILLER_3_2063 ();
 sg13g2_decap_4 FILLER_3_2068 ();
 sg13g2_fill_2 FILLER_3_2072 ();
 sg13g2_fill_2 FILLER_3_2096 ();
 sg13g2_fill_2 FILLER_3_2103 ();
 sg13g2_fill_2 FILLER_3_2141 ();
 sg13g2_fill_2 FILLER_3_2169 ();
 sg13g2_fill_2 FILLER_3_2176 ();
 sg13g2_fill_1 FILLER_3_2182 ();
 sg13g2_decap_8 FILLER_3_2274 ();
 sg13g2_decap_8 FILLER_3_2281 ();
 sg13g2_decap_8 FILLER_3_2288 ();
 sg13g2_decap_8 FILLER_3_2295 ();
 sg13g2_decap_8 FILLER_3_2302 ();
 sg13g2_decap_8 FILLER_3_2309 ();
 sg13g2_decap_8 FILLER_3_2316 ();
 sg13g2_decap_8 FILLER_3_2323 ();
 sg13g2_decap_8 FILLER_3_2330 ();
 sg13g2_decap_8 FILLER_3_2337 ();
 sg13g2_decap_8 FILLER_3_2344 ();
 sg13g2_decap_8 FILLER_3_2351 ();
 sg13g2_decap_8 FILLER_3_2358 ();
 sg13g2_decap_8 FILLER_3_2365 ();
 sg13g2_decap_8 FILLER_3_2372 ();
 sg13g2_decap_8 FILLER_3_2379 ();
 sg13g2_decap_8 FILLER_3_2386 ();
 sg13g2_decap_8 FILLER_3_2393 ();
 sg13g2_decap_8 FILLER_3_2400 ();
 sg13g2_decap_8 FILLER_3_2407 ();
 sg13g2_decap_8 FILLER_3_2414 ();
 sg13g2_decap_8 FILLER_3_2421 ();
 sg13g2_decap_8 FILLER_3_2428 ();
 sg13g2_decap_8 FILLER_3_2435 ();
 sg13g2_decap_8 FILLER_3_2442 ();
 sg13g2_decap_8 FILLER_3_2449 ();
 sg13g2_decap_8 FILLER_3_2456 ();
 sg13g2_decap_8 FILLER_3_2463 ();
 sg13g2_decap_8 FILLER_3_2470 ();
 sg13g2_decap_8 FILLER_3_2477 ();
 sg13g2_decap_8 FILLER_3_2484 ();
 sg13g2_decap_8 FILLER_3_2491 ();
 sg13g2_decap_8 FILLER_3_2498 ();
 sg13g2_decap_8 FILLER_3_2505 ();
 sg13g2_decap_8 FILLER_3_2512 ();
 sg13g2_decap_8 FILLER_3_2519 ();
 sg13g2_decap_8 FILLER_3_2526 ();
 sg13g2_decap_8 FILLER_3_2533 ();
 sg13g2_decap_8 FILLER_3_2540 ();
 sg13g2_decap_8 FILLER_3_2547 ();
 sg13g2_decap_8 FILLER_3_2554 ();
 sg13g2_decap_8 FILLER_3_2561 ();
 sg13g2_decap_8 FILLER_3_2568 ();
 sg13g2_decap_8 FILLER_3_2575 ();
 sg13g2_decap_8 FILLER_3_2582 ();
 sg13g2_decap_8 FILLER_3_2589 ();
 sg13g2_decap_8 FILLER_3_2596 ();
 sg13g2_decap_8 FILLER_3_2603 ();
 sg13g2_decap_8 FILLER_3_2610 ();
 sg13g2_decap_8 FILLER_3_2617 ();
 sg13g2_decap_8 FILLER_3_2624 ();
 sg13g2_decap_8 FILLER_3_2631 ();
 sg13g2_decap_8 FILLER_3_2638 ();
 sg13g2_decap_8 FILLER_3_2645 ();
 sg13g2_decap_8 FILLER_3_2652 ();
 sg13g2_decap_8 FILLER_3_2659 ();
 sg13g2_decap_8 FILLER_3_2666 ();
 sg13g2_fill_1 FILLER_3_2673 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_4 FILLER_4_441 ();
 sg13g2_fill_2 FILLER_4_445 ();
 sg13g2_decap_4 FILLER_4_499 ();
 sg13g2_fill_2 FILLER_4_507 ();
 sg13g2_fill_2 FILLER_4_549 ();
 sg13g2_fill_1 FILLER_4_556 ();
 sg13g2_fill_1 FILLER_4_562 ();
 sg13g2_fill_2 FILLER_4_572 ();
 sg13g2_fill_1 FILLER_4_656 ();
 sg13g2_fill_2 FILLER_4_684 ();
 sg13g2_fill_1 FILLER_4_695 ();
 sg13g2_decap_8 FILLER_4_713 ();
 sg13g2_fill_1 FILLER_4_760 ();
 sg13g2_fill_2 FILLER_4_827 ();
 sg13g2_fill_1 FILLER_4_834 ();
 sg13g2_fill_2 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_856 ();
 sg13g2_fill_1 FILLER_4_871 ();
 sg13g2_decap_8 FILLER_4_911 ();
 sg13g2_fill_1 FILLER_4_918 ();
 sg13g2_decap_8 FILLER_4_923 ();
 sg13g2_decap_4 FILLER_4_930 ();
 sg13g2_decap_8 FILLER_4_960 ();
 sg13g2_decap_8 FILLER_4_967 ();
 sg13g2_fill_2 FILLER_4_974 ();
 sg13g2_decap_8 FILLER_4_980 ();
 sg13g2_fill_1 FILLER_4_987 ();
 sg13g2_decap_4 FILLER_4_997 ();
 sg13g2_fill_1 FILLER_4_1001 ();
 sg13g2_fill_2 FILLER_4_1075 ();
 sg13g2_fill_1 FILLER_4_1077 ();
 sg13g2_fill_2 FILLER_4_1182 ();
 sg13g2_fill_1 FILLER_4_1193 ();
 sg13g2_fill_1 FILLER_4_1220 ();
 sg13g2_fill_2 FILLER_4_1291 ();
 sg13g2_decap_4 FILLER_4_1407 ();
 sg13g2_fill_1 FILLER_4_1411 ();
 sg13g2_fill_2 FILLER_4_1456 ();
 sg13g2_fill_1 FILLER_4_1458 ();
 sg13g2_fill_2 FILLER_4_1485 ();
 sg13g2_fill_2 FILLER_4_1501 ();
 sg13g2_fill_1 FILLER_4_1503 ();
 sg13g2_fill_2 FILLER_4_1508 ();
 sg13g2_fill_1 FILLER_4_1510 ();
 sg13g2_fill_1 FILLER_4_1515 ();
 sg13g2_decap_8 FILLER_4_1569 ();
 sg13g2_decap_4 FILLER_4_1593 ();
 sg13g2_fill_1 FILLER_4_1597 ();
 sg13g2_fill_1 FILLER_4_1632 ();
 sg13g2_fill_2 FILLER_4_1694 ();
 sg13g2_fill_2 FILLER_4_1749 ();
 sg13g2_fill_2 FILLER_4_1833 ();
 sg13g2_fill_1 FILLER_4_1835 ();
 sg13g2_decap_4 FILLER_4_1891 ();
 sg13g2_fill_2 FILLER_4_1895 ();
 sg13g2_fill_1 FILLER_4_1910 ();
 sg13g2_fill_2 FILLER_4_1928 ();
 sg13g2_decap_8 FILLER_4_1996 ();
 sg13g2_decap_4 FILLER_4_2003 ();
 sg13g2_fill_2 FILLER_4_2097 ();
 sg13g2_fill_2 FILLER_4_2160 ();
 sg13g2_fill_2 FILLER_4_2206 ();
 sg13g2_fill_1 FILLER_4_2208 ();
 sg13g2_decap_8 FILLER_4_2218 ();
 sg13g2_fill_2 FILLER_4_2225 ();
 sg13g2_fill_2 FILLER_4_2231 ();
 sg13g2_fill_1 FILLER_4_2233 ();
 sg13g2_decap_8 FILLER_4_2278 ();
 sg13g2_decap_8 FILLER_4_2285 ();
 sg13g2_decap_8 FILLER_4_2292 ();
 sg13g2_fill_1 FILLER_4_2299 ();
 sg13g2_decap_8 FILLER_4_2305 ();
 sg13g2_decap_8 FILLER_4_2312 ();
 sg13g2_decap_8 FILLER_4_2319 ();
 sg13g2_decap_8 FILLER_4_2326 ();
 sg13g2_decap_8 FILLER_4_2333 ();
 sg13g2_decap_8 FILLER_4_2340 ();
 sg13g2_decap_8 FILLER_4_2347 ();
 sg13g2_decap_8 FILLER_4_2354 ();
 sg13g2_decap_8 FILLER_4_2361 ();
 sg13g2_decap_8 FILLER_4_2368 ();
 sg13g2_decap_8 FILLER_4_2375 ();
 sg13g2_decap_8 FILLER_4_2382 ();
 sg13g2_decap_8 FILLER_4_2389 ();
 sg13g2_decap_8 FILLER_4_2396 ();
 sg13g2_decap_8 FILLER_4_2403 ();
 sg13g2_decap_8 FILLER_4_2410 ();
 sg13g2_decap_8 FILLER_4_2417 ();
 sg13g2_decap_8 FILLER_4_2424 ();
 sg13g2_decap_8 FILLER_4_2431 ();
 sg13g2_decap_8 FILLER_4_2438 ();
 sg13g2_decap_8 FILLER_4_2445 ();
 sg13g2_decap_8 FILLER_4_2452 ();
 sg13g2_decap_8 FILLER_4_2459 ();
 sg13g2_decap_8 FILLER_4_2466 ();
 sg13g2_decap_8 FILLER_4_2473 ();
 sg13g2_decap_8 FILLER_4_2480 ();
 sg13g2_decap_8 FILLER_4_2487 ();
 sg13g2_decap_8 FILLER_4_2494 ();
 sg13g2_decap_8 FILLER_4_2501 ();
 sg13g2_decap_8 FILLER_4_2508 ();
 sg13g2_decap_8 FILLER_4_2515 ();
 sg13g2_decap_8 FILLER_4_2522 ();
 sg13g2_decap_8 FILLER_4_2529 ();
 sg13g2_decap_8 FILLER_4_2536 ();
 sg13g2_decap_8 FILLER_4_2543 ();
 sg13g2_decap_8 FILLER_4_2550 ();
 sg13g2_decap_8 FILLER_4_2557 ();
 sg13g2_decap_8 FILLER_4_2564 ();
 sg13g2_decap_8 FILLER_4_2571 ();
 sg13g2_decap_8 FILLER_4_2578 ();
 sg13g2_decap_8 FILLER_4_2585 ();
 sg13g2_decap_8 FILLER_4_2592 ();
 sg13g2_decap_8 FILLER_4_2599 ();
 sg13g2_decap_8 FILLER_4_2606 ();
 sg13g2_decap_8 FILLER_4_2613 ();
 sg13g2_decap_8 FILLER_4_2620 ();
 sg13g2_decap_8 FILLER_4_2627 ();
 sg13g2_decap_8 FILLER_4_2634 ();
 sg13g2_decap_8 FILLER_4_2641 ();
 sg13g2_decap_8 FILLER_4_2648 ();
 sg13g2_decap_8 FILLER_4_2655 ();
 sg13g2_decap_8 FILLER_4_2662 ();
 sg13g2_decap_4 FILLER_4_2669 ();
 sg13g2_fill_1 FILLER_4_2673 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_fill_1 FILLER_5_441 ();
 sg13g2_fill_1 FILLER_5_464 ();
 sg13g2_fill_1 FILLER_5_494 ();
 sg13g2_fill_2 FILLER_5_521 ();
 sg13g2_fill_1 FILLER_5_549 ();
 sg13g2_fill_2 FILLER_5_584 ();
 sg13g2_fill_1 FILLER_5_586 ();
 sg13g2_decap_4 FILLER_5_618 ();
 sg13g2_fill_1 FILLER_5_622 ();
 sg13g2_fill_2 FILLER_5_628 ();
 sg13g2_fill_1 FILLER_5_630 ();
 sg13g2_decap_4 FILLER_5_636 ();
 sg13g2_fill_1 FILLER_5_640 ();
 sg13g2_fill_2 FILLER_5_649 ();
 sg13g2_fill_1 FILLER_5_677 ();
 sg13g2_fill_1 FILLER_5_713 ();
 sg13g2_decap_4 FILLER_5_731 ();
 sg13g2_fill_2 FILLER_5_739 ();
 sg13g2_fill_1 FILLER_5_741 ();
 sg13g2_fill_2 FILLER_5_783 ();
 sg13g2_fill_2 FILLER_5_809 ();
 sg13g2_fill_1 FILLER_5_811 ();
 sg13g2_decap_8 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_823 ();
 sg13g2_fill_2 FILLER_5_838 ();
 sg13g2_fill_2 FILLER_5_878 ();
 sg13g2_fill_1 FILLER_5_885 ();
 sg13g2_fill_1 FILLER_5_944 ();
 sg13g2_fill_2 FILLER_5_953 ();
 sg13g2_decap_8 FILLER_5_1004 ();
 sg13g2_fill_2 FILLER_5_1011 ();
 sg13g2_fill_2 FILLER_5_1035 ();
 sg13g2_fill_1 FILLER_5_1037 ();
 sg13g2_fill_2 FILLER_5_1064 ();
 sg13g2_fill_1 FILLER_5_1066 ();
 sg13g2_decap_8 FILLER_5_1103 ();
 sg13g2_fill_2 FILLER_5_1110 ();
 sg13g2_fill_1 FILLER_5_1112 ();
 sg13g2_fill_2 FILLER_5_1152 ();
 sg13g2_fill_1 FILLER_5_1154 ();
 sg13g2_fill_2 FILLER_5_1207 ();
 sg13g2_fill_1 FILLER_5_1214 ();
 sg13g2_decap_8 FILLER_5_1237 ();
 sg13g2_decap_4 FILLER_5_1244 ();
 sg13g2_fill_2 FILLER_5_1262 ();
 sg13g2_fill_2 FILLER_5_1286 ();
 sg13g2_fill_1 FILLER_5_1296 ();
 sg13g2_fill_1 FILLER_5_1315 ();
 sg13g2_fill_2 FILLER_5_1326 ();
 sg13g2_fill_1 FILLER_5_1328 ();
 sg13g2_fill_2 FILLER_5_1347 ();
 sg13g2_fill_1 FILLER_5_1349 ();
 sg13g2_fill_2 FILLER_5_1384 ();
 sg13g2_fill_1 FILLER_5_1386 ();
 sg13g2_fill_2 FILLER_5_1452 ();
 sg13g2_fill_1 FILLER_5_1454 ();
 sg13g2_fill_2 FILLER_5_1464 ();
 sg13g2_fill_1 FILLER_5_1466 ();
 sg13g2_fill_2 FILLER_5_1493 ();
 sg13g2_fill_2 FILLER_5_1535 ();
 sg13g2_fill_2 FILLER_5_1547 ();
 sg13g2_fill_1 FILLER_5_1549 ();
 sg13g2_fill_2 FILLER_5_1554 ();
 sg13g2_fill_2 FILLER_5_1561 ();
 sg13g2_fill_1 FILLER_5_1563 ();
 sg13g2_fill_1 FILLER_5_1582 ();
 sg13g2_fill_2 FILLER_5_1618 ();
 sg13g2_fill_1 FILLER_5_1620 ();
 sg13g2_fill_2 FILLER_5_1644 ();
 sg13g2_fill_2 FILLER_5_1676 ();
 sg13g2_fill_1 FILLER_5_1678 ();
 sg13g2_decap_8 FILLER_5_1683 ();
 sg13g2_fill_2 FILLER_5_1690 ();
 sg13g2_fill_2 FILLER_5_1701 ();
 sg13g2_fill_1 FILLER_5_1703 ();
 sg13g2_fill_1 FILLER_5_1708 ();
 sg13g2_fill_1 FILLER_5_1718 ();
 sg13g2_fill_2 FILLER_5_1723 ();
 sg13g2_fill_1 FILLER_5_1725 ();
 sg13g2_decap_4 FILLER_5_1760 ();
 sg13g2_fill_1 FILLER_5_1764 ();
 sg13g2_fill_2 FILLER_5_1774 ();
 sg13g2_fill_1 FILLER_5_1776 ();
 sg13g2_fill_2 FILLER_5_1785 ();
 sg13g2_fill_2 FILLER_5_1806 ();
 sg13g2_fill_2 FILLER_5_1847 ();
 sg13g2_fill_2 FILLER_5_1854 ();
 sg13g2_fill_2 FILLER_5_1861 ();
 sg13g2_fill_1 FILLER_5_1863 ();
 sg13g2_decap_4 FILLER_5_1877 ();
 sg13g2_fill_2 FILLER_5_1881 ();
 sg13g2_fill_2 FILLER_5_1949 ();
 sg13g2_fill_1 FILLER_5_1951 ();
 sg13g2_fill_2 FILLER_5_2004 ();
 sg13g2_fill_2 FILLER_5_2037 ();
 sg13g2_fill_1 FILLER_5_2039 ();
 sg13g2_decap_8 FILLER_5_2062 ();
 sg13g2_fill_1 FILLER_5_2069 ();
 sg13g2_decap_4 FILLER_5_2074 ();
 sg13g2_fill_2 FILLER_5_2088 ();
 sg13g2_fill_2 FILLER_5_2130 ();
 sg13g2_fill_1 FILLER_5_2132 ();
 sg13g2_decap_8 FILLER_5_2180 ();
 sg13g2_fill_2 FILLER_5_2187 ();
 sg13g2_fill_1 FILLER_5_2189 ();
 sg13g2_fill_2 FILLER_5_2206 ();
 sg13g2_fill_2 FILLER_5_2216 ();
 sg13g2_decap_4 FILLER_5_2231 ();
 sg13g2_fill_2 FILLER_5_2235 ();
 sg13g2_decap_4 FILLER_5_2246 ();
 sg13g2_fill_1 FILLER_5_2250 ();
 sg13g2_fill_2 FILLER_5_2268 ();
 sg13g2_fill_1 FILLER_5_2270 ();
 sg13g2_decap_8 FILLER_5_2284 ();
 sg13g2_decap_8 FILLER_5_2321 ();
 sg13g2_decap_8 FILLER_5_2328 ();
 sg13g2_decap_8 FILLER_5_2335 ();
 sg13g2_decap_8 FILLER_5_2342 ();
 sg13g2_decap_8 FILLER_5_2349 ();
 sg13g2_decap_8 FILLER_5_2356 ();
 sg13g2_decap_8 FILLER_5_2363 ();
 sg13g2_decap_8 FILLER_5_2370 ();
 sg13g2_decap_8 FILLER_5_2377 ();
 sg13g2_decap_8 FILLER_5_2384 ();
 sg13g2_decap_8 FILLER_5_2391 ();
 sg13g2_decap_8 FILLER_5_2398 ();
 sg13g2_decap_8 FILLER_5_2405 ();
 sg13g2_decap_8 FILLER_5_2412 ();
 sg13g2_decap_8 FILLER_5_2419 ();
 sg13g2_decap_8 FILLER_5_2426 ();
 sg13g2_decap_8 FILLER_5_2433 ();
 sg13g2_decap_8 FILLER_5_2440 ();
 sg13g2_decap_8 FILLER_5_2447 ();
 sg13g2_decap_8 FILLER_5_2454 ();
 sg13g2_decap_8 FILLER_5_2461 ();
 sg13g2_decap_8 FILLER_5_2468 ();
 sg13g2_decap_8 FILLER_5_2475 ();
 sg13g2_decap_8 FILLER_5_2482 ();
 sg13g2_decap_8 FILLER_5_2489 ();
 sg13g2_decap_8 FILLER_5_2496 ();
 sg13g2_decap_8 FILLER_5_2503 ();
 sg13g2_decap_8 FILLER_5_2510 ();
 sg13g2_decap_8 FILLER_5_2517 ();
 sg13g2_decap_8 FILLER_5_2524 ();
 sg13g2_decap_8 FILLER_5_2531 ();
 sg13g2_decap_8 FILLER_5_2538 ();
 sg13g2_decap_8 FILLER_5_2545 ();
 sg13g2_decap_8 FILLER_5_2552 ();
 sg13g2_decap_8 FILLER_5_2559 ();
 sg13g2_decap_8 FILLER_5_2566 ();
 sg13g2_decap_8 FILLER_5_2573 ();
 sg13g2_decap_8 FILLER_5_2580 ();
 sg13g2_decap_8 FILLER_5_2587 ();
 sg13g2_decap_8 FILLER_5_2594 ();
 sg13g2_decap_8 FILLER_5_2601 ();
 sg13g2_decap_8 FILLER_5_2608 ();
 sg13g2_decap_8 FILLER_5_2615 ();
 sg13g2_decap_8 FILLER_5_2622 ();
 sg13g2_decap_8 FILLER_5_2629 ();
 sg13g2_decap_8 FILLER_5_2636 ();
 sg13g2_decap_8 FILLER_5_2643 ();
 sg13g2_decap_8 FILLER_5_2650 ();
 sg13g2_decap_8 FILLER_5_2657 ();
 sg13g2_decap_8 FILLER_5_2664 ();
 sg13g2_fill_2 FILLER_5_2671 ();
 sg13g2_fill_1 FILLER_5_2673 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_fill_2 FILLER_6_467 ();
 sg13g2_fill_1 FILLER_6_469 ();
 sg13g2_fill_1 FILLER_6_491 ();
 sg13g2_fill_1 FILLER_6_501 ();
 sg13g2_decap_4 FILLER_6_546 ();
 sg13g2_fill_1 FILLER_6_575 ();
 sg13g2_decap_4 FILLER_6_658 ();
 sg13g2_fill_2 FILLER_6_667 ();
 sg13g2_fill_1 FILLER_6_679 ();
 sg13g2_fill_1 FILLER_6_684 ();
 sg13g2_fill_2 FILLER_6_729 ();
 sg13g2_decap_4 FILLER_6_744 ();
 sg13g2_fill_1 FILLER_6_748 ();
 sg13g2_fill_1 FILLER_6_754 ();
 sg13g2_fill_2 FILLER_6_786 ();
 sg13g2_fill_1 FILLER_6_788 ();
 sg13g2_fill_2 FILLER_6_910 ();
 sg13g2_fill_1 FILLER_6_912 ();
 sg13g2_fill_2 FILLER_6_963 ();
 sg13g2_fill_1 FILLER_6_965 ();
 sg13g2_fill_2 FILLER_6_979 ();
 sg13g2_fill_1 FILLER_6_981 ();
 sg13g2_fill_2 FILLER_6_1000 ();
 sg13g2_decap_4 FILLER_6_1046 ();
 sg13g2_fill_2 FILLER_6_1050 ();
 sg13g2_fill_2 FILLER_6_1086 ();
 sg13g2_decap_4 FILLER_6_1101 ();
 sg13g2_fill_1 FILLER_6_1123 ();
 sg13g2_fill_2 FILLER_6_1128 ();
 sg13g2_fill_1 FILLER_6_1130 ();
 sg13g2_fill_1 FILLER_6_1167 ();
 sg13g2_fill_2 FILLER_6_1275 ();
 sg13g2_fill_1 FILLER_6_1303 ();
 sg13g2_fill_1 FILLER_6_1330 ();
 sg13g2_fill_2 FILLER_6_1357 ();
 sg13g2_fill_1 FILLER_6_1359 ();
 sg13g2_fill_2 FILLER_6_1391 ();
 sg13g2_fill_1 FILLER_6_1393 ();
 sg13g2_decap_4 FILLER_6_1408 ();
 sg13g2_fill_1 FILLER_6_1412 ();
 sg13g2_decap_4 FILLER_6_1431 ();
 sg13g2_fill_1 FILLER_6_1435 ();
 sg13g2_fill_2 FILLER_6_1467 ();
 sg13g2_fill_2 FILLER_6_1474 ();
 sg13g2_decap_8 FILLER_6_1506 ();
 sg13g2_fill_2 FILLER_6_1560 ();
 sg13g2_fill_1 FILLER_6_1562 ();
 sg13g2_fill_2 FILLER_6_1603 ();
 sg13g2_fill_1 FILLER_6_1631 ();
 sg13g2_decap_4 FILLER_6_1680 ();
 sg13g2_fill_2 FILLER_6_1684 ();
 sg13g2_fill_2 FILLER_6_1738 ();
 sg13g2_fill_2 FILLER_6_1792 ();
 sg13g2_fill_1 FILLER_6_1794 ();
 sg13g2_fill_2 FILLER_6_1835 ();
 sg13g2_fill_2 FILLER_6_1851 ();
 sg13g2_fill_1 FILLER_6_1853 ();
 sg13g2_fill_2 FILLER_6_1889 ();
 sg13g2_fill_2 FILLER_6_1918 ();
 sg13g2_fill_1 FILLER_6_1920 ();
 sg13g2_fill_2 FILLER_6_1965 ();
 sg13g2_fill_2 FILLER_6_1993 ();
 sg13g2_fill_2 FILLER_6_2026 ();
 sg13g2_fill_1 FILLER_6_2028 ();
 sg13g2_decap_8 FILLER_6_2056 ();
 sg13g2_decap_8 FILLER_6_2063 ();
 sg13g2_fill_2 FILLER_6_2070 ();
 sg13g2_fill_2 FILLER_6_2076 ();
 sg13g2_fill_1 FILLER_6_2078 ();
 sg13g2_fill_2 FILLER_6_2092 ();
 sg13g2_fill_2 FILLER_6_2188 ();
 sg13g2_fill_1 FILLER_6_2190 ();
 sg13g2_decap_8 FILLER_6_2334 ();
 sg13g2_decap_8 FILLER_6_2341 ();
 sg13g2_decap_8 FILLER_6_2348 ();
 sg13g2_decap_8 FILLER_6_2355 ();
 sg13g2_decap_8 FILLER_6_2362 ();
 sg13g2_decap_8 FILLER_6_2369 ();
 sg13g2_decap_8 FILLER_6_2376 ();
 sg13g2_decap_8 FILLER_6_2383 ();
 sg13g2_decap_8 FILLER_6_2390 ();
 sg13g2_decap_8 FILLER_6_2397 ();
 sg13g2_decap_8 FILLER_6_2404 ();
 sg13g2_decap_8 FILLER_6_2411 ();
 sg13g2_decap_8 FILLER_6_2418 ();
 sg13g2_decap_8 FILLER_6_2425 ();
 sg13g2_decap_8 FILLER_6_2432 ();
 sg13g2_decap_8 FILLER_6_2439 ();
 sg13g2_decap_8 FILLER_6_2446 ();
 sg13g2_decap_8 FILLER_6_2453 ();
 sg13g2_decap_8 FILLER_6_2460 ();
 sg13g2_decap_8 FILLER_6_2467 ();
 sg13g2_decap_8 FILLER_6_2474 ();
 sg13g2_decap_8 FILLER_6_2481 ();
 sg13g2_decap_8 FILLER_6_2488 ();
 sg13g2_decap_8 FILLER_6_2495 ();
 sg13g2_decap_8 FILLER_6_2502 ();
 sg13g2_decap_8 FILLER_6_2509 ();
 sg13g2_decap_8 FILLER_6_2516 ();
 sg13g2_decap_8 FILLER_6_2523 ();
 sg13g2_decap_8 FILLER_6_2530 ();
 sg13g2_decap_8 FILLER_6_2537 ();
 sg13g2_decap_8 FILLER_6_2544 ();
 sg13g2_decap_8 FILLER_6_2551 ();
 sg13g2_decap_8 FILLER_6_2558 ();
 sg13g2_decap_8 FILLER_6_2565 ();
 sg13g2_decap_8 FILLER_6_2572 ();
 sg13g2_decap_8 FILLER_6_2579 ();
 sg13g2_decap_8 FILLER_6_2586 ();
 sg13g2_decap_8 FILLER_6_2593 ();
 sg13g2_decap_8 FILLER_6_2600 ();
 sg13g2_decap_8 FILLER_6_2607 ();
 sg13g2_decap_8 FILLER_6_2614 ();
 sg13g2_decap_8 FILLER_6_2621 ();
 sg13g2_decap_8 FILLER_6_2628 ();
 sg13g2_decap_8 FILLER_6_2635 ();
 sg13g2_decap_8 FILLER_6_2642 ();
 sg13g2_decap_8 FILLER_6_2649 ();
 sg13g2_decap_8 FILLER_6_2656 ();
 sg13g2_decap_8 FILLER_6_2663 ();
 sg13g2_decap_4 FILLER_6_2670 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_1 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_459 ();
 sg13g2_fill_2 FILLER_7_495 ();
 sg13g2_decap_8 FILLER_7_506 ();
 sg13g2_decap_8 FILLER_7_513 ();
 sg13g2_decap_4 FILLER_7_520 ();
 sg13g2_fill_2 FILLER_7_524 ();
 sg13g2_fill_1 FILLER_7_530 ();
 sg13g2_fill_1 FILLER_7_593 ();
 sg13g2_fill_2 FILLER_7_625 ();
 sg13g2_fill_1 FILLER_7_627 ();
 sg13g2_decap_4 FILLER_7_632 ();
 sg13g2_fill_1 FILLER_7_636 ();
 sg13g2_fill_2 FILLER_7_681 ();
 sg13g2_fill_2 FILLER_7_688 ();
 sg13g2_fill_2 FILLER_7_716 ();
 sg13g2_fill_1 FILLER_7_718 ();
 sg13g2_fill_1 FILLER_7_753 ();
 sg13g2_fill_1 FILLER_7_759 ();
 sg13g2_fill_2 FILLER_7_791 ();
 sg13g2_fill_2 FILLER_7_817 ();
 sg13g2_fill_2 FILLER_7_858 ();
 sg13g2_fill_1 FILLER_7_860 ();
 sg13g2_fill_2 FILLER_7_866 ();
 sg13g2_fill_1 FILLER_7_868 ();
 sg13g2_fill_1 FILLER_7_913 ();
 sg13g2_fill_1 FILLER_7_948 ();
 sg13g2_fill_1 FILLER_7_1062 ();
 sg13g2_fill_2 FILLER_7_1071 ();
 sg13g2_fill_1 FILLER_7_1073 ();
 sg13g2_fill_1 FILLER_7_1090 ();
 sg13g2_fill_2 FILLER_7_1100 ();
 sg13g2_fill_1 FILLER_7_1137 ();
 sg13g2_decap_4 FILLER_7_1143 ();
 sg13g2_decap_4 FILLER_7_1166 ();
 sg13g2_fill_1 FILLER_7_1170 ();
 sg13g2_fill_2 FILLER_7_1211 ();
 sg13g2_fill_1 FILLER_7_1213 ();
 sg13g2_fill_1 FILLER_7_1240 ();
 sg13g2_fill_1 FILLER_7_1309 ();
 sg13g2_fill_1 FILLER_7_1315 ();
 sg13g2_fill_2 FILLER_7_1320 ();
 sg13g2_fill_1 FILLER_7_1322 ();
 sg13g2_fill_1 FILLER_7_1327 ();
 sg13g2_decap_4 FILLER_7_1337 ();
 sg13g2_fill_1 FILLER_7_1341 ();
 sg13g2_fill_2 FILLER_7_1408 ();
 sg13g2_fill_1 FILLER_7_1410 ();
 sg13g2_decap_4 FILLER_7_1464 ();
 sg13g2_fill_1 FILLER_7_1468 ();
 sg13g2_fill_2 FILLER_7_1500 ();
 sg13g2_fill_2 FILLER_7_1549 ();
 sg13g2_fill_1 FILLER_7_1573 ();
 sg13g2_fill_2 FILLER_7_1588 ();
 sg13g2_fill_2 FILLER_7_1616 ();
 sg13g2_fill_1 FILLER_7_1623 ();
 sg13g2_fill_1 FILLER_7_1646 ();
 sg13g2_fill_2 FILLER_7_1661 ();
 sg13g2_decap_8 FILLER_7_1689 ();
 sg13g2_fill_1 FILLER_7_1696 ();
 sg13g2_decap_4 FILLER_7_1701 ();
 sg13g2_fill_2 FILLER_7_1714 ();
 sg13g2_fill_2 FILLER_7_1741 ();
 sg13g2_fill_1 FILLER_7_1743 ();
 sg13g2_fill_1 FILLER_7_1776 ();
 sg13g2_fill_1 FILLER_7_1790 ();
 sg13g2_fill_2 FILLER_7_1825 ();
 sg13g2_fill_2 FILLER_7_1867 ();
 sg13g2_fill_2 FILLER_7_1899 ();
 sg13g2_fill_1 FILLER_7_1901 ();
 sg13g2_fill_2 FILLER_7_1927 ();
 sg13g2_fill_1 FILLER_7_1929 ();
 sg13g2_decap_8 FILLER_7_1935 ();
 sg13g2_fill_1 FILLER_7_1942 ();
 sg13g2_fill_1 FILLER_7_1997 ();
 sg13g2_fill_2 FILLER_7_2007 ();
 sg13g2_fill_1 FILLER_7_2009 ();
 sg13g2_fill_1 FILLER_7_2019 ();
 sg13g2_fill_2 FILLER_7_2029 ();
 sg13g2_fill_2 FILLER_7_2112 ();
 sg13g2_fill_1 FILLER_7_2119 ();
 sg13g2_fill_2 FILLER_7_2133 ();
 sg13g2_fill_1 FILLER_7_2135 ();
 sg13g2_fill_2 FILLER_7_2149 ();
 sg13g2_fill_1 FILLER_7_2151 ();
 sg13g2_fill_2 FILLER_7_2209 ();
 sg13g2_fill_2 FILLER_7_2232 ();
 sg13g2_fill_1 FILLER_7_2234 ();
 sg13g2_fill_1 FILLER_7_2250 ();
 sg13g2_decap_8 FILLER_7_2255 ();
 sg13g2_fill_2 FILLER_7_2262 ();
 sg13g2_fill_1 FILLER_7_2264 ();
 sg13g2_fill_2 FILLER_7_2269 ();
 sg13g2_fill_2 FILLER_7_2276 ();
 sg13g2_fill_1 FILLER_7_2278 ();
 sg13g2_fill_2 FILLER_7_2283 ();
 sg13g2_fill_1 FILLER_7_2321 ();
 sg13g2_fill_2 FILLER_7_2327 ();
 sg13g2_decap_8 FILLER_7_2338 ();
 sg13g2_decap_8 FILLER_7_2345 ();
 sg13g2_decap_8 FILLER_7_2352 ();
 sg13g2_decap_8 FILLER_7_2359 ();
 sg13g2_decap_8 FILLER_7_2366 ();
 sg13g2_decap_8 FILLER_7_2373 ();
 sg13g2_decap_8 FILLER_7_2380 ();
 sg13g2_decap_8 FILLER_7_2387 ();
 sg13g2_decap_8 FILLER_7_2394 ();
 sg13g2_decap_8 FILLER_7_2401 ();
 sg13g2_decap_8 FILLER_7_2408 ();
 sg13g2_decap_8 FILLER_7_2415 ();
 sg13g2_decap_8 FILLER_7_2422 ();
 sg13g2_decap_8 FILLER_7_2429 ();
 sg13g2_decap_8 FILLER_7_2436 ();
 sg13g2_decap_8 FILLER_7_2443 ();
 sg13g2_decap_8 FILLER_7_2450 ();
 sg13g2_decap_8 FILLER_7_2457 ();
 sg13g2_decap_8 FILLER_7_2464 ();
 sg13g2_decap_8 FILLER_7_2471 ();
 sg13g2_decap_8 FILLER_7_2478 ();
 sg13g2_decap_8 FILLER_7_2485 ();
 sg13g2_decap_8 FILLER_7_2492 ();
 sg13g2_decap_8 FILLER_7_2499 ();
 sg13g2_decap_8 FILLER_7_2506 ();
 sg13g2_decap_8 FILLER_7_2513 ();
 sg13g2_decap_8 FILLER_7_2520 ();
 sg13g2_decap_8 FILLER_7_2527 ();
 sg13g2_decap_8 FILLER_7_2534 ();
 sg13g2_decap_8 FILLER_7_2541 ();
 sg13g2_decap_8 FILLER_7_2548 ();
 sg13g2_decap_8 FILLER_7_2555 ();
 sg13g2_decap_8 FILLER_7_2562 ();
 sg13g2_decap_8 FILLER_7_2569 ();
 sg13g2_decap_8 FILLER_7_2576 ();
 sg13g2_decap_8 FILLER_7_2583 ();
 sg13g2_decap_8 FILLER_7_2590 ();
 sg13g2_decap_8 FILLER_7_2597 ();
 sg13g2_decap_8 FILLER_7_2604 ();
 sg13g2_decap_8 FILLER_7_2611 ();
 sg13g2_decap_8 FILLER_7_2618 ();
 sg13g2_decap_8 FILLER_7_2625 ();
 sg13g2_decap_8 FILLER_7_2632 ();
 sg13g2_decap_8 FILLER_7_2639 ();
 sg13g2_decap_8 FILLER_7_2646 ();
 sg13g2_decap_8 FILLER_7_2653 ();
 sg13g2_decap_8 FILLER_7_2660 ();
 sg13g2_decap_8 FILLER_7_2667 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_451 ();
 sg13g2_fill_2 FILLER_8_461 ();
 sg13g2_fill_1 FILLER_8_480 ();
 sg13g2_fill_2 FILLER_8_490 ();
 sg13g2_fill_2 FILLER_8_588 ();
 sg13g2_fill_1 FILLER_8_590 ();
 sg13g2_decap_8 FILLER_8_638 ();
 sg13g2_fill_1 FILLER_8_645 ();
 sg13g2_fill_2 FILLER_8_650 ();
 sg13g2_fill_1 FILLER_8_656 ();
 sg13g2_fill_2 FILLER_8_683 ();
 sg13g2_fill_1 FILLER_8_685 ();
 sg13g2_fill_2 FILLER_8_720 ();
 sg13g2_fill_1 FILLER_8_722 ();
 sg13g2_fill_1 FILLER_8_728 ();
 sg13g2_fill_1 FILLER_8_743 ();
 sg13g2_fill_1 FILLER_8_762 ();
 sg13g2_fill_2 FILLER_8_802 ();
 sg13g2_fill_1 FILLER_8_804 ();
 sg13g2_fill_2 FILLER_8_819 ();
 sg13g2_fill_1 FILLER_8_821 ();
 sg13g2_fill_1 FILLER_8_848 ();
 sg13g2_fill_2 FILLER_8_892 ();
 sg13g2_fill_1 FILLER_8_894 ();
 sg13g2_fill_2 FILLER_8_930 ();
 sg13g2_fill_1 FILLER_8_932 ();
 sg13g2_decap_4 FILLER_8_980 ();
 sg13g2_fill_2 FILLER_8_984 ();
 sg13g2_fill_2 FILLER_8_995 ();
 sg13g2_fill_1 FILLER_8_1002 ();
 sg13g2_fill_2 FILLER_8_1008 ();
 sg13g2_fill_1 FILLER_8_1066 ();
 sg13g2_decap_4 FILLER_8_1110 ();
 sg13g2_fill_1 FILLER_8_1114 ();
 sg13g2_decap_4 FILLER_8_1170 ();
 sg13g2_fill_1 FILLER_8_1174 ();
 sg13g2_fill_2 FILLER_8_1192 ();
 sg13g2_fill_1 FILLER_8_1194 ();
 sg13g2_decap_8 FILLER_8_1229 ();
 sg13g2_fill_2 FILLER_8_1236 ();
 sg13g2_fill_1 FILLER_8_1238 ();
 sg13g2_fill_2 FILLER_8_1270 ();
 sg13g2_fill_1 FILLER_8_1272 ();
 sg13g2_fill_2 FILLER_8_1287 ();
 sg13g2_fill_2 FILLER_8_1303 ();
 sg13g2_fill_2 FILLER_8_1331 ();
 sg13g2_fill_1 FILLER_8_1333 ();
 sg13g2_fill_2 FILLER_8_1379 ();
 sg13g2_fill_1 FILLER_8_1402 ();
 sg13g2_decap_4 FILLER_8_1421 ();
 sg13g2_fill_2 FILLER_8_1425 ();
 sg13g2_fill_2 FILLER_8_1431 ();
 sg13g2_fill_2 FILLER_8_1442 ();
 sg13g2_fill_1 FILLER_8_1500 ();
 sg13g2_fill_2 FILLER_8_1521 ();
 sg13g2_fill_1 FILLER_8_1523 ();
 sg13g2_fill_1 FILLER_8_1591 ();
 sg13g2_fill_1 FILLER_8_1665 ();
 sg13g2_fill_2 FILLER_8_1670 ();
 sg13g2_fill_1 FILLER_8_1690 ();
 sg13g2_fill_1 FILLER_8_1717 ();
 sg13g2_fill_2 FILLER_8_1741 ();
 sg13g2_fill_1 FILLER_8_1743 ();
 sg13g2_fill_1 FILLER_8_1809 ();
 sg13g2_fill_2 FILLER_8_1844 ();
 sg13g2_fill_1 FILLER_8_1846 ();
 sg13g2_fill_2 FILLER_8_1852 ();
 sg13g2_fill_1 FILLER_8_1867 ();
 sg13g2_fill_2 FILLER_8_1894 ();
 sg13g2_fill_2 FILLER_8_1914 ();
 sg13g2_fill_1 FILLER_8_1916 ();
 sg13g2_fill_1 FILLER_8_1960 ();
 sg13g2_fill_1 FILLER_8_1997 ();
 sg13g2_fill_2 FILLER_8_2003 ();
 sg13g2_fill_2 FILLER_8_2031 ();
 sg13g2_fill_1 FILLER_8_2033 ();
 sg13g2_decap_8 FILLER_8_2055 ();
 sg13g2_decap_8 FILLER_8_2062 ();
 sg13g2_fill_1 FILLER_8_2069 ();
 sg13g2_fill_2 FILLER_8_2074 ();
 sg13g2_fill_1 FILLER_8_2076 ();
 sg13g2_fill_1 FILLER_8_2150 ();
 sg13g2_fill_1 FILLER_8_2170 ();
 sg13g2_decap_4 FILLER_8_2244 ();
 sg13g2_fill_1 FILLER_8_2248 ();
 sg13g2_decap_8 FILLER_8_2350 ();
 sg13g2_decap_8 FILLER_8_2357 ();
 sg13g2_decap_8 FILLER_8_2364 ();
 sg13g2_decap_8 FILLER_8_2371 ();
 sg13g2_decap_8 FILLER_8_2378 ();
 sg13g2_decap_8 FILLER_8_2385 ();
 sg13g2_decap_8 FILLER_8_2392 ();
 sg13g2_decap_8 FILLER_8_2399 ();
 sg13g2_decap_8 FILLER_8_2406 ();
 sg13g2_decap_8 FILLER_8_2413 ();
 sg13g2_decap_8 FILLER_8_2420 ();
 sg13g2_decap_8 FILLER_8_2427 ();
 sg13g2_decap_8 FILLER_8_2434 ();
 sg13g2_decap_8 FILLER_8_2441 ();
 sg13g2_decap_8 FILLER_8_2448 ();
 sg13g2_decap_8 FILLER_8_2455 ();
 sg13g2_decap_8 FILLER_8_2462 ();
 sg13g2_decap_8 FILLER_8_2469 ();
 sg13g2_decap_8 FILLER_8_2476 ();
 sg13g2_decap_8 FILLER_8_2483 ();
 sg13g2_decap_8 FILLER_8_2490 ();
 sg13g2_decap_8 FILLER_8_2497 ();
 sg13g2_decap_8 FILLER_8_2504 ();
 sg13g2_decap_8 FILLER_8_2511 ();
 sg13g2_decap_8 FILLER_8_2518 ();
 sg13g2_decap_8 FILLER_8_2525 ();
 sg13g2_decap_8 FILLER_8_2532 ();
 sg13g2_decap_8 FILLER_8_2539 ();
 sg13g2_decap_8 FILLER_8_2546 ();
 sg13g2_decap_8 FILLER_8_2553 ();
 sg13g2_decap_8 FILLER_8_2560 ();
 sg13g2_decap_8 FILLER_8_2567 ();
 sg13g2_decap_8 FILLER_8_2574 ();
 sg13g2_decap_8 FILLER_8_2581 ();
 sg13g2_decap_8 FILLER_8_2588 ();
 sg13g2_decap_8 FILLER_8_2595 ();
 sg13g2_decap_8 FILLER_8_2602 ();
 sg13g2_decap_8 FILLER_8_2609 ();
 sg13g2_decap_8 FILLER_8_2616 ();
 sg13g2_decap_8 FILLER_8_2623 ();
 sg13g2_decap_8 FILLER_8_2630 ();
 sg13g2_decap_8 FILLER_8_2637 ();
 sg13g2_decap_8 FILLER_8_2644 ();
 sg13g2_decap_8 FILLER_8_2651 ();
 sg13g2_decap_8 FILLER_8_2658 ();
 sg13g2_decap_8 FILLER_8_2665 ();
 sg13g2_fill_2 FILLER_8_2672 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_fill_2 FILLER_9_465 ();
 sg13g2_decap_4 FILLER_9_489 ();
 sg13g2_fill_1 FILLER_9_493 ();
 sg13g2_fill_2 FILLER_9_503 ();
 sg13g2_fill_1 FILLER_9_505 ();
 sg13g2_fill_1 FILLER_9_568 ();
 sg13g2_fill_2 FILLER_9_608 ();
 sg13g2_fill_2 FILLER_9_640 ();
 sg13g2_fill_2 FILLER_9_656 ();
 sg13g2_fill_1 FILLER_9_658 ();
 sg13g2_fill_2 FILLER_9_669 ();
 sg13g2_fill_1 FILLER_9_671 ();
 sg13g2_fill_1 FILLER_9_712 ();
 sg13g2_fill_2 FILLER_9_730 ();
 sg13g2_fill_1 FILLER_9_737 ();
 sg13g2_fill_1 FILLER_9_778 ();
 sg13g2_fill_2 FILLER_9_788 ();
 sg13g2_fill_1 FILLER_9_790 ();
 sg13g2_fill_2 FILLER_9_804 ();
 sg13g2_fill_2 FILLER_9_832 ();
 sg13g2_fill_1 FILLER_9_938 ();
 sg13g2_fill_2 FILLER_9_965 ();
 sg13g2_fill_1 FILLER_9_967 ();
 sg13g2_fill_2 FILLER_9_1020 ();
 sg13g2_fill_1 FILLER_9_1103 ();
 sg13g2_fill_2 FILLER_9_1130 ();
 sg13g2_fill_1 FILLER_9_1150 ();
 sg13g2_decap_4 FILLER_9_1155 ();
 sg13g2_fill_1 FILLER_9_1159 ();
 sg13g2_fill_2 FILLER_9_1169 ();
 sg13g2_fill_1 FILLER_9_1171 ();
 sg13g2_fill_1 FILLER_9_1206 ();
 sg13g2_fill_1 FILLER_9_1268 ();
 sg13g2_decap_8 FILLER_9_1342 ();
 sg13g2_decap_8 FILLER_9_1353 ();
 sg13g2_fill_2 FILLER_9_1360 ();
 sg13g2_fill_2 FILLER_9_1422 ();
 sg13g2_fill_2 FILLER_9_1432 ();
 sg13g2_fill_1 FILLER_9_1434 ();
 sg13g2_fill_2 FILLER_9_1456 ();
 sg13g2_fill_1 FILLER_9_1458 ();
 sg13g2_fill_2 FILLER_9_1538 ();
 sg13g2_fill_1 FILLER_9_1540 ();
 sg13g2_fill_2 FILLER_9_1550 ();
 sg13g2_fill_2 FILLER_9_1583 ();
 sg13g2_fill_1 FILLER_9_1585 ();
 sg13g2_decap_4 FILLER_9_1590 ();
 sg13g2_fill_1 FILLER_9_1594 ();
 sg13g2_fill_2 FILLER_9_1608 ();
 sg13g2_fill_2 FILLER_9_1649 ();
 sg13g2_fill_1 FILLER_9_1651 ();
 sg13g2_fill_1 FILLER_9_1761 ();
 sg13g2_fill_2 FILLER_9_1794 ();
 sg13g2_fill_1 FILLER_9_1817 ();
 sg13g2_fill_2 FILLER_9_1889 ();
 sg13g2_fill_1 FILLER_9_1922 ();
 sg13g2_fill_1 FILLER_9_1958 ();
 sg13g2_fill_2 FILLER_9_1987 ();
 sg13g2_fill_2 FILLER_9_2028 ();
 sg13g2_fill_1 FILLER_9_2030 ();
 sg13g2_fill_2 FILLER_9_2036 ();
 sg13g2_fill_2 FILLER_9_2123 ();
 sg13g2_fill_1 FILLER_9_2194 ();
 sg13g2_fill_2 FILLER_9_2200 ();
 sg13g2_fill_1 FILLER_9_2202 ();
 sg13g2_decap_4 FILLER_9_2273 ();
 sg13g2_fill_2 FILLER_9_2285 ();
 sg13g2_fill_1 FILLER_9_2287 ();
 sg13g2_fill_2 FILLER_9_2306 ();
 sg13g2_fill_1 FILLER_9_2308 ();
 sg13g2_fill_1 FILLER_9_2332 ();
 sg13g2_decap_8 FILLER_9_2368 ();
 sg13g2_decap_8 FILLER_9_2375 ();
 sg13g2_decap_8 FILLER_9_2382 ();
 sg13g2_decap_8 FILLER_9_2389 ();
 sg13g2_decap_8 FILLER_9_2396 ();
 sg13g2_decap_8 FILLER_9_2403 ();
 sg13g2_decap_8 FILLER_9_2410 ();
 sg13g2_decap_8 FILLER_9_2417 ();
 sg13g2_decap_8 FILLER_9_2424 ();
 sg13g2_decap_8 FILLER_9_2431 ();
 sg13g2_decap_8 FILLER_9_2438 ();
 sg13g2_decap_8 FILLER_9_2445 ();
 sg13g2_decap_8 FILLER_9_2452 ();
 sg13g2_decap_8 FILLER_9_2459 ();
 sg13g2_decap_8 FILLER_9_2466 ();
 sg13g2_decap_8 FILLER_9_2473 ();
 sg13g2_decap_8 FILLER_9_2480 ();
 sg13g2_decap_8 FILLER_9_2487 ();
 sg13g2_decap_8 FILLER_9_2494 ();
 sg13g2_decap_8 FILLER_9_2501 ();
 sg13g2_decap_8 FILLER_9_2508 ();
 sg13g2_decap_8 FILLER_9_2515 ();
 sg13g2_decap_8 FILLER_9_2522 ();
 sg13g2_decap_8 FILLER_9_2529 ();
 sg13g2_decap_8 FILLER_9_2536 ();
 sg13g2_decap_8 FILLER_9_2543 ();
 sg13g2_decap_8 FILLER_9_2550 ();
 sg13g2_decap_8 FILLER_9_2557 ();
 sg13g2_decap_8 FILLER_9_2564 ();
 sg13g2_decap_8 FILLER_9_2571 ();
 sg13g2_decap_8 FILLER_9_2578 ();
 sg13g2_decap_8 FILLER_9_2585 ();
 sg13g2_decap_8 FILLER_9_2592 ();
 sg13g2_decap_8 FILLER_9_2599 ();
 sg13g2_decap_8 FILLER_9_2606 ();
 sg13g2_decap_8 FILLER_9_2613 ();
 sg13g2_decap_8 FILLER_9_2620 ();
 sg13g2_decap_8 FILLER_9_2627 ();
 sg13g2_decap_8 FILLER_9_2634 ();
 sg13g2_decap_8 FILLER_9_2641 ();
 sg13g2_decap_8 FILLER_9_2648 ();
 sg13g2_decap_8 FILLER_9_2655 ();
 sg13g2_decap_8 FILLER_9_2662 ();
 sg13g2_decap_4 FILLER_9_2669 ();
 sg13g2_fill_1 FILLER_9_2673 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_4 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_424 ();
 sg13g2_fill_1 FILLER_10_466 ();
 sg13g2_decap_8 FILLER_10_519 ();
 sg13g2_fill_1 FILLER_10_526 ();
 sg13g2_fill_2 FILLER_10_535 ();
 sg13g2_fill_2 FILLER_10_558 ();
 sg13g2_decap_8 FILLER_10_582 ();
 sg13g2_fill_2 FILLER_10_589 ();
 sg13g2_fill_1 FILLER_10_604 ();
 sg13g2_fill_1 FILLER_10_628 ();
 sg13g2_fill_1 FILLER_10_650 ();
 sg13g2_fill_1 FILLER_10_670 ();
 sg13g2_fill_2 FILLER_10_702 ();
 sg13g2_fill_1 FILLER_10_704 ();
 sg13g2_fill_1 FILLER_10_722 ();
 sg13g2_fill_2 FILLER_10_737 ();
 sg13g2_fill_1 FILLER_10_744 ();
 sg13g2_fill_1 FILLER_10_758 ();
 sg13g2_fill_2 FILLER_10_816 ();
 sg13g2_fill_1 FILLER_10_818 ();
 sg13g2_fill_2 FILLER_10_839 ();
 sg13g2_fill_1 FILLER_10_841 ();
 sg13g2_fill_1 FILLER_10_864 ();
 sg13g2_fill_2 FILLER_10_899 ();
 sg13g2_fill_1 FILLER_10_901 ();
 sg13g2_fill_2 FILLER_10_927 ();
 sg13g2_fill_1 FILLER_10_939 ();
 sg13g2_fill_1 FILLER_10_949 ();
 sg13g2_fill_2 FILLER_10_958 ();
 sg13g2_fill_2 FILLER_10_969 ();
 sg13g2_fill_1 FILLER_10_971 ();
 sg13g2_fill_1 FILLER_10_976 ();
 sg13g2_fill_2 FILLER_10_1026 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_fill_1 FILLER_10_1038 ();
 sg13g2_fill_2 FILLER_10_1043 ();
 sg13g2_fill_1 FILLER_10_1045 ();
 sg13g2_fill_1 FILLER_10_1070 ();
 sg13g2_fill_1 FILLER_10_1078 ();
 sg13g2_decap_4 FILLER_10_1125 ();
 sg13g2_fill_1 FILLER_10_1129 ();
 sg13g2_fill_1 FILLER_10_1143 ();
 sg13g2_fill_1 FILLER_10_1154 ();
 sg13g2_fill_1 FILLER_10_1190 ();
 sg13g2_fill_1 FILLER_10_1217 ();
 sg13g2_fill_1 FILLER_10_1227 ();
 sg13g2_fill_2 FILLER_10_1232 ();
 sg13g2_decap_4 FILLER_10_1239 ();
 sg13g2_fill_2 FILLER_10_1243 ();
 sg13g2_fill_2 FILLER_10_1250 ();
 sg13g2_fill_1 FILLER_10_1301 ();
 sg13g2_fill_2 FILLER_10_1312 ();
 sg13g2_decap_4 FILLER_10_1323 ();
 sg13g2_fill_1 FILLER_10_1327 ();
 sg13g2_fill_2 FILLER_10_1333 ();
 sg13g2_fill_1 FILLER_10_1335 ();
 sg13g2_fill_1 FILLER_10_1340 ();
 sg13g2_fill_2 FILLER_10_1387 ();
 sg13g2_fill_1 FILLER_10_1389 ();
 sg13g2_fill_1 FILLER_10_1409 ();
 sg13g2_fill_1 FILLER_10_1441 ();
 sg13g2_fill_2 FILLER_10_1447 ();
 sg13g2_fill_1 FILLER_10_1449 ();
 sg13g2_decap_4 FILLER_10_1454 ();
 sg13g2_fill_2 FILLER_10_1458 ();
 sg13g2_fill_2 FILLER_10_1474 ();
 sg13g2_fill_1 FILLER_10_1479 ();
 sg13g2_fill_1 FILLER_10_1502 ();
 sg13g2_fill_1 FILLER_10_1552 ();
 sg13g2_fill_1 FILLER_10_1562 ();
 sg13g2_decap_8 FILLER_10_1576 ();
 sg13g2_fill_1 FILLER_10_1587 ();
 sg13g2_fill_1 FILLER_10_1636 ();
 sg13g2_fill_2 FILLER_10_1701 ();
 sg13g2_fill_2 FILLER_10_1725 ();
 sg13g2_decap_4 FILLER_10_1834 ();
 sg13g2_fill_2 FILLER_10_1850 ();
 sg13g2_fill_2 FILLER_10_1871 ();
 sg13g2_fill_1 FILLER_10_1873 ();
 sg13g2_fill_2 FILLER_10_1892 ();
 sg13g2_fill_2 FILLER_10_1898 ();
 sg13g2_decap_4 FILLER_10_1913 ();
 sg13g2_fill_2 FILLER_10_1929 ();
 sg13g2_fill_2 FILLER_10_1940 ();
 sg13g2_decap_4 FILLER_10_1998 ();
 sg13g2_fill_1 FILLER_10_2023 ();
 sg13g2_fill_2 FILLER_10_2074 ();
 sg13g2_decap_4 FILLER_10_2110 ();
 sg13g2_decap_8 FILLER_10_2153 ();
 sg13g2_decap_4 FILLER_10_2160 ();
 sg13g2_fill_2 FILLER_10_2168 ();
 sg13g2_fill_2 FILLER_10_2179 ();
 sg13g2_fill_1 FILLER_10_2190 ();
 sg13g2_fill_2 FILLER_10_2201 ();
 sg13g2_fill_2 FILLER_10_2217 ();
 sg13g2_fill_1 FILLER_10_2219 ();
 sg13g2_fill_2 FILLER_10_2230 ();
 sg13g2_fill_2 FILLER_10_2266 ();
 sg13g2_decap_8 FILLER_10_2273 ();
 sg13g2_decap_4 FILLER_10_2280 ();
 sg13g2_fill_2 FILLER_10_2284 ();
 sg13g2_fill_1 FILLER_10_2295 ();
 sg13g2_fill_2 FILLER_10_2301 ();
 sg13g2_fill_1 FILLER_10_2303 ();
 sg13g2_fill_2 FILLER_10_2316 ();
 sg13g2_decap_8 FILLER_10_2352 ();
 sg13g2_decap_8 FILLER_10_2359 ();
 sg13g2_decap_8 FILLER_10_2366 ();
 sg13g2_decap_8 FILLER_10_2373 ();
 sg13g2_decap_8 FILLER_10_2380 ();
 sg13g2_decap_8 FILLER_10_2387 ();
 sg13g2_decap_8 FILLER_10_2394 ();
 sg13g2_decap_8 FILLER_10_2401 ();
 sg13g2_decap_8 FILLER_10_2408 ();
 sg13g2_decap_8 FILLER_10_2415 ();
 sg13g2_decap_8 FILLER_10_2422 ();
 sg13g2_decap_8 FILLER_10_2429 ();
 sg13g2_decap_8 FILLER_10_2436 ();
 sg13g2_decap_8 FILLER_10_2443 ();
 sg13g2_decap_8 FILLER_10_2450 ();
 sg13g2_decap_8 FILLER_10_2457 ();
 sg13g2_decap_8 FILLER_10_2464 ();
 sg13g2_decap_8 FILLER_10_2471 ();
 sg13g2_decap_8 FILLER_10_2478 ();
 sg13g2_decap_8 FILLER_10_2485 ();
 sg13g2_decap_8 FILLER_10_2492 ();
 sg13g2_decap_8 FILLER_10_2499 ();
 sg13g2_decap_8 FILLER_10_2506 ();
 sg13g2_decap_8 FILLER_10_2513 ();
 sg13g2_decap_8 FILLER_10_2520 ();
 sg13g2_decap_8 FILLER_10_2527 ();
 sg13g2_decap_8 FILLER_10_2534 ();
 sg13g2_decap_8 FILLER_10_2541 ();
 sg13g2_decap_8 FILLER_10_2548 ();
 sg13g2_decap_8 FILLER_10_2555 ();
 sg13g2_decap_8 FILLER_10_2562 ();
 sg13g2_decap_8 FILLER_10_2569 ();
 sg13g2_decap_8 FILLER_10_2576 ();
 sg13g2_decap_8 FILLER_10_2583 ();
 sg13g2_decap_8 FILLER_10_2590 ();
 sg13g2_decap_8 FILLER_10_2597 ();
 sg13g2_decap_8 FILLER_10_2604 ();
 sg13g2_decap_8 FILLER_10_2611 ();
 sg13g2_decap_8 FILLER_10_2618 ();
 sg13g2_decap_8 FILLER_10_2625 ();
 sg13g2_decap_8 FILLER_10_2632 ();
 sg13g2_decap_8 FILLER_10_2639 ();
 sg13g2_decap_8 FILLER_10_2646 ();
 sg13g2_decap_8 FILLER_10_2653 ();
 sg13g2_decap_8 FILLER_10_2660 ();
 sg13g2_decap_8 FILLER_10_2667 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_4 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_431 ();
 sg13g2_fill_1 FILLER_11_449 ();
 sg13g2_fill_2 FILLER_11_485 ();
 sg13g2_fill_1 FILLER_11_487 ();
 sg13g2_fill_2 FILLER_11_493 ();
 sg13g2_fill_2 FILLER_11_512 ();
 sg13g2_fill_1 FILLER_11_559 ();
 sg13g2_fill_1 FILLER_11_660 ();
 sg13g2_fill_1 FILLER_11_666 ();
 sg13g2_decap_4 FILLER_11_676 ();
 sg13g2_fill_2 FILLER_11_680 ();
 sg13g2_fill_2 FILLER_11_695 ();
 sg13g2_fill_1 FILLER_11_707 ();
 sg13g2_fill_2 FILLER_11_769 ();
 sg13g2_fill_1 FILLER_11_781 ();
 sg13g2_fill_2 FILLER_11_801 ();
 sg13g2_decap_8 FILLER_11_834 ();
 sg13g2_decap_4 FILLER_11_841 ();
 sg13g2_fill_1 FILLER_11_885 ();
 sg13g2_fill_2 FILLER_11_895 ();
 sg13g2_fill_1 FILLER_11_907 ();
 sg13g2_fill_1 FILLER_11_965 ();
 sg13g2_fill_1 FILLER_11_997 ();
 sg13g2_fill_1 FILLER_11_1067 ();
 sg13g2_fill_2 FILLER_11_1094 ();
 sg13g2_fill_2 FILLER_11_1153 ();
 sg13g2_fill_2 FILLER_11_1188 ();
 sg13g2_fill_1 FILLER_11_1190 ();
 sg13g2_fill_2 FILLER_11_1200 ();
 sg13g2_fill_1 FILLER_11_1202 ();
 sg13g2_decap_4 FILLER_11_1277 ();
 sg13g2_fill_2 FILLER_11_1293 ();
 sg13g2_fill_1 FILLER_11_1295 ();
 sg13g2_fill_1 FILLER_11_1300 ();
 sg13g2_fill_2 FILLER_11_1310 ();
 sg13g2_fill_1 FILLER_11_1312 ();
 sg13g2_fill_1 FILLER_11_1387 ();
 sg13g2_fill_2 FILLER_11_1428 ();
 sg13g2_fill_1 FILLER_11_1465 ();
 sg13g2_fill_1 FILLER_11_1475 ();
 sg13g2_fill_2 FILLER_11_1487 ();
 sg13g2_fill_1 FILLER_11_1515 ();
 sg13g2_fill_2 FILLER_11_1536 ();
 sg13g2_fill_1 FILLER_11_1538 ();
 sg13g2_decap_8 FILLER_11_1586 ();
 sg13g2_decap_4 FILLER_11_1593 ();
 sg13g2_fill_1 FILLER_11_1597 ();
 sg13g2_decap_8 FILLER_11_1606 ();
 sg13g2_fill_2 FILLER_11_1613 ();
 sg13g2_fill_2 FILLER_11_1668 ();
 sg13g2_fill_2 FILLER_11_1679 ();
 sg13g2_fill_1 FILLER_11_1681 ();
 sg13g2_decap_8 FILLER_11_1695 ();
 sg13g2_fill_2 FILLER_11_1702 ();
 sg13g2_fill_1 FILLER_11_1704 ();
 sg13g2_decap_8 FILLER_11_1770 ();
 sg13g2_fill_2 FILLER_11_1782 ();
 sg13g2_fill_2 FILLER_11_1792 ();
 sg13g2_fill_1 FILLER_11_1794 ();
 sg13g2_fill_1 FILLER_11_1834 ();
 sg13g2_fill_1 FILLER_11_1854 ();
 sg13g2_fill_1 FILLER_11_1872 ();
 sg13g2_fill_1 FILLER_11_1913 ();
 sg13g2_fill_2 FILLER_11_1945 ();
 sg13g2_decap_4 FILLER_11_1951 ();
 sg13g2_fill_1 FILLER_11_1973 ();
 sg13g2_fill_2 FILLER_11_2005 ();
 sg13g2_fill_1 FILLER_11_2007 ();
 sg13g2_fill_1 FILLER_11_2018 ();
 sg13g2_fill_1 FILLER_11_2058 ();
 sg13g2_fill_2 FILLER_11_2085 ();
 sg13g2_fill_1 FILLER_11_2087 ();
 sg13g2_fill_1 FILLER_11_2097 ();
 sg13g2_fill_1 FILLER_11_2232 ();
 sg13g2_fill_2 FILLER_11_2247 ();
 sg13g2_fill_1 FILLER_11_2249 ();
 sg13g2_decap_8 FILLER_11_2351 ();
 sg13g2_decap_8 FILLER_11_2358 ();
 sg13g2_decap_8 FILLER_11_2365 ();
 sg13g2_decap_8 FILLER_11_2372 ();
 sg13g2_decap_8 FILLER_11_2379 ();
 sg13g2_decap_8 FILLER_11_2386 ();
 sg13g2_decap_8 FILLER_11_2393 ();
 sg13g2_decap_8 FILLER_11_2400 ();
 sg13g2_decap_8 FILLER_11_2407 ();
 sg13g2_decap_8 FILLER_11_2414 ();
 sg13g2_decap_8 FILLER_11_2421 ();
 sg13g2_decap_8 FILLER_11_2428 ();
 sg13g2_decap_8 FILLER_11_2435 ();
 sg13g2_decap_8 FILLER_11_2442 ();
 sg13g2_decap_8 FILLER_11_2449 ();
 sg13g2_decap_8 FILLER_11_2456 ();
 sg13g2_decap_8 FILLER_11_2463 ();
 sg13g2_decap_8 FILLER_11_2470 ();
 sg13g2_decap_8 FILLER_11_2477 ();
 sg13g2_decap_8 FILLER_11_2484 ();
 sg13g2_decap_8 FILLER_11_2491 ();
 sg13g2_decap_8 FILLER_11_2498 ();
 sg13g2_decap_8 FILLER_11_2505 ();
 sg13g2_decap_8 FILLER_11_2512 ();
 sg13g2_decap_8 FILLER_11_2519 ();
 sg13g2_decap_8 FILLER_11_2526 ();
 sg13g2_decap_8 FILLER_11_2533 ();
 sg13g2_decap_8 FILLER_11_2540 ();
 sg13g2_decap_8 FILLER_11_2547 ();
 sg13g2_decap_8 FILLER_11_2554 ();
 sg13g2_decap_8 FILLER_11_2561 ();
 sg13g2_decap_8 FILLER_11_2568 ();
 sg13g2_decap_8 FILLER_11_2575 ();
 sg13g2_decap_8 FILLER_11_2582 ();
 sg13g2_decap_8 FILLER_11_2589 ();
 sg13g2_decap_8 FILLER_11_2596 ();
 sg13g2_decap_8 FILLER_11_2603 ();
 sg13g2_decap_8 FILLER_11_2610 ();
 sg13g2_decap_8 FILLER_11_2617 ();
 sg13g2_decap_8 FILLER_11_2624 ();
 sg13g2_decap_8 FILLER_11_2631 ();
 sg13g2_decap_8 FILLER_11_2638 ();
 sg13g2_decap_8 FILLER_11_2645 ();
 sg13g2_decap_8 FILLER_11_2652 ();
 sg13g2_decap_8 FILLER_11_2659 ();
 sg13g2_decap_8 FILLER_11_2666 ();
 sg13g2_fill_1 FILLER_11_2673 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_4 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_424 ();
 sg13g2_fill_1 FILLER_12_505 ();
 sg13g2_fill_1 FILLER_12_520 ();
 sg13g2_decap_4 FILLER_12_543 ();
 sg13g2_decap_8 FILLER_12_590 ();
 sg13g2_fill_2 FILLER_12_597 ();
 sg13g2_fill_2 FILLER_12_607 ();
 sg13g2_fill_1 FILLER_12_609 ();
 sg13g2_fill_2 FILLER_12_614 ();
 sg13g2_fill_1 FILLER_12_616 ();
 sg13g2_decap_4 FILLER_12_621 ();
 sg13g2_fill_1 FILLER_12_625 ();
 sg13g2_fill_2 FILLER_12_643 ();
 sg13g2_fill_1 FILLER_12_645 ();
 sg13g2_fill_2 FILLER_12_681 ();
 sg13g2_fill_1 FILLER_12_683 ();
 sg13g2_decap_4 FILLER_12_702 ();
 sg13g2_fill_1 FILLER_12_706 ();
 sg13g2_decap_8 FILLER_12_724 ();
 sg13g2_fill_1 FILLER_12_731 ();
 sg13g2_fill_1 FILLER_12_736 ();
 sg13g2_fill_1 FILLER_12_745 ();
 sg13g2_decap_4 FILLER_12_754 ();
 sg13g2_fill_1 FILLER_12_758 ();
 sg13g2_fill_1 FILLER_12_822 ();
 sg13g2_fill_2 FILLER_12_872 ();
 sg13g2_fill_1 FILLER_12_919 ();
 sg13g2_fill_2 FILLER_12_970 ();
 sg13g2_decap_4 FILLER_12_981 ();
 sg13g2_decap_4 FILLER_12_989 ();
 sg13g2_fill_2 FILLER_12_993 ();
 sg13g2_fill_2 FILLER_12_1005 ();
 sg13g2_fill_1 FILLER_12_1017 ();
 sg13g2_decap_8 FILLER_12_1026 ();
 sg13g2_decap_8 FILLER_12_1033 ();
 sg13g2_decap_4 FILLER_12_1046 ();
 sg13g2_fill_2 FILLER_12_1050 ();
 sg13g2_fill_2 FILLER_12_1066 ();
 sg13g2_fill_1 FILLER_12_1068 ();
 sg13g2_fill_1 FILLER_12_1078 ();
 sg13g2_fill_1 FILLER_12_1093 ();
 sg13g2_fill_1 FILLER_12_1099 ();
 sg13g2_fill_2 FILLER_12_1109 ();
 sg13g2_fill_1 FILLER_12_1111 ();
 sg13g2_fill_1 FILLER_12_1125 ();
 sg13g2_fill_2 FILLER_12_1148 ();
 sg13g2_fill_1 FILLER_12_1150 ();
 sg13g2_fill_1 FILLER_12_1167 ();
 sg13g2_fill_2 FILLER_12_1194 ();
 sg13g2_fill_2 FILLER_12_1242 ();
 sg13g2_fill_1 FILLER_12_1279 ();
 sg13g2_decap_8 FILLER_12_1311 ();
 sg13g2_fill_2 FILLER_12_1318 ();
 sg13g2_fill_1 FILLER_12_1320 ();
 sg13g2_fill_2 FILLER_12_1369 ();
 sg13g2_decap_8 FILLER_12_1406 ();
 sg13g2_decap_4 FILLER_12_1439 ();
 sg13g2_fill_2 FILLER_12_1443 ();
 sg13g2_fill_1 FILLER_12_1479 ();
 sg13g2_fill_2 FILLER_12_1561 ();
 sg13g2_fill_2 FILLER_12_1577 ();
 sg13g2_fill_2 FILLER_12_1603 ();
 sg13g2_fill_1 FILLER_12_1631 ();
 sg13g2_fill_2 FILLER_12_1637 ();
 sg13g2_fill_2 FILLER_12_1649 ();
 sg13g2_fill_2 FILLER_12_1693 ();
 sg13g2_fill_1 FILLER_12_1695 ();
 sg13g2_fill_2 FILLER_12_1706 ();
 sg13g2_fill_1 FILLER_12_1708 ();
 sg13g2_fill_2 FILLER_12_1735 ();
 sg13g2_fill_2 FILLER_12_1754 ();
 sg13g2_fill_1 FILLER_12_1756 ();
 sg13g2_decap_4 FILLER_12_1766 ();
 sg13g2_fill_1 FILLER_12_1770 ();
 sg13g2_fill_2 FILLER_12_1811 ();
 sg13g2_fill_1 FILLER_12_1822 ();
 sg13g2_decap_8 FILLER_12_1885 ();
 sg13g2_decap_4 FILLER_12_1892 ();
 sg13g2_fill_2 FILLER_12_1896 ();
 sg13g2_fill_2 FILLER_12_1924 ();
 sg13g2_fill_1 FILLER_12_1926 ();
 sg13g2_fill_2 FILLER_12_1988 ();
 sg13g2_fill_1 FILLER_12_1990 ();
 sg13g2_fill_2 FILLER_12_2043 ();
 sg13g2_fill_1 FILLER_12_2045 ();
 sg13g2_fill_1 FILLER_12_2063 ();
 sg13g2_fill_1 FILLER_12_2068 ();
 sg13g2_fill_1 FILLER_12_2109 ();
 sg13g2_fill_2 FILLER_12_2158 ();
 sg13g2_fill_1 FILLER_12_2178 ();
 sg13g2_fill_2 FILLER_12_2188 ();
 sg13g2_fill_1 FILLER_12_2195 ();
 sg13g2_fill_2 FILLER_12_2209 ();
 sg13g2_fill_2 FILLER_12_2225 ();
 sg13g2_fill_1 FILLER_12_2253 ();
 sg13g2_fill_2 FILLER_12_2266 ();
 sg13g2_fill_1 FILLER_12_2268 ();
 sg13g2_fill_2 FILLER_12_2310 ();
 sg13g2_fill_1 FILLER_12_2333 ();
 sg13g2_decap_8 FILLER_12_2360 ();
 sg13g2_decap_8 FILLER_12_2367 ();
 sg13g2_decap_8 FILLER_12_2374 ();
 sg13g2_decap_8 FILLER_12_2381 ();
 sg13g2_decap_8 FILLER_12_2388 ();
 sg13g2_decap_8 FILLER_12_2395 ();
 sg13g2_decap_8 FILLER_12_2402 ();
 sg13g2_decap_8 FILLER_12_2409 ();
 sg13g2_decap_8 FILLER_12_2416 ();
 sg13g2_decap_8 FILLER_12_2423 ();
 sg13g2_decap_8 FILLER_12_2430 ();
 sg13g2_decap_8 FILLER_12_2437 ();
 sg13g2_decap_8 FILLER_12_2444 ();
 sg13g2_decap_8 FILLER_12_2451 ();
 sg13g2_decap_8 FILLER_12_2458 ();
 sg13g2_decap_8 FILLER_12_2465 ();
 sg13g2_decap_8 FILLER_12_2472 ();
 sg13g2_decap_8 FILLER_12_2479 ();
 sg13g2_decap_8 FILLER_12_2486 ();
 sg13g2_decap_8 FILLER_12_2493 ();
 sg13g2_decap_8 FILLER_12_2500 ();
 sg13g2_decap_8 FILLER_12_2507 ();
 sg13g2_decap_8 FILLER_12_2514 ();
 sg13g2_decap_8 FILLER_12_2521 ();
 sg13g2_decap_8 FILLER_12_2528 ();
 sg13g2_decap_8 FILLER_12_2535 ();
 sg13g2_decap_8 FILLER_12_2542 ();
 sg13g2_decap_8 FILLER_12_2549 ();
 sg13g2_decap_8 FILLER_12_2556 ();
 sg13g2_decap_8 FILLER_12_2563 ();
 sg13g2_decap_8 FILLER_12_2570 ();
 sg13g2_decap_8 FILLER_12_2577 ();
 sg13g2_decap_8 FILLER_12_2584 ();
 sg13g2_decap_8 FILLER_12_2591 ();
 sg13g2_decap_8 FILLER_12_2598 ();
 sg13g2_decap_8 FILLER_12_2605 ();
 sg13g2_decap_8 FILLER_12_2612 ();
 sg13g2_decap_8 FILLER_12_2619 ();
 sg13g2_decap_8 FILLER_12_2626 ();
 sg13g2_decap_8 FILLER_12_2633 ();
 sg13g2_decap_8 FILLER_12_2640 ();
 sg13g2_decap_8 FILLER_12_2647 ();
 sg13g2_decap_8 FILLER_12_2654 ();
 sg13g2_decap_8 FILLER_12_2661 ();
 sg13g2_decap_4 FILLER_12_2668 ();
 sg13g2_fill_2 FILLER_12_2672 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_1 FILLER_13_427 ();
 sg13g2_fill_2 FILLER_13_445 ();
 sg13g2_fill_1 FILLER_13_447 ();
 sg13g2_fill_2 FILLER_13_500 ();
 sg13g2_fill_1 FILLER_13_528 ();
 sg13g2_fill_2 FILLER_13_574 ();
 sg13g2_decap_4 FILLER_13_602 ();
 sg13g2_fill_1 FILLER_13_606 ();
 sg13g2_fill_1 FILLER_13_620 ();
 sg13g2_fill_2 FILLER_13_626 ();
 sg13g2_fill_1 FILLER_13_628 ();
 sg13g2_fill_2 FILLER_13_668 ();
 sg13g2_fill_2 FILLER_13_675 ();
 sg13g2_fill_1 FILLER_13_703 ();
 sg13g2_decap_4 FILLER_13_709 ();
 sg13g2_fill_1 FILLER_13_757 ();
 sg13g2_fill_1 FILLER_13_767 ();
 sg13g2_fill_1 FILLER_13_795 ();
 sg13g2_fill_2 FILLER_13_801 ();
 sg13g2_fill_2 FILLER_13_821 ();
 sg13g2_fill_1 FILLER_13_827 ();
 sg13g2_fill_2 FILLER_13_841 ();
 sg13g2_fill_1 FILLER_13_843 ();
 sg13g2_fill_2 FILLER_13_857 ();
 sg13g2_fill_1 FILLER_13_859 ();
 sg13g2_fill_2 FILLER_13_900 ();
 sg13g2_fill_1 FILLER_13_915 ();
 sg13g2_fill_1 FILLER_13_938 ();
 sg13g2_fill_1 FILLER_13_1039 ();
 sg13g2_fill_2 FILLER_13_1053 ();
 sg13g2_fill_1 FILLER_13_1060 ();
 sg13g2_fill_1 FILLER_13_1165 ();
 sg13g2_fill_1 FILLER_13_1249 ();
 sg13g2_fill_1 FILLER_13_1286 ();
 sg13g2_fill_2 FILLER_13_1345 ();
 sg13g2_decap_4 FILLER_13_1416 ();
 sg13g2_fill_1 FILLER_13_1420 ();
 sg13g2_fill_2 FILLER_13_1429 ();
 sg13g2_fill_1 FILLER_13_1440 ();
 sg13g2_fill_2 FILLER_13_1485 ();
 sg13g2_fill_1 FILLER_13_1547 ();
 sg13g2_fill_1 FILLER_13_1566 ();
 sg13g2_fill_1 FILLER_13_1603 ();
 sg13g2_fill_2 FILLER_13_1664 ();
 sg13g2_fill_1 FILLER_13_1666 ();
 sg13g2_fill_1 FILLER_13_1671 ();
 sg13g2_fill_2 FILLER_13_1681 ();
 sg13g2_fill_1 FILLER_13_1683 ();
 sg13g2_fill_2 FILLER_13_1755 ();
 sg13g2_fill_1 FILLER_13_1757 ();
 sg13g2_fill_2 FILLER_13_1784 ();
 sg13g2_fill_2 FILLER_13_1790 ();
 sg13g2_fill_2 FILLER_13_1831 ();
 sg13g2_fill_1 FILLER_13_1833 ();
 sg13g2_fill_1 FILLER_13_1838 ();
 sg13g2_fill_2 FILLER_13_1844 ();
 sg13g2_fill_1 FILLER_13_1846 ();
 sg13g2_fill_2 FILLER_13_1870 ();
 sg13g2_fill_1 FILLER_13_1872 ();
 sg13g2_fill_2 FILLER_13_1887 ();
 sg13g2_fill_1 FILLER_13_1889 ();
 sg13g2_decap_4 FILLER_13_1942 ();
 sg13g2_fill_1 FILLER_13_1946 ();
 sg13g2_decap_4 FILLER_13_1951 ();
 sg13g2_fill_1 FILLER_13_1955 ();
 sg13g2_fill_2 FILLER_13_1981 ();
 sg13g2_fill_2 FILLER_13_1987 ();
 sg13g2_fill_1 FILLER_13_1989 ();
 sg13g2_fill_2 FILLER_13_2007 ();
 sg13g2_fill_2 FILLER_13_2028 ();
 sg13g2_fill_1 FILLER_13_2030 ();
 sg13g2_fill_2 FILLER_13_2041 ();
 sg13g2_fill_1 FILLER_13_2052 ();
 sg13g2_fill_2 FILLER_13_2083 ();
 sg13g2_decap_4 FILLER_13_2098 ();
 sg13g2_fill_2 FILLER_13_2111 ();
 sg13g2_fill_1 FILLER_13_2129 ();
 sg13g2_fill_1 FILLER_13_2183 ();
 sg13g2_fill_2 FILLER_13_2189 ();
 sg13g2_fill_1 FILLER_13_2191 ();
 sg13g2_fill_2 FILLER_13_2205 ();
 sg13g2_fill_1 FILLER_13_2216 ();
 sg13g2_fill_1 FILLER_13_2222 ();
 sg13g2_fill_2 FILLER_13_2228 ();
 sg13g2_fill_2 FILLER_13_2247 ();
 sg13g2_fill_2 FILLER_13_2291 ();
 sg13g2_fill_2 FILLER_13_2342 ();
 sg13g2_fill_1 FILLER_13_2344 ();
 sg13g2_decap_8 FILLER_13_2367 ();
 sg13g2_decap_8 FILLER_13_2374 ();
 sg13g2_decap_8 FILLER_13_2381 ();
 sg13g2_decap_8 FILLER_13_2388 ();
 sg13g2_decap_8 FILLER_13_2395 ();
 sg13g2_decap_8 FILLER_13_2402 ();
 sg13g2_decap_8 FILLER_13_2409 ();
 sg13g2_decap_8 FILLER_13_2416 ();
 sg13g2_decap_8 FILLER_13_2423 ();
 sg13g2_decap_8 FILLER_13_2430 ();
 sg13g2_decap_8 FILLER_13_2437 ();
 sg13g2_decap_8 FILLER_13_2444 ();
 sg13g2_decap_8 FILLER_13_2451 ();
 sg13g2_decap_8 FILLER_13_2458 ();
 sg13g2_decap_8 FILLER_13_2465 ();
 sg13g2_decap_8 FILLER_13_2472 ();
 sg13g2_decap_8 FILLER_13_2479 ();
 sg13g2_decap_8 FILLER_13_2486 ();
 sg13g2_decap_8 FILLER_13_2493 ();
 sg13g2_decap_8 FILLER_13_2500 ();
 sg13g2_decap_8 FILLER_13_2507 ();
 sg13g2_decap_8 FILLER_13_2514 ();
 sg13g2_decap_8 FILLER_13_2521 ();
 sg13g2_decap_8 FILLER_13_2528 ();
 sg13g2_decap_8 FILLER_13_2535 ();
 sg13g2_decap_8 FILLER_13_2542 ();
 sg13g2_decap_8 FILLER_13_2549 ();
 sg13g2_decap_8 FILLER_13_2556 ();
 sg13g2_decap_8 FILLER_13_2563 ();
 sg13g2_decap_8 FILLER_13_2570 ();
 sg13g2_decap_8 FILLER_13_2577 ();
 sg13g2_decap_8 FILLER_13_2584 ();
 sg13g2_decap_8 FILLER_13_2591 ();
 sg13g2_decap_8 FILLER_13_2598 ();
 sg13g2_decap_8 FILLER_13_2605 ();
 sg13g2_decap_8 FILLER_13_2612 ();
 sg13g2_decap_8 FILLER_13_2619 ();
 sg13g2_decap_8 FILLER_13_2626 ();
 sg13g2_decap_8 FILLER_13_2633 ();
 sg13g2_decap_8 FILLER_13_2640 ();
 sg13g2_decap_8 FILLER_13_2647 ();
 sg13g2_decap_8 FILLER_13_2654 ();
 sg13g2_decap_8 FILLER_13_2661 ();
 sg13g2_decap_4 FILLER_13_2668 ();
 sg13g2_fill_2 FILLER_13_2672 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_4 FILLER_14_420 ();
 sg13g2_fill_1 FILLER_14_424 ();
 sg13g2_fill_1 FILLER_14_468 ();
 sg13g2_decap_8 FILLER_14_478 ();
 sg13g2_decap_8 FILLER_14_485 ();
 sg13g2_decap_8 FILLER_14_501 ();
 sg13g2_fill_2 FILLER_14_508 ();
 sg13g2_fill_1 FILLER_14_515 ();
 sg13g2_fill_2 FILLER_14_537 ();
 sg13g2_fill_2 FILLER_14_544 ();
 sg13g2_fill_1 FILLER_14_546 ();
 sg13g2_fill_1 FILLER_14_586 ();
 sg13g2_fill_1 FILLER_14_591 ();
 sg13g2_fill_2 FILLER_14_636 ();
 sg13g2_decap_4 FILLER_14_673 ();
 sg13g2_fill_2 FILLER_14_686 ();
 sg13g2_fill_1 FILLER_14_688 ();
 sg13g2_fill_1 FILLER_14_737 ();
 sg13g2_fill_2 FILLER_14_747 ();
 sg13g2_fill_1 FILLER_14_749 ();
 sg13g2_fill_2 FILLER_14_758 ();
 sg13g2_fill_1 FILLER_14_863 ();
 sg13g2_decap_4 FILLER_14_890 ();
 sg13g2_fill_1 FILLER_14_923 ();
 sg13g2_fill_2 FILLER_14_929 ();
 sg13g2_fill_1 FILLER_14_945 ();
 sg13g2_fill_2 FILLER_14_972 ();
 sg13g2_fill_1 FILLER_14_1017 ();
 sg13g2_fill_2 FILLER_14_1043 ();
 sg13g2_fill_2 FILLER_14_1100 ();
 sg13g2_fill_1 FILLER_14_1102 ();
 sg13g2_decap_8 FILLER_14_1124 ();
 sg13g2_decap_4 FILLER_14_1131 ();
 sg13g2_fill_2 FILLER_14_1183 ();
 sg13g2_fill_2 FILLER_14_1190 ();
 sg13g2_fill_1 FILLER_14_1192 ();
 sg13g2_fill_1 FILLER_14_1198 ();
 sg13g2_fill_2 FILLER_14_1212 ();
 sg13g2_fill_1 FILLER_14_1214 ();
 sg13g2_decap_4 FILLER_14_1238 ();
 sg13g2_fill_1 FILLER_14_1242 ();
 sg13g2_fill_2 FILLER_14_1287 ();
 sg13g2_fill_1 FILLER_14_1289 ();
 sg13g2_decap_4 FILLER_14_1317 ();
 sg13g2_fill_1 FILLER_14_1321 ();
 sg13g2_fill_2 FILLER_14_1373 ();
 sg13g2_fill_1 FILLER_14_1375 ();
 sg13g2_fill_2 FILLER_14_1429 ();
 sg13g2_fill_1 FILLER_14_1431 ();
 sg13g2_fill_1 FILLER_14_1467 ();
 sg13g2_fill_1 FILLER_14_1481 ();
 sg13g2_fill_1 FILLER_14_1487 ();
 sg13g2_fill_2 FILLER_14_1498 ();
 sg13g2_fill_2 FILLER_14_1509 ();
 sg13g2_fill_1 FILLER_14_1516 ();
 sg13g2_decap_4 FILLER_14_1545 ();
 sg13g2_decap_4 FILLER_14_1558 ();
 sg13g2_fill_1 FILLER_14_1562 ();
 sg13g2_fill_2 FILLER_14_1590 ();
 sg13g2_fill_1 FILLER_14_1592 ();
 sg13g2_fill_1 FILLER_14_1602 ();
 sg13g2_fill_2 FILLER_14_1613 ();
 sg13g2_fill_2 FILLER_14_1629 ();
 sg13g2_fill_1 FILLER_14_1648 ();
 sg13g2_fill_1 FILLER_14_1672 ();
 sg13g2_fill_1 FILLER_14_1683 ();
 sg13g2_fill_1 FILLER_14_1706 ();
 sg13g2_decap_4 FILLER_14_1732 ();
 sg13g2_fill_2 FILLER_14_1746 ();
 sg13g2_fill_1 FILLER_14_1748 ();
 sg13g2_fill_1 FILLER_14_1754 ();
 sg13g2_decap_4 FILLER_14_1760 ();
 sg13g2_fill_1 FILLER_14_1764 ();
 sg13g2_fill_2 FILLER_14_1773 ();
 sg13g2_fill_1 FILLER_14_1804 ();
 sg13g2_fill_1 FILLER_14_1809 ();
 sg13g2_fill_1 FILLER_14_1849 ();
 sg13g2_fill_2 FILLER_14_1959 ();
 sg13g2_fill_1 FILLER_14_1961 ();
 sg13g2_decap_4 FILLER_14_1993 ();
 sg13g2_fill_1 FILLER_14_2018 ();
 sg13g2_fill_2 FILLER_14_2062 ();
 sg13g2_fill_2 FILLER_14_2099 ();
 sg13g2_fill_1 FILLER_14_2101 ();
 sg13g2_fill_2 FILLER_14_2111 ();
 sg13g2_fill_1 FILLER_14_2129 ();
 sg13g2_fill_1 FILLER_14_2161 ();
 sg13g2_fill_2 FILLER_14_2167 ();
 sg13g2_fill_1 FILLER_14_2169 ();
 sg13g2_decap_8 FILLER_14_2182 ();
 sg13g2_fill_2 FILLER_14_2269 ();
 sg13g2_fill_1 FILLER_14_2271 ();
 sg13g2_fill_2 FILLER_14_2298 ();
 sg13g2_decap_8 FILLER_14_2313 ();
 sg13g2_fill_1 FILLER_14_2320 ();
 sg13g2_fill_1 FILLER_14_2337 ();
 sg13g2_decap_8 FILLER_14_2364 ();
 sg13g2_decap_8 FILLER_14_2371 ();
 sg13g2_decap_8 FILLER_14_2378 ();
 sg13g2_decap_8 FILLER_14_2385 ();
 sg13g2_decap_8 FILLER_14_2392 ();
 sg13g2_decap_8 FILLER_14_2399 ();
 sg13g2_decap_8 FILLER_14_2406 ();
 sg13g2_decap_8 FILLER_14_2413 ();
 sg13g2_decap_8 FILLER_14_2420 ();
 sg13g2_decap_8 FILLER_14_2427 ();
 sg13g2_decap_8 FILLER_14_2434 ();
 sg13g2_decap_8 FILLER_14_2441 ();
 sg13g2_decap_8 FILLER_14_2448 ();
 sg13g2_decap_8 FILLER_14_2455 ();
 sg13g2_decap_8 FILLER_14_2462 ();
 sg13g2_decap_8 FILLER_14_2469 ();
 sg13g2_decap_8 FILLER_14_2476 ();
 sg13g2_decap_8 FILLER_14_2483 ();
 sg13g2_decap_8 FILLER_14_2490 ();
 sg13g2_decap_8 FILLER_14_2497 ();
 sg13g2_decap_8 FILLER_14_2504 ();
 sg13g2_decap_8 FILLER_14_2511 ();
 sg13g2_decap_8 FILLER_14_2518 ();
 sg13g2_decap_8 FILLER_14_2525 ();
 sg13g2_decap_8 FILLER_14_2532 ();
 sg13g2_decap_8 FILLER_14_2539 ();
 sg13g2_decap_8 FILLER_14_2546 ();
 sg13g2_decap_8 FILLER_14_2553 ();
 sg13g2_decap_8 FILLER_14_2560 ();
 sg13g2_decap_8 FILLER_14_2567 ();
 sg13g2_decap_8 FILLER_14_2574 ();
 sg13g2_decap_8 FILLER_14_2581 ();
 sg13g2_decap_8 FILLER_14_2588 ();
 sg13g2_decap_8 FILLER_14_2595 ();
 sg13g2_decap_8 FILLER_14_2602 ();
 sg13g2_decap_8 FILLER_14_2609 ();
 sg13g2_decap_8 FILLER_14_2616 ();
 sg13g2_decap_8 FILLER_14_2623 ();
 sg13g2_decap_8 FILLER_14_2630 ();
 sg13g2_decap_8 FILLER_14_2637 ();
 sg13g2_decap_8 FILLER_14_2644 ();
 sg13g2_decap_8 FILLER_14_2651 ();
 sg13g2_decap_8 FILLER_14_2658 ();
 sg13g2_decap_8 FILLER_14_2665 ();
 sg13g2_fill_2 FILLER_14_2672 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_fill_2 FILLER_15_459 ();
 sg13g2_fill_1 FILLER_15_475 ();
 sg13g2_fill_2 FILLER_15_551 ();
 sg13g2_fill_1 FILLER_15_553 ();
 sg13g2_fill_1 FILLER_15_567 ();
 sg13g2_fill_2 FILLER_15_582 ();
 sg13g2_decap_4 FILLER_15_605 ();
 sg13g2_fill_1 FILLER_15_645 ();
 sg13g2_decap_8 FILLER_15_668 ();
 sg13g2_fill_1 FILLER_15_675 ();
 sg13g2_fill_2 FILLER_15_723 ();
 sg13g2_fill_2 FILLER_15_739 ();
 sg13g2_fill_1 FILLER_15_741 ();
 sg13g2_fill_2 FILLER_15_750 ();
 sg13g2_fill_2 FILLER_15_757 ();
 sg13g2_fill_2 FILLER_15_764 ();
 sg13g2_fill_1 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_779 ();
 sg13g2_decap_4 FILLER_15_786 ();
 sg13g2_decap_4 FILLER_15_798 ();
 sg13g2_fill_1 FILLER_15_802 ();
 sg13g2_fill_2 FILLER_15_834 ();
 sg13g2_fill_2 FILLER_15_849 ();
 sg13g2_decap_8 FILLER_15_856 ();
 sg13g2_fill_2 FILLER_15_863 ();
 sg13g2_fill_2 FILLER_15_883 ();
 sg13g2_fill_1 FILLER_15_894 ();
 sg13g2_decap_4 FILLER_15_920 ();
 sg13g2_decap_4 FILLER_15_954 ();
 sg13g2_fill_2 FILLER_15_958 ();
 sg13g2_fill_2 FILLER_15_1048 ();
 sg13g2_fill_1 FILLER_15_1050 ();
 sg13g2_fill_2 FILLER_15_1060 ();
 sg13g2_fill_1 FILLER_15_1062 ();
 sg13g2_fill_1 FILLER_15_1070 ();
 sg13g2_fill_2 FILLER_15_1102 ();
 sg13g2_fill_1 FILLER_15_1104 ();
 sg13g2_decap_4 FILLER_15_1118 ();
 sg13g2_fill_2 FILLER_15_1156 ();
 sg13g2_decap_4 FILLER_15_1220 ();
 sg13g2_fill_2 FILLER_15_1224 ();
 sg13g2_fill_2 FILLER_15_1252 ();
 sg13g2_fill_1 FILLER_15_1254 ();
 sg13g2_fill_1 FILLER_15_1281 ();
 sg13g2_fill_1 FILLER_15_1322 ();
 sg13g2_fill_1 FILLER_15_1331 ();
 sg13g2_decap_8 FILLER_15_1336 ();
 sg13g2_fill_2 FILLER_15_1343 ();
 sg13g2_fill_1 FILLER_15_1350 ();
 sg13g2_fill_1 FILLER_15_1399 ();
 sg13g2_decap_4 FILLER_15_1450 ();
 sg13g2_fill_1 FILLER_15_1466 ();
 sg13g2_fill_2 FILLER_15_1489 ();
 sg13g2_fill_2 FILLER_15_1529 ();
 sg13g2_fill_1 FILLER_15_1531 ();
 sg13g2_fill_2 FILLER_15_1614 ();
 sg13g2_fill_1 FILLER_15_1616 ();
 sg13g2_fill_2 FILLER_15_1648 ();
 sg13g2_fill_1 FILLER_15_1650 ();
 sg13g2_fill_1 FILLER_15_1706 ();
 sg13g2_fill_2 FILLER_15_1725 ();
 sg13g2_fill_2 FILLER_15_1732 ();
 sg13g2_fill_1 FILLER_15_1734 ();
 sg13g2_fill_2 FILLER_15_1757 ();
 sg13g2_fill_2 FILLER_15_1772 ();
 sg13g2_fill_1 FILLER_15_1774 ();
 sg13g2_fill_2 FILLER_15_1790 ();
 sg13g2_decap_4 FILLER_15_1827 ();
 sg13g2_fill_1 FILLER_15_1838 ();
 sg13g2_fill_2 FILLER_15_1864 ();
 sg13g2_fill_2 FILLER_15_1870 ();
 sg13g2_fill_1 FILLER_15_1872 ();
 sg13g2_decap_4 FILLER_15_1933 ();
 sg13g2_fill_1 FILLER_15_1990 ();
 sg13g2_fill_1 FILLER_15_1996 ();
 sg13g2_decap_8 FILLER_15_2049 ();
 sg13g2_fill_1 FILLER_15_2056 ();
 sg13g2_fill_2 FILLER_15_2118 ();
 sg13g2_decap_8 FILLER_15_2124 ();
 sg13g2_fill_2 FILLER_15_2131 ();
 sg13g2_fill_2 FILLER_15_2211 ();
 sg13g2_fill_1 FILLER_15_2213 ();
 sg13g2_fill_2 FILLER_15_2223 ();
 sg13g2_fill_2 FILLER_15_2243 ();
 sg13g2_fill_2 FILLER_15_2249 ();
 sg13g2_fill_2 FILLER_15_2265 ();
 sg13g2_fill_1 FILLER_15_2267 ();
 sg13g2_fill_2 FILLER_15_2282 ();
 sg13g2_fill_1 FILLER_15_2284 ();
 sg13g2_fill_2 FILLER_15_2308 ();
 sg13g2_fill_1 FILLER_15_2310 ();
 sg13g2_fill_2 FILLER_15_2319 ();
 sg13g2_fill_1 FILLER_15_2321 ();
 sg13g2_decap_8 FILLER_15_2335 ();
 sg13g2_fill_1 FILLER_15_2342 ();
 sg13g2_decap_8 FILLER_15_2360 ();
 sg13g2_decap_8 FILLER_15_2367 ();
 sg13g2_decap_8 FILLER_15_2374 ();
 sg13g2_decap_8 FILLER_15_2381 ();
 sg13g2_decap_8 FILLER_15_2388 ();
 sg13g2_decap_8 FILLER_15_2395 ();
 sg13g2_decap_8 FILLER_15_2402 ();
 sg13g2_decap_8 FILLER_15_2409 ();
 sg13g2_decap_8 FILLER_15_2416 ();
 sg13g2_decap_8 FILLER_15_2423 ();
 sg13g2_decap_8 FILLER_15_2430 ();
 sg13g2_decap_8 FILLER_15_2437 ();
 sg13g2_decap_8 FILLER_15_2444 ();
 sg13g2_decap_8 FILLER_15_2451 ();
 sg13g2_decap_8 FILLER_15_2458 ();
 sg13g2_decap_8 FILLER_15_2465 ();
 sg13g2_decap_8 FILLER_15_2472 ();
 sg13g2_decap_8 FILLER_15_2479 ();
 sg13g2_decap_8 FILLER_15_2486 ();
 sg13g2_decap_8 FILLER_15_2493 ();
 sg13g2_decap_8 FILLER_15_2500 ();
 sg13g2_decap_8 FILLER_15_2507 ();
 sg13g2_decap_8 FILLER_15_2514 ();
 sg13g2_decap_8 FILLER_15_2521 ();
 sg13g2_decap_8 FILLER_15_2528 ();
 sg13g2_decap_8 FILLER_15_2535 ();
 sg13g2_decap_8 FILLER_15_2542 ();
 sg13g2_decap_8 FILLER_15_2549 ();
 sg13g2_decap_8 FILLER_15_2556 ();
 sg13g2_decap_8 FILLER_15_2563 ();
 sg13g2_decap_8 FILLER_15_2570 ();
 sg13g2_decap_8 FILLER_15_2577 ();
 sg13g2_decap_8 FILLER_15_2584 ();
 sg13g2_decap_8 FILLER_15_2591 ();
 sg13g2_decap_8 FILLER_15_2598 ();
 sg13g2_decap_8 FILLER_15_2605 ();
 sg13g2_decap_8 FILLER_15_2612 ();
 sg13g2_decap_8 FILLER_15_2619 ();
 sg13g2_decap_8 FILLER_15_2626 ();
 sg13g2_decap_8 FILLER_15_2633 ();
 sg13g2_decap_8 FILLER_15_2640 ();
 sg13g2_decap_8 FILLER_15_2647 ();
 sg13g2_decap_8 FILLER_15_2654 ();
 sg13g2_decap_8 FILLER_15_2661 ();
 sg13g2_decap_4 FILLER_15_2668 ();
 sg13g2_fill_2 FILLER_15_2672 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_fill_2 FILLER_16_460 ();
 sg13g2_fill_2 FILLER_16_497 ();
 sg13g2_fill_1 FILLER_16_508 ();
 sg13g2_fill_2 FILLER_16_535 ();
 sg13g2_fill_1 FILLER_16_537 ();
 sg13g2_fill_1 FILLER_16_547 ();
 sg13g2_fill_2 FILLER_16_605 ();
 sg13g2_fill_2 FILLER_16_613 ();
 sg13g2_fill_2 FILLER_16_632 ();
 sg13g2_fill_1 FILLER_16_634 ();
 sg13g2_fill_1 FILLER_16_692 ();
 sg13g2_fill_2 FILLER_16_711 ();
 sg13g2_fill_1 FILLER_16_713 ();
 sg13g2_fill_2 FILLER_16_752 ();
 sg13g2_fill_2 FILLER_16_797 ();
 sg13g2_fill_2 FILLER_16_804 ();
 sg13g2_fill_1 FILLER_16_818 ();
 sg13g2_decap_4 FILLER_16_900 ();
 sg13g2_decap_8 FILLER_16_913 ();
 sg13g2_decap_8 FILLER_16_924 ();
 sg13g2_fill_2 FILLER_16_931 ();
 sg13g2_fill_2 FILLER_16_938 ();
 sg13g2_decap_4 FILLER_16_976 ();
 sg13g2_fill_1 FILLER_16_980 ();
 sg13g2_fill_2 FILLER_16_985 ();
 sg13g2_fill_1 FILLER_16_987 ();
 sg13g2_fill_2 FILLER_16_1028 ();
 sg13g2_fill_1 FILLER_16_1043 ();
 sg13g2_fill_1 FILLER_16_1140 ();
 sg13g2_fill_2 FILLER_16_1149 ();
 sg13g2_fill_2 FILLER_16_1160 ();
 sg13g2_fill_1 FILLER_16_1162 ();
 sg13g2_decap_8 FILLER_16_1193 ();
 sg13g2_decap_4 FILLER_16_1200 ();
 sg13g2_fill_1 FILLER_16_1225 ();
 sg13g2_fill_1 FILLER_16_1265 ();
 sg13g2_fill_1 FILLER_16_1270 ();
 sg13g2_fill_2 FILLER_16_1276 ();
 sg13g2_decap_4 FILLER_16_1287 ();
 sg13g2_fill_2 FILLER_16_1295 ();
 sg13g2_fill_1 FILLER_16_1297 ();
 sg13g2_fill_1 FILLER_16_1302 ();
 sg13g2_decap_8 FILLER_16_1319 ();
 sg13g2_decap_4 FILLER_16_1335 ();
 sg13g2_fill_2 FILLER_16_1339 ();
 sg13g2_fill_2 FILLER_16_1381 ();
 sg13g2_fill_1 FILLER_16_1383 ();
 sg13g2_fill_2 FILLER_16_1435 ();
 sg13g2_fill_2 FILLER_16_1472 ();
 sg13g2_fill_1 FILLER_16_1474 ();
 sg13g2_fill_1 FILLER_16_1505 ();
 sg13g2_decap_4 FILLER_16_1523 ();
 sg13g2_fill_2 FILLER_16_1527 ();
 sg13g2_fill_2 FILLER_16_1534 ();
 sg13g2_fill_2 FILLER_16_1540 ();
 sg13g2_fill_1 FILLER_16_1542 ();
 sg13g2_fill_2 FILLER_16_1556 ();
 sg13g2_fill_1 FILLER_16_1558 ();
 sg13g2_decap_8 FILLER_16_1577 ();
 sg13g2_fill_2 FILLER_16_1584 ();
 sg13g2_fill_2 FILLER_16_1599 ();
 sg13g2_fill_1 FILLER_16_1601 ();
 sg13g2_fill_2 FILLER_16_1625 ();
 sg13g2_decap_8 FILLER_16_1637 ();
 sg13g2_decap_4 FILLER_16_1644 ();
 sg13g2_fill_1 FILLER_16_1648 ();
 sg13g2_fill_2 FILLER_16_1658 ();
 sg13g2_fill_1 FILLER_16_1660 ();
 sg13g2_fill_2 FILLER_16_1683 ();
 sg13g2_fill_1 FILLER_16_1685 ();
 sg13g2_decap_8 FILLER_16_1691 ();
 sg13g2_fill_2 FILLER_16_1698 ();
 sg13g2_fill_1 FILLER_16_1700 ();
 sg13g2_fill_1 FILLER_16_1792 ();
 sg13g2_fill_2 FILLER_16_1807 ();
 sg13g2_fill_2 FILLER_16_1813 ();
 sg13g2_fill_1 FILLER_16_1815 ();
 sg13g2_fill_1 FILLER_16_1837 ();
 sg13g2_fill_2 FILLER_16_1845 ();
 sg13g2_fill_2 FILLER_16_1852 ();
 sg13g2_fill_2 FILLER_16_1885 ();
 sg13g2_fill_2 FILLER_16_1895 ();
 sg13g2_fill_2 FILLER_16_1911 ();
 sg13g2_fill_1 FILLER_16_1927 ();
 sg13g2_fill_2 FILLER_16_1937 ();
 sg13g2_fill_1 FILLER_16_1939 ();
 sg13g2_decap_8 FILLER_16_1945 ();
 sg13g2_decap_8 FILLER_16_1952 ();
 sg13g2_fill_2 FILLER_16_1959 ();
 sg13g2_decap_8 FILLER_16_1981 ();
 sg13g2_decap_4 FILLER_16_1988 ();
 sg13g2_fill_2 FILLER_16_2000 ();
 sg13g2_fill_2 FILLER_16_2006 ();
 sg13g2_decap_4 FILLER_16_2012 ();
 sg13g2_fill_1 FILLER_16_2030 ();
 sg13g2_fill_1 FILLER_16_2057 ();
 sg13g2_fill_1 FILLER_16_2066 ();
 sg13g2_fill_2 FILLER_16_2076 ();
 sg13g2_fill_1 FILLER_16_2078 ();
 sg13g2_fill_2 FILLER_16_2092 ();
 sg13g2_fill_2 FILLER_16_2111 ();
 sg13g2_fill_1 FILLER_16_2113 ();
 sg13g2_fill_2 FILLER_16_2119 ();
 sg13g2_fill_2 FILLER_16_2178 ();
 sg13g2_fill_1 FILLER_16_2194 ();
 sg13g2_fill_2 FILLER_16_2221 ();
 sg13g2_fill_1 FILLER_16_2223 ();
 sg13g2_decap_4 FILLER_16_2250 ();
 sg13g2_fill_1 FILLER_16_2269 ();
 sg13g2_decap_8 FILLER_16_2301 ();
 sg13g2_decap_4 FILLER_16_2312 ();
 sg13g2_fill_1 FILLER_16_2316 ();
 sg13g2_fill_2 FILLER_16_2325 ();
 sg13g2_fill_1 FILLER_16_2327 ();
 sg13g2_decap_8 FILLER_16_2363 ();
 sg13g2_decap_8 FILLER_16_2370 ();
 sg13g2_decap_8 FILLER_16_2377 ();
 sg13g2_decap_8 FILLER_16_2384 ();
 sg13g2_decap_8 FILLER_16_2391 ();
 sg13g2_decap_8 FILLER_16_2398 ();
 sg13g2_decap_8 FILLER_16_2405 ();
 sg13g2_decap_8 FILLER_16_2412 ();
 sg13g2_decap_8 FILLER_16_2419 ();
 sg13g2_decap_8 FILLER_16_2426 ();
 sg13g2_decap_8 FILLER_16_2433 ();
 sg13g2_decap_8 FILLER_16_2440 ();
 sg13g2_decap_8 FILLER_16_2447 ();
 sg13g2_decap_8 FILLER_16_2454 ();
 sg13g2_decap_8 FILLER_16_2461 ();
 sg13g2_decap_8 FILLER_16_2468 ();
 sg13g2_decap_8 FILLER_16_2475 ();
 sg13g2_decap_8 FILLER_16_2482 ();
 sg13g2_decap_8 FILLER_16_2489 ();
 sg13g2_decap_8 FILLER_16_2496 ();
 sg13g2_decap_8 FILLER_16_2503 ();
 sg13g2_decap_8 FILLER_16_2510 ();
 sg13g2_decap_8 FILLER_16_2517 ();
 sg13g2_decap_8 FILLER_16_2524 ();
 sg13g2_decap_8 FILLER_16_2531 ();
 sg13g2_decap_8 FILLER_16_2538 ();
 sg13g2_decap_8 FILLER_16_2545 ();
 sg13g2_decap_8 FILLER_16_2552 ();
 sg13g2_decap_8 FILLER_16_2559 ();
 sg13g2_decap_8 FILLER_16_2566 ();
 sg13g2_decap_8 FILLER_16_2573 ();
 sg13g2_decap_8 FILLER_16_2580 ();
 sg13g2_decap_8 FILLER_16_2587 ();
 sg13g2_decap_8 FILLER_16_2594 ();
 sg13g2_decap_8 FILLER_16_2601 ();
 sg13g2_decap_8 FILLER_16_2608 ();
 sg13g2_decap_8 FILLER_16_2615 ();
 sg13g2_decap_8 FILLER_16_2622 ();
 sg13g2_decap_8 FILLER_16_2629 ();
 sg13g2_decap_8 FILLER_16_2636 ();
 sg13g2_decap_8 FILLER_16_2643 ();
 sg13g2_decap_8 FILLER_16_2650 ();
 sg13g2_decap_8 FILLER_16_2657 ();
 sg13g2_decap_8 FILLER_16_2664 ();
 sg13g2_fill_2 FILLER_16_2671 ();
 sg13g2_fill_1 FILLER_16_2673 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_4 FILLER_17_420 ();
 sg13g2_fill_1 FILLER_17_480 ();
 sg13g2_fill_2 FILLER_17_485 ();
 sg13g2_fill_2 FILLER_17_496 ();
 sg13g2_fill_1 FILLER_17_498 ();
 sg13g2_fill_1 FILLER_17_547 ();
 sg13g2_fill_2 FILLER_17_552 ();
 sg13g2_fill_1 FILLER_17_554 ();
 sg13g2_fill_2 FILLER_17_563 ();
 sg13g2_decap_4 FILLER_17_569 ();
 sg13g2_decap_4 FILLER_17_582 ();
 sg13g2_fill_2 FILLER_17_586 ();
 sg13g2_decap_4 FILLER_17_601 ();
 sg13g2_fill_2 FILLER_17_605 ();
 sg13g2_fill_2 FILLER_17_619 ();
 sg13g2_fill_1 FILLER_17_621 ();
 sg13g2_fill_2 FILLER_17_635 ();
 sg13g2_fill_1 FILLER_17_637 ();
 sg13g2_fill_2 FILLER_17_651 ();
 sg13g2_decap_4 FILLER_17_717 ();
 sg13g2_fill_1 FILLER_17_721 ();
 sg13g2_decap_4 FILLER_17_727 ();
 sg13g2_fill_1 FILLER_17_731 ();
 sg13g2_fill_2 FILLER_17_740 ();
 sg13g2_decap_4 FILLER_17_747 ();
 sg13g2_fill_1 FILLER_17_751 ();
 sg13g2_fill_1 FILLER_17_761 ();
 sg13g2_fill_2 FILLER_17_786 ();
 sg13g2_fill_1 FILLER_17_788 ();
 sg13g2_fill_1 FILLER_17_799 ();
 sg13g2_fill_2 FILLER_17_808 ();
 sg13g2_decap_4 FILLER_17_825 ();
 sg13g2_fill_1 FILLER_17_829 ();
 sg13g2_fill_1 FILLER_17_844 ();
 sg13g2_fill_1 FILLER_17_857 ();
 sg13g2_fill_2 FILLER_17_867 ();
 sg13g2_fill_1 FILLER_17_883 ();
 sg13g2_fill_2 FILLER_17_935 ();
 sg13g2_fill_2 FILLER_17_946 ();
 sg13g2_decap_8 FILLER_17_1005 ();
 sg13g2_fill_1 FILLER_17_1012 ();
 sg13g2_decap_4 FILLER_17_1017 ();
 sg13g2_fill_1 FILLER_17_1021 ();
 sg13g2_fill_2 FILLER_17_1075 ();
 sg13g2_fill_1 FILLER_17_1077 ();
 sg13g2_decap_4 FILLER_17_1090 ();
 sg13g2_decap_4 FILLER_17_1103 ();
 sg13g2_fill_1 FILLER_17_1107 ();
 sg13g2_fill_1 FILLER_17_1173 ();
 sg13g2_fill_1 FILLER_17_1183 ();
 sg13g2_fill_2 FILLER_17_1224 ();
 sg13g2_fill_1 FILLER_17_1270 ();
 sg13g2_fill_1 FILLER_17_1314 ();
 sg13g2_fill_2 FILLER_17_1350 ();
 sg13g2_decap_4 FILLER_17_1356 ();
 sg13g2_fill_2 FILLER_17_1360 ();
 sg13g2_fill_1 FILLER_17_1382 ();
 sg13g2_decap_8 FILLER_17_1401 ();
 sg13g2_fill_1 FILLER_17_1408 ();
 sg13g2_decap_4 FILLER_17_1422 ();
 sg13g2_fill_1 FILLER_17_1430 ();
 sg13g2_fill_1 FILLER_17_1471 ();
 sg13g2_fill_1 FILLER_17_1486 ();
 sg13g2_fill_2 FILLER_17_1558 ();
 sg13g2_fill_1 FILLER_17_1560 ();
 sg13g2_fill_2 FILLER_17_1634 ();
 sg13g2_fill_1 FILLER_17_1636 ();
 sg13g2_fill_2 FILLER_17_1663 ();
 sg13g2_fill_1 FILLER_17_1665 ();
 sg13g2_fill_2 FILLER_17_1736 ();
 sg13g2_fill_1 FILLER_17_1738 ();
 sg13g2_decap_8 FILLER_17_1765 ();
 sg13g2_fill_1 FILLER_17_1781 ();
 sg13g2_fill_2 FILLER_17_1809 ();
 sg13g2_fill_1 FILLER_17_1811 ();
 sg13g2_fill_2 FILLER_17_1841 ();
 sg13g2_decap_8 FILLER_17_1861 ();
 sg13g2_fill_2 FILLER_17_1868 ();
 sg13g2_decap_8 FILLER_17_1973 ();
 sg13g2_decap_8 FILLER_17_1980 ();
 sg13g2_decap_8 FILLER_17_1991 ();
 sg13g2_fill_1 FILLER_17_2034 ();
 sg13g2_fill_2 FILLER_17_2107 ();
 sg13g2_fill_1 FILLER_17_2109 ();
 sg13g2_fill_1 FILLER_17_2140 ();
 sg13g2_fill_2 FILLER_17_2206 ();
 sg13g2_fill_2 FILLER_17_2213 ();
 sg13g2_fill_1 FILLER_17_2241 ();
 sg13g2_fill_2 FILLER_17_2251 ();
 sg13g2_fill_1 FILLER_17_2253 ();
 sg13g2_fill_2 FILLER_17_2262 ();
 sg13g2_fill_1 FILLER_17_2281 ();
 sg13g2_fill_2 FILLER_17_2290 ();
 sg13g2_fill_2 FILLER_17_2323 ();
 sg13g2_fill_1 FILLER_17_2325 ();
 sg13g2_fill_2 FILLER_17_2331 ();
 sg13g2_fill_1 FILLER_17_2333 ();
 sg13g2_decap_8 FILLER_17_2365 ();
 sg13g2_decap_8 FILLER_17_2372 ();
 sg13g2_decap_8 FILLER_17_2379 ();
 sg13g2_decap_8 FILLER_17_2386 ();
 sg13g2_decap_8 FILLER_17_2393 ();
 sg13g2_decap_8 FILLER_17_2400 ();
 sg13g2_decap_8 FILLER_17_2407 ();
 sg13g2_decap_8 FILLER_17_2414 ();
 sg13g2_decap_8 FILLER_17_2421 ();
 sg13g2_decap_8 FILLER_17_2428 ();
 sg13g2_decap_8 FILLER_17_2435 ();
 sg13g2_decap_8 FILLER_17_2442 ();
 sg13g2_decap_8 FILLER_17_2449 ();
 sg13g2_decap_8 FILLER_17_2456 ();
 sg13g2_decap_8 FILLER_17_2463 ();
 sg13g2_decap_8 FILLER_17_2470 ();
 sg13g2_decap_8 FILLER_17_2477 ();
 sg13g2_decap_8 FILLER_17_2484 ();
 sg13g2_decap_8 FILLER_17_2491 ();
 sg13g2_decap_8 FILLER_17_2498 ();
 sg13g2_decap_8 FILLER_17_2505 ();
 sg13g2_decap_8 FILLER_17_2512 ();
 sg13g2_decap_8 FILLER_17_2519 ();
 sg13g2_decap_8 FILLER_17_2526 ();
 sg13g2_decap_8 FILLER_17_2533 ();
 sg13g2_decap_8 FILLER_17_2540 ();
 sg13g2_decap_8 FILLER_17_2547 ();
 sg13g2_decap_8 FILLER_17_2554 ();
 sg13g2_decap_8 FILLER_17_2561 ();
 sg13g2_decap_8 FILLER_17_2568 ();
 sg13g2_decap_8 FILLER_17_2575 ();
 sg13g2_decap_8 FILLER_17_2582 ();
 sg13g2_decap_8 FILLER_17_2589 ();
 sg13g2_decap_8 FILLER_17_2596 ();
 sg13g2_decap_8 FILLER_17_2603 ();
 sg13g2_decap_8 FILLER_17_2610 ();
 sg13g2_decap_8 FILLER_17_2617 ();
 sg13g2_decap_8 FILLER_17_2624 ();
 sg13g2_decap_8 FILLER_17_2631 ();
 sg13g2_decap_8 FILLER_17_2638 ();
 sg13g2_decap_8 FILLER_17_2645 ();
 sg13g2_decap_8 FILLER_17_2652 ();
 sg13g2_decap_8 FILLER_17_2659 ();
 sg13g2_decap_8 FILLER_17_2666 ();
 sg13g2_fill_1 FILLER_17_2673 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_fill_2 FILLER_18_434 ();
 sg13g2_fill_2 FILLER_18_467 ();
 sg13g2_fill_2 FILLER_18_482 ();
 sg13g2_fill_1 FILLER_18_484 ();
 sg13g2_fill_2 FILLER_18_501 ();
 sg13g2_fill_1 FILLER_18_503 ();
 sg13g2_fill_2 FILLER_18_508 ();
 sg13g2_fill_1 FILLER_18_523 ();
 sg13g2_fill_2 FILLER_18_602 ();
 sg13g2_fill_2 FILLER_18_644 ();
 sg13g2_fill_1 FILLER_18_646 ();
 sg13g2_fill_2 FILLER_18_659 ();
 sg13g2_fill_2 FILLER_18_717 ();
 sg13g2_fill_1 FILLER_18_719 ();
 sg13g2_fill_1 FILLER_18_746 ();
 sg13g2_decap_4 FILLER_18_782 ();
 sg13g2_fill_2 FILLER_18_804 ();
 sg13g2_fill_1 FILLER_18_818 ();
 sg13g2_fill_2 FILLER_18_845 ();
 sg13g2_fill_2 FILLER_18_859 ();
 sg13g2_fill_1 FILLER_18_874 ();
 sg13g2_decap_4 FILLER_18_937 ();
 sg13g2_fill_2 FILLER_18_941 ();
 sg13g2_decap_4 FILLER_18_974 ();
 sg13g2_fill_2 FILLER_18_989 ();
 sg13g2_fill_2 FILLER_18_1030 ();
 sg13g2_fill_2 FILLER_18_1067 ();
 sg13g2_fill_1 FILLER_18_1069 ();
 sg13g2_fill_1 FILLER_18_1122 ();
 sg13g2_fill_2 FILLER_18_1140 ();
 sg13g2_fill_2 FILLER_18_1147 ();
 sg13g2_fill_1 FILLER_18_1157 ();
 sg13g2_fill_1 FILLER_18_1171 ();
 sg13g2_fill_2 FILLER_18_1181 ();
 sg13g2_fill_1 FILLER_18_1183 ();
 sg13g2_fill_1 FILLER_18_1201 ();
 sg13g2_fill_2 FILLER_18_1207 ();
 sg13g2_fill_1 FILLER_18_1209 ();
 sg13g2_fill_2 FILLER_18_1214 ();
 sg13g2_decap_8 FILLER_18_1225 ();
 sg13g2_fill_1 FILLER_18_1232 ();
 sg13g2_decap_4 FILLER_18_1242 ();
 sg13g2_fill_1 FILLER_18_1246 ();
 sg13g2_decap_8 FILLER_18_1287 ();
 sg13g2_fill_2 FILLER_18_1298 ();
 sg13g2_decap_4 FILLER_18_1309 ();
 sg13g2_fill_1 FILLER_18_1318 ();
 sg13g2_decap_8 FILLER_18_1331 ();
 sg13g2_fill_1 FILLER_18_1343 ();
 sg13g2_decap_8 FILLER_18_1357 ();
 sg13g2_fill_1 FILLER_18_1364 ();
 sg13g2_decap_4 FILLER_18_1374 ();
 sg13g2_fill_1 FILLER_18_1378 ();
 sg13g2_fill_2 FILLER_18_1405 ();
 sg13g2_fill_2 FILLER_18_1498 ();
 sg13g2_fill_1 FILLER_18_1500 ();
 sg13g2_decap_8 FILLER_18_1524 ();
 sg13g2_fill_1 FILLER_18_1531 ();
 sg13g2_decap_8 FILLER_18_1536 ();
 sg13g2_fill_2 FILLER_18_1565 ();
 sg13g2_fill_1 FILLER_18_1567 ();
 sg13g2_fill_1 FILLER_18_1592 ();
 sg13g2_fill_1 FILLER_18_1602 ();
 sg13g2_fill_1 FILLER_18_1611 ();
 sg13g2_decap_4 FILLER_18_1677 ();
 sg13g2_fill_2 FILLER_18_1681 ();
 sg13g2_decap_4 FILLER_18_1692 ();
 sg13g2_fill_2 FILLER_18_1696 ();
 sg13g2_fill_1 FILLER_18_1707 ();
 sg13g2_fill_2 FILLER_18_1734 ();
 sg13g2_fill_1 FILLER_18_1754 ();
 sg13g2_decap_4 FILLER_18_1772 ();
 sg13g2_fill_1 FILLER_18_1776 ();
 sg13g2_decap_4 FILLER_18_1786 ();
 sg13g2_fill_1 FILLER_18_1790 ();
 sg13g2_fill_2 FILLER_18_1821 ();
 sg13g2_fill_1 FILLER_18_1831 ();
 sg13g2_decap_8 FILLER_18_1870 ();
 sg13g2_fill_2 FILLER_18_1889 ();
 sg13g2_fill_1 FILLER_18_1891 ();
 sg13g2_decap_4 FILLER_18_1921 ();
 sg13g2_fill_1 FILLER_18_1942 ();
 sg13g2_fill_2 FILLER_18_1947 ();
 sg13g2_fill_1 FILLER_18_2012 ();
 sg13g2_fill_2 FILLER_18_2017 ();
 sg13g2_decap_8 FILLER_18_2060 ();
 sg13g2_decap_4 FILLER_18_2067 ();
 sg13g2_fill_2 FILLER_18_2071 ();
 sg13g2_decap_4 FILLER_18_2077 ();
 sg13g2_fill_2 FILLER_18_2081 ();
 sg13g2_decap_4 FILLER_18_2118 ();
 sg13g2_fill_2 FILLER_18_2122 ();
 sg13g2_fill_1 FILLER_18_2167 ();
 sg13g2_fill_2 FILLER_18_2206 ();
 sg13g2_fill_1 FILLER_18_2216 ();
 sg13g2_fill_1 FILLER_18_2247 ();
 sg13g2_fill_2 FILLER_18_2263 ();
 sg13g2_fill_1 FILLER_18_2265 ();
 sg13g2_decap_8 FILLER_18_2297 ();
 sg13g2_fill_2 FILLER_18_2304 ();
 sg13g2_fill_1 FILLER_18_2306 ();
 sg13g2_fill_2 FILLER_18_2347 ();
 sg13g2_fill_1 FILLER_18_2349 ();
 sg13g2_decap_8 FILLER_18_2376 ();
 sg13g2_decap_8 FILLER_18_2383 ();
 sg13g2_decap_8 FILLER_18_2390 ();
 sg13g2_decap_8 FILLER_18_2397 ();
 sg13g2_decap_8 FILLER_18_2404 ();
 sg13g2_decap_8 FILLER_18_2411 ();
 sg13g2_decap_8 FILLER_18_2418 ();
 sg13g2_decap_8 FILLER_18_2425 ();
 sg13g2_decap_8 FILLER_18_2432 ();
 sg13g2_decap_8 FILLER_18_2439 ();
 sg13g2_decap_8 FILLER_18_2446 ();
 sg13g2_decap_8 FILLER_18_2453 ();
 sg13g2_decap_8 FILLER_18_2460 ();
 sg13g2_decap_8 FILLER_18_2467 ();
 sg13g2_decap_8 FILLER_18_2474 ();
 sg13g2_decap_8 FILLER_18_2481 ();
 sg13g2_decap_8 FILLER_18_2488 ();
 sg13g2_decap_8 FILLER_18_2495 ();
 sg13g2_decap_8 FILLER_18_2502 ();
 sg13g2_decap_8 FILLER_18_2509 ();
 sg13g2_decap_8 FILLER_18_2516 ();
 sg13g2_decap_8 FILLER_18_2523 ();
 sg13g2_decap_8 FILLER_18_2530 ();
 sg13g2_decap_8 FILLER_18_2537 ();
 sg13g2_decap_8 FILLER_18_2544 ();
 sg13g2_decap_8 FILLER_18_2551 ();
 sg13g2_decap_8 FILLER_18_2558 ();
 sg13g2_decap_8 FILLER_18_2565 ();
 sg13g2_decap_8 FILLER_18_2572 ();
 sg13g2_decap_8 FILLER_18_2579 ();
 sg13g2_decap_8 FILLER_18_2586 ();
 sg13g2_decap_8 FILLER_18_2593 ();
 sg13g2_decap_8 FILLER_18_2600 ();
 sg13g2_decap_8 FILLER_18_2607 ();
 sg13g2_decap_8 FILLER_18_2614 ();
 sg13g2_decap_8 FILLER_18_2621 ();
 sg13g2_decap_8 FILLER_18_2628 ();
 sg13g2_decap_8 FILLER_18_2635 ();
 sg13g2_decap_8 FILLER_18_2642 ();
 sg13g2_decap_8 FILLER_18_2649 ();
 sg13g2_decap_8 FILLER_18_2656 ();
 sg13g2_decap_8 FILLER_18_2663 ();
 sg13g2_decap_4 FILLER_18_2670 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_fill_2 FILLER_19_441 ();
 sg13g2_fill_1 FILLER_19_443 ();
 sg13g2_fill_1 FILLER_19_461 ();
 sg13g2_fill_1 FILLER_19_537 ();
 sg13g2_fill_2 FILLER_19_585 ();
 sg13g2_fill_1 FILLER_19_613 ();
 sg13g2_fill_1 FILLER_19_639 ();
 sg13g2_fill_2 FILLER_19_666 ();
 sg13g2_fill_1 FILLER_19_668 ();
 sg13g2_fill_2 FILLER_19_673 ();
 sg13g2_fill_1 FILLER_19_675 ();
 sg13g2_fill_2 FILLER_19_716 ();
 sg13g2_decap_4 FILLER_19_753 ();
 sg13g2_fill_1 FILLER_19_757 ();
 sg13g2_decap_4 FILLER_19_762 ();
 sg13g2_fill_2 FILLER_19_766 ();
 sg13g2_fill_1 FILLER_19_794 ();
 sg13g2_fill_1 FILLER_19_821 ();
 sg13g2_decap_8 FILLER_19_825 ();
 sg13g2_fill_2 FILLER_19_832 ();
 sg13g2_decap_4 FILLER_19_893 ();
 sg13g2_fill_1 FILLER_19_897 ();
 sg13g2_decap_4 FILLER_19_912 ();
 sg13g2_fill_2 FILLER_19_916 ();
 sg13g2_decap_8 FILLER_19_965 ();
 sg13g2_fill_1 FILLER_19_972 ();
 sg13g2_fill_2 FILLER_19_981 ();
 sg13g2_fill_2 FILLER_19_991 ();
 sg13g2_fill_2 FILLER_19_1006 ();
 sg13g2_fill_1 FILLER_19_1008 ();
 sg13g2_fill_1 FILLER_19_1026 ();
 sg13g2_fill_1 FILLER_19_1036 ();
 sg13g2_decap_8 FILLER_19_1125 ();
 sg13g2_fill_2 FILLER_19_1153 ();
 sg13g2_fill_1 FILLER_19_1155 ();
 sg13g2_fill_2 FILLER_19_1160 ();
 sg13g2_fill_1 FILLER_19_1162 ();
 sg13g2_fill_2 FILLER_19_1189 ();
 sg13g2_fill_2 FILLER_19_1260 ();
 sg13g2_fill_1 FILLER_19_1262 ();
 sg13g2_fill_2 FILLER_19_1277 ();
 sg13g2_fill_2 FILLER_19_1292 ();
 sg13g2_fill_2 FILLER_19_1303 ();
 sg13g2_fill_1 FILLER_19_1305 ();
 sg13g2_fill_1 FILLER_19_1326 ();
 sg13g2_fill_1 FILLER_19_1335 ();
 sg13g2_fill_2 FILLER_19_1379 ();
 sg13g2_fill_2 FILLER_19_1394 ();
 sg13g2_fill_1 FILLER_19_1441 ();
 sg13g2_fill_1 FILLER_19_1452 ();
 sg13g2_fill_1 FILLER_19_1462 ();
 sg13g2_decap_4 FILLER_19_1471 ();
 sg13g2_fill_2 FILLER_19_1475 ();
 sg13g2_fill_2 FILLER_19_1491 ();
 sg13g2_fill_1 FILLER_19_1493 ();
 sg13g2_decap_8 FILLER_19_1534 ();
 sg13g2_fill_2 FILLER_19_1593 ();
 sg13g2_fill_2 FILLER_19_1603 ();
 sg13g2_fill_2 FILLER_19_1663 ();
 sg13g2_decap_4 FILLER_19_1691 ();
 sg13g2_fill_1 FILLER_19_1695 ();
 sg13g2_fill_2 FILLER_19_1704 ();
 sg13g2_fill_1 FILLER_19_1711 ();
 sg13g2_fill_2 FILLER_19_1717 ();
 sg13g2_fill_2 FILLER_19_1723 ();
 sg13g2_fill_1 FILLER_19_1725 ();
 sg13g2_decap_4 FILLER_19_1767 ();
 sg13g2_fill_2 FILLER_19_1786 ();
 sg13g2_fill_1 FILLER_19_1837 ();
 sg13g2_fill_1 FILLER_19_1894 ();
 sg13g2_decap_4 FILLER_19_1917 ();
 sg13g2_decap_8 FILLER_19_1978 ();
 sg13g2_fill_2 FILLER_19_1985 ();
 sg13g2_fill_1 FILLER_19_2008 ();
 sg13g2_decap_4 FILLER_19_2022 ();
 sg13g2_fill_2 FILLER_19_2026 ();
 sg13g2_fill_2 FILLER_19_2036 ();
 sg13g2_fill_2 FILLER_19_2047 ();
 sg13g2_fill_1 FILLER_19_2058 ();
 sg13g2_fill_2 FILLER_19_2067 ();
 sg13g2_decap_8 FILLER_19_2086 ();
 sg13g2_fill_1 FILLER_19_2093 ();
 sg13g2_fill_1 FILLER_19_2098 ();
 sg13g2_decap_8 FILLER_19_2104 ();
 sg13g2_fill_1 FILLER_19_2115 ();
 sg13g2_fill_1 FILLER_19_2126 ();
 sg13g2_fill_2 FILLER_19_2131 ();
 sg13g2_fill_2 FILLER_19_2207 ();
 sg13g2_fill_1 FILLER_19_2209 ();
 sg13g2_decap_4 FILLER_19_2223 ();
 sg13g2_fill_1 FILLER_19_2227 ();
 sg13g2_fill_2 FILLER_19_2237 ();
 sg13g2_decap_8 FILLER_19_2280 ();
 sg13g2_fill_2 FILLER_19_2287 ();
 sg13g2_fill_1 FILLER_19_2289 ();
 sg13g2_decap_8 FILLER_19_2298 ();
 sg13g2_decap_4 FILLER_19_2305 ();
 sg13g2_decap_4 FILLER_19_2314 ();
 sg13g2_fill_1 FILLER_19_2331 ();
 sg13g2_fill_1 FILLER_19_2337 ();
 sg13g2_decap_8 FILLER_19_2368 ();
 sg13g2_decap_8 FILLER_19_2375 ();
 sg13g2_decap_8 FILLER_19_2382 ();
 sg13g2_decap_8 FILLER_19_2389 ();
 sg13g2_decap_8 FILLER_19_2396 ();
 sg13g2_decap_8 FILLER_19_2403 ();
 sg13g2_decap_8 FILLER_19_2410 ();
 sg13g2_decap_8 FILLER_19_2417 ();
 sg13g2_decap_8 FILLER_19_2424 ();
 sg13g2_decap_8 FILLER_19_2431 ();
 sg13g2_decap_8 FILLER_19_2438 ();
 sg13g2_decap_8 FILLER_19_2445 ();
 sg13g2_decap_8 FILLER_19_2452 ();
 sg13g2_decap_8 FILLER_19_2459 ();
 sg13g2_decap_8 FILLER_19_2466 ();
 sg13g2_decap_8 FILLER_19_2473 ();
 sg13g2_decap_8 FILLER_19_2480 ();
 sg13g2_decap_8 FILLER_19_2487 ();
 sg13g2_decap_8 FILLER_19_2494 ();
 sg13g2_decap_8 FILLER_19_2501 ();
 sg13g2_decap_8 FILLER_19_2508 ();
 sg13g2_decap_8 FILLER_19_2515 ();
 sg13g2_decap_8 FILLER_19_2522 ();
 sg13g2_decap_8 FILLER_19_2529 ();
 sg13g2_decap_8 FILLER_19_2536 ();
 sg13g2_decap_8 FILLER_19_2543 ();
 sg13g2_decap_8 FILLER_19_2550 ();
 sg13g2_decap_8 FILLER_19_2557 ();
 sg13g2_decap_8 FILLER_19_2564 ();
 sg13g2_decap_8 FILLER_19_2571 ();
 sg13g2_decap_8 FILLER_19_2578 ();
 sg13g2_decap_8 FILLER_19_2585 ();
 sg13g2_decap_8 FILLER_19_2592 ();
 sg13g2_decap_8 FILLER_19_2599 ();
 sg13g2_decap_8 FILLER_19_2606 ();
 sg13g2_decap_8 FILLER_19_2613 ();
 sg13g2_decap_8 FILLER_19_2620 ();
 sg13g2_decap_8 FILLER_19_2627 ();
 sg13g2_decap_8 FILLER_19_2634 ();
 sg13g2_decap_8 FILLER_19_2641 ();
 sg13g2_decap_8 FILLER_19_2648 ();
 sg13g2_decap_8 FILLER_19_2655 ();
 sg13g2_decap_8 FILLER_19_2662 ();
 sg13g2_decap_4 FILLER_19_2669 ();
 sg13g2_fill_1 FILLER_19_2673 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_4 FILLER_20_441 ();
 sg13g2_fill_2 FILLER_20_445 ();
 sg13g2_fill_1 FILLER_20_452 ();
 sg13g2_fill_2 FILLER_20_504 ();
 sg13g2_fill_1 FILLER_20_506 ();
 sg13g2_fill_2 FILLER_20_511 ();
 sg13g2_fill_1 FILLER_20_518 ();
 sg13g2_fill_2 FILLER_20_523 ();
 sg13g2_fill_1 FILLER_20_534 ();
 sg13g2_decap_8 FILLER_20_575 ();
 sg13g2_fill_1 FILLER_20_582 ();
 sg13g2_fill_1 FILLER_20_599 ();
 sg13g2_fill_1 FILLER_20_635 ();
 sg13g2_fill_1 FILLER_20_641 ();
 sg13g2_fill_2 FILLER_20_659 ();
 sg13g2_fill_2 FILLER_20_682 ();
 sg13g2_fill_2 FILLER_20_731 ();
 sg13g2_fill_2 FILLER_20_759 ();
 sg13g2_fill_1 FILLER_20_774 ();
 sg13g2_fill_2 FILLER_20_810 ();
 sg13g2_fill_1 FILLER_20_821 ();
 sg13g2_fill_2 FILLER_20_848 ();
 sg13g2_fill_1 FILLER_20_850 ();
 sg13g2_fill_2 FILLER_20_860 ();
 sg13g2_decap_8 FILLER_20_894 ();
 sg13g2_decap_4 FILLER_20_901 ();
 sg13g2_decap_8 FILLER_20_910 ();
 sg13g2_fill_1 FILLER_20_917 ();
 sg13g2_decap_4 FILLER_20_922 ();
 sg13g2_fill_2 FILLER_20_931 ();
 sg13g2_decap_8 FILLER_20_938 ();
 sg13g2_decap_4 FILLER_20_945 ();
 sg13g2_fill_1 FILLER_20_949 ();
 sg13g2_fill_2 FILLER_20_954 ();
 sg13g2_fill_1 FILLER_20_961 ();
 sg13g2_fill_1 FILLER_20_1002 ();
 sg13g2_fill_2 FILLER_20_1008 ();
 sg13g2_fill_1 FILLER_20_1010 ();
 sg13g2_fill_1 FILLER_20_1072 ();
 sg13g2_fill_1 FILLER_20_1108 ();
 sg13g2_fill_1 FILLER_20_1140 ();
 sg13g2_fill_2 FILLER_20_1166 ();
 sg13g2_fill_2 FILLER_20_1172 ();
 sg13g2_decap_4 FILLER_20_1178 ();
 sg13g2_fill_1 FILLER_20_1182 ();
 sg13g2_fill_2 FILLER_20_1195 ();
 sg13g2_fill_1 FILLER_20_1206 ();
 sg13g2_fill_1 FILLER_20_1216 ();
 sg13g2_decap_4 FILLER_20_1225 ();
 sg13g2_fill_1 FILLER_20_1229 ();
 sg13g2_fill_2 FILLER_20_1243 ();
 sg13g2_fill_1 FILLER_20_1245 ();
 sg13g2_fill_2 FILLER_20_1281 ();
 sg13g2_decap_4 FILLER_20_1309 ();
 sg13g2_fill_1 FILLER_20_1335 ();
 sg13g2_decap_4 FILLER_20_1341 ();
 sg13g2_fill_1 FILLER_20_1345 ();
 sg13g2_fill_2 FILLER_20_1367 ();
 sg13g2_fill_2 FILLER_20_1421 ();
 sg13g2_fill_2 FILLER_20_1449 ();
 sg13g2_fill_1 FILLER_20_1451 ();
 sg13g2_fill_2 FILLER_20_1557 ();
 sg13g2_fill_1 FILLER_20_1559 ();
 sg13g2_fill_1 FILLER_20_1567 ();
 sg13g2_decap_4 FILLER_20_1572 ();
 sg13g2_fill_2 FILLER_20_1576 ();
 sg13g2_fill_2 FILLER_20_1605 ();
 sg13g2_fill_2 FILLER_20_1630 ();
 sg13g2_fill_1 FILLER_20_1632 ();
 sg13g2_fill_1 FILLER_20_1647 ();
 sg13g2_decap_8 FILLER_20_1682 ();
 sg13g2_decap_4 FILLER_20_1689 ();
 sg13g2_fill_2 FILLER_20_1693 ();
 sg13g2_decap_4 FILLER_20_1700 ();
 sg13g2_fill_1 FILLER_20_1739 ();
 sg13g2_fill_2 FILLER_20_1775 ();
 sg13g2_fill_1 FILLER_20_1777 ();
 sg13g2_fill_1 FILLER_20_1786 ();
 sg13g2_decap_8 FILLER_20_1870 ();
 sg13g2_fill_1 FILLER_20_1877 ();
 sg13g2_fill_2 FILLER_20_1913 ();
 sg13g2_fill_2 FILLER_20_1936 ();
 sg13g2_fill_1 FILLER_20_1938 ();
 sg13g2_fill_2 FILLER_20_1943 ();
 sg13g2_fill_1 FILLER_20_1945 ();
 sg13g2_decap_4 FILLER_20_1950 ();
 sg13g2_fill_2 FILLER_20_1992 ();
 sg13g2_fill_1 FILLER_20_1994 ();
 sg13g2_fill_2 FILLER_20_2000 ();
 sg13g2_fill_2 FILLER_20_2063 ();
 sg13g2_fill_1 FILLER_20_2091 ();
 sg13g2_fill_2 FILLER_20_2110 ();
 sg13g2_fill_1 FILLER_20_2161 ();
 sg13g2_fill_1 FILLER_20_2181 ();
 sg13g2_decap_4 FILLER_20_2198 ();
 sg13g2_fill_1 FILLER_20_2206 ();
 sg13g2_fill_1 FILLER_20_2212 ();
 sg13g2_fill_1 FILLER_20_2217 ();
 sg13g2_fill_1 FILLER_20_2227 ();
 sg13g2_fill_1 FILLER_20_2259 ();
 sg13g2_fill_2 FILLER_20_2352 ();
 sg13g2_decap_8 FILLER_20_2367 ();
 sg13g2_decap_8 FILLER_20_2374 ();
 sg13g2_decap_8 FILLER_20_2381 ();
 sg13g2_decap_8 FILLER_20_2388 ();
 sg13g2_decap_8 FILLER_20_2395 ();
 sg13g2_decap_8 FILLER_20_2402 ();
 sg13g2_decap_8 FILLER_20_2409 ();
 sg13g2_decap_8 FILLER_20_2416 ();
 sg13g2_decap_8 FILLER_20_2423 ();
 sg13g2_decap_8 FILLER_20_2430 ();
 sg13g2_decap_8 FILLER_20_2437 ();
 sg13g2_decap_8 FILLER_20_2444 ();
 sg13g2_decap_8 FILLER_20_2451 ();
 sg13g2_decap_8 FILLER_20_2458 ();
 sg13g2_decap_8 FILLER_20_2465 ();
 sg13g2_decap_8 FILLER_20_2472 ();
 sg13g2_decap_8 FILLER_20_2479 ();
 sg13g2_decap_8 FILLER_20_2486 ();
 sg13g2_decap_8 FILLER_20_2493 ();
 sg13g2_decap_8 FILLER_20_2500 ();
 sg13g2_decap_8 FILLER_20_2507 ();
 sg13g2_decap_8 FILLER_20_2514 ();
 sg13g2_decap_8 FILLER_20_2521 ();
 sg13g2_decap_8 FILLER_20_2528 ();
 sg13g2_decap_8 FILLER_20_2535 ();
 sg13g2_decap_8 FILLER_20_2542 ();
 sg13g2_decap_8 FILLER_20_2549 ();
 sg13g2_decap_8 FILLER_20_2556 ();
 sg13g2_decap_8 FILLER_20_2563 ();
 sg13g2_decap_8 FILLER_20_2570 ();
 sg13g2_decap_8 FILLER_20_2577 ();
 sg13g2_decap_8 FILLER_20_2584 ();
 sg13g2_decap_8 FILLER_20_2591 ();
 sg13g2_decap_8 FILLER_20_2598 ();
 sg13g2_decap_8 FILLER_20_2605 ();
 sg13g2_decap_8 FILLER_20_2612 ();
 sg13g2_decap_8 FILLER_20_2619 ();
 sg13g2_decap_8 FILLER_20_2626 ();
 sg13g2_decap_8 FILLER_20_2633 ();
 sg13g2_decap_8 FILLER_20_2640 ();
 sg13g2_decap_8 FILLER_20_2647 ();
 sg13g2_decap_8 FILLER_20_2654 ();
 sg13g2_decap_8 FILLER_20_2661 ();
 sg13g2_decap_4 FILLER_20_2668 ();
 sg13g2_fill_2 FILLER_20_2672 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_fill_2 FILLER_21_427 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_fill_1 FILLER_21_456 ();
 sg13g2_fill_2 FILLER_21_502 ();
 sg13g2_fill_2 FILLER_21_556 ();
 sg13g2_fill_1 FILLER_21_593 ();
 sg13g2_fill_2 FILLER_21_599 ();
 sg13g2_fill_2 FILLER_21_702 ();
 sg13g2_fill_2 FILLER_21_709 ();
 sg13g2_fill_1 FILLER_21_729 ();
 sg13g2_fill_2 FILLER_21_743 ();
 sg13g2_fill_1 FILLER_21_785 ();
 sg13g2_fill_1 FILLER_21_817 ();
 sg13g2_fill_2 FILLER_21_840 ();
 sg13g2_fill_2 FILLER_21_933 ();
 sg13g2_decap_4 FILLER_21_940 ();
 sg13g2_decap_4 FILLER_21_949 ();
 sg13g2_fill_1 FILLER_21_961 ();
 sg13g2_fill_2 FILLER_21_992 ();
 sg13g2_fill_1 FILLER_21_994 ();
 sg13g2_fill_2 FILLER_21_1021 ();
 sg13g2_fill_1 FILLER_21_1023 ();
 sg13g2_fill_2 FILLER_21_1041 ();
 sg13g2_fill_2 FILLER_21_1061 ();
 sg13g2_fill_1 FILLER_21_1063 ();
 sg13g2_fill_2 FILLER_21_1073 ();
 sg13g2_fill_2 FILLER_21_1080 ();
 sg13g2_fill_1 FILLER_21_1082 ();
 sg13g2_fill_2 FILLER_21_1087 ();
 sg13g2_fill_1 FILLER_21_1089 ();
 sg13g2_fill_2 FILLER_21_1107 ();
 sg13g2_fill_1 FILLER_21_1109 ();
 sg13g2_decap_8 FILLER_21_1144 ();
 sg13g2_decap_4 FILLER_21_1151 ();
 sg13g2_fill_2 FILLER_21_1155 ();
 sg13g2_decap_4 FILLER_21_1192 ();
 sg13g2_fill_1 FILLER_21_1196 ();
 sg13g2_decap_8 FILLER_21_1242 ();
 sg13g2_fill_2 FILLER_21_1249 ();
 sg13g2_fill_2 FILLER_21_1285 ();
 sg13g2_fill_1 FILLER_21_1292 ();
 sg13g2_fill_2 FILLER_21_1320 ();
 sg13g2_fill_1 FILLER_21_1322 ();
 sg13g2_fill_2 FILLER_21_1349 ();
 sg13g2_fill_1 FILLER_21_1351 ();
 sg13g2_fill_2 FILLER_21_1356 ();
 sg13g2_fill_2 FILLER_21_1363 ();
 sg13g2_fill_1 FILLER_21_1365 ();
 sg13g2_fill_2 FILLER_21_1375 ();
 sg13g2_decap_4 FILLER_21_1407 ();
 sg13g2_fill_1 FILLER_21_1411 ();
 sg13g2_decap_4 FILLER_21_1421 ();
 sg13g2_decap_8 FILLER_21_1452 ();
 sg13g2_fill_1 FILLER_21_1459 ();
 sg13g2_fill_1 FILLER_21_1506 ();
 sg13g2_decap_4 FILLER_21_1534 ();
 sg13g2_fill_1 FILLER_21_1538 ();
 sg13g2_fill_2 FILLER_21_1547 ();
 sg13g2_decap_4 FILLER_21_1625 ();
 sg13g2_fill_1 FILLER_21_1629 ();
 sg13g2_fill_2 FILLER_21_1640 ();
 sg13g2_fill_2 FILLER_21_1673 ();
 sg13g2_decap_4 FILLER_21_1696 ();
 sg13g2_fill_1 FILLER_21_1704 ();
 sg13g2_decap_4 FILLER_21_1709 ();
 sg13g2_fill_1 FILLER_21_1713 ();
 sg13g2_fill_2 FILLER_21_1735 ();
 sg13g2_fill_1 FILLER_21_1737 ();
 sg13g2_fill_1 FILLER_21_1789 ();
 sg13g2_fill_1 FILLER_21_1803 ();
 sg13g2_decap_8 FILLER_21_1816 ();
 sg13g2_decap_4 FILLER_21_1823 ();
 sg13g2_fill_2 FILLER_21_1827 ();
 sg13g2_fill_2 FILLER_21_1851 ();
 sg13g2_fill_1 FILLER_21_1883 ();
 sg13g2_decap_4 FILLER_21_1892 ();
 sg13g2_fill_2 FILLER_21_1896 ();
 sg13g2_fill_2 FILLER_21_1919 ();
 sg13g2_decap_4 FILLER_21_1929 ();
 sg13g2_fill_2 FILLER_21_1933 ();
 sg13g2_fill_1 FILLER_21_1969 ();
 sg13g2_fill_2 FILLER_21_2000 ();
 sg13g2_fill_2 FILLER_21_2007 ();
 sg13g2_fill_1 FILLER_21_2009 ();
 sg13g2_decap_8 FILLER_21_2018 ();
 sg13g2_fill_1 FILLER_21_2074 ();
 sg13g2_fill_1 FILLER_21_2084 ();
 sg13g2_fill_2 FILLER_21_2094 ();
 sg13g2_fill_1 FILLER_21_2109 ();
 sg13g2_fill_2 FILLER_21_2130 ();
 sg13g2_fill_1 FILLER_21_2132 ();
 sg13g2_fill_2 FILLER_21_2142 ();
 sg13g2_fill_2 FILLER_21_2188 ();
 sg13g2_fill_1 FILLER_21_2190 ();
 sg13g2_fill_2 FILLER_21_2196 ();
 sg13g2_fill_1 FILLER_21_2237 ();
 sg13g2_fill_2 FILLER_21_2261 ();
 sg13g2_fill_2 FILLER_21_2281 ();
 sg13g2_fill_1 FILLER_21_2283 ();
 sg13g2_fill_1 FILLER_21_2289 ();
 sg13g2_decap_4 FILLER_21_2298 ();
 sg13g2_fill_2 FILLER_21_2315 ();
 sg13g2_decap_8 FILLER_21_2365 ();
 sg13g2_decap_8 FILLER_21_2372 ();
 sg13g2_decap_8 FILLER_21_2379 ();
 sg13g2_decap_8 FILLER_21_2386 ();
 sg13g2_decap_8 FILLER_21_2393 ();
 sg13g2_decap_8 FILLER_21_2400 ();
 sg13g2_decap_8 FILLER_21_2407 ();
 sg13g2_decap_8 FILLER_21_2414 ();
 sg13g2_decap_8 FILLER_21_2421 ();
 sg13g2_decap_8 FILLER_21_2428 ();
 sg13g2_decap_8 FILLER_21_2435 ();
 sg13g2_decap_8 FILLER_21_2442 ();
 sg13g2_decap_8 FILLER_21_2449 ();
 sg13g2_decap_8 FILLER_21_2456 ();
 sg13g2_decap_8 FILLER_21_2463 ();
 sg13g2_decap_8 FILLER_21_2470 ();
 sg13g2_decap_8 FILLER_21_2477 ();
 sg13g2_decap_8 FILLER_21_2484 ();
 sg13g2_decap_8 FILLER_21_2491 ();
 sg13g2_decap_8 FILLER_21_2498 ();
 sg13g2_decap_8 FILLER_21_2505 ();
 sg13g2_decap_8 FILLER_21_2512 ();
 sg13g2_decap_8 FILLER_21_2519 ();
 sg13g2_decap_8 FILLER_21_2526 ();
 sg13g2_decap_8 FILLER_21_2533 ();
 sg13g2_decap_8 FILLER_21_2540 ();
 sg13g2_decap_8 FILLER_21_2547 ();
 sg13g2_decap_8 FILLER_21_2554 ();
 sg13g2_decap_8 FILLER_21_2561 ();
 sg13g2_decap_8 FILLER_21_2568 ();
 sg13g2_decap_8 FILLER_21_2575 ();
 sg13g2_decap_8 FILLER_21_2582 ();
 sg13g2_decap_8 FILLER_21_2589 ();
 sg13g2_decap_8 FILLER_21_2596 ();
 sg13g2_decap_8 FILLER_21_2603 ();
 sg13g2_decap_8 FILLER_21_2610 ();
 sg13g2_decap_8 FILLER_21_2617 ();
 sg13g2_decap_8 FILLER_21_2624 ();
 sg13g2_decap_8 FILLER_21_2631 ();
 sg13g2_decap_8 FILLER_21_2638 ();
 sg13g2_decap_8 FILLER_21_2645 ();
 sg13g2_decap_8 FILLER_21_2652 ();
 sg13g2_decap_8 FILLER_21_2659 ();
 sg13g2_decap_8 FILLER_21_2666 ();
 sg13g2_fill_1 FILLER_21_2673 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_4 FILLER_22_427 ();
 sg13g2_fill_2 FILLER_22_431 ();
 sg13g2_fill_2 FILLER_22_459 ();
 sg13g2_fill_1 FILLER_22_496 ();
 sg13g2_fill_2 FILLER_22_506 ();
 sg13g2_fill_1 FILLER_22_516 ();
 sg13g2_fill_1 FILLER_22_542 ();
 sg13g2_fill_1 FILLER_22_561 ();
 sg13g2_fill_2 FILLER_22_567 ();
 sg13g2_fill_2 FILLER_22_577 ();
 sg13g2_fill_2 FILLER_22_618 ();
 sg13g2_fill_1 FILLER_22_620 ();
 sg13g2_fill_2 FILLER_22_654 ();
 sg13g2_fill_2 FILLER_22_660 ();
 sg13g2_fill_2 FILLER_22_688 ();
 sg13g2_fill_2 FILLER_22_735 ();
 sg13g2_fill_1 FILLER_22_775 ();
 sg13g2_decap_8 FILLER_22_786 ();
 sg13g2_fill_2 FILLER_22_793 ();
 sg13g2_fill_2 FILLER_22_806 ();
 sg13g2_fill_2 FILLER_22_816 ();
 sg13g2_fill_1 FILLER_22_826 ();
 sg13g2_fill_2 FILLER_22_853 ();
 sg13g2_fill_2 FILLER_22_901 ();
 sg13g2_fill_1 FILLER_22_903 ();
 sg13g2_fill_1 FILLER_22_917 ();
 sg13g2_fill_2 FILLER_22_948 ();
 sg13g2_fill_1 FILLER_22_958 ();
 sg13g2_fill_2 FILLER_22_985 ();
 sg13g2_fill_1 FILLER_22_997 ();
 sg13g2_fill_2 FILLER_22_1019 ();
 sg13g2_fill_2 FILLER_22_1066 ();
 sg13g2_fill_1 FILLER_22_1068 ();
 sg13g2_fill_1 FILLER_22_1125 ();
 sg13g2_fill_1 FILLER_22_1135 ();
 sg13g2_fill_2 FILLER_22_1231 ();
 sg13g2_fill_1 FILLER_22_1250 ();
 sg13g2_fill_1 FILLER_22_1292 ();
 sg13g2_fill_2 FILLER_22_1302 ();
 sg13g2_fill_1 FILLER_22_1320 ();
 sg13g2_fill_2 FILLER_22_1357 ();
 sg13g2_fill_2 FILLER_22_1377 ();
 sg13g2_fill_1 FILLER_22_1379 ();
 sg13g2_fill_1 FILLER_22_1385 ();
 sg13g2_fill_2 FILLER_22_1403 ();
 sg13g2_fill_1 FILLER_22_1405 ();
 sg13g2_fill_1 FILLER_22_1490 ();
 sg13g2_decap_8 FILLER_22_1552 ();
 sg13g2_fill_1 FILLER_22_1559 ();
 sg13g2_decap_8 FILLER_22_1568 ();
 sg13g2_fill_2 FILLER_22_1578 ();
 sg13g2_fill_1 FILLER_22_1590 ();
 sg13g2_fill_2 FILLER_22_1596 ();
 sg13g2_fill_2 FILLER_22_1653 ();
 sg13g2_fill_1 FILLER_22_1655 ();
 sg13g2_fill_2 FILLER_22_1696 ();
 sg13g2_fill_1 FILLER_22_1729 ();
 sg13g2_fill_2 FILLER_22_1740 ();
 sg13g2_fill_2 FILLER_22_1755 ();
 sg13g2_fill_1 FILLER_22_1757 ();
 sg13g2_fill_2 FILLER_22_1794 ();
 sg13g2_fill_1 FILLER_22_1796 ();
 sg13g2_decap_8 FILLER_22_1852 ();
 sg13g2_decap_4 FILLER_22_1859 ();
 sg13g2_fill_1 FILLER_22_1863 ();
 sg13g2_fill_2 FILLER_22_1868 ();
 sg13g2_fill_1 FILLER_22_1879 ();
 sg13g2_fill_1 FILLER_22_1941 ();
 sg13g2_fill_2 FILLER_22_1951 ();
 sg13g2_fill_1 FILLER_22_1958 ();
 sg13g2_fill_1 FILLER_22_1978 ();
 sg13g2_fill_2 FILLER_22_2045 ();
 sg13g2_fill_1 FILLER_22_2057 ();
 sg13g2_fill_2 FILLER_22_2174 ();
 sg13g2_fill_1 FILLER_22_2176 ();
 sg13g2_fill_1 FILLER_22_2203 ();
 sg13g2_fill_2 FILLER_22_2254 ();
 sg13g2_decap_4 FILLER_22_2282 ();
 sg13g2_fill_1 FILLER_22_2325 ();
 sg13g2_fill_1 FILLER_22_2331 ();
 sg13g2_decap_4 FILLER_22_2349 ();
 sg13g2_fill_1 FILLER_22_2353 ();
 sg13g2_decap_8 FILLER_22_2367 ();
 sg13g2_decap_8 FILLER_22_2374 ();
 sg13g2_decap_8 FILLER_22_2381 ();
 sg13g2_decap_8 FILLER_22_2388 ();
 sg13g2_decap_8 FILLER_22_2395 ();
 sg13g2_decap_8 FILLER_22_2402 ();
 sg13g2_decap_8 FILLER_22_2409 ();
 sg13g2_decap_8 FILLER_22_2416 ();
 sg13g2_decap_8 FILLER_22_2423 ();
 sg13g2_decap_8 FILLER_22_2430 ();
 sg13g2_decap_8 FILLER_22_2437 ();
 sg13g2_decap_8 FILLER_22_2444 ();
 sg13g2_decap_8 FILLER_22_2451 ();
 sg13g2_decap_8 FILLER_22_2458 ();
 sg13g2_decap_8 FILLER_22_2465 ();
 sg13g2_decap_8 FILLER_22_2472 ();
 sg13g2_decap_8 FILLER_22_2479 ();
 sg13g2_decap_8 FILLER_22_2486 ();
 sg13g2_decap_8 FILLER_22_2493 ();
 sg13g2_decap_8 FILLER_22_2500 ();
 sg13g2_decap_8 FILLER_22_2507 ();
 sg13g2_decap_8 FILLER_22_2514 ();
 sg13g2_decap_8 FILLER_22_2521 ();
 sg13g2_decap_8 FILLER_22_2528 ();
 sg13g2_decap_8 FILLER_22_2535 ();
 sg13g2_decap_8 FILLER_22_2542 ();
 sg13g2_decap_8 FILLER_22_2549 ();
 sg13g2_decap_8 FILLER_22_2556 ();
 sg13g2_decap_8 FILLER_22_2563 ();
 sg13g2_decap_8 FILLER_22_2570 ();
 sg13g2_decap_8 FILLER_22_2577 ();
 sg13g2_decap_8 FILLER_22_2584 ();
 sg13g2_decap_8 FILLER_22_2591 ();
 sg13g2_decap_8 FILLER_22_2598 ();
 sg13g2_decap_8 FILLER_22_2605 ();
 sg13g2_decap_8 FILLER_22_2612 ();
 sg13g2_decap_8 FILLER_22_2619 ();
 sg13g2_decap_8 FILLER_22_2626 ();
 sg13g2_decap_8 FILLER_22_2633 ();
 sg13g2_decap_8 FILLER_22_2640 ();
 sg13g2_decap_8 FILLER_22_2647 ();
 sg13g2_decap_8 FILLER_22_2654 ();
 sg13g2_decap_8 FILLER_22_2661 ();
 sg13g2_decap_4 FILLER_22_2668 ();
 sg13g2_fill_2 FILLER_22_2672 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_fill_2 FILLER_23_491 ();
 sg13g2_fill_1 FILLER_23_493 ();
 sg13g2_fill_2 FILLER_23_524 ();
 sg13g2_fill_1 FILLER_23_552 ();
 sg13g2_fill_1 FILLER_23_556 ();
 sg13g2_fill_2 FILLER_23_607 ();
 sg13g2_fill_1 FILLER_23_609 ();
 sg13g2_fill_1 FILLER_23_624 ();
 sg13g2_fill_2 FILLER_23_635 ();
 sg13g2_decap_8 FILLER_23_663 ();
 sg13g2_fill_2 FILLER_23_670 ();
 sg13g2_fill_2 FILLER_23_676 ();
 sg13g2_fill_1 FILLER_23_678 ();
 sg13g2_decap_4 FILLER_23_688 ();
 sg13g2_fill_1 FILLER_23_705 ();
 sg13g2_fill_1 FILLER_23_710 ();
 sg13g2_fill_1 FILLER_23_763 ();
 sg13g2_fill_1 FILLER_23_773 ();
 sg13g2_fill_2 FILLER_23_779 ();
 sg13g2_fill_1 FILLER_23_781 ();
 sg13g2_fill_1 FILLER_23_790 ();
 sg13g2_fill_2 FILLER_23_808 ();
 sg13g2_fill_1 FILLER_23_810 ();
 sg13g2_fill_2 FILLER_23_815 ();
 sg13g2_fill_2 FILLER_23_827 ();
 sg13g2_fill_1 FILLER_23_829 ();
 sg13g2_fill_2 FILLER_23_873 ();
 sg13g2_fill_1 FILLER_23_875 ();
 sg13g2_fill_2 FILLER_23_894 ();
 sg13g2_fill_2 FILLER_23_904 ();
 sg13g2_fill_1 FILLER_23_918 ();
 sg13g2_fill_2 FILLER_23_928 ();
 sg13g2_fill_1 FILLER_23_930 ();
 sg13g2_fill_1 FILLER_23_958 ();
 sg13g2_fill_2 FILLER_23_985 ();
 sg13g2_fill_1 FILLER_23_997 ();
 sg13g2_decap_4 FILLER_23_1037 ();
 sg13g2_fill_2 FILLER_23_1049 ();
 sg13g2_fill_1 FILLER_23_1051 ();
 sg13g2_fill_2 FILLER_23_1088 ();
 sg13g2_fill_1 FILLER_23_1090 ();
 sg13g2_fill_2 FILLER_23_1104 ();
 sg13g2_fill_1 FILLER_23_1106 ();
 sg13g2_fill_2 FILLER_23_1121 ();
 sg13g2_fill_1 FILLER_23_1136 ();
 sg13g2_fill_1 FILLER_23_1162 ();
 sg13g2_fill_1 FILLER_23_1171 ();
 sg13g2_fill_2 FILLER_23_1211 ();
 sg13g2_fill_1 FILLER_23_1213 ();
 sg13g2_fill_2 FILLER_23_1219 ();
 sg13g2_fill_1 FILLER_23_1221 ();
 sg13g2_decap_8 FILLER_23_1226 ();
 sg13g2_decap_4 FILLER_23_1233 ();
 sg13g2_decap_8 FILLER_23_1247 ();
 sg13g2_decap_8 FILLER_23_1254 ();
 sg13g2_fill_2 FILLER_23_1261 ();
 sg13g2_fill_1 FILLER_23_1311 ();
 sg13g2_fill_1 FILLER_23_1359 ();
 sg13g2_fill_1 FILLER_23_1381 ();
 sg13g2_fill_1 FILLER_23_1408 ();
 sg13g2_fill_1 FILLER_23_1425 ();
 sg13g2_fill_2 FILLER_23_1430 ();
 sg13g2_fill_1 FILLER_23_1432 ();
 sg13g2_decap_4 FILLER_23_1438 ();
 sg13g2_fill_2 FILLER_23_1442 ();
 sg13g2_fill_1 FILLER_23_1502 ();
 sg13g2_decap_8 FILLER_23_1516 ();
 sg13g2_fill_1 FILLER_23_1523 ();
 sg13g2_fill_2 FILLER_23_1541 ();
 sg13g2_fill_1 FILLER_23_1543 ();
 sg13g2_fill_2 FILLER_23_1663 ();
 sg13g2_fill_1 FILLER_23_1704 ();
 sg13g2_fill_1 FILLER_23_1748 ();
 sg13g2_fill_1 FILLER_23_1780 ();
 sg13g2_fill_2 FILLER_23_1811 ();
 sg13g2_fill_1 FILLER_23_1813 ();
 sg13g2_fill_2 FILLER_23_1832 ();
 sg13g2_fill_2 FILLER_23_1866 ();
 sg13g2_fill_1 FILLER_23_1912 ();
 sg13g2_fill_2 FILLER_23_1921 ();
 sg13g2_fill_1 FILLER_23_1923 ();
 sg13g2_fill_2 FILLER_23_1938 ();
 sg13g2_fill_1 FILLER_23_1940 ();
 sg13g2_fill_2 FILLER_23_1989 ();
 sg13g2_fill_1 FILLER_23_2008 ();
 sg13g2_fill_1 FILLER_23_2026 ();
 sg13g2_fill_2 FILLER_23_2078 ();
 sg13g2_fill_2 FILLER_23_2094 ();
 sg13g2_fill_1 FILLER_23_2096 ();
 sg13g2_fill_2 FILLER_23_2114 ();
 sg13g2_fill_1 FILLER_23_2116 ();
 sg13g2_decap_4 FILLER_23_2123 ();
 sg13g2_decap_8 FILLER_23_2131 ();
 sg13g2_fill_2 FILLER_23_2138 ();
 sg13g2_fill_2 FILLER_23_2192 ();
 sg13g2_fill_1 FILLER_23_2208 ();
 sg13g2_decap_4 FILLER_23_2235 ();
 sg13g2_decap_4 FILLER_23_2247 ();
 sg13g2_decap_4 FILLER_23_2276 ();
 sg13g2_fill_1 FILLER_23_2284 ();
 sg13g2_fill_2 FILLER_23_2317 ();
 sg13g2_decap_8 FILLER_23_2371 ();
 sg13g2_decap_8 FILLER_23_2378 ();
 sg13g2_decap_8 FILLER_23_2385 ();
 sg13g2_decap_8 FILLER_23_2392 ();
 sg13g2_decap_8 FILLER_23_2399 ();
 sg13g2_decap_8 FILLER_23_2406 ();
 sg13g2_decap_8 FILLER_23_2413 ();
 sg13g2_decap_8 FILLER_23_2420 ();
 sg13g2_decap_8 FILLER_23_2427 ();
 sg13g2_decap_8 FILLER_23_2434 ();
 sg13g2_decap_8 FILLER_23_2441 ();
 sg13g2_decap_8 FILLER_23_2448 ();
 sg13g2_decap_8 FILLER_23_2455 ();
 sg13g2_decap_8 FILLER_23_2462 ();
 sg13g2_decap_8 FILLER_23_2469 ();
 sg13g2_decap_8 FILLER_23_2476 ();
 sg13g2_decap_8 FILLER_23_2483 ();
 sg13g2_decap_8 FILLER_23_2490 ();
 sg13g2_decap_8 FILLER_23_2497 ();
 sg13g2_decap_8 FILLER_23_2504 ();
 sg13g2_decap_8 FILLER_23_2511 ();
 sg13g2_decap_8 FILLER_23_2518 ();
 sg13g2_decap_8 FILLER_23_2525 ();
 sg13g2_decap_8 FILLER_23_2532 ();
 sg13g2_decap_8 FILLER_23_2539 ();
 sg13g2_decap_8 FILLER_23_2546 ();
 sg13g2_decap_8 FILLER_23_2553 ();
 sg13g2_decap_8 FILLER_23_2560 ();
 sg13g2_decap_8 FILLER_23_2567 ();
 sg13g2_decap_8 FILLER_23_2574 ();
 sg13g2_decap_8 FILLER_23_2581 ();
 sg13g2_decap_8 FILLER_23_2588 ();
 sg13g2_decap_8 FILLER_23_2595 ();
 sg13g2_decap_8 FILLER_23_2602 ();
 sg13g2_decap_8 FILLER_23_2609 ();
 sg13g2_decap_8 FILLER_23_2616 ();
 sg13g2_decap_8 FILLER_23_2623 ();
 sg13g2_decap_8 FILLER_23_2630 ();
 sg13g2_decap_8 FILLER_23_2637 ();
 sg13g2_decap_8 FILLER_23_2644 ();
 sg13g2_decap_8 FILLER_23_2651 ();
 sg13g2_decap_8 FILLER_23_2658 ();
 sg13g2_decap_8 FILLER_23_2665 ();
 sg13g2_fill_2 FILLER_23_2672 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_4 FILLER_24_434 ();
 sg13g2_fill_2 FILLER_24_438 ();
 sg13g2_decap_4 FILLER_24_444 ();
 sg13g2_fill_1 FILLER_24_448 ();
 sg13g2_fill_2 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_477 ();
 sg13g2_fill_1 FILLER_24_484 ();
 sg13g2_decap_4 FILLER_24_490 ();
 sg13g2_fill_2 FILLER_24_494 ();
 sg13g2_fill_2 FILLER_24_532 ();
 sg13g2_fill_1 FILLER_24_534 ();
 sg13g2_fill_2 FILLER_24_569 ();
 sg13g2_fill_1 FILLER_24_571 ();
 sg13g2_fill_2 FILLER_24_585 ();
 sg13g2_fill_1 FILLER_24_587 ();
 sg13g2_fill_1 FILLER_24_601 ();
 sg13g2_fill_2 FILLER_24_637 ();
 sg13g2_fill_1 FILLER_24_639 ();
 sg13g2_fill_1 FILLER_24_662 ();
 sg13g2_fill_2 FILLER_24_698 ();
 sg13g2_fill_1 FILLER_24_700 ();
 sg13g2_fill_1 FILLER_24_714 ();
 sg13g2_fill_2 FILLER_24_747 ();
 sg13g2_fill_1 FILLER_24_749 ();
 sg13g2_decap_4 FILLER_24_768 ();
 sg13g2_fill_2 FILLER_24_772 ();
 sg13g2_decap_4 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_800 ();
 sg13g2_fill_1 FILLER_24_807 ();
 sg13g2_fill_2 FILLER_24_818 ();
 sg13g2_fill_2 FILLER_24_824 ();
 sg13g2_fill_1 FILLER_24_826 ();
 sg13g2_fill_1 FILLER_24_839 ();
 sg13g2_fill_2 FILLER_24_907 ();
 sg13g2_fill_2 FILLER_24_950 ();
 sg13g2_fill_2 FILLER_24_1019 ();
 sg13g2_fill_1 FILLER_24_1021 ();
 sg13g2_fill_1 FILLER_24_1025 ();
 sg13g2_decap_4 FILLER_24_1034 ();
 sg13g2_fill_2 FILLER_24_1051 ();
 sg13g2_fill_1 FILLER_24_1062 ();
 sg13g2_fill_2 FILLER_24_1093 ();
 sg13g2_fill_2 FILLER_24_1113 ();
 sg13g2_fill_1 FILLER_24_1150 ();
 sg13g2_fill_1 FILLER_24_1159 ();
 sg13g2_fill_1 FILLER_24_1177 ();
 sg13g2_fill_2 FILLER_24_1204 ();
 sg13g2_fill_1 FILLER_24_1206 ();
 sg13g2_fill_1 FILLER_24_1216 ();
 sg13g2_fill_1 FILLER_24_1233 ();
 sg13g2_fill_2 FILLER_24_1305 ();
 sg13g2_fill_1 FILLER_24_1312 ();
 sg13g2_fill_1 FILLER_24_1324 ();
 sg13g2_decap_8 FILLER_24_1329 ();
 sg13g2_decap_4 FILLER_24_1336 ();
 sg13g2_fill_1 FILLER_24_1340 ();
 sg13g2_fill_2 FILLER_24_1367 ();
 sg13g2_fill_1 FILLER_24_1369 ();
 sg13g2_decap_8 FILLER_24_1422 ();
 sg13g2_decap_4 FILLER_24_1429 ();
 sg13g2_fill_2 FILLER_24_1433 ();
 sg13g2_decap_8 FILLER_24_1439 ();
 sg13g2_fill_1 FILLER_24_1446 ();
 sg13g2_fill_1 FILLER_24_1452 ();
 sg13g2_decap_8 FILLER_24_1458 ();
 sg13g2_fill_2 FILLER_24_1473 ();
 sg13g2_decap_8 FILLER_24_1506 ();
 sg13g2_fill_2 FILLER_24_1513 ();
 sg13g2_fill_1 FILLER_24_1515 ();
 sg13g2_fill_1 FILLER_24_1562 ();
 sg13g2_fill_2 FILLER_24_1572 ();
 sg13g2_fill_1 FILLER_24_1582 ();
 sg13g2_fill_2 FILLER_24_1612 ();
 sg13g2_fill_2 FILLER_24_1674 ();
 sg13g2_fill_2 FILLER_24_1684 ();
 sg13g2_fill_1 FILLER_24_1718 ();
 sg13g2_fill_2 FILLER_24_1769 ();
 sg13g2_fill_2 FILLER_24_1799 ();
 sg13g2_fill_2 FILLER_24_1839 ();
 sg13g2_fill_2 FILLER_24_1903 ();
 sg13g2_fill_2 FILLER_24_1949 ();
 sg13g2_fill_1 FILLER_24_1955 ();
 sg13g2_decap_4 FILLER_24_2028 ();
 sg13g2_fill_1 FILLER_24_2032 ();
 sg13g2_fill_1 FILLER_24_2066 ();
 sg13g2_decap_8 FILLER_24_2135 ();
 sg13g2_fill_1 FILLER_24_2142 ();
 sg13g2_decap_8 FILLER_24_2156 ();
 sg13g2_fill_1 FILLER_24_2163 ();
 sg13g2_fill_1 FILLER_24_2168 ();
 sg13g2_fill_2 FILLER_24_2179 ();
 sg13g2_fill_2 FILLER_24_2185 ();
 sg13g2_fill_1 FILLER_24_2187 ();
 sg13g2_fill_1 FILLER_24_2201 ();
 sg13g2_decap_4 FILLER_24_2233 ();
 sg13g2_fill_1 FILLER_24_2237 ();
 sg13g2_fill_2 FILLER_24_2243 ();
 sg13g2_fill_1 FILLER_24_2266 ();
 sg13g2_fill_2 FILLER_24_2308 ();
 sg13g2_fill_1 FILLER_24_2346 ();
 sg13g2_decap_8 FILLER_24_2373 ();
 sg13g2_decap_8 FILLER_24_2380 ();
 sg13g2_decap_8 FILLER_24_2387 ();
 sg13g2_decap_8 FILLER_24_2394 ();
 sg13g2_decap_8 FILLER_24_2401 ();
 sg13g2_decap_8 FILLER_24_2408 ();
 sg13g2_decap_8 FILLER_24_2415 ();
 sg13g2_decap_8 FILLER_24_2422 ();
 sg13g2_decap_8 FILLER_24_2429 ();
 sg13g2_decap_8 FILLER_24_2436 ();
 sg13g2_decap_8 FILLER_24_2443 ();
 sg13g2_decap_8 FILLER_24_2450 ();
 sg13g2_decap_8 FILLER_24_2457 ();
 sg13g2_decap_8 FILLER_24_2464 ();
 sg13g2_decap_8 FILLER_24_2471 ();
 sg13g2_decap_8 FILLER_24_2478 ();
 sg13g2_decap_8 FILLER_24_2485 ();
 sg13g2_decap_8 FILLER_24_2492 ();
 sg13g2_decap_8 FILLER_24_2499 ();
 sg13g2_decap_8 FILLER_24_2506 ();
 sg13g2_decap_8 FILLER_24_2513 ();
 sg13g2_decap_8 FILLER_24_2520 ();
 sg13g2_decap_8 FILLER_24_2527 ();
 sg13g2_decap_8 FILLER_24_2534 ();
 sg13g2_decap_8 FILLER_24_2541 ();
 sg13g2_decap_8 FILLER_24_2548 ();
 sg13g2_decap_8 FILLER_24_2555 ();
 sg13g2_decap_8 FILLER_24_2562 ();
 sg13g2_decap_8 FILLER_24_2569 ();
 sg13g2_decap_8 FILLER_24_2576 ();
 sg13g2_decap_8 FILLER_24_2583 ();
 sg13g2_decap_8 FILLER_24_2590 ();
 sg13g2_decap_8 FILLER_24_2597 ();
 sg13g2_decap_8 FILLER_24_2604 ();
 sg13g2_decap_8 FILLER_24_2611 ();
 sg13g2_decap_8 FILLER_24_2618 ();
 sg13g2_decap_8 FILLER_24_2625 ();
 sg13g2_decap_8 FILLER_24_2632 ();
 sg13g2_decap_8 FILLER_24_2639 ();
 sg13g2_decap_8 FILLER_24_2646 ();
 sg13g2_decap_8 FILLER_24_2653 ();
 sg13g2_decap_8 FILLER_24_2660 ();
 sg13g2_decap_8 FILLER_24_2667 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_decap_8 FILLER_25_427 ();
 sg13g2_decap_4 FILLER_25_434 ();
 sg13g2_fill_1 FILLER_25_438 ();
 sg13g2_fill_1 FILLER_25_496 ();
 sg13g2_fill_2 FILLER_25_501 ();
 sg13g2_fill_1 FILLER_25_503 ();
 sg13g2_fill_1 FILLER_25_514 ();
 sg13g2_fill_2 FILLER_25_525 ();
 sg13g2_fill_1 FILLER_25_556 ();
 sg13g2_fill_2 FILLER_25_566 ();
 sg13g2_fill_1 FILLER_25_568 ();
 sg13g2_fill_2 FILLER_25_595 ();
 sg13g2_fill_2 FILLER_25_614 ();
 sg13g2_fill_2 FILLER_25_681 ();
 sg13g2_fill_2 FILLER_25_740 ();
 sg13g2_fill_2 FILLER_25_821 ();
 sg13g2_fill_1 FILLER_25_871 ();
 sg13g2_fill_1 FILLER_25_893 ();
 sg13g2_fill_2 FILLER_25_904 ();
 sg13g2_fill_1 FILLER_25_906 ();
 sg13g2_fill_2 FILLER_25_912 ();
 sg13g2_decap_4 FILLER_25_918 ();
 sg13g2_fill_2 FILLER_25_922 ();
 sg13g2_fill_2 FILLER_25_933 ();
 sg13g2_fill_2 FILLER_25_939 ();
 sg13g2_fill_1 FILLER_25_941 ();
 sg13g2_decap_4 FILLER_25_972 ();
 sg13g2_fill_2 FILLER_25_993 ();
 sg13g2_fill_1 FILLER_25_995 ();
 sg13g2_fill_2 FILLER_25_1000 ();
 sg13g2_fill_1 FILLER_25_1002 ();
 sg13g2_fill_1 FILLER_25_1008 ();
 sg13g2_fill_2 FILLER_25_1145 ();
 sg13g2_fill_2 FILLER_25_1171 ();
 sg13g2_fill_1 FILLER_25_1218 ();
 sg13g2_decap_8 FILLER_25_1232 ();
 sg13g2_fill_1 FILLER_25_1239 ();
 sg13g2_fill_1 FILLER_25_1313 ();
 sg13g2_fill_1 FILLER_25_1328 ();
 sg13g2_decap_8 FILLER_25_1338 ();
 sg13g2_decap_4 FILLER_25_1345 ();
 sg13g2_fill_1 FILLER_25_1349 ();
 sg13g2_fill_1 FILLER_25_1359 ();
 sg13g2_fill_2 FILLER_25_1365 ();
 sg13g2_fill_2 FILLER_25_1372 ();
 sg13g2_fill_2 FILLER_25_1413 ();
 sg13g2_fill_2 FILLER_25_1451 ();
 sg13g2_fill_1 FILLER_25_1453 ();
 sg13g2_decap_8 FILLER_25_1527 ();
 sg13g2_fill_2 FILLER_25_1620 ();
 sg13g2_fill_1 FILLER_25_1683 ();
 sg13g2_decap_8 FILLER_25_1719 ();
 sg13g2_decap_8 FILLER_25_1738 ();
 sg13g2_fill_2 FILLER_25_1771 ();
 sg13g2_fill_1 FILLER_25_1773 ();
 sg13g2_decap_8 FILLER_25_1804 ();
 sg13g2_decap_4 FILLER_25_1815 ();
 sg13g2_decap_8 FILLER_25_1860 ();
 sg13g2_fill_1 FILLER_25_1867 ();
 sg13g2_fill_2 FILLER_25_1894 ();
 sg13g2_fill_1 FILLER_25_1896 ();
 sg13g2_fill_2 FILLER_25_1905 ();
 sg13g2_fill_1 FILLER_25_1907 ();
 sg13g2_fill_1 FILLER_25_1913 ();
 sg13g2_fill_2 FILLER_25_1923 ();
 sg13g2_fill_1 FILLER_25_1925 ();
 sg13g2_fill_1 FILLER_25_1939 ();
 sg13g2_decap_4 FILLER_25_1966 ();
 sg13g2_fill_2 FILLER_25_1974 ();
 sg13g2_fill_1 FILLER_25_1976 ();
 sg13g2_fill_2 FILLER_25_1982 ();
 sg13g2_fill_1 FILLER_25_1993 ();
 sg13g2_fill_2 FILLER_25_1999 ();
 sg13g2_fill_1 FILLER_25_2041 ();
 sg13g2_fill_2 FILLER_25_2060 ();
 sg13g2_fill_1 FILLER_25_2062 ();
 sg13g2_fill_2 FILLER_25_2075 ();
 sg13g2_fill_1 FILLER_25_2077 ();
 sg13g2_decap_4 FILLER_25_2082 ();
 sg13g2_fill_2 FILLER_25_2108 ();
 sg13g2_fill_2 FILLER_25_2142 ();
 sg13g2_fill_2 FILLER_25_2179 ();
 sg13g2_fill_1 FILLER_25_2212 ();
 sg13g2_fill_1 FILLER_25_2234 ();
 sg13g2_decap_4 FILLER_25_2275 ();
 sg13g2_fill_2 FILLER_25_2279 ();
 sg13g2_fill_2 FILLER_25_2290 ();
 sg13g2_fill_1 FILLER_25_2292 ();
 sg13g2_decap_8 FILLER_25_2297 ();
 sg13g2_fill_2 FILLER_25_2304 ();
 sg13g2_decap_8 FILLER_25_2315 ();
 sg13g2_decap_4 FILLER_25_2322 ();
 sg13g2_fill_2 FILLER_25_2326 ();
 sg13g2_fill_2 FILLER_25_2341 ();
 sg13g2_decap_4 FILLER_25_2352 ();
 sg13g2_decap_8 FILLER_25_2378 ();
 sg13g2_decap_8 FILLER_25_2385 ();
 sg13g2_decap_8 FILLER_25_2392 ();
 sg13g2_decap_8 FILLER_25_2399 ();
 sg13g2_decap_8 FILLER_25_2406 ();
 sg13g2_decap_8 FILLER_25_2413 ();
 sg13g2_decap_8 FILLER_25_2420 ();
 sg13g2_decap_8 FILLER_25_2427 ();
 sg13g2_decap_8 FILLER_25_2434 ();
 sg13g2_decap_8 FILLER_25_2441 ();
 sg13g2_decap_8 FILLER_25_2448 ();
 sg13g2_decap_8 FILLER_25_2455 ();
 sg13g2_decap_8 FILLER_25_2462 ();
 sg13g2_decap_8 FILLER_25_2469 ();
 sg13g2_decap_8 FILLER_25_2476 ();
 sg13g2_decap_8 FILLER_25_2483 ();
 sg13g2_decap_8 FILLER_25_2490 ();
 sg13g2_decap_8 FILLER_25_2497 ();
 sg13g2_decap_8 FILLER_25_2504 ();
 sg13g2_decap_8 FILLER_25_2511 ();
 sg13g2_decap_8 FILLER_25_2518 ();
 sg13g2_decap_8 FILLER_25_2525 ();
 sg13g2_decap_8 FILLER_25_2532 ();
 sg13g2_decap_8 FILLER_25_2539 ();
 sg13g2_decap_8 FILLER_25_2546 ();
 sg13g2_decap_8 FILLER_25_2553 ();
 sg13g2_decap_8 FILLER_25_2560 ();
 sg13g2_decap_8 FILLER_25_2567 ();
 sg13g2_decap_8 FILLER_25_2574 ();
 sg13g2_decap_8 FILLER_25_2581 ();
 sg13g2_decap_8 FILLER_25_2588 ();
 sg13g2_decap_8 FILLER_25_2595 ();
 sg13g2_decap_8 FILLER_25_2602 ();
 sg13g2_decap_8 FILLER_25_2609 ();
 sg13g2_decap_8 FILLER_25_2616 ();
 sg13g2_decap_8 FILLER_25_2623 ();
 sg13g2_decap_8 FILLER_25_2630 ();
 sg13g2_decap_8 FILLER_25_2637 ();
 sg13g2_decap_8 FILLER_25_2644 ();
 sg13g2_decap_8 FILLER_25_2651 ();
 sg13g2_decap_8 FILLER_25_2658 ();
 sg13g2_decap_8 FILLER_25_2665 ();
 sg13g2_fill_2 FILLER_25_2672 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_decap_8 FILLER_26_427 ();
 sg13g2_decap_8 FILLER_26_434 ();
 sg13g2_decap_4 FILLER_26_441 ();
 sg13g2_fill_1 FILLER_26_445 ();
 sg13g2_fill_1 FILLER_26_477 ();
 sg13g2_decap_8 FILLER_26_527 ();
 sg13g2_fill_2 FILLER_26_534 ();
 sg13g2_fill_1 FILLER_26_536 ();
 sg13g2_fill_1 FILLER_26_541 ();
 sg13g2_fill_2 FILLER_26_550 ();
 sg13g2_fill_2 FILLER_26_583 ();
 sg13g2_fill_2 FILLER_26_647 ();
 sg13g2_fill_1 FILLER_26_649 ();
 sg13g2_fill_2 FILLER_26_660 ();
 sg13g2_fill_1 FILLER_26_662 ();
 sg13g2_fill_2 FILLER_26_766 ();
 sg13g2_fill_1 FILLER_26_768 ();
 sg13g2_fill_2 FILLER_26_793 ();
 sg13g2_fill_1 FILLER_26_795 ();
 sg13g2_fill_2 FILLER_26_813 ();
 sg13g2_fill_1 FILLER_26_815 ();
 sg13g2_fill_2 FILLER_26_852 ();
 sg13g2_fill_1 FILLER_26_854 ();
 sg13g2_fill_1 FILLER_26_908 ();
 sg13g2_decap_4 FILLER_26_925 ();
 sg13g2_fill_1 FILLER_26_929 ();
 sg13g2_decap_4 FILLER_26_934 ();
 sg13g2_fill_2 FILLER_26_938 ();
 sg13g2_fill_1 FILLER_26_946 ();
 sg13g2_fill_1 FILLER_26_957 ();
 sg13g2_fill_2 FILLER_26_967 ();
 sg13g2_fill_1 FILLER_26_1009 ();
 sg13g2_fill_2 FILLER_26_1036 ();
 sg13g2_fill_1 FILLER_26_1038 ();
 sg13g2_fill_2 FILLER_26_1064 ();
 sg13g2_fill_1 FILLER_26_1066 ();
 sg13g2_fill_1 FILLER_26_1076 ();
 sg13g2_fill_2 FILLER_26_1086 ();
 sg13g2_fill_2 FILLER_26_1115 ();
 sg13g2_fill_1 FILLER_26_1122 ();
 sg13g2_decap_8 FILLER_26_1145 ();
 sg13g2_fill_2 FILLER_26_1157 ();
 sg13g2_decap_4 FILLER_26_1236 ();
 sg13g2_fill_1 FILLER_26_1266 ();
 sg13g2_fill_2 FILLER_26_1301 ();
 sg13g2_fill_1 FILLER_26_1303 ();
 sg13g2_fill_2 FILLER_26_1318 ();
 sg13g2_fill_1 FILLER_26_1320 ();
 sg13g2_decap_8 FILLER_26_1324 ();
 sg13g2_fill_2 FILLER_26_1331 ();
 sg13g2_fill_1 FILLER_26_1333 ();
 sg13g2_fill_2 FILLER_26_1338 ();
 sg13g2_fill_1 FILLER_26_1391 ();
 sg13g2_fill_2 FILLER_26_1396 ();
 sg13g2_fill_1 FILLER_26_1398 ();
 sg13g2_fill_1 FILLER_26_1417 ();
 sg13g2_fill_1 FILLER_26_1491 ();
 sg13g2_fill_1 FILLER_26_1541 ();
 sg13g2_fill_1 FILLER_26_1568 ();
 sg13g2_decap_4 FILLER_26_1595 ();
 sg13g2_decap_4 FILLER_26_1635 ();
 sg13g2_fill_1 FILLER_26_1685 ();
 sg13g2_fill_2 FILLER_26_1709 ();
 sg13g2_fill_1 FILLER_26_1720 ();
 sg13g2_fill_2 FILLER_26_1738 ();
 sg13g2_fill_2 FILLER_26_1759 ();
 sg13g2_fill_1 FILLER_26_1761 ();
 sg13g2_fill_2 FILLER_26_1781 ();
 sg13g2_fill_2 FILLER_26_1835 ();
 sg13g2_fill_2 FILLER_26_1876 ();
 sg13g2_fill_2 FILLER_26_1896 ();
 sg13g2_fill_1 FILLER_26_1898 ();
 sg13g2_fill_1 FILLER_26_1921 ();
 sg13g2_fill_1 FILLER_26_1931 ();
 sg13g2_fill_1 FILLER_26_1941 ();
 sg13g2_decap_8 FILLER_26_1951 ();
 sg13g2_fill_2 FILLER_26_1958 ();
 sg13g2_fill_2 FILLER_26_2007 ();
 sg13g2_fill_1 FILLER_26_2009 ();
 sg13g2_decap_8 FILLER_26_2071 ();
 sg13g2_fill_1 FILLER_26_2078 ();
 sg13g2_decap_4 FILLER_26_2105 ();
 sg13g2_fill_1 FILLER_26_2109 ();
 sg13g2_decap_8 FILLER_26_2113 ();
 sg13g2_decap_8 FILLER_26_2120 ();
 sg13g2_fill_2 FILLER_26_2127 ();
 sg13g2_fill_1 FILLER_26_2129 ();
 sg13g2_fill_2 FILLER_26_2139 ();
 sg13g2_fill_1 FILLER_26_2141 ();
 sg13g2_decap_4 FILLER_26_2151 ();
 sg13g2_fill_2 FILLER_26_2198 ();
 sg13g2_fill_1 FILLER_26_2200 ();
 sg13g2_fill_1 FILLER_26_2227 ();
 sg13g2_decap_4 FILLER_26_2237 ();
 sg13g2_fill_2 FILLER_26_2241 ();
 sg13g2_fill_2 FILLER_26_2279 ();
 sg13g2_fill_1 FILLER_26_2281 ();
 sg13g2_fill_2 FILLER_26_2308 ();
 sg13g2_fill_1 FILLER_26_2320 ();
 sg13g2_decap_8 FILLER_26_2374 ();
 sg13g2_decap_8 FILLER_26_2381 ();
 sg13g2_decap_8 FILLER_26_2388 ();
 sg13g2_decap_8 FILLER_26_2395 ();
 sg13g2_decap_8 FILLER_26_2402 ();
 sg13g2_decap_8 FILLER_26_2409 ();
 sg13g2_decap_8 FILLER_26_2416 ();
 sg13g2_decap_8 FILLER_26_2423 ();
 sg13g2_decap_8 FILLER_26_2430 ();
 sg13g2_decap_8 FILLER_26_2437 ();
 sg13g2_decap_8 FILLER_26_2444 ();
 sg13g2_decap_8 FILLER_26_2451 ();
 sg13g2_decap_8 FILLER_26_2458 ();
 sg13g2_decap_8 FILLER_26_2465 ();
 sg13g2_decap_8 FILLER_26_2472 ();
 sg13g2_decap_8 FILLER_26_2479 ();
 sg13g2_decap_8 FILLER_26_2486 ();
 sg13g2_decap_8 FILLER_26_2493 ();
 sg13g2_decap_8 FILLER_26_2500 ();
 sg13g2_decap_8 FILLER_26_2507 ();
 sg13g2_decap_8 FILLER_26_2514 ();
 sg13g2_decap_8 FILLER_26_2521 ();
 sg13g2_decap_8 FILLER_26_2528 ();
 sg13g2_decap_8 FILLER_26_2535 ();
 sg13g2_decap_8 FILLER_26_2542 ();
 sg13g2_decap_8 FILLER_26_2549 ();
 sg13g2_decap_8 FILLER_26_2556 ();
 sg13g2_decap_8 FILLER_26_2563 ();
 sg13g2_decap_8 FILLER_26_2570 ();
 sg13g2_decap_8 FILLER_26_2577 ();
 sg13g2_decap_8 FILLER_26_2584 ();
 sg13g2_decap_8 FILLER_26_2591 ();
 sg13g2_decap_8 FILLER_26_2598 ();
 sg13g2_decap_8 FILLER_26_2605 ();
 sg13g2_decap_8 FILLER_26_2612 ();
 sg13g2_decap_8 FILLER_26_2619 ();
 sg13g2_decap_8 FILLER_26_2626 ();
 sg13g2_decap_8 FILLER_26_2633 ();
 sg13g2_decap_8 FILLER_26_2640 ();
 sg13g2_decap_8 FILLER_26_2647 ();
 sg13g2_decap_8 FILLER_26_2654 ();
 sg13g2_decap_8 FILLER_26_2661 ();
 sg13g2_decap_4 FILLER_26_2668 ();
 sg13g2_fill_2 FILLER_26_2672 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_fill_2 FILLER_27_427 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_fill_2 FILLER_27_456 ();
 sg13g2_fill_1 FILLER_27_488 ();
 sg13g2_decap_4 FILLER_27_507 ();
 sg13g2_fill_2 FILLER_27_532 ();
 sg13g2_fill_1 FILLER_27_543 ();
 sg13g2_decap_4 FILLER_27_548 ();
 sg13g2_decap_4 FILLER_27_567 ();
 sg13g2_fill_1 FILLER_27_580 ();
 sg13g2_decap_4 FILLER_27_589 ();
 sg13g2_fill_1 FILLER_27_598 ();
 sg13g2_fill_1 FILLER_27_603 ();
 sg13g2_decap_8 FILLER_27_612 ();
 sg13g2_fill_2 FILLER_27_619 ();
 sg13g2_fill_1 FILLER_27_621 ();
 sg13g2_fill_2 FILLER_27_627 ();
 sg13g2_fill_2 FILLER_27_637 ();
 sg13g2_fill_2 FILLER_27_647 ();
 sg13g2_fill_1 FILLER_27_649 ();
 sg13g2_fill_2 FILLER_27_655 ();
 sg13g2_fill_1 FILLER_27_657 ();
 sg13g2_fill_1 FILLER_27_663 ();
 sg13g2_fill_2 FILLER_27_673 ();
 sg13g2_fill_2 FILLER_27_679 ();
 sg13g2_fill_1 FILLER_27_681 ();
 sg13g2_fill_1 FILLER_27_713 ();
 sg13g2_fill_2 FILLER_27_745 ();
 sg13g2_fill_2 FILLER_27_759 ();
 sg13g2_fill_1 FILLER_27_778 ();
 sg13g2_fill_2 FILLER_27_815 ();
 sg13g2_fill_2 FILLER_27_827 ();
 sg13g2_fill_1 FILLER_27_829 ();
 sg13g2_fill_1 FILLER_27_835 ();
 sg13g2_fill_2 FILLER_27_855 ();
 sg13g2_fill_1 FILLER_27_870 ();
 sg13g2_fill_2 FILLER_27_884 ();
 sg13g2_decap_4 FILLER_27_895 ();
 sg13g2_decap_4 FILLER_27_913 ();
 sg13g2_fill_2 FILLER_27_948 ();
 sg13g2_fill_1 FILLER_27_950 ();
 sg13g2_fill_1 FILLER_27_990 ();
 sg13g2_fill_1 FILLER_27_996 ();
 sg13g2_fill_1 FILLER_27_1020 ();
 sg13g2_fill_2 FILLER_27_1046 ();
 sg13g2_fill_2 FILLER_27_1078 ();
 sg13g2_fill_1 FILLER_27_1080 ();
 sg13g2_fill_2 FILLER_27_1168 ();
 sg13g2_fill_1 FILLER_27_1170 ();
 sg13g2_fill_1 FILLER_27_1202 ();
 sg13g2_fill_2 FILLER_27_1312 ();
 sg13g2_fill_2 FILLER_27_1357 ();
 sg13g2_fill_2 FILLER_27_1378 ();
 sg13g2_fill_1 FILLER_27_1380 ();
 sg13g2_fill_1 FILLER_27_1416 ();
 sg13g2_fill_1 FILLER_27_1421 ();
 sg13g2_fill_2 FILLER_27_1445 ();
 sg13g2_fill_1 FILLER_27_1447 ();
 sg13g2_fill_2 FILLER_27_1524 ();
 sg13g2_decap_8 FILLER_27_1596 ();
 sg13g2_decap_8 FILLER_27_1603 ();
 sg13g2_decap_4 FILLER_27_1614 ();
 sg13g2_decap_8 FILLER_27_1622 ();
 sg13g2_fill_2 FILLER_27_1629 ();
 sg13g2_decap_4 FILLER_27_1644 ();
 sg13g2_fill_2 FILLER_27_1648 ();
 sg13g2_fill_2 FILLER_27_1654 ();
 sg13g2_fill_1 FILLER_27_1697 ();
 sg13g2_fill_2 FILLER_27_1743 ();
 sg13g2_fill_2 FILLER_27_1753 ();
 sg13g2_fill_1 FILLER_27_1755 ();
 sg13g2_fill_1 FILLER_27_1800 ();
 sg13g2_fill_1 FILLER_27_1856 ();
 sg13g2_fill_1 FILLER_27_1960 ();
 sg13g2_fill_1 FILLER_27_1970 ();
 sg13g2_decap_8 FILLER_27_1976 ();
 sg13g2_fill_2 FILLER_27_1983 ();
 sg13g2_fill_1 FILLER_27_1985 ();
 sg13g2_fill_2 FILLER_27_1990 ();
 sg13g2_fill_1 FILLER_27_1992 ();
 sg13g2_decap_8 FILLER_27_2062 ();
 sg13g2_fill_1 FILLER_27_2069 ();
 sg13g2_fill_2 FILLER_27_2104 ();
 sg13g2_fill_1 FILLER_27_2106 ();
 sg13g2_fill_1 FILLER_27_2130 ();
 sg13g2_fill_2 FILLER_27_2141 ();
 sg13g2_fill_1 FILLER_27_2143 ();
 sg13g2_fill_2 FILLER_27_2149 ();
 sg13g2_fill_2 FILLER_27_2156 ();
 sg13g2_fill_2 FILLER_27_2172 ();
 sg13g2_fill_1 FILLER_27_2196 ();
 sg13g2_fill_2 FILLER_27_2211 ();
 sg13g2_fill_1 FILLER_27_2213 ();
 sg13g2_fill_2 FILLER_27_2249 ();
 sg13g2_decap_4 FILLER_27_2255 ();
 sg13g2_fill_1 FILLER_27_2281 ();
 sg13g2_fill_1 FILLER_27_2304 ();
 sg13g2_decap_8 FILLER_27_2349 ();
 sg13g2_decap_8 FILLER_27_2373 ();
 sg13g2_decap_8 FILLER_27_2380 ();
 sg13g2_decap_8 FILLER_27_2387 ();
 sg13g2_decap_8 FILLER_27_2394 ();
 sg13g2_decap_8 FILLER_27_2401 ();
 sg13g2_decap_8 FILLER_27_2408 ();
 sg13g2_decap_8 FILLER_27_2415 ();
 sg13g2_decap_8 FILLER_27_2422 ();
 sg13g2_decap_8 FILLER_27_2429 ();
 sg13g2_decap_8 FILLER_27_2436 ();
 sg13g2_decap_8 FILLER_27_2443 ();
 sg13g2_decap_8 FILLER_27_2450 ();
 sg13g2_decap_8 FILLER_27_2457 ();
 sg13g2_decap_8 FILLER_27_2464 ();
 sg13g2_decap_8 FILLER_27_2471 ();
 sg13g2_decap_8 FILLER_27_2478 ();
 sg13g2_decap_8 FILLER_27_2485 ();
 sg13g2_decap_8 FILLER_27_2492 ();
 sg13g2_decap_8 FILLER_27_2499 ();
 sg13g2_decap_8 FILLER_27_2506 ();
 sg13g2_decap_8 FILLER_27_2513 ();
 sg13g2_decap_8 FILLER_27_2520 ();
 sg13g2_decap_8 FILLER_27_2527 ();
 sg13g2_decap_8 FILLER_27_2534 ();
 sg13g2_decap_8 FILLER_27_2541 ();
 sg13g2_decap_8 FILLER_27_2548 ();
 sg13g2_decap_8 FILLER_27_2555 ();
 sg13g2_decap_8 FILLER_27_2562 ();
 sg13g2_decap_8 FILLER_27_2569 ();
 sg13g2_decap_8 FILLER_27_2576 ();
 sg13g2_decap_8 FILLER_27_2583 ();
 sg13g2_decap_8 FILLER_27_2590 ();
 sg13g2_decap_8 FILLER_27_2597 ();
 sg13g2_decap_8 FILLER_27_2604 ();
 sg13g2_decap_8 FILLER_27_2611 ();
 sg13g2_decap_8 FILLER_27_2618 ();
 sg13g2_decap_8 FILLER_27_2625 ();
 sg13g2_decap_8 FILLER_27_2632 ();
 sg13g2_decap_8 FILLER_27_2639 ();
 sg13g2_decap_8 FILLER_27_2646 ();
 sg13g2_decap_8 FILLER_27_2653 ();
 sg13g2_decap_8 FILLER_27_2660 ();
 sg13g2_decap_8 FILLER_27_2667 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_420 ();
 sg13g2_fill_2 FILLER_28_427 ();
 sg13g2_fill_1 FILLER_28_465 ();
 sg13g2_fill_2 FILLER_28_475 ();
 sg13g2_fill_2 FILLER_28_482 ();
 sg13g2_fill_1 FILLER_28_501 ();
 sg13g2_fill_2 FILLER_28_507 ();
 sg13g2_fill_1 FILLER_28_509 ();
 sg13g2_fill_2 FILLER_28_519 ();
 sg13g2_decap_4 FILLER_28_529 ();
 sg13g2_fill_1 FILLER_28_587 ();
 sg13g2_decap_4 FILLER_28_598 ();
 sg13g2_decap_4 FILLER_28_610 ();
 sg13g2_fill_2 FILLER_28_614 ();
 sg13g2_decap_4 FILLER_28_651 ();
 sg13g2_fill_2 FILLER_28_700 ();
 sg13g2_fill_1 FILLER_28_716 ();
 sg13g2_fill_1 FILLER_28_740 ();
 sg13g2_fill_2 FILLER_28_816 ();
 sg13g2_fill_1 FILLER_28_818 ();
 sg13g2_fill_1 FILLER_28_845 ();
 sg13g2_fill_2 FILLER_28_881 ();
 sg13g2_fill_1 FILLER_28_883 ();
 sg13g2_fill_1 FILLER_28_928 ();
 sg13g2_fill_2 FILLER_28_991 ();
 sg13g2_fill_1 FILLER_28_993 ();
 sg13g2_decap_4 FILLER_28_1024 ();
 sg13g2_fill_1 FILLER_28_1028 ();
 sg13g2_decap_8 FILLER_28_1037 ();
 sg13g2_fill_2 FILLER_28_1053 ();
 sg13g2_fill_1 FILLER_28_1055 ();
 sg13g2_fill_2 FILLER_28_1095 ();
 sg13g2_fill_1 FILLER_28_1097 ();
 sg13g2_fill_2 FILLER_28_1113 ();
 sg13g2_fill_1 FILLER_28_1115 ();
 sg13g2_decap_4 FILLER_28_1158 ();
 sg13g2_fill_1 FILLER_28_1162 ();
 sg13g2_fill_2 FILLER_28_1215 ();
 sg13g2_fill_2 FILLER_28_1245 ();
 sg13g2_decap_8 FILLER_28_1255 ();
 sg13g2_decap_4 FILLER_28_1262 ();
 sg13g2_decap_4 FILLER_28_1271 ();
 sg13g2_fill_1 FILLER_28_1349 ();
 sg13g2_decap_8 FILLER_28_1401 ();
 sg13g2_fill_1 FILLER_28_1416 ();
 sg13g2_fill_2 FILLER_28_1464 ();
 sg13g2_fill_1 FILLER_28_1466 ();
 sg13g2_fill_2 FILLER_28_1484 ();
 sg13g2_fill_1 FILLER_28_1486 ();
 sg13g2_fill_2 FILLER_28_1500 ();
 sg13g2_fill_1 FILLER_28_1502 ();
 sg13g2_fill_2 FILLER_28_1524 ();
 sg13g2_fill_1 FILLER_28_1526 ();
 sg13g2_fill_2 FILLER_28_1576 ();
 sg13g2_fill_1 FILLER_28_1578 ();
 sg13g2_fill_1 FILLER_28_1614 ();
 sg13g2_fill_2 FILLER_28_1633 ();
 sg13g2_decap_8 FILLER_28_1639 ();
 sg13g2_decap_8 FILLER_28_1646 ();
 sg13g2_decap_4 FILLER_28_1653 ();
 sg13g2_decap_8 FILLER_28_1661 ();
 sg13g2_decap_4 FILLER_28_1676 ();
 sg13g2_fill_2 FILLER_28_1680 ();
 sg13g2_decap_4 FILLER_28_1686 ();
 sg13g2_fill_2 FILLER_28_1707 ();
 sg13g2_decap_8 FILLER_28_1718 ();
 sg13g2_fill_2 FILLER_28_1761 ();
 sg13g2_fill_1 FILLER_28_1763 ();
 sg13g2_fill_2 FILLER_28_1769 ();
 sg13g2_fill_1 FILLER_28_1771 ();
 sg13g2_decap_4 FILLER_28_1811 ();
 sg13g2_fill_1 FILLER_28_1815 ();
 sg13g2_fill_2 FILLER_28_1833 ();
 sg13g2_fill_1 FILLER_28_1835 ();
 sg13g2_fill_1 FILLER_28_1841 ();
 sg13g2_fill_2 FILLER_28_1855 ();
 sg13g2_fill_2 FILLER_28_1866 ();
 sg13g2_fill_2 FILLER_28_1894 ();
 sg13g2_fill_1 FILLER_28_1896 ();
 sg13g2_fill_1 FILLER_28_1910 ();
 sg13g2_fill_1 FILLER_28_1916 ();
 sg13g2_fill_1 FILLER_28_1940 ();
 sg13g2_fill_2 FILLER_28_1972 ();
 sg13g2_fill_2 FILLER_28_1978 ();
 sg13g2_fill_1 FILLER_28_1980 ();
 sg13g2_fill_2 FILLER_28_2012 ();
 sg13g2_fill_1 FILLER_28_2014 ();
 sg13g2_fill_2 FILLER_28_2024 ();
 sg13g2_fill_1 FILLER_28_2026 ();
 sg13g2_fill_2 FILLER_28_2036 ();
 sg13g2_fill_2 FILLER_28_2074 ();
 sg13g2_fill_1 FILLER_28_2076 ();
 sg13g2_decap_8 FILLER_28_2096 ();
 sg13g2_fill_2 FILLER_28_2103 ();
 sg13g2_fill_1 FILLER_28_2105 ();
 sg13g2_fill_2 FILLER_28_2113 ();
 sg13g2_decap_4 FILLER_28_2123 ();
 sg13g2_fill_1 FILLER_28_2127 ();
 sg13g2_fill_2 FILLER_28_2154 ();
 sg13g2_fill_1 FILLER_28_2182 ();
 sg13g2_fill_1 FILLER_28_2226 ();
 sg13g2_fill_1 FILLER_28_2240 ();
 sg13g2_fill_1 FILLER_28_2246 ();
 sg13g2_fill_1 FILLER_28_2299 ();
 sg13g2_fill_2 FILLER_28_2305 ();
 sg13g2_fill_2 FILLER_28_2321 ();
 sg13g2_fill_1 FILLER_28_2323 ();
 sg13g2_decap_8 FILLER_28_2373 ();
 sg13g2_decap_8 FILLER_28_2380 ();
 sg13g2_decap_8 FILLER_28_2387 ();
 sg13g2_decap_8 FILLER_28_2394 ();
 sg13g2_decap_8 FILLER_28_2401 ();
 sg13g2_decap_8 FILLER_28_2408 ();
 sg13g2_decap_8 FILLER_28_2415 ();
 sg13g2_decap_8 FILLER_28_2422 ();
 sg13g2_decap_8 FILLER_28_2429 ();
 sg13g2_decap_8 FILLER_28_2436 ();
 sg13g2_decap_8 FILLER_28_2443 ();
 sg13g2_decap_8 FILLER_28_2450 ();
 sg13g2_decap_8 FILLER_28_2457 ();
 sg13g2_decap_8 FILLER_28_2464 ();
 sg13g2_decap_8 FILLER_28_2471 ();
 sg13g2_decap_8 FILLER_28_2478 ();
 sg13g2_decap_8 FILLER_28_2485 ();
 sg13g2_decap_8 FILLER_28_2492 ();
 sg13g2_decap_8 FILLER_28_2499 ();
 sg13g2_decap_8 FILLER_28_2506 ();
 sg13g2_decap_8 FILLER_28_2513 ();
 sg13g2_decap_8 FILLER_28_2520 ();
 sg13g2_decap_8 FILLER_28_2527 ();
 sg13g2_decap_8 FILLER_28_2534 ();
 sg13g2_decap_8 FILLER_28_2541 ();
 sg13g2_decap_8 FILLER_28_2548 ();
 sg13g2_decap_8 FILLER_28_2555 ();
 sg13g2_decap_8 FILLER_28_2562 ();
 sg13g2_decap_8 FILLER_28_2569 ();
 sg13g2_decap_8 FILLER_28_2576 ();
 sg13g2_decap_8 FILLER_28_2583 ();
 sg13g2_decap_8 FILLER_28_2590 ();
 sg13g2_decap_8 FILLER_28_2597 ();
 sg13g2_decap_8 FILLER_28_2604 ();
 sg13g2_decap_8 FILLER_28_2611 ();
 sg13g2_decap_8 FILLER_28_2618 ();
 sg13g2_decap_8 FILLER_28_2625 ();
 sg13g2_decap_8 FILLER_28_2632 ();
 sg13g2_decap_8 FILLER_28_2639 ();
 sg13g2_decap_8 FILLER_28_2646 ();
 sg13g2_decap_8 FILLER_28_2653 ();
 sg13g2_decap_8 FILLER_28_2660 ();
 sg13g2_decap_8 FILLER_28_2667 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_decap_8 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_fill_2 FILLER_29_420 ();
 sg13g2_fill_2 FILLER_29_462 ();
 sg13g2_fill_1 FILLER_29_499 ();
 sg13g2_fill_1 FILLER_29_508 ();
 sg13g2_fill_2 FILLER_29_544 ();
 sg13g2_fill_2 FILLER_29_555 ();
 sg13g2_fill_1 FILLER_29_557 ();
 sg13g2_decap_4 FILLER_29_631 ();
 sg13g2_fill_2 FILLER_29_635 ();
 sg13g2_decap_4 FILLER_29_658 ();
 sg13g2_fill_1 FILLER_29_667 ();
 sg13g2_fill_1 FILLER_29_756 ();
 sg13g2_fill_2 FILLER_29_766 ();
 sg13g2_fill_1 FILLER_29_768 ();
 sg13g2_fill_2 FILLER_29_820 ();
 sg13g2_fill_2 FILLER_29_827 ();
 sg13g2_fill_2 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_843 ();
 sg13g2_fill_1 FILLER_29_855 ();
 sg13g2_fill_1 FILLER_29_864 ();
 sg13g2_fill_2 FILLER_29_870 ();
 sg13g2_fill_1 FILLER_29_887 ();
 sg13g2_decap_8 FILLER_29_892 ();
 sg13g2_fill_1 FILLER_29_899 ();
 sg13g2_fill_1 FILLER_29_904 ();
 sg13g2_fill_1 FILLER_29_910 ();
 sg13g2_fill_2 FILLER_29_915 ();
 sg13g2_fill_1 FILLER_29_921 ();
 sg13g2_fill_2 FILLER_29_927 ();
 sg13g2_fill_1 FILLER_29_929 ();
 sg13g2_fill_2 FILLER_29_994 ();
 sg13g2_fill_1 FILLER_29_1001 ();
 sg13g2_decap_4 FILLER_29_1016 ();
 sg13g2_fill_1 FILLER_29_1020 ();
 sg13g2_fill_2 FILLER_29_1034 ();
 sg13g2_fill_1 FILLER_29_1036 ();
 sg13g2_decap_4 FILLER_29_1090 ();
 sg13g2_fill_2 FILLER_29_1094 ();
 sg13g2_fill_2 FILLER_29_1139 ();
 sg13g2_fill_1 FILLER_29_1141 ();
 sg13g2_fill_1 FILLER_29_1168 ();
 sg13g2_fill_2 FILLER_29_1187 ();
 sg13g2_fill_1 FILLER_29_1189 ();
 sg13g2_fill_2 FILLER_29_1233 ();
 sg13g2_fill_1 FILLER_29_1235 ();
 sg13g2_fill_2 FILLER_29_1266 ();
 sg13g2_fill_1 FILLER_29_1268 ();
 sg13g2_fill_1 FILLER_29_1289 ();
 sg13g2_fill_2 FILLER_29_1302 ();
 sg13g2_fill_1 FILLER_29_1304 ();
 sg13g2_fill_2 FILLER_29_1331 ();
 sg13g2_fill_2 FILLER_29_1358 ();
 sg13g2_fill_1 FILLER_29_1360 ();
 sg13g2_decap_4 FILLER_29_1369 ();
 sg13g2_fill_1 FILLER_29_1408 ();
 sg13g2_fill_2 FILLER_29_1418 ();
 sg13g2_fill_1 FILLER_29_1424 ();
 sg13g2_decap_4 FILLER_29_1438 ();
 sg13g2_fill_1 FILLER_29_1442 ();
 sg13g2_decap_8 FILLER_29_1448 ();
 sg13g2_decap_4 FILLER_29_1455 ();
 sg13g2_fill_1 FILLER_29_1459 ();
 sg13g2_fill_1 FILLER_29_1468 ();
 sg13g2_fill_1 FILLER_29_1473 ();
 sg13g2_fill_2 FILLER_29_1544 ();
 sg13g2_fill_1 FILLER_29_1546 ();
 sg13g2_fill_2 FILLER_29_1582 ();
 sg13g2_fill_1 FILLER_29_1584 ();
 sg13g2_fill_2 FILLER_29_1610 ();
 sg13g2_fill_1 FILLER_29_1623 ();
 sg13g2_fill_1 FILLER_29_1664 ();
 sg13g2_fill_2 FILLER_29_1673 ();
 sg13g2_decap_4 FILLER_29_1716 ();
 sg13g2_decap_4 FILLER_29_1733 ();
 sg13g2_fill_1 FILLER_29_1737 ();
 sg13g2_fill_2 FILLER_29_1795 ();
 sg13g2_fill_1 FILLER_29_1836 ();
 sg13g2_fill_1 FILLER_29_1842 ();
 sg13g2_fill_1 FILLER_29_1962 ();
 sg13g2_fill_2 FILLER_29_2004 ();
 sg13g2_fill_1 FILLER_29_2040 ();
 sg13g2_fill_2 FILLER_29_2050 ();
 sg13g2_fill_1 FILLER_29_2052 ();
 sg13g2_decap_8 FILLER_29_2082 ();
 sg13g2_decap_8 FILLER_29_2089 ();
 sg13g2_fill_1 FILLER_29_2101 ();
 sg13g2_fill_1 FILLER_29_2146 ();
 sg13g2_fill_2 FILLER_29_2170 ();
 sg13g2_fill_2 FILLER_29_2176 ();
 sg13g2_fill_1 FILLER_29_2178 ();
 sg13g2_fill_1 FILLER_29_2198 ();
 sg13g2_fill_2 FILLER_29_2203 ();
 sg13g2_fill_2 FILLER_29_2225 ();
 sg13g2_fill_1 FILLER_29_2227 ();
 sg13g2_fill_1 FILLER_29_2233 ();
 sg13g2_decap_4 FILLER_29_2282 ();
 sg13g2_fill_1 FILLER_29_2286 ();
 sg13g2_fill_1 FILLER_29_2322 ();
 sg13g2_decap_8 FILLER_29_2361 ();
 sg13g2_decap_8 FILLER_29_2368 ();
 sg13g2_decap_8 FILLER_29_2375 ();
 sg13g2_decap_8 FILLER_29_2382 ();
 sg13g2_decap_8 FILLER_29_2389 ();
 sg13g2_decap_8 FILLER_29_2396 ();
 sg13g2_decap_8 FILLER_29_2403 ();
 sg13g2_decap_8 FILLER_29_2410 ();
 sg13g2_decap_8 FILLER_29_2417 ();
 sg13g2_decap_8 FILLER_29_2424 ();
 sg13g2_decap_8 FILLER_29_2431 ();
 sg13g2_decap_8 FILLER_29_2438 ();
 sg13g2_decap_8 FILLER_29_2445 ();
 sg13g2_decap_8 FILLER_29_2452 ();
 sg13g2_decap_8 FILLER_29_2459 ();
 sg13g2_decap_8 FILLER_29_2466 ();
 sg13g2_decap_8 FILLER_29_2473 ();
 sg13g2_decap_8 FILLER_29_2480 ();
 sg13g2_decap_8 FILLER_29_2487 ();
 sg13g2_decap_8 FILLER_29_2494 ();
 sg13g2_decap_8 FILLER_29_2501 ();
 sg13g2_decap_8 FILLER_29_2508 ();
 sg13g2_decap_8 FILLER_29_2515 ();
 sg13g2_decap_8 FILLER_29_2522 ();
 sg13g2_decap_8 FILLER_29_2529 ();
 sg13g2_decap_8 FILLER_29_2536 ();
 sg13g2_decap_8 FILLER_29_2543 ();
 sg13g2_decap_8 FILLER_29_2550 ();
 sg13g2_decap_8 FILLER_29_2557 ();
 sg13g2_decap_8 FILLER_29_2564 ();
 sg13g2_decap_8 FILLER_29_2571 ();
 sg13g2_decap_8 FILLER_29_2578 ();
 sg13g2_decap_8 FILLER_29_2585 ();
 sg13g2_decap_8 FILLER_29_2592 ();
 sg13g2_decap_8 FILLER_29_2599 ();
 sg13g2_decap_8 FILLER_29_2606 ();
 sg13g2_decap_8 FILLER_29_2613 ();
 sg13g2_decap_8 FILLER_29_2620 ();
 sg13g2_decap_8 FILLER_29_2627 ();
 sg13g2_decap_8 FILLER_29_2634 ();
 sg13g2_decap_8 FILLER_29_2641 ();
 sg13g2_decap_8 FILLER_29_2648 ();
 sg13g2_decap_8 FILLER_29_2655 ();
 sg13g2_decap_8 FILLER_29_2662 ();
 sg13g2_decap_4 FILLER_29_2669 ();
 sg13g2_fill_1 FILLER_29_2673 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_decap_8 FILLER_30_427 ();
 sg13g2_decap_4 FILLER_30_434 ();
 sg13g2_fill_1 FILLER_30_438 ();
 sg13g2_decap_4 FILLER_30_443 ();
 sg13g2_fill_1 FILLER_30_447 ();
 sg13g2_fill_2 FILLER_30_453 ();
 sg13g2_fill_1 FILLER_30_455 ();
 sg13g2_fill_2 FILLER_30_465 ();
 sg13g2_fill_2 FILLER_30_471 ();
 sg13g2_fill_1 FILLER_30_473 ();
 sg13g2_fill_2 FILLER_30_509 ();
 sg13g2_fill_1 FILLER_30_511 ();
 sg13g2_fill_2 FILLER_30_586 ();
 sg13g2_fill_2 FILLER_30_628 ();
 sg13g2_fill_1 FILLER_30_630 ();
 sg13g2_fill_2 FILLER_30_639 ();
 sg13g2_fill_1 FILLER_30_706 ();
 sg13g2_fill_2 FILLER_30_711 ();
 sg13g2_fill_2 FILLER_30_737 ();
 sg13g2_fill_1 FILLER_30_739 ();
 sg13g2_fill_1 FILLER_30_846 ();
 sg13g2_fill_2 FILLER_30_904 ();
 sg13g2_fill_2 FILLER_30_954 ();
 sg13g2_fill_1 FILLER_30_956 ();
 sg13g2_fill_2 FILLER_30_966 ();
 sg13g2_fill_1 FILLER_30_968 ();
 sg13g2_fill_1 FILLER_30_1038 ();
 sg13g2_decap_4 FILLER_30_1044 ();
 sg13g2_decap_8 FILLER_30_1095 ();
 sg13g2_fill_1 FILLER_30_1102 ();
 sg13g2_fill_1 FILLER_30_1108 ();
 sg13g2_fill_2 FILLER_30_1118 ();
 sg13g2_fill_1 FILLER_30_1120 ();
 sg13g2_fill_1 FILLER_30_1125 ();
 sg13g2_fill_2 FILLER_30_1154 ();
 sg13g2_fill_2 FILLER_30_1168 ();
 sg13g2_fill_1 FILLER_30_1170 ();
 sg13g2_fill_1 FILLER_30_1185 ();
 sg13g2_fill_1 FILLER_30_1190 ();
 sg13g2_fill_2 FILLER_30_1209 ();
 sg13g2_fill_1 FILLER_30_1211 ();
 sg13g2_fill_2 FILLER_30_1230 ();
 sg13g2_fill_1 FILLER_30_1232 ();
 sg13g2_fill_1 FILLER_30_1251 ();
 sg13g2_fill_1 FILLER_30_1278 ();
 sg13g2_fill_1 FILLER_30_1305 ();
 sg13g2_fill_1 FILLER_30_1320 ();
 sg13g2_decap_4 FILLER_30_1364 ();
 sg13g2_fill_2 FILLER_30_1368 ();
 sg13g2_decap_8 FILLER_30_1398 ();
 sg13g2_decap_4 FILLER_30_1405 ();
 sg13g2_decap_4 FILLER_30_1439 ();
 sg13g2_fill_1 FILLER_30_1443 ();
 sg13g2_fill_2 FILLER_30_1484 ();
 sg13g2_fill_1 FILLER_30_1486 ();
 sg13g2_fill_2 FILLER_30_1492 ();
 sg13g2_decap_4 FILLER_30_1499 ();
 sg13g2_fill_1 FILLER_30_1503 ();
 sg13g2_decap_8 FILLER_30_1518 ();
 sg13g2_fill_2 FILLER_30_1525 ();
 sg13g2_fill_1 FILLER_30_1588 ();
 sg13g2_fill_2 FILLER_30_1631 ();
 sg13g2_decap_8 FILLER_30_1672 ();
 sg13g2_fill_1 FILLER_30_1679 ();
 sg13g2_decap_4 FILLER_30_1711 ();
 sg13g2_fill_2 FILLER_30_1760 ();
 sg13g2_fill_2 FILLER_30_1771 ();
 sg13g2_fill_1 FILLER_30_1773 ();
 sg13g2_decap_4 FILLER_30_1814 ();
 sg13g2_fill_2 FILLER_30_1866 ();
 sg13g2_fill_2 FILLER_30_1872 ();
 sg13g2_decap_4 FILLER_30_1878 ();
 sg13g2_fill_2 FILLER_30_1913 ();
 sg13g2_fill_1 FILLER_30_1933 ();
 sg13g2_fill_2 FILLER_30_1964 ();
 sg13g2_fill_1 FILLER_30_1974 ();
 sg13g2_fill_2 FILLER_30_1997 ();
 sg13g2_fill_1 FILLER_30_1999 ();
 sg13g2_fill_2 FILLER_30_2008 ();
 sg13g2_fill_1 FILLER_30_2010 ();
 sg13g2_fill_2 FILLER_30_2026 ();
 sg13g2_fill_1 FILLER_30_2044 ();
 sg13g2_decap_8 FILLER_30_2080 ();
 sg13g2_fill_2 FILLER_30_2087 ();
 sg13g2_fill_1 FILLER_30_2089 ();
 sg13g2_fill_2 FILLER_30_2116 ();
 sg13g2_decap_4 FILLER_30_2158 ();
 sg13g2_fill_1 FILLER_30_2162 ();
 sg13g2_fill_1 FILLER_30_2198 ();
 sg13g2_fill_1 FILLER_30_2256 ();
 sg13g2_fill_1 FILLER_30_2262 ();
 sg13g2_fill_2 FILLER_30_2272 ();
 sg13g2_decap_4 FILLER_30_2290 ();
 sg13g2_fill_2 FILLER_30_2324 ();
 sg13g2_fill_1 FILLER_30_2326 ();
 sg13g2_decap_8 FILLER_30_2362 ();
 sg13g2_decap_8 FILLER_30_2369 ();
 sg13g2_decap_8 FILLER_30_2376 ();
 sg13g2_decap_8 FILLER_30_2383 ();
 sg13g2_decap_8 FILLER_30_2390 ();
 sg13g2_decap_8 FILLER_30_2397 ();
 sg13g2_decap_8 FILLER_30_2404 ();
 sg13g2_decap_8 FILLER_30_2411 ();
 sg13g2_decap_8 FILLER_30_2418 ();
 sg13g2_decap_8 FILLER_30_2425 ();
 sg13g2_decap_8 FILLER_30_2432 ();
 sg13g2_decap_8 FILLER_30_2439 ();
 sg13g2_decap_8 FILLER_30_2446 ();
 sg13g2_decap_8 FILLER_30_2453 ();
 sg13g2_decap_8 FILLER_30_2460 ();
 sg13g2_decap_8 FILLER_30_2467 ();
 sg13g2_decap_8 FILLER_30_2474 ();
 sg13g2_decap_8 FILLER_30_2481 ();
 sg13g2_decap_8 FILLER_30_2488 ();
 sg13g2_decap_8 FILLER_30_2495 ();
 sg13g2_decap_8 FILLER_30_2502 ();
 sg13g2_decap_8 FILLER_30_2509 ();
 sg13g2_decap_8 FILLER_30_2516 ();
 sg13g2_decap_8 FILLER_30_2523 ();
 sg13g2_decap_8 FILLER_30_2530 ();
 sg13g2_decap_8 FILLER_30_2537 ();
 sg13g2_decap_8 FILLER_30_2544 ();
 sg13g2_decap_8 FILLER_30_2551 ();
 sg13g2_decap_8 FILLER_30_2558 ();
 sg13g2_decap_8 FILLER_30_2565 ();
 sg13g2_decap_8 FILLER_30_2572 ();
 sg13g2_decap_8 FILLER_30_2579 ();
 sg13g2_decap_8 FILLER_30_2586 ();
 sg13g2_decap_8 FILLER_30_2593 ();
 sg13g2_decap_8 FILLER_30_2600 ();
 sg13g2_decap_8 FILLER_30_2607 ();
 sg13g2_decap_8 FILLER_30_2614 ();
 sg13g2_decap_8 FILLER_30_2621 ();
 sg13g2_decap_8 FILLER_30_2628 ();
 sg13g2_decap_8 FILLER_30_2635 ();
 sg13g2_decap_8 FILLER_30_2642 ();
 sg13g2_decap_8 FILLER_30_2649 ();
 sg13g2_decap_8 FILLER_30_2656 ();
 sg13g2_decap_8 FILLER_30_2663 ();
 sg13g2_decap_4 FILLER_30_2670 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_406 ();
 sg13g2_decap_8 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_fill_1 FILLER_31_427 ();
 sg13g2_fill_2 FILLER_31_454 ();
 sg13g2_fill_2 FILLER_31_470 ();
 sg13g2_fill_1 FILLER_31_472 ();
 sg13g2_fill_1 FILLER_31_478 ();
 sg13g2_fill_2 FILLER_31_497 ();
 sg13g2_fill_1 FILLER_31_499 ();
 sg13g2_fill_1 FILLER_31_514 ();
 sg13g2_fill_2 FILLER_31_524 ();
 sg13g2_fill_2 FILLER_31_540 ();
 sg13g2_fill_1 FILLER_31_651 ();
 sg13g2_fill_2 FILLER_31_657 ();
 sg13g2_fill_2 FILLER_31_674 ();
 sg13g2_fill_2 FILLER_31_684 ();
 sg13g2_fill_2 FILLER_31_700 ();
 sg13g2_fill_1 FILLER_31_757 ();
 sg13g2_fill_1 FILLER_31_775 ();
 sg13g2_fill_2 FILLER_31_780 ();
 sg13g2_fill_1 FILLER_31_782 ();
 sg13g2_fill_2 FILLER_31_793 ();
 sg13g2_fill_2 FILLER_31_826 ();
 sg13g2_fill_2 FILLER_31_854 ();
 sg13g2_fill_2 FILLER_31_868 ();
 sg13g2_fill_1 FILLER_31_870 ();
 sg13g2_fill_1 FILLER_31_937 ();
 sg13g2_fill_2 FILLER_31_973 ();
 sg13g2_fill_2 FILLER_31_1000 ();
 sg13g2_decap_8 FILLER_31_1006 ();
 sg13g2_decap_8 FILLER_31_1013 ();
 sg13g2_decap_8 FILLER_31_1020 ();
 sg13g2_decap_4 FILLER_31_1027 ();
 sg13g2_fill_1 FILLER_31_1031 ();
 sg13g2_fill_2 FILLER_31_1058 ();
 sg13g2_fill_1 FILLER_31_1060 ();
 sg13g2_fill_2 FILLER_31_1071 ();
 sg13g2_fill_1 FILLER_31_1073 ();
 sg13g2_fill_2 FILLER_31_1158 ();
 sg13g2_fill_1 FILLER_31_1164 ();
 sg13g2_decap_8 FILLER_31_1186 ();
 sg13g2_fill_2 FILLER_31_1193 ();
 sg13g2_fill_1 FILLER_31_1195 ();
 sg13g2_fill_1 FILLER_31_1252 ();
 sg13g2_fill_2 FILLER_31_1301 ();
 sg13g2_fill_2 FILLER_31_1352 ();
 sg13g2_fill_1 FILLER_31_1363 ();
 sg13g2_fill_2 FILLER_31_1377 ();
 sg13g2_fill_1 FILLER_31_1409 ();
 sg13g2_fill_1 FILLER_31_1415 ();
 sg13g2_decap_4 FILLER_31_1421 ();
 sg13g2_fill_2 FILLER_31_1425 ();
 sg13g2_fill_2 FILLER_31_1471 ();
 sg13g2_fill_2 FILLER_31_1542 ();
 sg13g2_fill_1 FILLER_31_1554 ();
 sg13g2_fill_2 FILLER_31_1568 ();
 sg13g2_fill_1 FILLER_31_1570 ();
 sg13g2_fill_2 FILLER_31_1593 ();
 sg13g2_fill_1 FILLER_31_1595 ();
 sg13g2_decap_4 FILLER_31_1636 ();
 sg13g2_fill_1 FILLER_31_1640 ();
 sg13g2_fill_1 FILLER_31_1650 ();
 sg13g2_decap_8 FILLER_31_1677 ();
 sg13g2_fill_2 FILLER_31_1696 ();
 sg13g2_fill_1 FILLER_31_1698 ();
 sg13g2_fill_1 FILLER_31_1704 ();
 sg13g2_fill_2 FILLER_31_1714 ();
 sg13g2_fill_2 FILLER_31_1738 ();
 sg13g2_fill_1 FILLER_31_1740 ();
 sg13g2_fill_1 FILLER_31_1758 ();
 sg13g2_fill_2 FILLER_31_1794 ();
 sg13g2_fill_1 FILLER_31_1796 ();
 sg13g2_fill_1 FILLER_31_1828 ();
 sg13g2_fill_2 FILLER_31_1859 ();
 sg13g2_fill_1 FILLER_31_1861 ();
 sg13g2_fill_2 FILLER_31_1872 ();
 sg13g2_fill_2 FILLER_31_1879 ();
 sg13g2_fill_1 FILLER_31_1881 ();
 sg13g2_fill_2 FILLER_31_1891 ();
 sg13g2_fill_2 FILLER_31_1901 ();
 sg13g2_fill_1 FILLER_31_1935 ();
 sg13g2_fill_1 FILLER_31_1953 ();
 sg13g2_fill_1 FILLER_31_2043 ();
 sg13g2_fill_2 FILLER_31_2049 ();
 sg13g2_fill_2 FILLER_31_2108 ();
 sg13g2_fill_1 FILLER_31_2110 ();
 sg13g2_decap_4 FILLER_31_2128 ();
 sg13g2_fill_1 FILLER_31_2148 ();
 sg13g2_fill_2 FILLER_31_2162 ();
 sg13g2_fill_1 FILLER_31_2164 ();
 sg13g2_fill_1 FILLER_31_2191 ();
 sg13g2_fill_1 FILLER_31_2196 ();
 sg13g2_decap_4 FILLER_31_2201 ();
 sg13g2_fill_1 FILLER_31_2214 ();
 sg13g2_fill_2 FILLER_31_2219 ();
 sg13g2_fill_2 FILLER_31_2248 ();
 sg13g2_fill_1 FILLER_31_2250 ();
 sg13g2_fill_2 FILLER_31_2274 ();
 sg13g2_decap_8 FILLER_31_2280 ();
 sg13g2_fill_2 FILLER_31_2297 ();
 sg13g2_fill_2 FILLER_31_2325 ();
 sg13g2_fill_2 FILLER_31_2349 ();
 sg13g2_fill_1 FILLER_31_2351 ();
 sg13g2_decap_8 FILLER_31_2369 ();
 sg13g2_decap_8 FILLER_31_2376 ();
 sg13g2_decap_8 FILLER_31_2383 ();
 sg13g2_decap_8 FILLER_31_2390 ();
 sg13g2_decap_8 FILLER_31_2397 ();
 sg13g2_decap_8 FILLER_31_2404 ();
 sg13g2_decap_8 FILLER_31_2411 ();
 sg13g2_decap_8 FILLER_31_2418 ();
 sg13g2_decap_8 FILLER_31_2425 ();
 sg13g2_decap_8 FILLER_31_2432 ();
 sg13g2_decap_8 FILLER_31_2439 ();
 sg13g2_decap_8 FILLER_31_2446 ();
 sg13g2_decap_8 FILLER_31_2453 ();
 sg13g2_decap_8 FILLER_31_2460 ();
 sg13g2_decap_8 FILLER_31_2467 ();
 sg13g2_decap_8 FILLER_31_2474 ();
 sg13g2_decap_8 FILLER_31_2481 ();
 sg13g2_decap_8 FILLER_31_2488 ();
 sg13g2_decap_8 FILLER_31_2495 ();
 sg13g2_decap_8 FILLER_31_2502 ();
 sg13g2_decap_8 FILLER_31_2509 ();
 sg13g2_decap_8 FILLER_31_2516 ();
 sg13g2_decap_8 FILLER_31_2523 ();
 sg13g2_decap_8 FILLER_31_2530 ();
 sg13g2_decap_8 FILLER_31_2537 ();
 sg13g2_decap_8 FILLER_31_2544 ();
 sg13g2_decap_8 FILLER_31_2551 ();
 sg13g2_decap_8 FILLER_31_2558 ();
 sg13g2_decap_8 FILLER_31_2565 ();
 sg13g2_decap_8 FILLER_31_2572 ();
 sg13g2_decap_8 FILLER_31_2579 ();
 sg13g2_decap_8 FILLER_31_2586 ();
 sg13g2_decap_8 FILLER_31_2593 ();
 sg13g2_decap_8 FILLER_31_2600 ();
 sg13g2_decap_8 FILLER_31_2607 ();
 sg13g2_decap_8 FILLER_31_2614 ();
 sg13g2_decap_8 FILLER_31_2621 ();
 sg13g2_decap_8 FILLER_31_2628 ();
 sg13g2_decap_8 FILLER_31_2635 ();
 sg13g2_decap_8 FILLER_31_2642 ();
 sg13g2_decap_8 FILLER_31_2649 ();
 sg13g2_decap_8 FILLER_31_2656 ();
 sg13g2_decap_8 FILLER_31_2663 ();
 sg13g2_decap_4 FILLER_31_2670 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_413 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_decap_8 FILLER_32_427 ();
 sg13g2_decap_4 FILLER_32_434 ();
 sg13g2_fill_1 FILLER_32_584 ();
 sg13g2_fill_2 FILLER_32_590 ();
 sg13g2_fill_1 FILLER_32_592 ();
 sg13g2_fill_2 FILLER_32_621 ();
 sg13g2_fill_1 FILLER_32_623 ();
 sg13g2_fill_1 FILLER_32_641 ();
 sg13g2_fill_1 FILLER_32_659 ();
 sg13g2_fill_1 FILLER_32_695 ();
 sg13g2_fill_2 FILLER_32_722 ();
 sg13g2_fill_1 FILLER_32_724 ();
 sg13g2_fill_1 FILLER_32_739 ();
 sg13g2_fill_1 FILLER_32_781 ();
 sg13g2_fill_2 FILLER_32_791 ();
 sg13g2_decap_4 FILLER_32_807 ();
 sg13g2_decap_8 FILLER_32_815 ();
 sg13g2_fill_1 FILLER_32_822 ();
 sg13g2_decap_4 FILLER_32_827 ();
 sg13g2_fill_1 FILLER_32_862 ();
 sg13g2_fill_1 FILLER_32_894 ();
 sg13g2_fill_1 FILLER_32_921 ();
 sg13g2_decap_8 FILLER_32_957 ();
 sg13g2_fill_2 FILLER_32_990 ();
 sg13g2_fill_1 FILLER_32_1002 ();
 sg13g2_fill_2 FILLER_32_1022 ();
 sg13g2_fill_1 FILLER_32_1024 ();
 sg13g2_decap_4 FILLER_32_1038 ();
 sg13g2_fill_2 FILLER_32_1064 ();
 sg13g2_fill_2 FILLER_32_1141 ();
 sg13g2_fill_1 FILLER_32_1143 ();
 sg13g2_fill_2 FILLER_32_1230 ();
 sg13g2_fill_2 FILLER_32_1242 ();
 sg13g2_fill_2 FILLER_32_1258 ();
 sg13g2_fill_1 FILLER_32_1260 ();
 sg13g2_decap_8 FILLER_32_1266 ();
 sg13g2_fill_1 FILLER_32_1273 ();
 sg13g2_fill_1 FILLER_32_1288 ();
 sg13g2_fill_1 FILLER_32_1307 ();
 sg13g2_fill_1 FILLER_32_1312 ();
 sg13g2_fill_1 FILLER_32_1318 ();
 sg13g2_fill_2 FILLER_32_1366 ();
 sg13g2_fill_1 FILLER_32_1368 ();
 sg13g2_fill_2 FILLER_32_1373 ();
 sg13g2_fill_2 FILLER_32_1383 ();
 sg13g2_fill_1 FILLER_32_1385 ();
 sg13g2_fill_2 FILLER_32_1435 ();
 sg13g2_fill_1 FILLER_32_1437 ();
 sg13g2_fill_2 FILLER_32_1442 ();
 sg13g2_fill_1 FILLER_32_1448 ();
 sg13g2_decap_4 FILLER_32_1480 ();
 sg13g2_decap_4 FILLER_32_1501 ();
 sg13g2_fill_1 FILLER_32_1505 ();
 sg13g2_fill_2 FILLER_32_1515 ();
 sg13g2_fill_1 FILLER_32_1517 ();
 sg13g2_decap_8 FILLER_32_1522 ();
 sg13g2_fill_2 FILLER_32_1618 ();
 sg13g2_fill_1 FILLER_32_1620 ();
 sg13g2_fill_2 FILLER_32_1692 ();
 sg13g2_fill_1 FILLER_32_1694 ();
 sg13g2_fill_2 FILLER_32_1721 ();
 sg13g2_fill_1 FILLER_32_1723 ();
 sg13g2_fill_2 FILLER_32_1777 ();
 sg13g2_fill_2 FILLER_32_1797 ();
 sg13g2_fill_2 FILLER_32_1812 ();
 sg13g2_fill_2 FILLER_32_1819 ();
 sg13g2_fill_2 FILLER_32_1835 ();
 sg13g2_fill_1 FILLER_32_1837 ();
 sg13g2_decap_8 FILLER_32_1899 ();
 sg13g2_decap_4 FILLER_32_1970 ();
 sg13g2_fill_1 FILLER_32_1974 ();
 sg13g2_fill_2 FILLER_32_1987 ();
 sg13g2_fill_1 FILLER_32_1989 ();
 sg13g2_decap_8 FILLER_32_2016 ();
 sg13g2_decap_4 FILLER_32_2023 ();
 sg13g2_fill_2 FILLER_32_2031 ();
 sg13g2_fill_1 FILLER_32_2055 ();
 sg13g2_fill_2 FILLER_32_2096 ();
 sg13g2_decap_4 FILLER_32_2132 ();
 sg13g2_fill_1 FILLER_32_2136 ();
 sg13g2_decap_4 FILLER_32_2142 ();
 sg13g2_fill_1 FILLER_32_2212 ();
 sg13g2_decap_4 FILLER_32_2226 ();
 sg13g2_decap_8 FILLER_32_2291 ();
 sg13g2_decap_8 FILLER_32_2298 ();
 sg13g2_decap_4 FILLER_32_2305 ();
 sg13g2_fill_1 FILLER_32_2309 ();
 sg13g2_fill_1 FILLER_32_2324 ();
 sg13g2_fill_1 FILLER_32_2363 ();
 sg13g2_decap_8 FILLER_32_2373 ();
 sg13g2_decap_8 FILLER_32_2380 ();
 sg13g2_decap_8 FILLER_32_2387 ();
 sg13g2_decap_8 FILLER_32_2394 ();
 sg13g2_decap_8 FILLER_32_2401 ();
 sg13g2_decap_8 FILLER_32_2408 ();
 sg13g2_decap_8 FILLER_32_2415 ();
 sg13g2_decap_8 FILLER_32_2422 ();
 sg13g2_decap_8 FILLER_32_2429 ();
 sg13g2_decap_8 FILLER_32_2436 ();
 sg13g2_decap_8 FILLER_32_2443 ();
 sg13g2_decap_8 FILLER_32_2450 ();
 sg13g2_decap_8 FILLER_32_2457 ();
 sg13g2_decap_8 FILLER_32_2464 ();
 sg13g2_decap_8 FILLER_32_2471 ();
 sg13g2_decap_8 FILLER_32_2478 ();
 sg13g2_decap_8 FILLER_32_2485 ();
 sg13g2_decap_8 FILLER_32_2492 ();
 sg13g2_decap_8 FILLER_32_2499 ();
 sg13g2_decap_8 FILLER_32_2506 ();
 sg13g2_decap_8 FILLER_32_2513 ();
 sg13g2_decap_8 FILLER_32_2520 ();
 sg13g2_decap_8 FILLER_32_2527 ();
 sg13g2_decap_8 FILLER_32_2534 ();
 sg13g2_decap_8 FILLER_32_2541 ();
 sg13g2_decap_8 FILLER_32_2548 ();
 sg13g2_decap_8 FILLER_32_2555 ();
 sg13g2_decap_8 FILLER_32_2562 ();
 sg13g2_decap_8 FILLER_32_2569 ();
 sg13g2_decap_8 FILLER_32_2576 ();
 sg13g2_decap_8 FILLER_32_2583 ();
 sg13g2_decap_8 FILLER_32_2590 ();
 sg13g2_decap_8 FILLER_32_2597 ();
 sg13g2_decap_8 FILLER_32_2604 ();
 sg13g2_decap_8 FILLER_32_2611 ();
 sg13g2_decap_8 FILLER_32_2618 ();
 sg13g2_decap_8 FILLER_32_2625 ();
 sg13g2_decap_8 FILLER_32_2632 ();
 sg13g2_decap_8 FILLER_32_2639 ();
 sg13g2_decap_8 FILLER_32_2646 ();
 sg13g2_decap_8 FILLER_32_2653 ();
 sg13g2_decap_8 FILLER_32_2660 ();
 sg13g2_decap_8 FILLER_32_2667 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_decap_8 FILLER_33_406 ();
 sg13g2_decap_8 FILLER_33_413 ();
 sg13g2_decap_8 FILLER_33_420 ();
 sg13g2_decap_8 FILLER_33_427 ();
 sg13g2_decap_8 FILLER_33_434 ();
 sg13g2_decap_8 FILLER_33_441 ();
 sg13g2_fill_1 FILLER_33_448 ();
 sg13g2_decap_8 FILLER_33_475 ();
 sg13g2_decap_8 FILLER_33_482 ();
 sg13g2_fill_2 FILLER_33_489 ();
 sg13g2_fill_2 FILLER_33_495 ();
 sg13g2_fill_1 FILLER_33_497 ();
 sg13g2_fill_2 FILLER_33_503 ();
 sg13g2_fill_1 FILLER_33_505 ();
 sg13g2_decap_8 FILLER_33_519 ();
 sg13g2_fill_1 FILLER_33_526 ();
 sg13g2_fill_2 FILLER_33_540 ();
 sg13g2_fill_1 FILLER_33_568 ();
 sg13g2_fill_1 FILLER_33_595 ();
 sg13g2_fill_2 FILLER_33_626 ();
 sg13g2_fill_1 FILLER_33_628 ();
 sg13g2_fill_2 FILLER_33_664 ();
 sg13g2_fill_1 FILLER_33_666 ();
 sg13g2_fill_2 FILLER_33_672 ();
 sg13g2_fill_1 FILLER_33_674 ();
 sg13g2_fill_2 FILLER_33_688 ();
 sg13g2_fill_1 FILLER_33_690 ();
 sg13g2_fill_1 FILLER_33_708 ();
 sg13g2_fill_1 FILLER_33_717 ();
 sg13g2_fill_2 FILLER_33_732 ();
 sg13g2_fill_1 FILLER_33_734 ();
 sg13g2_fill_1 FILLER_33_749 ();
 sg13g2_fill_2 FILLER_33_758 ();
 sg13g2_fill_1 FILLER_33_760 ();
 sg13g2_fill_2 FILLER_33_778 ();
 sg13g2_fill_1 FILLER_33_780 ();
 sg13g2_decap_4 FILLER_33_807 ();
 sg13g2_fill_1 FILLER_33_887 ();
 sg13g2_decap_4 FILLER_33_892 ();
 sg13g2_fill_1 FILLER_33_896 ();
 sg13g2_fill_2 FILLER_33_901 ();
 sg13g2_fill_2 FILLER_33_915 ();
 sg13g2_fill_1 FILLER_33_926 ();
 sg13g2_fill_2 FILLER_33_941 ();
 sg13g2_fill_1 FILLER_33_960 ();
 sg13g2_fill_2 FILLER_33_974 ();
 sg13g2_fill_1 FILLER_33_976 ();
 sg13g2_fill_2 FILLER_33_987 ();
 sg13g2_fill_2 FILLER_33_1023 ();
 sg13g2_decap_4 FILLER_33_1033 ();
 sg13g2_decap_4 FILLER_33_1067 ();
 sg13g2_fill_2 FILLER_33_1080 ();
 sg13g2_fill_2 FILLER_33_1091 ();
 sg13g2_fill_2 FILLER_33_1102 ();
 sg13g2_fill_1 FILLER_33_1104 ();
 sg13g2_fill_2 FILLER_33_1113 ();
 sg13g2_fill_1 FILLER_33_1115 ();
 sg13g2_decap_8 FILLER_33_1142 ();
 sg13g2_decap_4 FILLER_33_1149 ();
 sg13g2_fill_2 FILLER_33_1153 ();
 sg13g2_fill_2 FILLER_33_1164 ();
 sg13g2_fill_2 FILLER_33_1197 ();
 sg13g2_fill_2 FILLER_33_1290 ();
 sg13g2_decap_8 FILLER_33_1336 ();
 sg13g2_fill_2 FILLER_33_1343 ();
 sg13g2_fill_1 FILLER_33_1345 ();
 sg13g2_decap_4 FILLER_33_1350 ();
 sg13g2_fill_2 FILLER_33_1354 ();
 sg13g2_decap_4 FILLER_33_1413 ();
 sg13g2_fill_2 FILLER_33_1417 ();
 sg13g2_fill_2 FILLER_33_1424 ();
 sg13g2_fill_1 FILLER_33_1426 ();
 sg13g2_fill_2 FILLER_33_1458 ();
 sg13g2_fill_2 FILLER_33_1477 ();
 sg13g2_fill_1 FILLER_33_1479 ();
 sg13g2_decap_8 FILLER_33_1489 ();
 sg13g2_fill_2 FILLER_33_1496 ();
 sg13g2_fill_1 FILLER_33_1538 ();
 sg13g2_fill_2 FILLER_33_1543 ();
 sg13g2_fill_1 FILLER_33_1589 ();
 sg13g2_fill_2 FILLER_33_1629 ();
 sg13g2_decap_4 FILLER_33_1649 ();
 sg13g2_fill_1 FILLER_33_1663 ();
 sg13g2_decap_8 FILLER_33_1690 ();
 sg13g2_decap_4 FILLER_33_1697 ();
 sg13g2_fill_2 FILLER_33_1706 ();
 sg13g2_fill_1 FILLER_33_1739 ();
 sg13g2_fill_2 FILLER_33_1750 ();
 sg13g2_fill_1 FILLER_33_1752 ();
 sg13g2_fill_1 FILLER_33_1789 ();
 sg13g2_fill_1 FILLER_33_1816 ();
 sg13g2_fill_1 FILLER_33_1825 ();
 sg13g2_fill_2 FILLER_33_1830 ();
 sg13g2_fill_2 FILLER_33_1837 ();
 sg13g2_fill_1 FILLER_33_1839 ();
 sg13g2_fill_2 FILLER_33_1850 ();
 sg13g2_decap_8 FILLER_33_1909 ();
 sg13g2_decap_8 FILLER_33_1916 ();
 sg13g2_fill_1 FILLER_33_1923 ();
 sg13g2_decap_8 FILLER_33_1934 ();
 sg13g2_fill_2 FILLER_33_1956 ();
 sg13g2_fill_1 FILLER_33_1958 ();
 sg13g2_decap_8 FILLER_33_1974 ();
 sg13g2_fill_1 FILLER_33_1985 ();
 sg13g2_fill_1 FILLER_33_1995 ();
 sg13g2_decap_8 FILLER_33_2009 ();
 sg13g2_fill_2 FILLER_33_2016 ();
 sg13g2_fill_1 FILLER_33_2018 ();
 sg13g2_fill_1 FILLER_33_2098 ();
 sg13g2_fill_1 FILLER_33_2108 ();
 sg13g2_decap_4 FILLER_33_2113 ();
 sg13g2_decap_4 FILLER_33_2121 ();
 sg13g2_fill_2 FILLER_33_2125 ();
 sg13g2_fill_2 FILLER_33_2148 ();
 sg13g2_fill_2 FILLER_33_2164 ();
 sg13g2_fill_2 FILLER_33_2205 ();
 sg13g2_fill_2 FILLER_33_2212 ();
 sg13g2_fill_1 FILLER_33_2214 ();
 sg13g2_fill_2 FILLER_33_2326 ();
 sg13g2_decap_8 FILLER_33_2375 ();
 sg13g2_decap_8 FILLER_33_2382 ();
 sg13g2_decap_8 FILLER_33_2389 ();
 sg13g2_decap_8 FILLER_33_2396 ();
 sg13g2_decap_8 FILLER_33_2403 ();
 sg13g2_decap_8 FILLER_33_2410 ();
 sg13g2_decap_8 FILLER_33_2417 ();
 sg13g2_decap_8 FILLER_33_2424 ();
 sg13g2_decap_8 FILLER_33_2431 ();
 sg13g2_decap_8 FILLER_33_2438 ();
 sg13g2_decap_8 FILLER_33_2445 ();
 sg13g2_decap_8 FILLER_33_2452 ();
 sg13g2_decap_8 FILLER_33_2459 ();
 sg13g2_decap_8 FILLER_33_2466 ();
 sg13g2_decap_8 FILLER_33_2473 ();
 sg13g2_decap_8 FILLER_33_2480 ();
 sg13g2_decap_8 FILLER_33_2487 ();
 sg13g2_decap_8 FILLER_33_2494 ();
 sg13g2_decap_8 FILLER_33_2501 ();
 sg13g2_decap_8 FILLER_33_2508 ();
 sg13g2_decap_8 FILLER_33_2515 ();
 sg13g2_decap_8 FILLER_33_2522 ();
 sg13g2_decap_8 FILLER_33_2529 ();
 sg13g2_decap_8 FILLER_33_2536 ();
 sg13g2_decap_8 FILLER_33_2543 ();
 sg13g2_decap_8 FILLER_33_2550 ();
 sg13g2_decap_8 FILLER_33_2557 ();
 sg13g2_decap_8 FILLER_33_2564 ();
 sg13g2_decap_8 FILLER_33_2571 ();
 sg13g2_decap_8 FILLER_33_2578 ();
 sg13g2_decap_8 FILLER_33_2585 ();
 sg13g2_decap_8 FILLER_33_2592 ();
 sg13g2_decap_8 FILLER_33_2599 ();
 sg13g2_decap_8 FILLER_33_2606 ();
 sg13g2_decap_8 FILLER_33_2613 ();
 sg13g2_decap_8 FILLER_33_2620 ();
 sg13g2_decap_8 FILLER_33_2627 ();
 sg13g2_decap_8 FILLER_33_2634 ();
 sg13g2_decap_8 FILLER_33_2641 ();
 sg13g2_decap_8 FILLER_33_2648 ();
 sg13g2_decap_8 FILLER_33_2655 ();
 sg13g2_decap_8 FILLER_33_2662 ();
 sg13g2_decap_4 FILLER_33_2669 ();
 sg13g2_fill_1 FILLER_33_2673 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_34_406 ();
 sg13g2_decap_8 FILLER_34_413 ();
 sg13g2_decap_8 FILLER_34_420 ();
 sg13g2_decap_8 FILLER_34_427 ();
 sg13g2_decap_8 FILLER_34_434 ();
 sg13g2_decap_8 FILLER_34_441 ();
 sg13g2_decap_8 FILLER_34_448 ();
 sg13g2_decap_8 FILLER_34_455 ();
 sg13g2_fill_1 FILLER_34_462 ();
 sg13g2_decap_4 FILLER_34_468 ();
 sg13g2_fill_2 FILLER_34_551 ();
 sg13g2_fill_1 FILLER_34_562 ();
 sg13g2_fill_1 FILLER_34_576 ();
 sg13g2_fill_1 FILLER_34_586 ();
 sg13g2_decap_4 FILLER_34_591 ();
 sg13g2_fill_2 FILLER_34_595 ();
 sg13g2_fill_2 FILLER_34_629 ();
 sg13g2_fill_2 FILLER_34_650 ();
 sg13g2_fill_2 FILLER_34_754 ();
 sg13g2_fill_1 FILLER_34_756 ();
 sg13g2_fill_1 FILLER_34_766 ();
 sg13g2_fill_1 FILLER_34_808 ();
 sg13g2_fill_2 FILLER_34_884 ();
 sg13g2_decap_4 FILLER_34_952 ();
 sg13g2_fill_2 FILLER_34_991 ();
 sg13g2_fill_2 FILLER_34_1012 ();
 sg13g2_fill_1 FILLER_34_1014 ();
 sg13g2_fill_1 FILLER_34_1049 ();
 sg13g2_decap_4 FILLER_34_1114 ();
 sg13g2_fill_2 FILLER_34_1118 ();
 sg13g2_fill_1 FILLER_34_1129 ();
 sg13g2_decap_4 FILLER_34_1143 ();
 sg13g2_decap_4 FILLER_34_1182 ();
 sg13g2_fill_1 FILLER_34_1244 ();
 sg13g2_decap_8 FILLER_34_1261 ();
 sg13g2_decap_8 FILLER_34_1268 ();
 sg13g2_fill_2 FILLER_34_1301 ();
 sg13g2_fill_1 FILLER_34_1303 ();
 sg13g2_fill_2 FILLER_34_1382 ();
 sg13g2_fill_1 FILLER_34_1384 ();
 sg13g2_fill_2 FILLER_34_1446 ();
 sg13g2_fill_1 FILLER_34_1448 ();
 sg13g2_fill_1 FILLER_34_1541 ();
 sg13g2_decap_4 FILLER_34_1555 ();
 sg13g2_fill_2 FILLER_34_1559 ();
 sg13g2_fill_1 FILLER_34_1592 ();
 sg13g2_decap_4 FILLER_34_1610 ();
 sg13g2_fill_2 FILLER_34_1678 ();
 sg13g2_decap_4 FILLER_34_1700 ();
 sg13g2_fill_2 FILLER_34_1704 ();
 sg13g2_fill_1 FILLER_34_1710 ();
 sg13g2_fill_2 FILLER_34_1723 ();
 sg13g2_decap_8 FILLER_34_1755 ();
 sg13g2_fill_2 FILLER_34_1762 ();
 sg13g2_fill_2 FILLER_34_1779 ();
 sg13g2_fill_2 FILLER_34_1830 ();
 sg13g2_fill_2 FILLER_34_1842 ();
 sg13g2_fill_1 FILLER_34_1844 ();
 sg13g2_fill_2 FILLER_34_1871 ();
 sg13g2_fill_1 FILLER_34_1873 ();
 sg13g2_fill_2 FILLER_34_1883 ();
 sg13g2_fill_1 FILLER_34_1885 ();
 sg13g2_fill_2 FILLER_34_1942 ();
 sg13g2_fill_1 FILLER_34_1944 ();
 sg13g2_fill_2 FILLER_34_2038 ();
 sg13g2_fill_1 FILLER_34_2040 ();
 sg13g2_fill_2 FILLER_34_2144 ();
 sg13g2_fill_1 FILLER_34_2146 ();
 sg13g2_decap_4 FILLER_34_2177 ();
 sg13g2_decap_4 FILLER_34_2220 ();
 sg13g2_fill_1 FILLER_34_2224 ();
 sg13g2_fill_1 FILLER_34_2243 ();
 sg13g2_fill_2 FILLER_34_2248 ();
 sg13g2_fill_2 FILLER_34_2259 ();
 sg13g2_decap_4 FILLER_34_2265 ();
 sg13g2_fill_2 FILLER_34_2292 ();
 sg13g2_fill_2 FILLER_34_2307 ();
 sg13g2_fill_2 FILLER_34_2339 ();
 sg13g2_fill_1 FILLER_34_2341 ();
 sg13g2_decap_8 FILLER_34_2373 ();
 sg13g2_decap_8 FILLER_34_2380 ();
 sg13g2_decap_8 FILLER_34_2387 ();
 sg13g2_decap_8 FILLER_34_2394 ();
 sg13g2_decap_8 FILLER_34_2401 ();
 sg13g2_decap_8 FILLER_34_2408 ();
 sg13g2_decap_8 FILLER_34_2415 ();
 sg13g2_decap_8 FILLER_34_2422 ();
 sg13g2_decap_8 FILLER_34_2429 ();
 sg13g2_decap_8 FILLER_34_2436 ();
 sg13g2_decap_8 FILLER_34_2443 ();
 sg13g2_decap_8 FILLER_34_2450 ();
 sg13g2_decap_8 FILLER_34_2457 ();
 sg13g2_decap_8 FILLER_34_2464 ();
 sg13g2_decap_8 FILLER_34_2471 ();
 sg13g2_decap_8 FILLER_34_2478 ();
 sg13g2_decap_8 FILLER_34_2485 ();
 sg13g2_decap_8 FILLER_34_2492 ();
 sg13g2_decap_8 FILLER_34_2499 ();
 sg13g2_decap_8 FILLER_34_2506 ();
 sg13g2_decap_8 FILLER_34_2513 ();
 sg13g2_decap_8 FILLER_34_2520 ();
 sg13g2_decap_8 FILLER_34_2527 ();
 sg13g2_decap_8 FILLER_34_2534 ();
 sg13g2_decap_8 FILLER_34_2541 ();
 sg13g2_decap_8 FILLER_34_2548 ();
 sg13g2_decap_8 FILLER_34_2555 ();
 sg13g2_decap_8 FILLER_34_2562 ();
 sg13g2_decap_8 FILLER_34_2569 ();
 sg13g2_decap_8 FILLER_34_2576 ();
 sg13g2_decap_8 FILLER_34_2583 ();
 sg13g2_decap_8 FILLER_34_2590 ();
 sg13g2_decap_8 FILLER_34_2597 ();
 sg13g2_decap_8 FILLER_34_2604 ();
 sg13g2_decap_8 FILLER_34_2611 ();
 sg13g2_decap_8 FILLER_34_2618 ();
 sg13g2_decap_8 FILLER_34_2625 ();
 sg13g2_decap_8 FILLER_34_2632 ();
 sg13g2_decap_8 FILLER_34_2639 ();
 sg13g2_decap_8 FILLER_34_2646 ();
 sg13g2_decap_8 FILLER_34_2653 ();
 sg13g2_decap_8 FILLER_34_2660 ();
 sg13g2_decap_8 FILLER_34_2667 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_decap_8 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_413 ();
 sg13g2_decap_8 FILLER_35_420 ();
 sg13g2_decap_8 FILLER_35_427 ();
 sg13g2_decap_8 FILLER_35_434 ();
 sg13g2_decap_8 FILLER_35_441 ();
 sg13g2_decap_8 FILLER_35_448 ();
 sg13g2_decap_4 FILLER_35_455 ();
 sg13g2_fill_2 FILLER_35_459 ();
 sg13g2_fill_1 FILLER_35_474 ();
 sg13g2_fill_2 FILLER_35_514 ();
 sg13g2_fill_1 FILLER_35_516 ();
 sg13g2_fill_1 FILLER_35_538 ();
 sg13g2_fill_2 FILLER_35_573 ();
 sg13g2_fill_1 FILLER_35_575 ();
 sg13g2_fill_2 FILLER_35_611 ();
 sg13g2_fill_2 FILLER_35_648 ();
 sg13g2_decap_4 FILLER_35_682 ();
 sg13g2_fill_2 FILLER_35_736 ();
 sg13g2_fill_1 FILLER_35_738 ();
 sg13g2_fill_1 FILLER_35_765 ();
 sg13g2_fill_2 FILLER_35_823 ();
 sg13g2_fill_1 FILLER_35_825 ();
 sg13g2_fill_2 FILLER_35_864 ();
 sg13g2_fill_1 FILLER_35_866 ();
 sg13g2_fill_2 FILLER_35_881 ();
 sg13g2_decap_4 FILLER_35_919 ();
 sg13g2_fill_1 FILLER_35_923 ();
 sg13g2_fill_1 FILLER_35_932 ();
 sg13g2_decap_8 FILLER_35_937 ();
 sg13g2_fill_1 FILLER_35_944 ();
 sg13g2_fill_2 FILLER_35_950 ();
 sg13g2_fill_1 FILLER_35_957 ();
 sg13g2_decap_4 FILLER_35_963 ();
 sg13g2_decap_4 FILLER_35_1027 ();
 sg13g2_fill_1 FILLER_35_1031 ();
 sg13g2_fill_1 FILLER_35_1041 ();
 sg13g2_fill_2 FILLER_35_1077 ();
 sg13g2_decap_4 FILLER_35_1110 ();
 sg13g2_decap_8 FILLER_35_1122 ();
 sg13g2_fill_2 FILLER_35_1155 ();
 sg13g2_fill_1 FILLER_35_1157 ();
 sg13g2_decap_8 FILLER_35_1162 ();
 sg13g2_decap_4 FILLER_35_1169 ();
 sg13g2_fill_1 FILLER_35_1204 ();
 sg13g2_decap_8 FILLER_35_1221 ();
 sg13g2_fill_2 FILLER_35_1228 ();
 sg13g2_fill_1 FILLER_35_1256 ();
 sg13g2_fill_1 FILLER_35_1306 ();
 sg13g2_fill_2 FILLER_35_1316 ();
 sg13g2_fill_1 FILLER_35_1318 ();
 sg13g2_fill_1 FILLER_35_1364 ();
 sg13g2_fill_2 FILLER_35_1390 ();
 sg13g2_decap_4 FILLER_35_1401 ();
 sg13g2_fill_1 FILLER_35_1405 ();
 sg13g2_decap_4 FILLER_35_1410 ();
 sg13g2_fill_2 FILLER_35_1414 ();
 sg13g2_fill_2 FILLER_35_1438 ();
 sg13g2_fill_1 FILLER_35_1440 ();
 sg13g2_decap_8 FILLER_35_1481 ();
 sg13g2_decap_4 FILLER_35_1488 ();
 sg13g2_fill_1 FILLER_35_1492 ();
 sg13g2_fill_1 FILLER_35_1511 ();
 sg13g2_decap_4 FILLER_35_1533 ();
 sg13g2_fill_1 FILLER_35_1537 ();
 sg13g2_fill_2 FILLER_35_1552 ();
 sg13g2_fill_1 FILLER_35_1554 ();
 sg13g2_fill_1 FILLER_35_1573 ();
 sg13g2_fill_2 FILLER_35_1580 ();
 sg13g2_fill_1 FILLER_35_1582 ();
 sg13g2_fill_2 FILLER_35_1586 ();
 sg13g2_fill_2 FILLER_35_1597 ();
 sg13g2_fill_1 FILLER_35_1599 ();
 sg13g2_decap_4 FILLER_35_1610 ();
 sg13g2_fill_2 FILLER_35_1614 ();
 sg13g2_fill_2 FILLER_35_1647 ();
 sg13g2_fill_1 FILLER_35_1649 ();
 sg13g2_fill_2 FILLER_35_1654 ();
 sg13g2_fill_1 FILLER_35_1656 ();
 sg13g2_fill_1 FILLER_35_1672 ();
 sg13g2_fill_1 FILLER_35_1718 ();
 sg13g2_decap_4 FILLER_35_1732 ();
 sg13g2_fill_1 FILLER_35_1736 ();
 sg13g2_decap_8 FILLER_35_1742 ();
 sg13g2_decap_8 FILLER_35_1749 ();
 sg13g2_fill_1 FILLER_35_1756 ();
 sg13g2_decap_8 FILLER_35_1762 ();
 sg13g2_decap_8 FILLER_35_1769 ();
 sg13g2_decap_4 FILLER_35_1784 ();
 sg13g2_fill_2 FILLER_35_1788 ();
 sg13g2_fill_1 FILLER_35_1808 ();
 sg13g2_fill_1 FILLER_35_1814 ();
 sg13g2_fill_1 FILLER_35_1824 ();
 sg13g2_decap_8 FILLER_35_1838 ();
 sg13g2_fill_2 FILLER_35_1845 ();
 sg13g2_fill_1 FILLER_35_1847 ();
 sg13g2_fill_2 FILLER_35_1869 ();
 sg13g2_fill_1 FILLER_35_1871 ();
 sg13g2_decap_4 FILLER_35_1920 ();
 sg13g2_decap_4 FILLER_35_1946 ();
 sg13g2_fill_1 FILLER_35_1966 ();
 sg13g2_decap_8 FILLER_35_1976 ();
 sg13g2_fill_1 FILLER_35_1983 ();
 sg13g2_fill_2 FILLER_35_1992 ();
 sg13g2_fill_1 FILLER_35_1994 ();
 sg13g2_fill_2 FILLER_35_2004 ();
 sg13g2_fill_2 FILLER_35_2064 ();
 sg13g2_fill_1 FILLER_35_2066 ();
 sg13g2_fill_2 FILLER_35_2089 ();
 sg13g2_fill_2 FILLER_35_2096 ();
 sg13g2_decap_4 FILLER_35_2124 ();
 sg13g2_fill_1 FILLER_35_2128 ();
 sg13g2_decap_8 FILLER_35_2141 ();
 sg13g2_fill_1 FILLER_35_2148 ();
 sg13g2_fill_2 FILLER_35_2166 ();
 sg13g2_fill_1 FILLER_35_2168 ();
 sg13g2_decap_8 FILLER_35_2221 ();
 sg13g2_fill_2 FILLER_35_2228 ();
 sg13g2_fill_1 FILLER_35_2266 ();
 sg13g2_fill_1 FILLER_35_2307 ();
 sg13g2_decap_4 FILLER_35_2349 ();
 sg13g2_decap_8 FILLER_35_2375 ();
 sg13g2_decap_8 FILLER_35_2382 ();
 sg13g2_decap_8 FILLER_35_2389 ();
 sg13g2_decap_8 FILLER_35_2396 ();
 sg13g2_decap_8 FILLER_35_2403 ();
 sg13g2_decap_8 FILLER_35_2410 ();
 sg13g2_decap_8 FILLER_35_2417 ();
 sg13g2_decap_8 FILLER_35_2424 ();
 sg13g2_decap_8 FILLER_35_2431 ();
 sg13g2_decap_8 FILLER_35_2438 ();
 sg13g2_decap_8 FILLER_35_2445 ();
 sg13g2_decap_8 FILLER_35_2452 ();
 sg13g2_decap_8 FILLER_35_2459 ();
 sg13g2_decap_8 FILLER_35_2466 ();
 sg13g2_decap_8 FILLER_35_2473 ();
 sg13g2_decap_8 FILLER_35_2480 ();
 sg13g2_decap_8 FILLER_35_2487 ();
 sg13g2_decap_8 FILLER_35_2494 ();
 sg13g2_decap_8 FILLER_35_2501 ();
 sg13g2_decap_8 FILLER_35_2508 ();
 sg13g2_decap_8 FILLER_35_2515 ();
 sg13g2_decap_8 FILLER_35_2522 ();
 sg13g2_decap_8 FILLER_35_2529 ();
 sg13g2_decap_8 FILLER_35_2536 ();
 sg13g2_decap_8 FILLER_35_2543 ();
 sg13g2_decap_8 FILLER_35_2550 ();
 sg13g2_decap_8 FILLER_35_2557 ();
 sg13g2_decap_8 FILLER_35_2564 ();
 sg13g2_decap_8 FILLER_35_2571 ();
 sg13g2_decap_8 FILLER_35_2578 ();
 sg13g2_decap_8 FILLER_35_2585 ();
 sg13g2_decap_8 FILLER_35_2592 ();
 sg13g2_decap_8 FILLER_35_2599 ();
 sg13g2_decap_8 FILLER_35_2606 ();
 sg13g2_decap_8 FILLER_35_2613 ();
 sg13g2_decap_8 FILLER_35_2620 ();
 sg13g2_decap_8 FILLER_35_2627 ();
 sg13g2_decap_8 FILLER_35_2634 ();
 sg13g2_decap_8 FILLER_35_2641 ();
 sg13g2_decap_8 FILLER_35_2648 ();
 sg13g2_decap_8 FILLER_35_2655 ();
 sg13g2_decap_8 FILLER_35_2662 ();
 sg13g2_decap_4 FILLER_35_2669 ();
 sg13g2_fill_1 FILLER_35_2673 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_36_406 ();
 sg13g2_decap_8 FILLER_36_413 ();
 sg13g2_decap_8 FILLER_36_420 ();
 sg13g2_decap_8 FILLER_36_427 ();
 sg13g2_decap_8 FILLER_36_434 ();
 sg13g2_decap_8 FILLER_36_441 ();
 sg13g2_decap_4 FILLER_36_448 ();
 sg13g2_fill_2 FILLER_36_452 ();
 sg13g2_fill_2 FILLER_36_519 ();
 sg13g2_fill_1 FILLER_36_521 ();
 sg13g2_fill_2 FILLER_36_557 ();
 sg13g2_decap_4 FILLER_36_589 ();
 sg13g2_fill_1 FILLER_36_593 ();
 sg13g2_fill_2 FILLER_36_608 ();
 sg13g2_fill_2 FILLER_36_614 ();
 sg13g2_fill_2 FILLER_36_629 ();
 sg13g2_fill_1 FILLER_36_631 ();
 sg13g2_fill_2 FILLER_36_649 ();
 sg13g2_fill_2 FILLER_36_668 ();
 sg13g2_fill_1 FILLER_36_670 ();
 sg13g2_fill_1 FILLER_36_680 ();
 sg13g2_decap_4 FILLER_36_691 ();
 sg13g2_fill_1 FILLER_36_695 ();
 sg13g2_fill_2 FILLER_36_700 ();
 sg13g2_fill_2 FILLER_36_728 ();
 sg13g2_fill_1 FILLER_36_730 ();
 sg13g2_fill_2 FILLER_36_746 ();
 sg13g2_fill_1 FILLER_36_748 ();
 sg13g2_fill_1 FILLER_36_785 ();
 sg13g2_fill_2 FILLER_36_838 ();
 sg13g2_fill_2 FILLER_36_849 ();
 sg13g2_fill_1 FILLER_36_851 ();
 sg13g2_fill_2 FILLER_36_878 ();
 sg13g2_fill_1 FILLER_36_880 ();
 sg13g2_decap_4 FILLER_36_921 ();
 sg13g2_fill_1 FILLER_36_925 ();
 sg13g2_decap_4 FILLER_36_956 ();
 sg13g2_decap_4 FILLER_36_968 ();
 sg13g2_fill_2 FILLER_36_972 ();
 sg13g2_fill_2 FILLER_36_979 ();
 sg13g2_fill_1 FILLER_36_981 ();
 sg13g2_fill_1 FILLER_36_986 ();
 sg13g2_decap_4 FILLER_36_991 ();
 sg13g2_fill_1 FILLER_36_995 ();
 sg13g2_fill_2 FILLER_36_1010 ();
 sg13g2_fill_2 FILLER_36_1030 ();
 sg13g2_fill_1 FILLER_36_1032 ();
 sg13g2_fill_2 FILLER_36_1064 ();
 sg13g2_fill_1 FILLER_36_1066 ();
 sg13g2_fill_2 FILLER_36_1098 ();
 sg13g2_fill_1 FILLER_36_1126 ();
 sg13g2_fill_1 FILLER_36_1134 ();
 sg13g2_decap_4 FILLER_36_1157 ();
 sg13g2_fill_2 FILLER_36_1161 ();
 sg13g2_fill_2 FILLER_36_1172 ();
 sg13g2_fill_1 FILLER_36_1200 ();
 sg13g2_fill_1 FILLER_36_1215 ();
 sg13g2_decap_8 FILLER_36_1220 ();
 sg13g2_decap_4 FILLER_36_1227 ();
 sg13g2_fill_2 FILLER_36_1231 ();
 sg13g2_fill_1 FILLER_36_1240 ();
 sg13g2_decap_4 FILLER_36_1245 ();
 sg13g2_fill_1 FILLER_36_1249 ();
 sg13g2_decap_8 FILLER_36_1266 ();
 sg13g2_decap_4 FILLER_36_1273 ();
 sg13g2_fill_2 FILLER_36_1277 ();
 sg13g2_fill_2 FILLER_36_1374 ();
 sg13g2_fill_1 FILLER_36_1376 ();
 sg13g2_fill_2 FILLER_36_1455 ();
 sg13g2_fill_1 FILLER_36_1457 ();
 sg13g2_decap_8 FILLER_36_1510 ();
 sg13g2_fill_2 FILLER_36_1517 ();
 sg13g2_decap_8 FILLER_36_1529 ();
 sg13g2_decap_4 FILLER_36_1536 ();
 sg13g2_fill_2 FILLER_36_1550 ();
 sg13g2_fill_1 FILLER_36_1552 ();
 sg13g2_fill_2 FILLER_36_1566 ();
 sg13g2_fill_1 FILLER_36_1568 ();
 sg13g2_fill_2 FILLER_36_1574 ();
 sg13g2_fill_1 FILLER_36_1599 ();
 sg13g2_decap_4 FILLER_36_1626 ();
 sg13g2_fill_1 FILLER_36_1630 ();
 sg13g2_decap_4 FILLER_36_1638 ();
 sg13g2_decap_4 FILLER_36_1682 ();
 sg13g2_decap_8 FILLER_36_1694 ();
 sg13g2_decap_8 FILLER_36_1741 ();
 sg13g2_fill_2 FILLER_36_1748 ();
 sg13g2_decap_4 FILLER_36_1771 ();
 sg13g2_fill_2 FILLER_36_1775 ();
 sg13g2_decap_4 FILLER_36_1895 ();
 sg13g2_fill_1 FILLER_36_1904 ();
 sg13g2_fill_2 FILLER_36_1940 ();
 sg13g2_fill_1 FILLER_36_1942 ();
 sg13g2_fill_2 FILLER_36_1951 ();
 sg13g2_fill_1 FILLER_36_1953 ();
 sg13g2_decap_8 FILLER_36_1980 ();
 sg13g2_fill_2 FILLER_36_1987 ();
 sg13g2_fill_2 FILLER_36_1997 ();
 sg13g2_fill_1 FILLER_36_1999 ();
 sg13g2_decap_4 FILLER_36_2032 ();
 sg13g2_fill_2 FILLER_36_2133 ();
 sg13g2_fill_1 FILLER_36_2171 ();
 sg13g2_fill_2 FILLER_36_2202 ();
 sg13g2_fill_1 FILLER_36_2204 ();
 sg13g2_fill_1 FILLER_36_2244 ();
 sg13g2_fill_1 FILLER_36_2249 ();
 sg13g2_fill_1 FILLER_36_2276 ();
 sg13g2_fill_2 FILLER_36_2290 ();
 sg13g2_fill_2 FILLER_36_2300 ();
 sg13g2_fill_1 FILLER_36_2341 ();
 sg13g2_fill_1 FILLER_36_2347 ();
 sg13g2_decap_8 FILLER_36_2374 ();
 sg13g2_decap_8 FILLER_36_2381 ();
 sg13g2_decap_8 FILLER_36_2388 ();
 sg13g2_decap_8 FILLER_36_2395 ();
 sg13g2_decap_8 FILLER_36_2402 ();
 sg13g2_decap_8 FILLER_36_2409 ();
 sg13g2_decap_8 FILLER_36_2416 ();
 sg13g2_decap_8 FILLER_36_2423 ();
 sg13g2_decap_8 FILLER_36_2430 ();
 sg13g2_decap_8 FILLER_36_2437 ();
 sg13g2_decap_8 FILLER_36_2444 ();
 sg13g2_decap_8 FILLER_36_2451 ();
 sg13g2_decap_8 FILLER_36_2458 ();
 sg13g2_decap_8 FILLER_36_2465 ();
 sg13g2_decap_8 FILLER_36_2472 ();
 sg13g2_decap_8 FILLER_36_2479 ();
 sg13g2_decap_8 FILLER_36_2486 ();
 sg13g2_decap_8 FILLER_36_2493 ();
 sg13g2_decap_8 FILLER_36_2500 ();
 sg13g2_decap_8 FILLER_36_2507 ();
 sg13g2_decap_8 FILLER_36_2514 ();
 sg13g2_decap_8 FILLER_36_2521 ();
 sg13g2_decap_8 FILLER_36_2528 ();
 sg13g2_decap_8 FILLER_36_2535 ();
 sg13g2_decap_8 FILLER_36_2542 ();
 sg13g2_decap_8 FILLER_36_2549 ();
 sg13g2_decap_8 FILLER_36_2556 ();
 sg13g2_decap_8 FILLER_36_2563 ();
 sg13g2_decap_8 FILLER_36_2570 ();
 sg13g2_decap_8 FILLER_36_2577 ();
 sg13g2_decap_8 FILLER_36_2584 ();
 sg13g2_decap_8 FILLER_36_2591 ();
 sg13g2_decap_8 FILLER_36_2598 ();
 sg13g2_decap_8 FILLER_36_2605 ();
 sg13g2_decap_8 FILLER_36_2612 ();
 sg13g2_decap_8 FILLER_36_2619 ();
 sg13g2_decap_8 FILLER_36_2626 ();
 sg13g2_decap_8 FILLER_36_2633 ();
 sg13g2_decap_8 FILLER_36_2640 ();
 sg13g2_decap_8 FILLER_36_2647 ();
 sg13g2_decap_8 FILLER_36_2654 ();
 sg13g2_decap_8 FILLER_36_2661 ();
 sg13g2_decap_4 FILLER_36_2668 ();
 sg13g2_fill_2 FILLER_36_2672 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_decap_8 FILLER_37_427 ();
 sg13g2_decap_8 FILLER_37_434 ();
 sg13g2_decap_8 FILLER_37_441 ();
 sg13g2_decap_8 FILLER_37_448 ();
 sg13g2_decap_8 FILLER_37_455 ();
 sg13g2_fill_1 FILLER_37_493 ();
 sg13g2_decap_8 FILLER_37_524 ();
 sg13g2_fill_2 FILLER_37_531 ();
 sg13g2_fill_2 FILLER_37_537 ();
 sg13g2_fill_1 FILLER_37_539 ();
 sg13g2_fill_2 FILLER_37_544 ();
 sg13g2_fill_2 FILLER_37_551 ();
 sg13g2_fill_1 FILLER_37_553 ();
 sg13g2_fill_2 FILLER_37_563 ();
 sg13g2_fill_1 FILLER_37_565 ();
 sg13g2_fill_2 FILLER_37_583 ();
 sg13g2_fill_2 FILLER_37_593 ();
 sg13g2_fill_2 FILLER_37_621 ();
 sg13g2_fill_1 FILLER_37_657 ();
 sg13g2_decap_4 FILLER_37_684 ();
 sg13g2_decap_8 FILLER_37_700 ();
 sg13g2_decap_8 FILLER_37_707 ();
 sg13g2_fill_1 FILLER_37_714 ();
 sg13g2_decap_4 FILLER_37_725 ();
 sg13g2_fill_1 FILLER_37_760 ();
 sg13g2_fill_1 FILLER_37_796 ();
 sg13g2_fill_2 FILLER_37_815 ();
 sg13g2_fill_1 FILLER_37_817 ();
 sg13g2_decap_4 FILLER_37_846 ();
 sg13g2_fill_1 FILLER_37_901 ();
 sg13g2_decap_4 FILLER_37_936 ();
 sg13g2_fill_1 FILLER_37_971 ();
 sg13g2_fill_1 FILLER_37_982 ();
 sg13g2_fill_1 FILLER_37_1014 ();
 sg13g2_fill_1 FILLER_37_1021 ();
 sg13g2_decap_4 FILLER_37_1040 ();
 sg13g2_fill_1 FILLER_37_1048 ();
 sg13g2_fill_2 FILLER_37_1053 ();
 sg13g2_fill_2 FILLER_37_1068 ();
 sg13g2_fill_1 FILLER_37_1110 ();
 sg13g2_fill_1 FILLER_37_1115 ();
 sg13g2_fill_2 FILLER_37_1138 ();
 sg13g2_fill_1 FILLER_37_1209 ();
 sg13g2_fill_1 FILLER_37_1226 ();
 sg13g2_fill_2 FILLER_37_1250 ();
 sg13g2_fill_1 FILLER_37_1258 ();
 sg13g2_decap_8 FILLER_37_1272 ();
 sg13g2_decap_8 FILLER_37_1279 ();
 sg13g2_decap_4 FILLER_37_1286 ();
 sg13g2_fill_1 FILLER_37_1290 ();
 sg13g2_decap_4 FILLER_37_1321 ();
 sg13g2_fill_1 FILLER_37_1325 ();
 sg13g2_decap_8 FILLER_37_1330 ();
 sg13g2_decap_8 FILLER_37_1342 ();
 sg13g2_fill_2 FILLER_37_1358 ();
 sg13g2_fill_1 FILLER_37_1381 ();
 sg13g2_fill_1 FILLER_37_1390 ();
 sg13g2_fill_1 FILLER_37_1426 ();
 sg13g2_fill_2 FILLER_37_1466 ();
 sg13g2_fill_1 FILLER_37_1468 ();
 sg13g2_fill_2 FILLER_37_1477 ();
 sg13g2_fill_1 FILLER_37_1505 ();
 sg13g2_fill_2 FILLER_37_1533 ();
 sg13g2_fill_2 FILLER_37_1562 ();
 sg13g2_fill_1 FILLER_37_1568 ();
 sg13g2_fill_1 FILLER_37_1573 ();
 sg13g2_decap_4 FILLER_37_1583 ();
 sg13g2_fill_2 FILLER_37_1596 ();
 sg13g2_fill_1 FILLER_37_1598 ();
 sg13g2_fill_1 FILLER_37_1631 ();
 sg13g2_decap_8 FILLER_37_1636 ();
 sg13g2_decap_8 FILLER_37_1643 ();
 sg13g2_fill_1 FILLER_37_1663 ();
 sg13g2_decap_4 FILLER_37_1720 ();
 sg13g2_fill_2 FILLER_37_1724 ();
 sg13g2_decap_4 FILLER_37_1753 ();
 sg13g2_fill_1 FILLER_37_1757 ();
 sg13g2_decap_8 FILLER_37_1766 ();
 sg13g2_decap_4 FILLER_37_1773 ();
 sg13g2_decap_4 FILLER_37_1785 ();
 sg13g2_fill_2 FILLER_37_1789 ();
 sg13g2_fill_1 FILLER_37_1804 ();
 sg13g2_decap_8 FILLER_37_1818 ();
 sg13g2_decap_4 FILLER_37_1825 ();
 sg13g2_fill_1 FILLER_37_1859 ();
 sg13g2_decap_4 FILLER_37_1864 ();
 sg13g2_fill_2 FILLER_37_1938 ();
 sg13g2_fill_1 FILLER_37_1940 ();
 sg13g2_fill_1 FILLER_37_1957 ();
 sg13g2_fill_1 FILLER_37_2041 ();
 sg13g2_fill_2 FILLER_37_2067 ();
 sg13g2_fill_1 FILLER_37_2119 ();
 sg13g2_fill_2 FILLER_37_2160 ();
 sg13g2_fill_1 FILLER_37_2162 ();
 sg13g2_fill_1 FILLER_37_2168 ();
 sg13g2_fill_1 FILLER_37_2184 ();
 sg13g2_fill_1 FILLER_37_2208 ();
 sg13g2_decap_4 FILLER_37_2214 ();
 sg13g2_fill_2 FILLER_37_2222 ();
 sg13g2_fill_1 FILLER_37_2224 ();
 sg13g2_fill_2 FILLER_37_2252 ();
 sg13g2_fill_2 FILLER_37_2325 ();
 sg13g2_fill_1 FILLER_37_2327 ();
 sg13g2_fill_2 FILLER_37_2337 ();
 sg13g2_fill_1 FILLER_37_2339 ();
 sg13g2_decap_8 FILLER_37_2371 ();
 sg13g2_decap_8 FILLER_37_2378 ();
 sg13g2_decap_8 FILLER_37_2385 ();
 sg13g2_decap_8 FILLER_37_2392 ();
 sg13g2_decap_8 FILLER_37_2399 ();
 sg13g2_decap_8 FILLER_37_2406 ();
 sg13g2_decap_8 FILLER_37_2413 ();
 sg13g2_decap_8 FILLER_37_2420 ();
 sg13g2_decap_8 FILLER_37_2427 ();
 sg13g2_decap_8 FILLER_37_2434 ();
 sg13g2_decap_8 FILLER_37_2441 ();
 sg13g2_decap_8 FILLER_37_2448 ();
 sg13g2_decap_8 FILLER_37_2455 ();
 sg13g2_decap_8 FILLER_37_2462 ();
 sg13g2_decap_8 FILLER_37_2469 ();
 sg13g2_decap_8 FILLER_37_2476 ();
 sg13g2_decap_8 FILLER_37_2483 ();
 sg13g2_decap_8 FILLER_37_2490 ();
 sg13g2_decap_8 FILLER_37_2497 ();
 sg13g2_decap_8 FILLER_37_2504 ();
 sg13g2_decap_8 FILLER_37_2511 ();
 sg13g2_decap_8 FILLER_37_2518 ();
 sg13g2_decap_8 FILLER_37_2525 ();
 sg13g2_decap_8 FILLER_37_2532 ();
 sg13g2_decap_8 FILLER_37_2539 ();
 sg13g2_decap_8 FILLER_37_2546 ();
 sg13g2_decap_8 FILLER_37_2553 ();
 sg13g2_decap_8 FILLER_37_2560 ();
 sg13g2_decap_8 FILLER_37_2567 ();
 sg13g2_decap_8 FILLER_37_2574 ();
 sg13g2_decap_8 FILLER_37_2581 ();
 sg13g2_decap_8 FILLER_37_2588 ();
 sg13g2_decap_8 FILLER_37_2595 ();
 sg13g2_decap_8 FILLER_37_2602 ();
 sg13g2_decap_8 FILLER_37_2609 ();
 sg13g2_decap_8 FILLER_37_2616 ();
 sg13g2_decap_8 FILLER_37_2623 ();
 sg13g2_decap_8 FILLER_37_2630 ();
 sg13g2_decap_8 FILLER_37_2637 ();
 sg13g2_decap_8 FILLER_37_2644 ();
 sg13g2_decap_8 FILLER_37_2651 ();
 sg13g2_decap_8 FILLER_37_2658 ();
 sg13g2_decap_8 FILLER_37_2665 ();
 sg13g2_fill_2 FILLER_37_2672 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_decap_8 FILLER_38_427 ();
 sg13g2_decap_8 FILLER_38_434 ();
 sg13g2_fill_2 FILLER_38_441 ();
 sg13g2_fill_1 FILLER_38_478 ();
 sg13g2_fill_1 FILLER_38_528 ();
 sg13g2_fill_1 FILLER_38_537 ();
 sg13g2_decap_4 FILLER_38_542 ();
 sg13g2_fill_2 FILLER_38_546 ();
 sg13g2_decap_4 FILLER_38_566 ();
 sg13g2_fill_1 FILLER_38_570 ();
 sg13g2_decap_8 FILLER_38_623 ();
 sg13g2_fill_2 FILLER_38_630 ();
 sg13g2_decap_8 FILLER_38_645 ();
 sg13g2_decap_8 FILLER_38_652 ();
 sg13g2_fill_2 FILLER_38_659 ();
 sg13g2_fill_1 FILLER_38_661 ();
 sg13g2_decap_8 FILLER_38_666 ();
 sg13g2_decap_4 FILLER_38_673 ();
 sg13g2_fill_1 FILLER_38_677 ();
 sg13g2_fill_2 FILLER_38_683 ();
 sg13g2_decap_8 FILLER_38_708 ();
 sg13g2_fill_1 FILLER_38_715 ();
 sg13g2_decap_8 FILLER_38_736 ();
 sg13g2_fill_1 FILLER_38_743 ();
 sg13g2_fill_2 FILLER_38_748 ();
 sg13g2_fill_1 FILLER_38_750 ();
 sg13g2_fill_2 FILLER_38_756 ();
 sg13g2_fill_1 FILLER_38_777 ();
 sg13g2_fill_1 FILLER_38_863 ();
 sg13g2_fill_2 FILLER_38_905 ();
 sg13g2_decap_4 FILLER_38_945 ();
 sg13g2_fill_2 FILLER_38_949 ();
 sg13g2_fill_2 FILLER_38_955 ();
 sg13g2_fill_2 FILLER_38_962 ();
 sg13g2_fill_1 FILLER_38_964 ();
 sg13g2_decap_8 FILLER_38_977 ();
 sg13g2_decap_4 FILLER_38_984 ();
 sg13g2_decap_4 FILLER_38_1009 ();
 sg13g2_fill_1 FILLER_38_1013 ();
 sg13g2_fill_2 FILLER_38_1026 ();
 sg13g2_fill_1 FILLER_38_1028 ();
 sg13g2_fill_2 FILLER_38_1052 ();
 sg13g2_fill_1 FILLER_38_1054 ();
 sg13g2_decap_4 FILLER_38_1068 ();
 sg13g2_fill_1 FILLER_38_1098 ();
 sg13g2_fill_2 FILLER_38_1130 ();
 sg13g2_fill_1 FILLER_38_1132 ();
 sg13g2_decap_8 FILLER_38_1163 ();
 sg13g2_fill_2 FILLER_38_1170 ();
 sg13g2_decap_8 FILLER_38_1180 ();
 sg13g2_fill_1 FILLER_38_1193 ();
 sg13g2_fill_1 FILLER_38_1224 ();
 sg13g2_decap_8 FILLER_38_1243 ();
 sg13g2_fill_2 FILLER_38_1250 ();
 sg13g2_decap_4 FILLER_38_1260 ();
 sg13g2_decap_8 FILLER_38_1320 ();
 sg13g2_fill_1 FILLER_38_1327 ();
 sg13g2_decap_4 FILLER_38_1345 ();
 sg13g2_fill_1 FILLER_38_1349 ();
 sg13g2_fill_2 FILLER_38_1390 ();
 sg13g2_fill_2 FILLER_38_1406 ();
 sg13g2_decap_8 FILLER_38_1480 ();
 sg13g2_fill_2 FILLER_38_1487 ();
 sg13g2_fill_1 FILLER_38_1489 ();
 sg13g2_fill_1 FILLER_38_1518 ();
 sg13g2_decap_8 FILLER_38_1523 ();
 sg13g2_decap_4 FILLER_38_1530 ();
 sg13g2_fill_1 FILLER_38_1534 ();
 sg13g2_decap_4 FILLER_38_1540 ();
 sg13g2_fill_2 FILLER_38_1594 ();
 sg13g2_fill_2 FILLER_38_1604 ();
 sg13g2_fill_1 FILLER_38_1606 ();
 sg13g2_fill_2 FILLER_38_1611 ();
 sg13g2_fill_1 FILLER_38_1613 ();
 sg13g2_fill_1 FILLER_38_1618 ();
 sg13g2_fill_2 FILLER_38_1671 ();
 sg13g2_fill_2 FILLER_38_1677 ();
 sg13g2_fill_1 FILLER_38_1679 ();
 sg13g2_fill_1 FILLER_38_1684 ();
 sg13g2_decap_4 FILLER_38_1694 ();
 sg13g2_decap_4 FILLER_38_1729 ();
 sg13g2_fill_2 FILLER_38_1733 ();
 sg13g2_decap_8 FILLER_38_1739 ();
 sg13g2_fill_2 FILLER_38_1746 ();
 sg13g2_fill_1 FILLER_38_1748 ();
 sg13g2_decap_4 FILLER_38_1777 ();
 sg13g2_fill_1 FILLER_38_1804 ();
 sg13g2_decap_4 FILLER_38_1835 ();
 sg13g2_fill_1 FILLER_38_1883 ();
 sg13g2_fill_2 FILLER_38_1910 ();
 sg13g2_decap_8 FILLER_38_1933 ();
 sg13g2_decap_8 FILLER_38_1940 ();
 sg13g2_fill_2 FILLER_38_1947 ();
 sg13g2_fill_1 FILLER_38_1949 ();
 sg13g2_fill_1 FILLER_38_1955 ();
 sg13g2_fill_1 FILLER_38_1960 ();
 sg13g2_fill_2 FILLER_38_2039 ();
 sg13g2_fill_1 FILLER_38_2041 ();
 sg13g2_fill_2 FILLER_38_2051 ();
 sg13g2_fill_1 FILLER_38_2101 ();
 sg13g2_fill_2 FILLER_38_2105 ();
 sg13g2_fill_2 FILLER_38_2115 ();
 sg13g2_fill_1 FILLER_38_2117 ();
 sg13g2_fill_1 FILLER_38_2169 ();
 sg13g2_fill_2 FILLER_38_2231 ();
 sg13g2_fill_1 FILLER_38_2233 ();
 sg13g2_decap_4 FILLER_38_2296 ();
 sg13g2_fill_1 FILLER_38_2300 ();
 sg13g2_fill_2 FILLER_38_2314 ();
 sg13g2_fill_2 FILLER_38_2326 ();
 sg13g2_decap_8 FILLER_38_2346 ();
 sg13g2_fill_1 FILLER_38_2353 ();
 sg13g2_decap_8 FILLER_38_2371 ();
 sg13g2_decap_8 FILLER_38_2378 ();
 sg13g2_decap_8 FILLER_38_2385 ();
 sg13g2_decap_8 FILLER_38_2392 ();
 sg13g2_decap_8 FILLER_38_2399 ();
 sg13g2_decap_8 FILLER_38_2406 ();
 sg13g2_decap_8 FILLER_38_2413 ();
 sg13g2_decap_8 FILLER_38_2420 ();
 sg13g2_decap_8 FILLER_38_2427 ();
 sg13g2_decap_8 FILLER_38_2434 ();
 sg13g2_decap_8 FILLER_38_2441 ();
 sg13g2_decap_8 FILLER_38_2448 ();
 sg13g2_decap_8 FILLER_38_2455 ();
 sg13g2_decap_8 FILLER_38_2462 ();
 sg13g2_decap_8 FILLER_38_2469 ();
 sg13g2_decap_8 FILLER_38_2476 ();
 sg13g2_decap_8 FILLER_38_2483 ();
 sg13g2_decap_8 FILLER_38_2490 ();
 sg13g2_decap_8 FILLER_38_2497 ();
 sg13g2_decap_8 FILLER_38_2504 ();
 sg13g2_decap_8 FILLER_38_2511 ();
 sg13g2_decap_8 FILLER_38_2518 ();
 sg13g2_decap_8 FILLER_38_2525 ();
 sg13g2_decap_8 FILLER_38_2532 ();
 sg13g2_decap_8 FILLER_38_2539 ();
 sg13g2_decap_8 FILLER_38_2546 ();
 sg13g2_decap_8 FILLER_38_2553 ();
 sg13g2_decap_8 FILLER_38_2560 ();
 sg13g2_decap_8 FILLER_38_2567 ();
 sg13g2_decap_8 FILLER_38_2574 ();
 sg13g2_decap_8 FILLER_38_2581 ();
 sg13g2_decap_8 FILLER_38_2588 ();
 sg13g2_decap_8 FILLER_38_2595 ();
 sg13g2_decap_8 FILLER_38_2602 ();
 sg13g2_decap_8 FILLER_38_2609 ();
 sg13g2_decap_8 FILLER_38_2616 ();
 sg13g2_decap_8 FILLER_38_2623 ();
 sg13g2_decap_8 FILLER_38_2630 ();
 sg13g2_decap_8 FILLER_38_2637 ();
 sg13g2_decap_8 FILLER_38_2644 ();
 sg13g2_decap_8 FILLER_38_2651 ();
 sg13g2_decap_8 FILLER_38_2658 ();
 sg13g2_decap_8 FILLER_38_2665 ();
 sg13g2_fill_2 FILLER_38_2672 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_decap_8 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_238 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_decap_8 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_decap_8 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_336 ();
 sg13g2_decap_8 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_378 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_decap_8 FILLER_39_406 ();
 sg13g2_decap_8 FILLER_39_413 ();
 sg13g2_decap_8 FILLER_39_420 ();
 sg13g2_decap_8 FILLER_39_427 ();
 sg13g2_decap_8 FILLER_39_434 ();
 sg13g2_decap_8 FILLER_39_441 ();
 sg13g2_decap_4 FILLER_39_448 ();
 sg13g2_fill_2 FILLER_39_452 ();
 sg13g2_decap_4 FILLER_39_458 ();
 sg13g2_fill_2 FILLER_39_462 ();
 sg13g2_fill_1 FILLER_39_504 ();
 sg13g2_fill_1 FILLER_39_518 ();
 sg13g2_fill_1 FILLER_39_588 ();
 sg13g2_fill_1 FILLER_39_620 ();
 sg13g2_fill_2 FILLER_39_627 ();
 sg13g2_fill_1 FILLER_39_629 ();
 sg13g2_decap_8 FILLER_39_638 ();
 sg13g2_fill_2 FILLER_39_645 ();
 sg13g2_fill_1 FILLER_39_678 ();
 sg13g2_fill_2 FILLER_39_684 ();
 sg13g2_fill_2 FILLER_39_699 ();
 sg13g2_fill_2 FILLER_39_711 ();
 sg13g2_fill_1 FILLER_39_713 ();
 sg13g2_fill_1 FILLER_39_722 ();
 sg13g2_fill_2 FILLER_39_739 ();
 sg13g2_fill_1 FILLER_39_741 ();
 sg13g2_fill_2 FILLER_39_777 ();
 sg13g2_fill_1 FILLER_39_802 ();
 sg13g2_fill_2 FILLER_39_843 ();
 sg13g2_fill_2 FILLER_39_874 ();
 sg13g2_fill_2 FILLER_39_931 ();
 sg13g2_fill_2 FILLER_39_959 ();
 sg13g2_fill_1 FILLER_39_961 ();
 sg13g2_decap_4 FILLER_39_970 ();
 sg13g2_fill_1 FILLER_39_974 ();
 sg13g2_fill_2 FILLER_39_989 ();
 sg13g2_fill_1 FILLER_39_991 ();
 sg13g2_decap_4 FILLER_39_1011 ();
 sg13g2_fill_2 FILLER_39_1015 ();
 sg13g2_decap_4 FILLER_39_1023 ();
 sg13g2_fill_2 FILLER_39_1045 ();
 sg13g2_fill_2 FILLER_39_1082 ();
 sg13g2_fill_2 FILLER_39_1093 ();
 sg13g2_fill_2 FILLER_39_1108 ();
 sg13g2_decap_8 FILLER_39_1155 ();
 sg13g2_fill_2 FILLER_39_1162 ();
 sg13g2_fill_1 FILLER_39_1164 ();
 sg13g2_fill_2 FILLER_39_1178 ();
 sg13g2_fill_1 FILLER_39_1180 ();
 sg13g2_fill_2 FILLER_39_1252 ();
 sg13g2_fill_1 FILLER_39_1254 ();
 sg13g2_decap_8 FILLER_39_1263 ();
 sg13g2_decap_4 FILLER_39_1270 ();
 sg13g2_fill_2 FILLER_39_1274 ();
 sg13g2_fill_2 FILLER_39_1285 ();
 sg13g2_fill_1 FILLER_39_1287 ();
 sg13g2_fill_1 FILLER_39_1352 ();
 sg13g2_fill_2 FILLER_39_1366 ();
 sg13g2_fill_1 FILLER_39_1368 ();
 sg13g2_fill_2 FILLER_39_1398 ();
 sg13g2_decap_8 FILLER_39_1435 ();
 sg13g2_fill_2 FILLER_39_1442 ();
 sg13g2_fill_1 FILLER_39_1444 ();
 sg13g2_fill_2 FILLER_39_1458 ();
 sg13g2_fill_1 FILLER_39_1534 ();
 sg13g2_fill_1 FILLER_39_1554 ();
 sg13g2_fill_2 FILLER_39_1589 ();
 sg13g2_fill_2 FILLER_39_1596 ();
 sg13g2_fill_1 FILLER_39_1633 ();
 sg13g2_fill_2 FILLER_39_1656 ();
 sg13g2_fill_1 FILLER_39_1658 ();
 sg13g2_fill_1 FILLER_39_1668 ();
 sg13g2_fill_2 FILLER_39_1700 ();
 sg13g2_fill_1 FILLER_39_1702 ();
 sg13g2_fill_2 FILLER_39_1708 ();
 sg13g2_decap_4 FILLER_39_1776 ();
 sg13g2_fill_2 FILLER_39_1780 ();
 sg13g2_fill_1 FILLER_39_1813 ();
 sg13g2_fill_2 FILLER_39_1818 ();
 sg13g2_decap_4 FILLER_39_1824 ();
 sg13g2_fill_2 FILLER_39_1891 ();
 sg13g2_fill_1 FILLER_39_1893 ();
 sg13g2_fill_1 FILLER_39_1985 ();
 sg13g2_fill_1 FILLER_39_2013 ();
 sg13g2_fill_2 FILLER_39_2022 ();
 sg13g2_fill_2 FILLER_39_2038 ();
 sg13g2_fill_1 FILLER_39_2045 ();
 sg13g2_fill_1 FILLER_39_2063 ();
 sg13g2_fill_2 FILLER_39_2072 ();
 sg13g2_fill_2 FILLER_39_2083 ();
 sg13g2_decap_4 FILLER_39_2090 ();
 sg13g2_fill_1 FILLER_39_2098 ();
 sg13g2_fill_1 FILLER_39_2106 ();
 sg13g2_decap_4 FILLER_39_2173 ();
 sg13g2_decap_4 FILLER_39_2190 ();
 sg13g2_fill_2 FILLER_39_2198 ();
 sg13g2_fill_2 FILLER_39_2218 ();
 sg13g2_decap_4 FILLER_39_2246 ();
 sg13g2_fill_1 FILLER_39_2250 ();
 sg13g2_fill_2 FILLER_39_2256 ();
 sg13g2_fill_1 FILLER_39_2258 ();
 sg13g2_fill_2 FILLER_39_2264 ();
 sg13g2_fill_1 FILLER_39_2266 ();
 sg13g2_fill_2 FILLER_39_2280 ();
 sg13g2_decap_8 FILLER_39_2351 ();
 sg13g2_decap_8 FILLER_39_2358 ();
 sg13g2_decap_8 FILLER_39_2365 ();
 sg13g2_decap_8 FILLER_39_2372 ();
 sg13g2_decap_8 FILLER_39_2379 ();
 sg13g2_decap_8 FILLER_39_2386 ();
 sg13g2_decap_8 FILLER_39_2393 ();
 sg13g2_decap_8 FILLER_39_2400 ();
 sg13g2_decap_8 FILLER_39_2407 ();
 sg13g2_decap_8 FILLER_39_2414 ();
 sg13g2_decap_8 FILLER_39_2421 ();
 sg13g2_decap_8 FILLER_39_2428 ();
 sg13g2_decap_8 FILLER_39_2435 ();
 sg13g2_decap_8 FILLER_39_2442 ();
 sg13g2_decap_8 FILLER_39_2449 ();
 sg13g2_decap_8 FILLER_39_2456 ();
 sg13g2_decap_8 FILLER_39_2463 ();
 sg13g2_decap_8 FILLER_39_2470 ();
 sg13g2_decap_8 FILLER_39_2477 ();
 sg13g2_decap_8 FILLER_39_2484 ();
 sg13g2_decap_8 FILLER_39_2491 ();
 sg13g2_decap_8 FILLER_39_2498 ();
 sg13g2_decap_8 FILLER_39_2505 ();
 sg13g2_decap_8 FILLER_39_2512 ();
 sg13g2_decap_8 FILLER_39_2519 ();
 sg13g2_decap_8 FILLER_39_2526 ();
 sg13g2_decap_8 FILLER_39_2533 ();
 sg13g2_decap_8 FILLER_39_2540 ();
 sg13g2_decap_8 FILLER_39_2547 ();
 sg13g2_decap_8 FILLER_39_2554 ();
 sg13g2_decap_8 FILLER_39_2561 ();
 sg13g2_decap_8 FILLER_39_2568 ();
 sg13g2_decap_8 FILLER_39_2575 ();
 sg13g2_decap_8 FILLER_39_2582 ();
 sg13g2_decap_8 FILLER_39_2589 ();
 sg13g2_decap_8 FILLER_39_2596 ();
 sg13g2_decap_8 FILLER_39_2603 ();
 sg13g2_decap_8 FILLER_39_2610 ();
 sg13g2_decap_8 FILLER_39_2617 ();
 sg13g2_decap_8 FILLER_39_2624 ();
 sg13g2_decap_8 FILLER_39_2631 ();
 sg13g2_decap_8 FILLER_39_2638 ();
 sg13g2_decap_8 FILLER_39_2645 ();
 sg13g2_decap_8 FILLER_39_2652 ();
 sg13g2_decap_8 FILLER_39_2659 ();
 sg13g2_decap_8 FILLER_39_2666 ();
 sg13g2_fill_1 FILLER_39_2673 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_decap_8 FILLER_40_315 ();
 sg13g2_decap_8 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_decap_8 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_434 ();
 sg13g2_decap_8 FILLER_40_441 ();
 sg13g2_decap_8 FILLER_40_448 ();
 sg13g2_decap_8 FILLER_40_455 ();
 sg13g2_decap_4 FILLER_40_462 ();
 sg13g2_fill_2 FILLER_40_466 ();
 sg13g2_fill_2 FILLER_40_473 ();
 sg13g2_fill_1 FILLER_40_475 ();
 sg13g2_fill_2 FILLER_40_488 ();
 sg13g2_fill_1 FILLER_40_490 ();
 sg13g2_fill_2 FILLER_40_496 ();
 sg13g2_fill_1 FILLER_40_498 ();
 sg13g2_fill_2 FILLER_40_503 ();
 sg13g2_fill_1 FILLER_40_522 ();
 sg13g2_fill_1 FILLER_40_528 ();
 sg13g2_fill_2 FILLER_40_552 ();
 sg13g2_fill_1 FILLER_40_554 ();
 sg13g2_fill_2 FILLER_40_564 ();
 sg13g2_fill_1 FILLER_40_585 ();
 sg13g2_fill_2 FILLER_40_609 ();
 sg13g2_decap_8 FILLER_40_635 ();
 sg13g2_fill_1 FILLER_40_650 ();
 sg13g2_fill_2 FILLER_40_677 ();
 sg13g2_fill_1 FILLER_40_679 ();
 sg13g2_decap_4 FILLER_40_703 ();
 sg13g2_fill_2 FILLER_40_707 ();
 sg13g2_fill_2 FILLER_40_723 ();
 sg13g2_fill_1 FILLER_40_725 ();
 sg13g2_decap_8 FILLER_40_736 ();
 sg13g2_fill_2 FILLER_40_770 ();
 sg13g2_fill_1 FILLER_40_772 ();
 sg13g2_fill_2 FILLER_40_816 ();
 sg13g2_fill_2 FILLER_40_828 ();
 sg13g2_fill_2 FILLER_40_835 ();
 sg13g2_fill_1 FILLER_40_837 ();
 sg13g2_decap_4 FILLER_40_897 ();
 sg13g2_fill_2 FILLER_40_914 ();
 sg13g2_fill_2 FILLER_40_920 ();
 sg13g2_fill_1 FILLER_40_922 ();
 sg13g2_fill_2 FILLER_40_942 ();
 sg13g2_decap_8 FILLER_40_948 ();
 sg13g2_fill_2 FILLER_40_955 ();
 sg13g2_fill_2 FILLER_40_965 ();
 sg13g2_fill_1 FILLER_40_967 ();
 sg13g2_decap_4 FILLER_40_981 ();
 sg13g2_fill_1 FILLER_40_985 ();
 sg13g2_fill_1 FILLER_40_993 ();
 sg13g2_fill_1 FILLER_40_1019 ();
 sg13g2_fill_2 FILLER_40_1075 ();
 sg13g2_fill_1 FILLER_40_1077 ();
 sg13g2_fill_2 FILLER_40_1104 ();
 sg13g2_fill_1 FILLER_40_1106 ();
 sg13g2_decap_8 FILLER_40_1152 ();
 sg13g2_fill_2 FILLER_40_1163 ();
 sg13g2_fill_1 FILLER_40_1165 ();
 sg13g2_fill_1 FILLER_40_1172 ();
 sg13g2_decap_4 FILLER_40_1179 ();
 sg13g2_fill_1 FILLER_40_1189 ();
 sg13g2_fill_2 FILLER_40_1203 ();
 sg13g2_fill_1 FILLER_40_1218 ();
 sg13g2_decap_4 FILLER_40_1270 ();
 sg13g2_fill_2 FILLER_40_1274 ();
 sg13g2_fill_1 FILLER_40_1288 ();
 sg13g2_fill_2 FILLER_40_1306 ();
 sg13g2_fill_1 FILLER_40_1308 ();
 sg13g2_fill_1 FILLER_40_1314 ();
 sg13g2_decap_8 FILLER_40_1329 ();
 sg13g2_fill_2 FILLER_40_1336 ();
 sg13g2_fill_2 FILLER_40_1343 ();
 sg13g2_fill_2 FILLER_40_1368 ();
 sg13g2_fill_1 FILLER_40_1370 ();
 sg13g2_fill_1 FILLER_40_1419 ();
 sg13g2_decap_4 FILLER_40_1459 ();
 sg13g2_decap_4 FILLER_40_1485 ();
 sg13g2_fill_2 FILLER_40_1489 ();
 sg13g2_fill_2 FILLER_40_1521 ();
 sg13g2_decap_4 FILLER_40_1543 ();
 sg13g2_fill_1 FILLER_40_1547 ();
 sg13g2_fill_1 FILLER_40_1590 ();
 sg13g2_fill_2 FILLER_40_1617 ();
 sg13g2_decap_4 FILLER_40_1632 ();
 sg13g2_fill_2 FILLER_40_1636 ();
 sg13g2_fill_2 FILLER_40_1690 ();
 sg13g2_fill_2 FILLER_40_1701 ();
 sg13g2_fill_1 FILLER_40_1703 ();
 sg13g2_fill_1 FILLER_40_1713 ();
 sg13g2_fill_1 FILLER_40_1722 ();
 sg13g2_fill_2 FILLER_40_1732 ();
 sg13g2_fill_2 FILLER_40_1738 ();
 sg13g2_fill_1 FILLER_40_1797 ();
 sg13g2_decap_8 FILLER_40_1834 ();
 sg13g2_decap_4 FILLER_40_1841 ();
 sg13g2_fill_1 FILLER_40_1845 ();
 sg13g2_decap_4 FILLER_40_1898 ();
 sg13g2_fill_1 FILLER_40_1902 ();
 sg13g2_decap_8 FILLER_40_1916 ();
 sg13g2_fill_1 FILLER_40_1935 ();
 sg13g2_fill_2 FILLER_40_1940 ();
 sg13g2_fill_1 FILLER_40_1951 ();
 sg13g2_fill_2 FILLER_40_2001 ();
 sg13g2_fill_2 FILLER_40_2086 ();
 sg13g2_fill_1 FILLER_40_2088 ();
 sg13g2_fill_2 FILLER_40_2098 ();
 sg13g2_fill_2 FILLER_40_2104 ();
 sg13g2_fill_1 FILLER_40_2106 ();
 sg13g2_fill_2 FILLER_40_2127 ();
 sg13g2_fill_1 FILLER_40_2129 ();
 sg13g2_fill_2 FILLER_40_2143 ();
 sg13g2_fill_1 FILLER_40_2145 ();
 sg13g2_fill_1 FILLER_40_2163 ();
 sg13g2_fill_2 FILLER_40_2178 ();
 sg13g2_fill_1 FILLER_40_2180 ();
 sg13g2_fill_1 FILLER_40_2210 ();
 sg13g2_fill_1 FILLER_40_2224 ();
 sg13g2_fill_1 FILLER_40_2234 ();
 sg13g2_decap_4 FILLER_40_2249 ();
 sg13g2_fill_1 FILLER_40_2253 ();
 sg13g2_fill_2 FILLER_40_2272 ();
 sg13g2_decap_4 FILLER_40_2283 ();
 sg13g2_fill_1 FILLER_40_2287 ();
 sg13g2_fill_2 FILLER_40_2297 ();
 sg13g2_decap_4 FILLER_40_2303 ();
 sg13g2_fill_2 FILLER_40_2321 ();
 sg13g2_fill_1 FILLER_40_2323 ();
 sg13g2_decap_8 FILLER_40_2347 ();
 sg13g2_decap_8 FILLER_40_2354 ();
 sg13g2_decap_8 FILLER_40_2361 ();
 sg13g2_decap_8 FILLER_40_2368 ();
 sg13g2_decap_8 FILLER_40_2375 ();
 sg13g2_decap_8 FILLER_40_2382 ();
 sg13g2_decap_8 FILLER_40_2389 ();
 sg13g2_decap_8 FILLER_40_2396 ();
 sg13g2_decap_8 FILLER_40_2403 ();
 sg13g2_decap_8 FILLER_40_2410 ();
 sg13g2_decap_8 FILLER_40_2417 ();
 sg13g2_decap_8 FILLER_40_2424 ();
 sg13g2_decap_8 FILLER_40_2431 ();
 sg13g2_decap_8 FILLER_40_2438 ();
 sg13g2_decap_8 FILLER_40_2445 ();
 sg13g2_decap_8 FILLER_40_2452 ();
 sg13g2_decap_8 FILLER_40_2459 ();
 sg13g2_decap_8 FILLER_40_2466 ();
 sg13g2_decap_8 FILLER_40_2473 ();
 sg13g2_decap_8 FILLER_40_2480 ();
 sg13g2_decap_8 FILLER_40_2487 ();
 sg13g2_decap_8 FILLER_40_2494 ();
 sg13g2_decap_8 FILLER_40_2501 ();
 sg13g2_decap_8 FILLER_40_2508 ();
 sg13g2_decap_8 FILLER_40_2515 ();
 sg13g2_decap_8 FILLER_40_2522 ();
 sg13g2_decap_8 FILLER_40_2529 ();
 sg13g2_decap_8 FILLER_40_2536 ();
 sg13g2_decap_8 FILLER_40_2543 ();
 sg13g2_decap_8 FILLER_40_2550 ();
 sg13g2_decap_8 FILLER_40_2557 ();
 sg13g2_decap_8 FILLER_40_2564 ();
 sg13g2_decap_8 FILLER_40_2571 ();
 sg13g2_decap_8 FILLER_40_2578 ();
 sg13g2_decap_8 FILLER_40_2585 ();
 sg13g2_decap_8 FILLER_40_2592 ();
 sg13g2_decap_8 FILLER_40_2599 ();
 sg13g2_decap_8 FILLER_40_2606 ();
 sg13g2_decap_8 FILLER_40_2613 ();
 sg13g2_decap_8 FILLER_40_2620 ();
 sg13g2_decap_8 FILLER_40_2627 ();
 sg13g2_decap_8 FILLER_40_2634 ();
 sg13g2_decap_8 FILLER_40_2641 ();
 sg13g2_decap_8 FILLER_40_2648 ();
 sg13g2_decap_8 FILLER_40_2655 ();
 sg13g2_decap_8 FILLER_40_2662 ();
 sg13g2_decap_4 FILLER_40_2669 ();
 sg13g2_fill_1 FILLER_40_2673 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_287 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_308 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_decap_8 FILLER_41_420 ();
 sg13g2_decap_8 FILLER_41_427 ();
 sg13g2_decap_8 FILLER_41_434 ();
 sg13g2_decap_8 FILLER_41_441 ();
 sg13g2_decap_8 FILLER_41_448 ();
 sg13g2_fill_1 FILLER_41_455 ();
 sg13g2_fill_2 FILLER_41_486 ();
 sg13g2_fill_2 FILLER_41_614 ();
 sg13g2_decap_8 FILLER_41_666 ();
 sg13g2_fill_2 FILLER_41_673 ();
 sg13g2_fill_1 FILLER_41_684 ();
 sg13g2_decap_4 FILLER_41_694 ();
 sg13g2_fill_2 FILLER_41_698 ();
 sg13g2_fill_2 FILLER_41_729 ();
 sg13g2_fill_1 FILLER_41_736 ();
 sg13g2_decap_4 FILLER_41_741 ();
 sg13g2_fill_2 FILLER_41_745 ();
 sg13g2_fill_2 FILLER_41_752 ();
 sg13g2_decap_4 FILLER_41_764 ();
 sg13g2_fill_2 FILLER_41_768 ();
 sg13g2_fill_2 FILLER_41_774 ();
 sg13g2_fill_2 FILLER_41_788 ();
 sg13g2_fill_2 FILLER_41_805 ();
 sg13g2_fill_1 FILLER_41_807 ();
 sg13g2_fill_1 FILLER_41_817 ();
 sg13g2_fill_1 FILLER_41_832 ();
 sg13g2_fill_1 FILLER_41_865 ();
 sg13g2_decap_4 FILLER_41_893 ();
 sg13g2_fill_1 FILLER_41_931 ();
 sg13g2_decap_4 FILLER_41_935 ();
 sg13g2_fill_1 FILLER_41_965 ();
 sg13g2_decap_8 FILLER_41_996 ();
 sg13g2_decap_4 FILLER_41_1003 ();
 sg13g2_decap_8 FILLER_41_1026 ();
 sg13g2_decap_8 FILLER_41_1033 ();
 sg13g2_decap_8 FILLER_41_1040 ();
 sg13g2_fill_1 FILLER_41_1047 ();
 sg13g2_fill_2 FILLER_41_1056 ();
 sg13g2_fill_2 FILLER_41_1102 ();
 sg13g2_fill_1 FILLER_41_1104 ();
 sg13g2_fill_2 FILLER_41_1123 ();
 sg13g2_fill_1 FILLER_41_1129 ();
 sg13g2_fill_1 FILLER_41_1139 ();
 sg13g2_fill_2 FILLER_41_1175 ();
 sg13g2_fill_1 FILLER_41_1177 ();
 sg13g2_decap_8 FILLER_41_1182 ();
 sg13g2_decap_8 FILLER_41_1189 ();
 sg13g2_decap_4 FILLER_41_1196 ();
 sg13g2_fill_2 FILLER_41_1200 ();
 sg13g2_fill_2 FILLER_41_1208 ();
 sg13g2_fill_1 FILLER_41_1210 ();
 sg13g2_fill_2 FILLER_41_1229 ();
 sg13g2_fill_1 FILLER_41_1231 ();
 sg13g2_fill_2 FILLER_41_1291 ();
 sg13g2_fill_1 FILLER_41_1319 ();
 sg13g2_decap_4 FILLER_41_1351 ();
 sg13g2_fill_2 FILLER_41_1360 ();
 sg13g2_fill_1 FILLER_41_1362 ();
 sg13g2_decap_4 FILLER_41_1374 ();
 sg13g2_fill_2 FILLER_41_1378 ();
 sg13g2_fill_2 FILLER_41_1411 ();
 sg13g2_fill_2 FILLER_41_1446 ();
 sg13g2_fill_2 FILLER_41_1454 ();
 sg13g2_fill_2 FILLER_41_1513 ();
 sg13g2_fill_1 FILLER_41_1519 ();
 sg13g2_fill_1 FILLER_41_1524 ();
 sg13g2_fill_2 FILLER_41_1530 ();
 sg13g2_fill_1 FILLER_41_1532 ();
 sg13g2_fill_2 FILLER_41_1552 ();
 sg13g2_fill_2 FILLER_41_1568 ();
 sg13g2_decap_8 FILLER_41_1646 ();
 sg13g2_fill_2 FILLER_41_1653 ();
 sg13g2_fill_2 FILLER_41_1660 ();
 sg13g2_fill_1 FILLER_41_1801 ();
 sg13g2_fill_2 FILLER_41_1815 ();
 sg13g2_fill_2 FILLER_41_1826 ();
 sg13g2_fill_1 FILLER_41_1828 ();
 sg13g2_fill_2 FILLER_41_1847 ();
 sg13g2_decap_4 FILLER_41_1854 ();
 sg13g2_fill_1 FILLER_41_1858 ();
 sg13g2_decap_4 FILLER_41_1867 ();
 sg13g2_fill_1 FILLER_41_1892 ();
 sg13g2_decap_4 FILLER_41_1902 ();
 sg13g2_fill_1 FILLER_41_1906 ();
 sg13g2_decap_4 FILLER_41_2002 ();
 sg13g2_fill_1 FILLER_41_2006 ();
 sg13g2_decap_4 FILLER_41_2011 ();
 sg13g2_decap_4 FILLER_41_2032 ();
 sg13g2_fill_1 FILLER_41_2036 ();
 sg13g2_fill_2 FILLER_41_2050 ();
 sg13g2_fill_1 FILLER_41_2052 ();
 sg13g2_decap_4 FILLER_41_2057 ();
 sg13g2_fill_1 FILLER_41_2061 ();
 sg13g2_fill_2 FILLER_41_2066 ();
 sg13g2_decap_4 FILLER_41_2077 ();
 sg13g2_fill_2 FILLER_41_2081 ();
 sg13g2_fill_1 FILLER_41_2088 ();
 sg13g2_decap_4 FILLER_41_2115 ();
 sg13g2_fill_2 FILLER_41_2119 ();
 sg13g2_decap_8 FILLER_41_2142 ();
 sg13g2_decap_8 FILLER_41_2149 ();
 sg13g2_fill_1 FILLER_41_2166 ();
 sg13g2_fill_2 FILLER_41_2193 ();
 sg13g2_fill_1 FILLER_41_2195 ();
 sg13g2_fill_2 FILLER_41_2227 ();
 sg13g2_fill_1 FILLER_41_2229 ();
 sg13g2_fill_1 FILLER_41_2313 ();
 sg13g2_decap_8 FILLER_41_2344 ();
 sg13g2_decap_8 FILLER_41_2351 ();
 sg13g2_decap_8 FILLER_41_2358 ();
 sg13g2_decap_8 FILLER_41_2365 ();
 sg13g2_decap_8 FILLER_41_2372 ();
 sg13g2_decap_8 FILLER_41_2379 ();
 sg13g2_decap_8 FILLER_41_2386 ();
 sg13g2_decap_8 FILLER_41_2393 ();
 sg13g2_decap_8 FILLER_41_2400 ();
 sg13g2_decap_8 FILLER_41_2407 ();
 sg13g2_decap_8 FILLER_41_2414 ();
 sg13g2_decap_8 FILLER_41_2421 ();
 sg13g2_decap_8 FILLER_41_2428 ();
 sg13g2_decap_8 FILLER_41_2435 ();
 sg13g2_decap_8 FILLER_41_2442 ();
 sg13g2_decap_8 FILLER_41_2449 ();
 sg13g2_decap_8 FILLER_41_2456 ();
 sg13g2_decap_8 FILLER_41_2463 ();
 sg13g2_decap_8 FILLER_41_2470 ();
 sg13g2_decap_8 FILLER_41_2477 ();
 sg13g2_decap_8 FILLER_41_2484 ();
 sg13g2_decap_8 FILLER_41_2491 ();
 sg13g2_decap_8 FILLER_41_2498 ();
 sg13g2_decap_8 FILLER_41_2505 ();
 sg13g2_decap_8 FILLER_41_2512 ();
 sg13g2_decap_8 FILLER_41_2519 ();
 sg13g2_decap_8 FILLER_41_2526 ();
 sg13g2_decap_8 FILLER_41_2533 ();
 sg13g2_decap_8 FILLER_41_2540 ();
 sg13g2_decap_8 FILLER_41_2547 ();
 sg13g2_decap_8 FILLER_41_2554 ();
 sg13g2_decap_8 FILLER_41_2561 ();
 sg13g2_decap_8 FILLER_41_2568 ();
 sg13g2_decap_8 FILLER_41_2575 ();
 sg13g2_decap_8 FILLER_41_2582 ();
 sg13g2_decap_8 FILLER_41_2589 ();
 sg13g2_decap_8 FILLER_41_2596 ();
 sg13g2_decap_8 FILLER_41_2603 ();
 sg13g2_decap_8 FILLER_41_2610 ();
 sg13g2_decap_8 FILLER_41_2617 ();
 sg13g2_decap_8 FILLER_41_2624 ();
 sg13g2_decap_8 FILLER_41_2631 ();
 sg13g2_decap_8 FILLER_41_2638 ();
 sg13g2_decap_8 FILLER_41_2645 ();
 sg13g2_decap_8 FILLER_41_2652 ();
 sg13g2_decap_8 FILLER_41_2659 ();
 sg13g2_decap_8 FILLER_41_2666 ();
 sg13g2_fill_1 FILLER_41_2673 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_196 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_decap_8 FILLER_42_273 ();
 sg13g2_decap_8 FILLER_42_280 ();
 sg13g2_decap_8 FILLER_42_287 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_decap_8 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_378 ();
 sg13g2_decap_8 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_decap_8 FILLER_42_406 ();
 sg13g2_decap_8 FILLER_42_413 ();
 sg13g2_decap_8 FILLER_42_420 ();
 sg13g2_decap_8 FILLER_42_427 ();
 sg13g2_decap_8 FILLER_42_434 ();
 sg13g2_decap_8 FILLER_42_441 ();
 sg13g2_decap_8 FILLER_42_448 ();
 sg13g2_decap_8 FILLER_42_455 ();
 sg13g2_decap_4 FILLER_42_462 ();
 sg13g2_fill_1 FILLER_42_466 ();
 sg13g2_decap_8 FILLER_42_471 ();
 sg13g2_decap_4 FILLER_42_504 ();
 sg13g2_fill_1 FILLER_42_508 ();
 sg13g2_fill_1 FILLER_42_540 ();
 sg13g2_decap_4 FILLER_42_546 ();
 sg13g2_fill_2 FILLER_42_559 ();
 sg13g2_fill_1 FILLER_42_561 ();
 sg13g2_fill_2 FILLER_42_566 ();
 sg13g2_decap_4 FILLER_42_573 ();
 sg13g2_fill_1 FILLER_42_577 ();
 sg13g2_fill_2 FILLER_42_587 ();
 sg13g2_fill_2 FILLER_42_619 ();
 sg13g2_fill_2 FILLER_42_634 ();
 sg13g2_fill_1 FILLER_42_636 ();
 sg13g2_decap_8 FILLER_42_645 ();
 sg13g2_fill_2 FILLER_42_652 ();
 sg13g2_fill_2 FILLER_42_680 ();
 sg13g2_fill_1 FILLER_42_682 ();
 sg13g2_fill_2 FILLER_42_688 ();
 sg13g2_fill_2 FILLER_42_811 ();
 sg13g2_fill_2 FILLER_42_823 ();
 sg13g2_decap_8 FILLER_42_860 ();
 sg13g2_decap_8 FILLER_42_867 ();
 sg13g2_fill_2 FILLER_42_874 ();
 sg13g2_decap_4 FILLER_42_880 ();
 sg13g2_decap_8 FILLER_42_904 ();
 sg13g2_decap_4 FILLER_42_911 ();
 sg13g2_fill_1 FILLER_42_915 ();
 sg13g2_decap_4 FILLER_42_920 ();
 sg13g2_fill_2 FILLER_42_924 ();
 sg13g2_fill_2 FILLER_42_929 ();
 sg13g2_fill_2 FILLER_42_950 ();
 sg13g2_fill_1 FILLER_42_952 ();
 sg13g2_decap_4 FILLER_42_962 ();
 sg13g2_decap_8 FILLER_42_971 ();
 sg13g2_fill_1 FILLER_42_978 ();
 sg13g2_decap_4 FILLER_42_1005 ();
 sg13g2_fill_2 FILLER_42_1009 ();
 sg13g2_fill_1 FILLER_42_1024 ();
 sg13g2_fill_2 FILLER_42_1030 ();
 sg13g2_fill_1 FILLER_42_1032 ();
 sg13g2_fill_2 FILLER_42_1058 ();
 sg13g2_fill_1 FILLER_42_1068 ();
 sg13g2_fill_1 FILLER_42_1074 ();
 sg13g2_decap_4 FILLER_42_1079 ();
 sg13g2_fill_1 FILLER_42_1083 ();
 sg13g2_fill_2 FILLER_42_1156 ();
 sg13g2_fill_1 FILLER_42_1238 ();
 sg13g2_decap_8 FILLER_42_1286 ();
 sg13g2_decap_8 FILLER_42_1293 ();
 sg13g2_decap_8 FILLER_42_1300 ();
 sg13g2_decap_4 FILLER_42_1307 ();
 sg13g2_fill_2 FILLER_42_1311 ();
 sg13g2_fill_1 FILLER_42_1330 ();
 sg13g2_decap_4 FILLER_42_1335 ();
 sg13g2_fill_1 FILLER_42_1339 ();
 sg13g2_fill_1 FILLER_42_1353 ();
 sg13g2_fill_2 FILLER_42_1397 ();
 sg13g2_fill_2 FILLER_42_1408 ();
 sg13g2_fill_2 FILLER_42_1427 ();
 sg13g2_fill_1 FILLER_42_1454 ();
 sg13g2_decap_4 FILLER_42_1468 ();
 sg13g2_fill_2 FILLER_42_1472 ();
 sg13g2_decap_8 FILLER_42_1479 ();
 sg13g2_decap_8 FILLER_42_1486 ();
 sg13g2_decap_8 FILLER_42_1497 ();
 sg13g2_fill_2 FILLER_42_1504 ();
 sg13g2_fill_2 FILLER_42_1511 ();
 sg13g2_decap_8 FILLER_42_1548 ();
 sg13g2_fill_2 FILLER_42_1555 ();
 sg13g2_fill_1 FILLER_42_1557 ();
 sg13g2_fill_2 FILLER_42_1563 ();
 sg13g2_fill_2 FILLER_42_1582 ();
 sg13g2_fill_1 FILLER_42_1584 ();
 sg13g2_fill_1 FILLER_42_1599 ();
 sg13g2_decap_8 FILLER_42_1613 ();
 sg13g2_fill_2 FILLER_42_1665 ();
 sg13g2_fill_1 FILLER_42_1706 ();
 sg13g2_fill_1 FILLER_42_1716 ();
 sg13g2_fill_1 FILLER_42_1721 ();
 sg13g2_decap_4 FILLER_42_1743 ();
 sg13g2_fill_2 FILLER_42_1751 ();
 sg13g2_fill_2 FILLER_42_1762 ();
 sg13g2_decap_4 FILLER_42_1777 ();
 sg13g2_fill_2 FILLER_42_1816 ();
 sg13g2_fill_1 FILLER_42_1818 ();
 sg13g2_fill_1 FILLER_42_1876 ();
 sg13g2_fill_1 FILLER_42_1893 ();
 sg13g2_decap_8 FILLER_42_1905 ();
 sg13g2_decap_8 FILLER_42_1912 ();
 sg13g2_fill_2 FILLER_42_1919 ();
 sg13g2_decap_8 FILLER_42_1925 ();
 sg13g2_decap_4 FILLER_42_1932 ();
 sg13g2_fill_2 FILLER_42_1936 ();
 sg13g2_fill_2 FILLER_42_1947 ();
 sg13g2_fill_2 FILLER_42_1966 ();
 sg13g2_fill_1 FILLER_42_1968 ();
 sg13g2_fill_1 FILLER_42_2052 ();
 sg13g2_fill_1 FILLER_42_2062 ();
 sg13g2_fill_2 FILLER_42_2067 ();
 sg13g2_fill_2 FILLER_42_2083 ();
 sg13g2_fill_1 FILLER_42_2085 ();
 sg13g2_decap_8 FILLER_42_2099 ();
 sg13g2_decap_4 FILLER_42_2171 ();
 sg13g2_fill_2 FILLER_42_2175 ();
 sg13g2_fill_2 FILLER_42_2185 ();
 sg13g2_fill_1 FILLER_42_2187 ();
 sg13g2_decap_4 FILLER_42_2232 ();
 sg13g2_fill_1 FILLER_42_2236 ();
 sg13g2_decap_4 FILLER_42_2241 ();
 sg13g2_fill_1 FILLER_42_2249 ();
 sg13g2_decap_8 FILLER_42_2259 ();
 sg13g2_fill_1 FILLER_42_2266 ();
 sg13g2_decap_4 FILLER_42_2271 ();
 sg13g2_decap_8 FILLER_42_2279 ();
 sg13g2_decap_8 FILLER_42_2286 ();
 sg13g2_fill_2 FILLER_42_2293 ();
 sg13g2_decap_8 FILLER_42_2304 ();
 sg13g2_decap_8 FILLER_42_2345 ();
 sg13g2_decap_8 FILLER_42_2352 ();
 sg13g2_decap_8 FILLER_42_2359 ();
 sg13g2_decap_8 FILLER_42_2366 ();
 sg13g2_decap_8 FILLER_42_2373 ();
 sg13g2_decap_8 FILLER_42_2380 ();
 sg13g2_decap_8 FILLER_42_2387 ();
 sg13g2_decap_8 FILLER_42_2394 ();
 sg13g2_decap_8 FILLER_42_2401 ();
 sg13g2_decap_8 FILLER_42_2408 ();
 sg13g2_decap_8 FILLER_42_2415 ();
 sg13g2_decap_8 FILLER_42_2422 ();
 sg13g2_decap_8 FILLER_42_2429 ();
 sg13g2_decap_8 FILLER_42_2436 ();
 sg13g2_decap_8 FILLER_42_2443 ();
 sg13g2_decap_8 FILLER_42_2450 ();
 sg13g2_decap_8 FILLER_42_2457 ();
 sg13g2_decap_8 FILLER_42_2464 ();
 sg13g2_decap_8 FILLER_42_2471 ();
 sg13g2_decap_8 FILLER_42_2478 ();
 sg13g2_decap_8 FILLER_42_2485 ();
 sg13g2_decap_8 FILLER_42_2492 ();
 sg13g2_decap_8 FILLER_42_2499 ();
 sg13g2_decap_8 FILLER_42_2506 ();
 sg13g2_decap_8 FILLER_42_2513 ();
 sg13g2_decap_8 FILLER_42_2520 ();
 sg13g2_decap_8 FILLER_42_2527 ();
 sg13g2_decap_8 FILLER_42_2534 ();
 sg13g2_decap_8 FILLER_42_2541 ();
 sg13g2_decap_8 FILLER_42_2548 ();
 sg13g2_decap_8 FILLER_42_2555 ();
 sg13g2_decap_8 FILLER_42_2562 ();
 sg13g2_decap_8 FILLER_42_2569 ();
 sg13g2_decap_8 FILLER_42_2576 ();
 sg13g2_decap_8 FILLER_42_2583 ();
 sg13g2_decap_8 FILLER_42_2590 ();
 sg13g2_decap_8 FILLER_42_2597 ();
 sg13g2_decap_8 FILLER_42_2604 ();
 sg13g2_decap_8 FILLER_42_2611 ();
 sg13g2_decap_8 FILLER_42_2618 ();
 sg13g2_decap_8 FILLER_42_2625 ();
 sg13g2_decap_8 FILLER_42_2632 ();
 sg13g2_decap_8 FILLER_42_2639 ();
 sg13g2_decap_8 FILLER_42_2646 ();
 sg13g2_decap_8 FILLER_42_2653 ();
 sg13g2_decap_8 FILLER_42_2660 ();
 sg13g2_decap_8 FILLER_42_2667 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_266 ();
 sg13g2_decap_8 FILLER_43_273 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_decap_8 FILLER_43_301 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_315 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_decap_8 FILLER_43_427 ();
 sg13g2_decap_8 FILLER_43_434 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_8 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_455 ();
 sg13g2_decap_8 FILLER_43_462 ();
 sg13g2_decap_8 FILLER_43_469 ();
 sg13g2_fill_2 FILLER_43_507 ();
 sg13g2_fill_1 FILLER_43_509 ();
 sg13g2_fill_1 FILLER_43_524 ();
 sg13g2_fill_2 FILLER_43_529 ();
 sg13g2_decap_8 FILLER_43_540 ();
 sg13g2_fill_1 FILLER_43_547 ();
 sg13g2_fill_1 FILLER_43_578 ();
 sg13g2_fill_2 FILLER_43_609 ();
 sg13g2_decap_4 FILLER_43_619 ();
 sg13g2_fill_2 FILLER_43_623 ();
 sg13g2_fill_2 FILLER_43_671 ();
 sg13g2_fill_2 FILLER_43_699 ();
 sg13g2_fill_1 FILLER_43_715 ();
 sg13g2_fill_2 FILLER_43_721 ();
 sg13g2_decap_8 FILLER_43_736 ();
 sg13g2_fill_2 FILLER_43_743 ();
 sg13g2_decap_8 FILLER_43_768 ();
 sg13g2_fill_1 FILLER_43_775 ();
 sg13g2_fill_2 FILLER_43_790 ();
 sg13g2_fill_2 FILLER_43_797 ();
 sg13g2_fill_2 FILLER_43_813 ();
 sg13g2_fill_1 FILLER_43_815 ();
 sg13g2_fill_2 FILLER_43_824 ();
 sg13g2_decap_4 FILLER_43_852 ();
 sg13g2_fill_2 FILLER_43_896 ();
 sg13g2_fill_1 FILLER_43_898 ();
 sg13g2_fill_1 FILLER_43_925 ();
 sg13g2_fill_2 FILLER_43_941 ();
 sg13g2_fill_2 FILLER_43_953 ();
 sg13g2_fill_1 FILLER_43_955 ();
 sg13g2_decap_8 FILLER_43_970 ();
 sg13g2_decap_4 FILLER_43_977 ();
 sg13g2_fill_2 FILLER_43_981 ();
 sg13g2_fill_1 FILLER_43_992 ();
 sg13g2_decap_8 FILLER_43_1000 ();
 sg13g2_fill_2 FILLER_43_1007 ();
 sg13g2_fill_2 FILLER_43_1048 ();
 sg13g2_decap_8 FILLER_43_1125 ();
 sg13g2_fill_2 FILLER_43_1203 ();
 sg13g2_fill_1 FILLER_43_1205 ();
 sg13g2_fill_2 FILLER_43_1211 ();
 sg13g2_decap_4 FILLER_43_1222 ();
 sg13g2_fill_2 FILLER_43_1226 ();
 sg13g2_fill_2 FILLER_43_1246 ();
 sg13g2_fill_1 FILLER_43_1248 ();
 sg13g2_decap_4 FILLER_43_1327 ();
 sg13g2_fill_2 FILLER_43_1357 ();
 sg13g2_fill_1 FILLER_43_1359 ();
 sg13g2_fill_2 FILLER_43_1392 ();
 sg13g2_fill_1 FILLER_43_1394 ();
 sg13g2_fill_1 FILLER_43_1412 ();
 sg13g2_fill_2 FILLER_43_1416 ();
 sg13g2_fill_1 FILLER_43_1423 ();
 sg13g2_fill_2 FILLER_43_1433 ();
 sg13g2_decap_4 FILLER_43_1476 ();
 sg13g2_fill_2 FILLER_43_1510 ();
 sg13g2_fill_1 FILLER_43_1512 ();
 sg13g2_decap_8 FILLER_43_1518 ();
 sg13g2_fill_2 FILLER_43_1525 ();
 sg13g2_fill_1 FILLER_43_1527 ();
 sg13g2_fill_1 FILLER_43_1532 ();
 sg13g2_fill_2 FILLER_43_1559 ();
 sg13g2_fill_2 FILLER_43_1579 ();
 sg13g2_fill_2 FILLER_43_1616 ();
 sg13g2_fill_1 FILLER_43_1618 ();
 sg13g2_decap_8 FILLER_43_1623 ();
 sg13g2_fill_2 FILLER_43_1630 ();
 sg13g2_fill_1 FILLER_43_1692 ();
 sg13g2_fill_2 FILLER_43_1703 ();
 sg13g2_fill_1 FILLER_43_1705 ();
 sg13g2_decap_8 FILLER_43_1736 ();
 sg13g2_decap_8 FILLER_43_1743 ();
 sg13g2_decap_4 FILLER_43_1788 ();
 sg13g2_fill_1 FILLER_43_1792 ();
 sg13g2_fill_2 FILLER_43_1806 ();
 sg13g2_fill_1 FILLER_43_1808 ();
 sg13g2_decap_8 FILLER_43_1839 ();
 sg13g2_fill_2 FILLER_43_1846 ();
 sg13g2_fill_2 FILLER_43_1857 ();
 sg13g2_fill_1 FILLER_43_1859 ();
 sg13g2_fill_1 FILLER_43_1864 ();
 sg13g2_decap_8 FILLER_43_1874 ();
 sg13g2_fill_2 FILLER_43_1881 ();
 sg13g2_fill_1 FILLER_43_1883 ();
 sg13g2_decap_8 FILLER_43_1901 ();
 sg13g2_decap_8 FILLER_43_1908 ();
 sg13g2_fill_1 FILLER_43_1915 ();
 sg13g2_decap_8 FILLER_43_1921 ();
 sg13g2_decap_4 FILLER_43_1928 ();
 sg13g2_fill_1 FILLER_43_1936 ();
 sg13g2_fill_2 FILLER_43_1942 ();
 sg13g2_fill_1 FILLER_43_1944 ();
 sg13g2_fill_2 FILLER_43_1967 ();
 sg13g2_fill_1 FILLER_43_1969 ();
 sg13g2_fill_2 FILLER_43_2009 ();
 sg13g2_fill_1 FILLER_43_2011 ();
 sg13g2_fill_2 FILLER_43_2021 ();
 sg13g2_fill_1 FILLER_43_2023 ();
 sg13g2_decap_4 FILLER_43_2033 ();
 sg13g2_decap_8 FILLER_43_2041 ();
 sg13g2_decap_4 FILLER_43_2079 ();
 sg13g2_fill_1 FILLER_43_2122 ();
 sg13g2_fill_2 FILLER_43_2142 ();
 sg13g2_fill_1 FILLER_43_2144 ();
 sg13g2_fill_2 FILLER_43_2167 ();
 sg13g2_fill_1 FILLER_43_2174 ();
 sg13g2_decap_4 FILLER_43_2230 ();
 sg13g2_fill_2 FILLER_43_2252 ();
 sg13g2_fill_1 FILLER_43_2254 ();
 sg13g2_decap_4 FILLER_43_2316 ();
 sg13g2_fill_1 FILLER_43_2324 ();
 sg13g2_decap_8 FILLER_43_2351 ();
 sg13g2_decap_8 FILLER_43_2358 ();
 sg13g2_decap_8 FILLER_43_2365 ();
 sg13g2_decap_8 FILLER_43_2372 ();
 sg13g2_decap_8 FILLER_43_2379 ();
 sg13g2_decap_8 FILLER_43_2386 ();
 sg13g2_decap_8 FILLER_43_2393 ();
 sg13g2_decap_8 FILLER_43_2400 ();
 sg13g2_decap_8 FILLER_43_2407 ();
 sg13g2_decap_8 FILLER_43_2414 ();
 sg13g2_decap_8 FILLER_43_2421 ();
 sg13g2_decap_8 FILLER_43_2428 ();
 sg13g2_decap_8 FILLER_43_2435 ();
 sg13g2_decap_8 FILLER_43_2442 ();
 sg13g2_decap_8 FILLER_43_2449 ();
 sg13g2_decap_8 FILLER_43_2456 ();
 sg13g2_decap_8 FILLER_43_2463 ();
 sg13g2_decap_8 FILLER_43_2470 ();
 sg13g2_decap_8 FILLER_43_2477 ();
 sg13g2_decap_8 FILLER_43_2484 ();
 sg13g2_decap_8 FILLER_43_2491 ();
 sg13g2_decap_8 FILLER_43_2498 ();
 sg13g2_decap_8 FILLER_43_2505 ();
 sg13g2_decap_8 FILLER_43_2512 ();
 sg13g2_decap_8 FILLER_43_2519 ();
 sg13g2_decap_8 FILLER_43_2526 ();
 sg13g2_decap_8 FILLER_43_2533 ();
 sg13g2_decap_8 FILLER_43_2540 ();
 sg13g2_decap_8 FILLER_43_2547 ();
 sg13g2_decap_8 FILLER_43_2554 ();
 sg13g2_decap_8 FILLER_43_2561 ();
 sg13g2_decap_8 FILLER_43_2568 ();
 sg13g2_decap_8 FILLER_43_2575 ();
 sg13g2_decap_8 FILLER_43_2582 ();
 sg13g2_decap_8 FILLER_43_2589 ();
 sg13g2_decap_8 FILLER_43_2596 ();
 sg13g2_decap_8 FILLER_43_2603 ();
 sg13g2_decap_8 FILLER_43_2610 ();
 sg13g2_decap_8 FILLER_43_2617 ();
 sg13g2_decap_8 FILLER_43_2624 ();
 sg13g2_decap_8 FILLER_43_2631 ();
 sg13g2_decap_8 FILLER_43_2638 ();
 sg13g2_decap_8 FILLER_43_2645 ();
 sg13g2_decap_8 FILLER_43_2652 ();
 sg13g2_decap_8 FILLER_43_2659 ();
 sg13g2_decap_8 FILLER_43_2666 ();
 sg13g2_fill_1 FILLER_43_2673 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_decap_8 FILLER_44_196 ();
 sg13g2_decap_8 FILLER_44_203 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_decap_8 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_224 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_decap_8 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_259 ();
 sg13g2_decap_8 FILLER_44_266 ();
 sg13g2_decap_8 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_280 ();
 sg13g2_decap_8 FILLER_44_287 ();
 sg13g2_decap_8 FILLER_44_294 ();
 sg13g2_decap_8 FILLER_44_301 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_315 ();
 sg13g2_decap_8 FILLER_44_322 ();
 sg13g2_decap_8 FILLER_44_329 ();
 sg13g2_decap_8 FILLER_44_336 ();
 sg13g2_decap_8 FILLER_44_343 ();
 sg13g2_decap_8 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_decap_8 FILLER_44_406 ();
 sg13g2_decap_8 FILLER_44_413 ();
 sg13g2_decap_8 FILLER_44_420 ();
 sg13g2_decap_8 FILLER_44_427 ();
 sg13g2_decap_8 FILLER_44_434 ();
 sg13g2_decap_8 FILLER_44_441 ();
 sg13g2_decap_8 FILLER_44_448 ();
 sg13g2_decap_8 FILLER_44_455 ();
 sg13g2_decap_8 FILLER_44_462 ();
 sg13g2_decap_8 FILLER_44_469 ();
 sg13g2_decap_8 FILLER_44_476 ();
 sg13g2_fill_2 FILLER_44_483 ();
 sg13g2_fill_1 FILLER_44_524 ();
 sg13g2_fill_2 FILLER_44_560 ();
 sg13g2_fill_1 FILLER_44_562 ();
 sg13g2_decap_4 FILLER_44_577 ();
 sg13g2_fill_1 FILLER_44_581 ();
 sg13g2_fill_2 FILLER_44_586 ();
 sg13g2_fill_1 FILLER_44_588 ();
 sg13g2_decap_8 FILLER_44_607 ();
 sg13g2_fill_2 FILLER_44_614 ();
 sg13g2_decap_8 FILLER_44_645 ();
 sg13g2_decap_4 FILLER_44_652 ();
 sg13g2_fill_1 FILLER_44_656 ();
 sg13g2_fill_2 FILLER_44_728 ();
 sg13g2_fill_1 FILLER_44_730 ();
 sg13g2_fill_2 FILLER_44_757 ();
 sg13g2_fill_1 FILLER_44_759 ();
 sg13g2_fill_2 FILLER_44_799 ();
 sg13g2_fill_1 FILLER_44_801 ();
 sg13g2_decap_4 FILLER_44_815 ();
 sg13g2_fill_1 FILLER_44_819 ();
 sg13g2_fill_1 FILLER_44_876 ();
 sg13g2_fill_1 FILLER_44_899 ();
 sg13g2_fill_1 FILLER_44_909 ();
 sg13g2_decap_4 FILLER_44_914 ();
 sg13g2_decap_4 FILLER_44_922 ();
 sg13g2_fill_2 FILLER_44_926 ();
 sg13g2_decap_4 FILLER_44_1005 ();
 sg13g2_fill_1 FILLER_44_1017 ();
 sg13g2_fill_2 FILLER_44_1022 ();
 sg13g2_decap_4 FILLER_44_1041 ();
 sg13g2_fill_2 FILLER_44_1045 ();
 sg13g2_fill_2 FILLER_44_1097 ();
 sg13g2_fill_1 FILLER_44_1112 ();
 sg13g2_decap_4 FILLER_44_1118 ();
 sg13g2_fill_2 FILLER_44_1158 ();
 sg13g2_fill_2 FILLER_44_1174 ();
 sg13g2_fill_2 FILLER_44_1210 ();
 sg13g2_fill_1 FILLER_44_1212 ();
 sg13g2_fill_2 FILLER_44_1244 ();
 sg13g2_fill_2 FILLER_44_1251 ();
 sg13g2_fill_1 FILLER_44_1253 ();
 sg13g2_fill_2 FILLER_44_1268 ();
 sg13g2_fill_1 FILLER_44_1270 ();
 sg13g2_fill_2 FILLER_44_1280 ();
 sg13g2_fill_2 FILLER_44_1287 ();
 sg13g2_fill_1 FILLER_44_1297 ();
 sg13g2_fill_1 FILLER_44_1312 ();
 sg13g2_fill_2 FILLER_44_1340 ();
 sg13g2_fill_1 FILLER_44_1342 ();
 sg13g2_fill_2 FILLER_44_1367 ();
 sg13g2_fill_1 FILLER_44_1369 ();
 sg13g2_fill_1 FILLER_44_1405 ();
 sg13g2_fill_2 FILLER_44_1446 ();
 sg13g2_fill_1 FILLER_44_1448 ();
 sg13g2_fill_1 FILLER_44_1535 ();
 sg13g2_fill_1 FILLER_44_1593 ();
 sg13g2_decap_8 FILLER_44_1634 ();
 sg13g2_fill_2 FILLER_44_1641 ();
 sg13g2_decap_8 FILLER_44_1647 ();
 sg13g2_fill_2 FILLER_44_1668 ();
 sg13g2_fill_1 FILLER_44_1728 ();
 sg13g2_fill_1 FILLER_44_1755 ();
 sg13g2_fill_2 FILLER_44_1765 ();
 sg13g2_fill_1 FILLER_44_1767 ();
 sg13g2_fill_2 FILLER_44_1812 ();
 sg13g2_fill_2 FILLER_44_1823 ();
 sg13g2_fill_1 FILLER_44_1825 ();
 sg13g2_fill_2 FILLER_44_1847 ();
 sg13g2_decap_8 FILLER_44_1875 ();
 sg13g2_fill_2 FILLER_44_1882 ();
 sg13g2_fill_2 FILLER_44_1992 ();
 sg13g2_fill_1 FILLER_44_1994 ();
 sg13g2_fill_1 FILLER_44_2035 ();
 sg13g2_decap_4 FILLER_44_2044 ();
 sg13g2_fill_1 FILLER_44_2048 ();
 sg13g2_decap_8 FILLER_44_2075 ();
 sg13g2_fill_1 FILLER_44_2082 ();
 sg13g2_fill_2 FILLER_44_2087 ();
 sg13g2_fill_1 FILLER_44_2089 ();
 sg13g2_fill_2 FILLER_44_2108 ();
 sg13g2_fill_2 FILLER_44_2114 ();
 sg13g2_fill_1 FILLER_44_2116 ();
 sg13g2_fill_2 FILLER_44_2152 ();
 sg13g2_fill_2 FILLER_44_2193 ();
 sg13g2_fill_2 FILLER_44_2204 ();
 sg13g2_decap_4 FILLER_44_2211 ();
 sg13g2_fill_2 FILLER_44_2215 ();
 sg13g2_fill_2 FILLER_44_2252 ();
 sg13g2_fill_1 FILLER_44_2254 ();
 sg13g2_fill_1 FILLER_44_2260 ();
 sg13g2_fill_2 FILLER_44_2270 ();
 sg13g2_fill_1 FILLER_44_2272 ();
 sg13g2_fill_1 FILLER_44_2282 ();
 sg13g2_fill_1 FILLER_44_2312 ();
 sg13g2_decap_8 FILLER_44_2349 ();
 sg13g2_decap_8 FILLER_44_2356 ();
 sg13g2_decap_8 FILLER_44_2363 ();
 sg13g2_decap_8 FILLER_44_2370 ();
 sg13g2_decap_8 FILLER_44_2377 ();
 sg13g2_decap_8 FILLER_44_2384 ();
 sg13g2_decap_8 FILLER_44_2391 ();
 sg13g2_decap_8 FILLER_44_2398 ();
 sg13g2_decap_8 FILLER_44_2405 ();
 sg13g2_decap_8 FILLER_44_2412 ();
 sg13g2_decap_8 FILLER_44_2419 ();
 sg13g2_decap_8 FILLER_44_2426 ();
 sg13g2_decap_8 FILLER_44_2433 ();
 sg13g2_decap_8 FILLER_44_2440 ();
 sg13g2_decap_8 FILLER_44_2447 ();
 sg13g2_decap_8 FILLER_44_2454 ();
 sg13g2_decap_8 FILLER_44_2461 ();
 sg13g2_decap_8 FILLER_44_2468 ();
 sg13g2_decap_8 FILLER_44_2475 ();
 sg13g2_decap_8 FILLER_44_2482 ();
 sg13g2_decap_8 FILLER_44_2489 ();
 sg13g2_decap_8 FILLER_44_2496 ();
 sg13g2_decap_8 FILLER_44_2503 ();
 sg13g2_decap_8 FILLER_44_2510 ();
 sg13g2_decap_8 FILLER_44_2517 ();
 sg13g2_decap_8 FILLER_44_2524 ();
 sg13g2_decap_8 FILLER_44_2531 ();
 sg13g2_decap_8 FILLER_44_2538 ();
 sg13g2_decap_8 FILLER_44_2545 ();
 sg13g2_decap_8 FILLER_44_2552 ();
 sg13g2_decap_8 FILLER_44_2559 ();
 sg13g2_decap_8 FILLER_44_2566 ();
 sg13g2_decap_8 FILLER_44_2573 ();
 sg13g2_decap_8 FILLER_44_2580 ();
 sg13g2_decap_8 FILLER_44_2587 ();
 sg13g2_decap_8 FILLER_44_2594 ();
 sg13g2_decap_8 FILLER_44_2601 ();
 sg13g2_decap_8 FILLER_44_2608 ();
 sg13g2_decap_8 FILLER_44_2615 ();
 sg13g2_decap_8 FILLER_44_2622 ();
 sg13g2_decap_8 FILLER_44_2629 ();
 sg13g2_decap_8 FILLER_44_2636 ();
 sg13g2_decap_8 FILLER_44_2643 ();
 sg13g2_decap_8 FILLER_44_2650 ();
 sg13g2_decap_8 FILLER_44_2657 ();
 sg13g2_decap_8 FILLER_44_2664 ();
 sg13g2_fill_2 FILLER_44_2671 ();
 sg13g2_fill_1 FILLER_44_2673 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_decap_8 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_245 ();
 sg13g2_decap_8 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_329 ();
 sg13g2_decap_8 FILLER_45_336 ();
 sg13g2_decap_8 FILLER_45_343 ();
 sg13g2_decap_8 FILLER_45_350 ();
 sg13g2_decap_8 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_decap_8 FILLER_45_413 ();
 sg13g2_decap_8 FILLER_45_420 ();
 sg13g2_decap_8 FILLER_45_427 ();
 sg13g2_decap_8 FILLER_45_434 ();
 sg13g2_decap_8 FILLER_45_441 ();
 sg13g2_decap_8 FILLER_45_448 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_decap_8 FILLER_45_462 ();
 sg13g2_decap_8 FILLER_45_469 ();
 sg13g2_decap_8 FILLER_45_476 ();
 sg13g2_decap_8 FILLER_45_483 ();
 sg13g2_fill_1 FILLER_45_490 ();
 sg13g2_fill_1 FILLER_45_500 ();
 sg13g2_decap_8 FILLER_45_509 ();
 sg13g2_fill_2 FILLER_45_525 ();
 sg13g2_fill_1 FILLER_45_527 ();
 sg13g2_decap_4 FILLER_45_642 ();
 sg13g2_fill_1 FILLER_45_658 ();
 sg13g2_fill_2 FILLER_45_721 ();
 sg13g2_fill_2 FILLER_45_738 ();
 sg13g2_fill_1 FILLER_45_740 ();
 sg13g2_fill_2 FILLER_45_759 ();
 sg13g2_fill_1 FILLER_45_804 ();
 sg13g2_fill_2 FILLER_45_824 ();
 sg13g2_fill_1 FILLER_45_826 ();
 sg13g2_fill_2 FILLER_45_836 ();
 sg13g2_fill_1 FILLER_45_838 ();
 sg13g2_fill_2 FILLER_45_867 ();
 sg13g2_fill_1 FILLER_45_869 ();
 sg13g2_fill_2 FILLER_45_884 ();
 sg13g2_fill_1 FILLER_45_886 ();
 sg13g2_fill_1 FILLER_45_893 ();
 sg13g2_fill_2 FILLER_45_904 ();
 sg13g2_fill_1 FILLER_45_906 ();
 sg13g2_decap_8 FILLER_45_937 ();
 sg13g2_fill_1 FILLER_45_944 ();
 sg13g2_decap_8 FILLER_45_987 ();
 sg13g2_decap_8 FILLER_45_994 ();
 sg13g2_fill_1 FILLER_45_1001 ();
 sg13g2_decap_4 FILLER_45_1037 ();
 sg13g2_fill_2 FILLER_45_1052 ();
 sg13g2_fill_2 FILLER_45_1098 ();
 sg13g2_fill_1 FILLER_45_1108 ();
 sg13g2_fill_2 FILLER_45_1135 ();
 sg13g2_fill_2 FILLER_45_1156 ();
 sg13g2_fill_1 FILLER_45_1163 ();
 sg13g2_fill_1 FILLER_45_1195 ();
 sg13g2_fill_2 FILLER_45_1276 ();
 sg13g2_fill_1 FILLER_45_1278 ();
 sg13g2_fill_2 FILLER_45_1306 ();
 sg13g2_fill_1 FILLER_45_1308 ();
 sg13g2_fill_2 FILLER_45_1326 ();
 sg13g2_fill_2 FILLER_45_1354 ();
 sg13g2_decap_8 FILLER_45_1401 ();
 sg13g2_fill_2 FILLER_45_1408 ();
 sg13g2_fill_1 FILLER_45_1410 ();
 sg13g2_fill_2 FILLER_45_1427 ();
 sg13g2_fill_2 FILLER_45_1484 ();
 sg13g2_fill_1 FILLER_45_1486 ();
 sg13g2_fill_1 FILLER_45_1519 ();
 sg13g2_fill_2 FILLER_45_1578 ();
 sg13g2_fill_1 FILLER_45_1580 ();
 sg13g2_decap_4 FILLER_45_1620 ();
 sg13g2_decap_4 FILLER_45_1654 ();
 sg13g2_decap_4 FILLER_45_1663 ();
 sg13g2_fill_2 FILLER_45_1692 ();
 sg13g2_fill_2 FILLER_45_1749 ();
 sg13g2_fill_1 FILLER_45_1790 ();
 sg13g2_fill_2 FILLER_45_1810 ();
 sg13g2_fill_1 FILLER_45_1812 ();
 sg13g2_fill_2 FILLER_45_1818 ();
 sg13g2_decap_4 FILLER_45_1824 ();
 sg13g2_fill_2 FILLER_45_1846 ();
 sg13g2_fill_2 FILLER_45_1862 ();
 sg13g2_fill_1 FILLER_45_1864 ();
 sg13g2_decap_4 FILLER_45_1878 ();
 sg13g2_fill_2 FILLER_45_1882 ();
 sg13g2_decap_8 FILLER_45_1897 ();
 sg13g2_fill_2 FILLER_45_1904 ();
 sg13g2_fill_1 FILLER_45_1906 ();
 sg13g2_decap_8 FILLER_45_1918 ();
 sg13g2_fill_1 FILLER_45_1925 ();
 sg13g2_decap_8 FILLER_45_1931 ();
 sg13g2_fill_2 FILLER_45_1938 ();
 sg13g2_fill_2 FILLER_45_1961 ();
 sg13g2_fill_1 FILLER_45_1963 ();
 sg13g2_fill_1 FILLER_45_2015 ();
 sg13g2_fill_1 FILLER_45_2045 ();
 sg13g2_fill_2 FILLER_45_2051 ();
 sg13g2_fill_1 FILLER_45_2053 ();
 sg13g2_fill_1 FILLER_45_2135 ();
 sg13g2_fill_1 FILLER_45_2145 ();
 sg13g2_fill_1 FILLER_45_2168 ();
 sg13g2_fill_2 FILLER_45_2232 ();
 sg13g2_fill_2 FILLER_45_2239 ();
 sg13g2_fill_2 FILLER_45_2250 ();
 sg13g2_fill_1 FILLER_45_2252 ();
 sg13g2_fill_2 FILLER_45_2296 ();
 sg13g2_decap_8 FILLER_45_2350 ();
 sg13g2_decap_8 FILLER_45_2357 ();
 sg13g2_decap_8 FILLER_45_2364 ();
 sg13g2_decap_8 FILLER_45_2371 ();
 sg13g2_decap_8 FILLER_45_2378 ();
 sg13g2_decap_8 FILLER_45_2385 ();
 sg13g2_decap_8 FILLER_45_2392 ();
 sg13g2_decap_8 FILLER_45_2399 ();
 sg13g2_decap_8 FILLER_45_2406 ();
 sg13g2_decap_8 FILLER_45_2413 ();
 sg13g2_decap_8 FILLER_45_2420 ();
 sg13g2_decap_8 FILLER_45_2427 ();
 sg13g2_decap_8 FILLER_45_2434 ();
 sg13g2_decap_8 FILLER_45_2441 ();
 sg13g2_decap_8 FILLER_45_2448 ();
 sg13g2_decap_8 FILLER_45_2455 ();
 sg13g2_decap_8 FILLER_45_2462 ();
 sg13g2_decap_8 FILLER_45_2469 ();
 sg13g2_decap_8 FILLER_45_2476 ();
 sg13g2_decap_8 FILLER_45_2483 ();
 sg13g2_decap_8 FILLER_45_2490 ();
 sg13g2_decap_8 FILLER_45_2497 ();
 sg13g2_decap_8 FILLER_45_2504 ();
 sg13g2_decap_8 FILLER_45_2511 ();
 sg13g2_decap_8 FILLER_45_2518 ();
 sg13g2_decap_8 FILLER_45_2525 ();
 sg13g2_decap_8 FILLER_45_2532 ();
 sg13g2_decap_8 FILLER_45_2539 ();
 sg13g2_decap_8 FILLER_45_2546 ();
 sg13g2_decap_8 FILLER_45_2553 ();
 sg13g2_decap_8 FILLER_45_2560 ();
 sg13g2_decap_8 FILLER_45_2567 ();
 sg13g2_decap_8 FILLER_45_2574 ();
 sg13g2_decap_8 FILLER_45_2581 ();
 sg13g2_decap_8 FILLER_45_2588 ();
 sg13g2_decap_8 FILLER_45_2595 ();
 sg13g2_decap_8 FILLER_45_2602 ();
 sg13g2_decap_8 FILLER_45_2609 ();
 sg13g2_decap_8 FILLER_45_2616 ();
 sg13g2_decap_8 FILLER_45_2623 ();
 sg13g2_decap_8 FILLER_45_2630 ();
 sg13g2_decap_8 FILLER_45_2637 ();
 sg13g2_decap_8 FILLER_45_2644 ();
 sg13g2_decap_8 FILLER_45_2651 ();
 sg13g2_decap_8 FILLER_45_2658 ();
 sg13g2_decap_8 FILLER_45_2665 ();
 sg13g2_fill_2 FILLER_45_2672 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_357 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_441 ();
 sg13g2_decap_8 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_455 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_497 ();
 sg13g2_fill_2 FILLER_46_504 ();
 sg13g2_fill_2 FILLER_46_541 ();
 sg13g2_fill_2 FILLER_46_552 ();
 sg13g2_fill_1 FILLER_46_554 ();
 sg13g2_fill_2 FILLER_46_581 ();
 sg13g2_fill_1 FILLER_46_583 ();
 sg13g2_fill_2 FILLER_46_605 ();
 sg13g2_fill_1 FILLER_46_607 ();
 sg13g2_fill_2 FILLER_46_621 ();
 sg13g2_fill_2 FILLER_46_628 ();
 sg13g2_fill_1 FILLER_46_630 ();
 sg13g2_fill_1 FILLER_46_647 ();
 sg13g2_fill_2 FILLER_46_680 ();
 sg13g2_fill_1 FILLER_46_760 ();
 sg13g2_fill_2 FILLER_46_771 ();
 sg13g2_fill_1 FILLER_46_773 ();
 sg13g2_fill_2 FILLER_46_798 ();
 sg13g2_fill_2 FILLER_46_842 ();
 sg13g2_fill_2 FILLER_46_913 ();
 sg13g2_fill_2 FILLER_46_928 ();
 sg13g2_fill_2 FILLER_46_947 ();
 sg13g2_decap_8 FILLER_46_953 ();
 sg13g2_fill_1 FILLER_46_972 ();
 sg13g2_fill_2 FILLER_46_990 ();
 sg13g2_fill_2 FILLER_46_1005 ();
 sg13g2_fill_1 FILLER_46_1007 ();
 sg13g2_fill_2 FILLER_46_1013 ();
 sg13g2_fill_1 FILLER_46_1015 ();
 sg13g2_fill_1 FILLER_46_1054 ();
 sg13g2_fill_2 FILLER_46_1116 ();
 sg13g2_fill_1 FILLER_46_1118 ();
 sg13g2_fill_2 FILLER_46_1167 ();
 sg13g2_fill_1 FILLER_46_1173 ();
 sg13g2_decap_8 FILLER_46_1196 ();
 sg13g2_fill_2 FILLER_46_1203 ();
 sg13g2_fill_2 FILLER_46_1218 ();
 sg13g2_fill_1 FILLER_46_1220 ();
 sg13g2_fill_2 FILLER_46_1230 ();
 sg13g2_fill_1 FILLER_46_1232 ();
 sg13g2_fill_2 FILLER_46_1259 ();
 sg13g2_fill_1 FILLER_46_1261 ();
 sg13g2_fill_1 FILLER_46_1293 ();
 sg13g2_decap_8 FILLER_46_1330 ();
 sg13g2_fill_2 FILLER_46_1337 ();
 sg13g2_fill_2 FILLER_46_1347 ();
 sg13g2_fill_2 FILLER_46_1378 ();
 sg13g2_fill_2 FILLER_46_1397 ();
 sg13g2_fill_1 FILLER_46_1452 ();
 sg13g2_decap_8 FILLER_46_1458 ();
 sg13g2_fill_2 FILLER_46_1465 ();
 sg13g2_fill_2 FILLER_46_1521 ();
 sg13g2_fill_1 FILLER_46_1523 ();
 sg13g2_fill_2 FILLER_46_1529 ();
 sg13g2_fill_1 FILLER_46_1531 ();
 sg13g2_fill_2 FILLER_46_1536 ();
 sg13g2_fill_1 FILLER_46_1538 ();
 sg13g2_fill_2 FILLER_46_1545 ();
 sg13g2_fill_1 FILLER_46_1547 ();
 sg13g2_fill_1 FILLER_46_1580 ();
 sg13g2_fill_1 FILLER_46_1592 ();
 sg13g2_fill_2 FILLER_46_1633 ();
 sg13g2_fill_1 FILLER_46_1635 ();
 sg13g2_decap_8 FILLER_46_1660 ();
 sg13g2_fill_1 FILLER_46_1676 ();
 sg13g2_decap_8 FILLER_46_1686 ();
 sg13g2_fill_1 FILLER_46_1693 ();
 sg13g2_fill_2 FILLER_46_1713 ();
 sg13g2_fill_1 FILLER_46_1715 ();
 sg13g2_decap_4 FILLER_46_1729 ();
 sg13g2_fill_2 FILLER_46_1733 ();
 sg13g2_fill_2 FILLER_46_1748 ();
 sg13g2_fill_1 FILLER_46_1768 ();
 sg13g2_fill_2 FILLER_46_1788 ();
 sg13g2_fill_1 FILLER_46_1790 ();
 sg13g2_fill_1 FILLER_46_1821 ();
 sg13g2_fill_1 FILLER_46_1857 ();
 sg13g2_decap_4 FILLER_46_1969 ();
 sg13g2_fill_2 FILLER_46_1986 ();
 sg13g2_fill_1 FILLER_46_1988 ();
 sg13g2_fill_2 FILLER_46_1998 ();
 sg13g2_decap_4 FILLER_46_2017 ();
 sg13g2_fill_2 FILLER_46_2021 ();
 sg13g2_fill_2 FILLER_46_2039 ();
 sg13g2_fill_1 FILLER_46_2041 ();
 sg13g2_fill_1 FILLER_46_2077 ();
 sg13g2_decap_8 FILLER_46_2096 ();
 sg13g2_fill_1 FILLER_46_2103 ();
 sg13g2_fill_2 FILLER_46_2169 ();
 sg13g2_fill_1 FILLER_46_2178 ();
 sg13g2_fill_2 FILLER_46_2205 ();
 sg13g2_fill_1 FILLER_46_2207 ();
 sg13g2_decap_4 FILLER_46_2212 ();
 sg13g2_fill_1 FILLER_46_2220 ();
 sg13g2_fill_2 FILLER_46_2268 ();
 sg13g2_fill_1 FILLER_46_2270 ();
 sg13g2_fill_2 FILLER_46_2280 ();
 sg13g2_fill_1 FILLER_46_2286 ();
 sg13g2_decap_4 FILLER_46_2291 ();
 sg13g2_fill_2 FILLER_46_2304 ();
 sg13g2_fill_1 FILLER_46_2306 ();
 sg13g2_fill_1 FILLER_46_2321 ();
 sg13g2_fill_2 FILLER_46_2331 ();
 sg13g2_fill_1 FILLER_46_2333 ();
 sg13g2_decap_8 FILLER_46_2347 ();
 sg13g2_decap_8 FILLER_46_2354 ();
 sg13g2_decap_8 FILLER_46_2361 ();
 sg13g2_decap_8 FILLER_46_2368 ();
 sg13g2_decap_8 FILLER_46_2375 ();
 sg13g2_decap_8 FILLER_46_2382 ();
 sg13g2_decap_8 FILLER_46_2389 ();
 sg13g2_decap_8 FILLER_46_2396 ();
 sg13g2_decap_8 FILLER_46_2403 ();
 sg13g2_decap_8 FILLER_46_2410 ();
 sg13g2_decap_8 FILLER_46_2417 ();
 sg13g2_decap_8 FILLER_46_2424 ();
 sg13g2_decap_8 FILLER_46_2431 ();
 sg13g2_decap_8 FILLER_46_2438 ();
 sg13g2_decap_8 FILLER_46_2445 ();
 sg13g2_decap_8 FILLER_46_2452 ();
 sg13g2_decap_8 FILLER_46_2459 ();
 sg13g2_decap_8 FILLER_46_2466 ();
 sg13g2_decap_8 FILLER_46_2473 ();
 sg13g2_decap_8 FILLER_46_2480 ();
 sg13g2_decap_8 FILLER_46_2487 ();
 sg13g2_decap_8 FILLER_46_2494 ();
 sg13g2_decap_8 FILLER_46_2501 ();
 sg13g2_decap_8 FILLER_46_2508 ();
 sg13g2_decap_8 FILLER_46_2515 ();
 sg13g2_decap_8 FILLER_46_2522 ();
 sg13g2_decap_8 FILLER_46_2529 ();
 sg13g2_decap_8 FILLER_46_2536 ();
 sg13g2_decap_8 FILLER_46_2543 ();
 sg13g2_decap_8 FILLER_46_2550 ();
 sg13g2_decap_8 FILLER_46_2557 ();
 sg13g2_decap_8 FILLER_46_2564 ();
 sg13g2_decap_8 FILLER_46_2571 ();
 sg13g2_decap_8 FILLER_46_2578 ();
 sg13g2_decap_8 FILLER_46_2585 ();
 sg13g2_decap_8 FILLER_46_2592 ();
 sg13g2_decap_8 FILLER_46_2599 ();
 sg13g2_decap_8 FILLER_46_2606 ();
 sg13g2_decap_8 FILLER_46_2613 ();
 sg13g2_decap_8 FILLER_46_2620 ();
 sg13g2_decap_8 FILLER_46_2627 ();
 sg13g2_decap_8 FILLER_46_2634 ();
 sg13g2_decap_8 FILLER_46_2641 ();
 sg13g2_decap_8 FILLER_46_2648 ();
 sg13g2_decap_8 FILLER_46_2655 ();
 sg13g2_decap_8 FILLER_46_2662 ();
 sg13g2_decap_4 FILLER_46_2669 ();
 sg13g2_fill_1 FILLER_46_2673 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_fill_2 FILLER_47_462 ();
 sg13g2_fill_2 FILLER_47_482 ();
 sg13g2_fill_1 FILLER_47_484 ();
 sg13g2_fill_1 FILLER_47_516 ();
 sg13g2_decap_8 FILLER_47_521 ();
 sg13g2_fill_1 FILLER_47_562 ();
 sg13g2_fill_1 FILLER_47_581 ();
 sg13g2_decap_4 FILLER_47_626 ();
 sg13g2_fill_2 FILLER_47_630 ();
 sg13g2_decap_8 FILLER_47_640 ();
 sg13g2_fill_2 FILLER_47_647 ();
 sg13g2_decap_4 FILLER_47_652 ();
 sg13g2_fill_1 FILLER_47_682 ();
 sg13g2_fill_1 FILLER_47_692 ();
 sg13g2_fill_1 FILLER_47_709 ();
 sg13g2_fill_1 FILLER_47_756 ();
 sg13g2_fill_1 FILLER_47_791 ();
 sg13g2_fill_2 FILLER_47_800 ();
 sg13g2_fill_2 FILLER_47_824 ();
 sg13g2_fill_1 FILLER_47_826 ();
 sg13g2_fill_1 FILLER_47_831 ();
 sg13g2_fill_1 FILLER_47_840 ();
 sg13g2_fill_2 FILLER_47_853 ();
 sg13g2_decap_4 FILLER_47_869 ();
 sg13g2_fill_2 FILLER_47_878 ();
 sg13g2_fill_1 FILLER_47_880 ();
 sg13g2_fill_2 FILLER_47_902 ();
 sg13g2_fill_1 FILLER_47_904 ();
 sg13g2_fill_1 FILLER_47_924 ();
 sg13g2_decap_4 FILLER_47_964 ();
 sg13g2_fill_2 FILLER_47_968 ();
 sg13g2_fill_2 FILLER_47_1047 ();
 sg13g2_fill_1 FILLER_47_1049 ();
 sg13g2_fill_2 FILLER_47_1077 ();
 sg13g2_fill_1 FILLER_47_1083 ();
 sg13g2_decap_4 FILLER_47_1093 ();
 sg13g2_fill_2 FILLER_47_1110 ();
 sg13g2_fill_1 FILLER_47_1119 ();
 sg13g2_fill_2 FILLER_47_1130 ();
 sg13g2_fill_1 FILLER_47_1132 ();
 sg13g2_fill_2 FILLER_47_1159 ();
 sg13g2_fill_2 FILLER_47_1191 ();
 sg13g2_decap_4 FILLER_47_1201 ();
 sg13g2_fill_2 FILLER_47_1205 ();
 sg13g2_fill_1 FILLER_47_1232 ();
 sg13g2_decap_4 FILLER_47_1238 ();
 sg13g2_fill_2 FILLER_47_1242 ();
 sg13g2_fill_2 FILLER_47_1252 ();
 sg13g2_fill_1 FILLER_47_1254 ();
 sg13g2_fill_2 FILLER_47_1286 ();
 sg13g2_fill_2 FILLER_47_1297 ();
 sg13g2_fill_1 FILLER_47_1299 ();
 sg13g2_fill_1 FILLER_47_1305 ();
 sg13g2_fill_1 FILLER_47_1311 ();
 sg13g2_fill_2 FILLER_47_1317 ();
 sg13g2_fill_2 FILLER_47_1366 ();
 sg13g2_fill_1 FILLER_47_1368 ();
 sg13g2_decap_4 FILLER_47_1400 ();
 sg13g2_fill_2 FILLER_47_1404 ();
 sg13g2_decap_4 FILLER_47_1411 ();
 sg13g2_fill_1 FILLER_47_1415 ();
 sg13g2_fill_2 FILLER_47_1425 ();
 sg13g2_fill_2 FILLER_47_1475 ();
 sg13g2_fill_1 FILLER_47_1477 ();
 sg13g2_decap_4 FILLER_47_1499 ();
 sg13g2_fill_2 FILLER_47_1503 ();
 sg13g2_decap_8 FILLER_47_1510 ();
 sg13g2_fill_1 FILLER_47_1517 ();
 sg13g2_fill_2 FILLER_47_1548 ();
 sg13g2_fill_2 FILLER_47_1559 ();
 sg13g2_fill_1 FILLER_47_1561 ();
 sg13g2_fill_2 FILLER_47_1571 ();
 sg13g2_fill_2 FILLER_47_1587 ();
 sg13g2_fill_2 FILLER_47_1624 ();
 sg13g2_fill_1 FILLER_47_1631 ();
 sg13g2_fill_2 FILLER_47_1653 ();
 sg13g2_fill_1 FILLER_47_1655 ();
 sg13g2_fill_2 FILLER_47_1661 ();
 sg13g2_decap_8 FILLER_47_1672 ();
 sg13g2_fill_1 FILLER_47_1679 ();
 sg13g2_fill_1 FILLER_47_1694 ();
 sg13g2_fill_2 FILLER_47_1736 ();
 sg13g2_fill_1 FILLER_47_1738 ();
 sg13g2_fill_2 FILLER_47_1756 ();
 sg13g2_fill_1 FILLER_47_1758 ();
 sg13g2_fill_2 FILLER_47_1773 ();
 sg13g2_fill_1 FILLER_47_1775 ();
 sg13g2_fill_2 FILLER_47_1792 ();
 sg13g2_fill_1 FILLER_47_1812 ();
 sg13g2_fill_2 FILLER_47_1840 ();
 sg13g2_fill_1 FILLER_47_1842 ();
 sg13g2_decap_4 FILLER_47_1891 ();
 sg13g2_fill_2 FILLER_47_1895 ();
 sg13g2_fill_2 FILLER_47_1919 ();
 sg13g2_decap_4 FILLER_47_1925 ();
 sg13g2_fill_1 FILLER_47_1933 ();
 sg13g2_fill_2 FILLER_47_1953 ();
 sg13g2_fill_1 FILLER_47_1955 ();
 sg13g2_fill_1 FILLER_47_1982 ();
 sg13g2_fill_1 FILLER_47_2040 ();
 sg13g2_fill_2 FILLER_47_2076 ();
 sg13g2_fill_1 FILLER_47_2078 ();
 sg13g2_fill_2 FILLER_47_2105 ();
 sg13g2_fill_2 FILLER_47_2120 ();
 sg13g2_decap_4 FILLER_47_2143 ();
 sg13g2_fill_2 FILLER_47_2147 ();
 sg13g2_fill_1 FILLER_47_2167 ();
 sg13g2_decap_8 FILLER_47_2189 ();
 sg13g2_decap_4 FILLER_47_2196 ();
 sg13g2_fill_2 FILLER_47_2200 ();
 sg13g2_fill_1 FILLER_47_2210 ();
 sg13g2_decap_8 FILLER_47_2215 ();
 sg13g2_decap_8 FILLER_47_2222 ();
 sg13g2_decap_4 FILLER_47_2229 ();
 sg13g2_fill_1 FILLER_47_2233 ();
 sg13g2_fill_2 FILLER_47_2255 ();
 sg13g2_fill_1 FILLER_47_2257 ();
 sg13g2_fill_2 FILLER_47_2311 ();
 sg13g2_fill_1 FILLER_47_2313 ();
 sg13g2_decap_8 FILLER_47_2340 ();
 sg13g2_decap_8 FILLER_47_2347 ();
 sg13g2_decap_8 FILLER_47_2354 ();
 sg13g2_decap_8 FILLER_47_2361 ();
 sg13g2_decap_8 FILLER_47_2368 ();
 sg13g2_decap_8 FILLER_47_2375 ();
 sg13g2_decap_8 FILLER_47_2382 ();
 sg13g2_decap_8 FILLER_47_2389 ();
 sg13g2_decap_8 FILLER_47_2396 ();
 sg13g2_decap_8 FILLER_47_2403 ();
 sg13g2_decap_8 FILLER_47_2410 ();
 sg13g2_decap_8 FILLER_47_2417 ();
 sg13g2_decap_8 FILLER_47_2424 ();
 sg13g2_decap_8 FILLER_47_2431 ();
 sg13g2_decap_8 FILLER_47_2438 ();
 sg13g2_decap_8 FILLER_47_2445 ();
 sg13g2_decap_8 FILLER_47_2452 ();
 sg13g2_decap_8 FILLER_47_2459 ();
 sg13g2_decap_8 FILLER_47_2466 ();
 sg13g2_decap_8 FILLER_47_2473 ();
 sg13g2_decap_8 FILLER_47_2480 ();
 sg13g2_decap_8 FILLER_47_2487 ();
 sg13g2_decap_8 FILLER_47_2494 ();
 sg13g2_decap_8 FILLER_47_2501 ();
 sg13g2_decap_8 FILLER_47_2508 ();
 sg13g2_decap_8 FILLER_47_2515 ();
 sg13g2_decap_8 FILLER_47_2522 ();
 sg13g2_decap_8 FILLER_47_2529 ();
 sg13g2_decap_8 FILLER_47_2536 ();
 sg13g2_decap_8 FILLER_47_2543 ();
 sg13g2_decap_8 FILLER_47_2550 ();
 sg13g2_decap_8 FILLER_47_2557 ();
 sg13g2_decap_8 FILLER_47_2564 ();
 sg13g2_decap_8 FILLER_47_2571 ();
 sg13g2_decap_8 FILLER_47_2578 ();
 sg13g2_decap_8 FILLER_47_2585 ();
 sg13g2_decap_8 FILLER_47_2592 ();
 sg13g2_decap_8 FILLER_47_2599 ();
 sg13g2_decap_8 FILLER_47_2606 ();
 sg13g2_decap_8 FILLER_47_2613 ();
 sg13g2_decap_8 FILLER_47_2620 ();
 sg13g2_decap_8 FILLER_47_2627 ();
 sg13g2_decap_8 FILLER_47_2634 ();
 sg13g2_decap_8 FILLER_47_2641 ();
 sg13g2_decap_8 FILLER_47_2648 ();
 sg13g2_decap_8 FILLER_47_2655 ();
 sg13g2_decap_8 FILLER_47_2662 ();
 sg13g2_decap_4 FILLER_47_2669 ();
 sg13g2_fill_1 FILLER_47_2673 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_fill_2 FILLER_48_455 ();
 sg13g2_fill_2 FILLER_48_488 ();
 sg13g2_fill_1 FILLER_48_490 ();
 sg13g2_fill_2 FILLER_48_591 ();
 sg13g2_fill_1 FILLER_48_593 ();
 sg13g2_decap_8 FILLER_48_613 ();
 sg13g2_decap_4 FILLER_48_620 ();
 sg13g2_fill_2 FILLER_48_642 ();
 sg13g2_fill_2 FILLER_48_675 ();
 sg13g2_fill_1 FILLER_48_687 ();
 sg13g2_fill_2 FILLER_48_696 ();
 sg13g2_fill_2 FILLER_48_788 ();
 sg13g2_fill_1 FILLER_48_832 ();
 sg13g2_fill_1 FILLER_48_842 ();
 sg13g2_fill_1 FILLER_48_854 ();
 sg13g2_fill_2 FILLER_48_886 ();
 sg13g2_fill_1 FILLER_48_888 ();
 sg13g2_fill_2 FILLER_48_923 ();
 sg13g2_fill_1 FILLER_48_925 ();
 sg13g2_fill_2 FILLER_48_933 ();
 sg13g2_fill_1 FILLER_48_947 ();
 sg13g2_decap_4 FILLER_48_953 ();
 sg13g2_fill_2 FILLER_48_957 ();
 sg13g2_decap_8 FILLER_48_963 ();
 sg13g2_fill_2 FILLER_48_979 ();
 sg13g2_fill_2 FILLER_48_986 ();
 sg13g2_fill_1 FILLER_48_988 ();
 sg13g2_fill_2 FILLER_48_1002 ();
 sg13g2_fill_2 FILLER_48_1088 ();
 sg13g2_fill_1 FILLER_48_1099 ();
 sg13g2_fill_1 FILLER_48_1124 ();
 sg13g2_fill_2 FILLER_48_1152 ();
 sg13g2_fill_2 FILLER_48_1169 ();
 sg13g2_fill_1 FILLER_48_1171 ();
 sg13g2_fill_2 FILLER_48_1198 ();
 sg13g2_fill_1 FILLER_48_1289 ();
 sg13g2_fill_2 FILLER_48_1369 ();
 sg13g2_fill_1 FILLER_48_1371 ();
 sg13g2_fill_2 FILLER_48_1390 ();
 sg13g2_fill_2 FILLER_48_1418 ();
 sg13g2_fill_1 FILLER_48_1420 ();
 sg13g2_fill_2 FILLER_48_1428 ();
 sg13g2_fill_1 FILLER_48_1430 ();
 sg13g2_fill_2 FILLER_48_1454 ();
 sg13g2_decap_4 FILLER_48_1469 ();
 sg13g2_fill_1 FILLER_48_1473 ();
 sg13g2_decap_4 FILLER_48_1486 ();
 sg13g2_fill_1 FILLER_48_1499 ();
 sg13g2_decap_4 FILLER_48_1504 ();
 sg13g2_fill_2 FILLER_48_1508 ();
 sg13g2_fill_2 FILLER_48_1543 ();
 sg13g2_fill_1 FILLER_48_1626 ();
 sg13g2_fill_2 FILLER_48_1636 ();
 sg13g2_decap_8 FILLER_48_1642 ();
 sg13g2_fill_2 FILLER_48_1649 ();
 sg13g2_fill_1 FILLER_48_1651 ();
 sg13g2_fill_1 FILLER_48_1678 ();
 sg13g2_fill_1 FILLER_48_1718 ();
 sg13g2_fill_2 FILLER_48_1754 ();
 sg13g2_fill_1 FILLER_48_1756 ();
 sg13g2_fill_2 FILLER_48_1801 ();
 sg13g2_fill_1 FILLER_48_1817 ();
 sg13g2_fill_2 FILLER_48_1853 ();
 sg13g2_decap_4 FILLER_48_1882 ();
 sg13g2_fill_2 FILLER_48_1890 ();
 sg13g2_fill_1 FILLER_48_1892 ();
 sg13g2_fill_2 FILLER_48_1920 ();
 sg13g2_fill_1 FILLER_48_1922 ();
 sg13g2_fill_2 FILLER_48_1936 ();
 sg13g2_fill_2 FILLER_48_1943 ();
 sg13g2_fill_1 FILLER_48_1949 ();
 sg13g2_fill_1 FILLER_48_1968 ();
 sg13g2_fill_2 FILLER_48_1984 ();
 sg13g2_fill_2 FILLER_48_1994 ();
 sg13g2_fill_1 FILLER_48_1996 ();
 sg13g2_fill_2 FILLER_48_2010 ();
 sg13g2_fill_1 FILLER_48_2012 ();
 sg13g2_fill_2 FILLER_48_2017 ();
 sg13g2_fill_2 FILLER_48_2047 ();
 sg13g2_fill_1 FILLER_48_2049 ();
 sg13g2_fill_1 FILLER_48_2076 ();
 sg13g2_fill_1 FILLER_48_2099 ();
 sg13g2_decap_4 FILLER_48_2140 ();
 sg13g2_fill_2 FILLER_48_2144 ();
 sg13g2_fill_1 FILLER_48_2151 ();
 sg13g2_fill_2 FILLER_48_2156 ();
 sg13g2_fill_1 FILLER_48_2174 ();
 sg13g2_fill_1 FILLER_48_2250 ();
 sg13g2_fill_1 FILLER_48_2290 ();
 sg13g2_decap_4 FILLER_48_2295 ();
 sg13g2_fill_2 FILLER_48_2303 ();
 sg13g2_fill_2 FILLER_48_2309 ();
 sg13g2_decap_8 FILLER_48_2336 ();
 sg13g2_decap_8 FILLER_48_2343 ();
 sg13g2_decap_8 FILLER_48_2350 ();
 sg13g2_decap_8 FILLER_48_2357 ();
 sg13g2_decap_8 FILLER_48_2364 ();
 sg13g2_decap_8 FILLER_48_2371 ();
 sg13g2_decap_8 FILLER_48_2378 ();
 sg13g2_decap_8 FILLER_48_2385 ();
 sg13g2_decap_8 FILLER_48_2392 ();
 sg13g2_decap_8 FILLER_48_2399 ();
 sg13g2_decap_8 FILLER_48_2406 ();
 sg13g2_decap_8 FILLER_48_2413 ();
 sg13g2_decap_8 FILLER_48_2420 ();
 sg13g2_decap_8 FILLER_48_2427 ();
 sg13g2_decap_8 FILLER_48_2434 ();
 sg13g2_decap_8 FILLER_48_2441 ();
 sg13g2_decap_8 FILLER_48_2448 ();
 sg13g2_decap_8 FILLER_48_2455 ();
 sg13g2_decap_8 FILLER_48_2462 ();
 sg13g2_decap_8 FILLER_48_2469 ();
 sg13g2_decap_8 FILLER_48_2476 ();
 sg13g2_decap_8 FILLER_48_2483 ();
 sg13g2_decap_8 FILLER_48_2490 ();
 sg13g2_decap_8 FILLER_48_2497 ();
 sg13g2_decap_8 FILLER_48_2504 ();
 sg13g2_decap_8 FILLER_48_2511 ();
 sg13g2_decap_8 FILLER_48_2518 ();
 sg13g2_decap_8 FILLER_48_2525 ();
 sg13g2_decap_8 FILLER_48_2532 ();
 sg13g2_decap_8 FILLER_48_2539 ();
 sg13g2_decap_8 FILLER_48_2546 ();
 sg13g2_decap_8 FILLER_48_2553 ();
 sg13g2_decap_8 FILLER_48_2560 ();
 sg13g2_decap_8 FILLER_48_2567 ();
 sg13g2_decap_8 FILLER_48_2574 ();
 sg13g2_decap_8 FILLER_48_2581 ();
 sg13g2_decap_8 FILLER_48_2588 ();
 sg13g2_decap_8 FILLER_48_2595 ();
 sg13g2_decap_8 FILLER_48_2602 ();
 sg13g2_decap_8 FILLER_48_2609 ();
 sg13g2_decap_8 FILLER_48_2616 ();
 sg13g2_decap_8 FILLER_48_2623 ();
 sg13g2_decap_8 FILLER_48_2630 ();
 sg13g2_decap_8 FILLER_48_2637 ();
 sg13g2_decap_8 FILLER_48_2644 ();
 sg13g2_decap_8 FILLER_48_2651 ();
 sg13g2_decap_8 FILLER_48_2658 ();
 sg13g2_decap_8 FILLER_48_2665 ();
 sg13g2_fill_2 FILLER_48_2672 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_8 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_210 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_decap_8 FILLER_49_224 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_decap_8 FILLER_49_238 ();
 sg13g2_decap_8 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_decap_8 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_decap_8 FILLER_49_315 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_decap_8 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_decap_8 FILLER_49_406 ();
 sg13g2_decap_8 FILLER_49_413 ();
 sg13g2_decap_8 FILLER_49_420 ();
 sg13g2_decap_8 FILLER_49_427 ();
 sg13g2_decap_8 FILLER_49_434 ();
 sg13g2_decap_8 FILLER_49_441 ();
 sg13g2_decap_8 FILLER_49_448 ();
 sg13g2_decap_8 FILLER_49_455 ();
 sg13g2_decap_4 FILLER_49_462 ();
 sg13g2_decap_8 FILLER_49_470 ();
 sg13g2_fill_2 FILLER_49_477 ();
 sg13g2_fill_1 FILLER_49_479 ();
 sg13g2_fill_2 FILLER_49_520 ();
 sg13g2_fill_2 FILLER_49_531 ();
 sg13g2_fill_2 FILLER_49_560 ();
 sg13g2_fill_1 FILLER_49_562 ();
 sg13g2_fill_2 FILLER_49_616 ();
 sg13g2_fill_2 FILLER_49_644 ();
 sg13g2_fill_1 FILLER_49_693 ();
 sg13g2_fill_2 FILLER_49_707 ();
 sg13g2_fill_1 FILLER_49_709 ();
 sg13g2_fill_2 FILLER_49_721 ();
 sg13g2_fill_1 FILLER_49_803 ();
 sg13g2_fill_1 FILLER_49_821 ();
 sg13g2_fill_2 FILLER_49_896 ();
 sg13g2_fill_2 FILLER_49_946 ();
 sg13g2_fill_1 FILLER_49_948 ();
 sg13g2_fill_2 FILLER_49_987 ();
 sg13g2_fill_1 FILLER_49_1041 ();
 sg13g2_fill_2 FILLER_49_1051 ();
 sg13g2_fill_2 FILLER_49_1071 ();
 sg13g2_fill_1 FILLER_49_1099 ();
 sg13g2_fill_2 FILLER_49_1105 ();
 sg13g2_fill_1 FILLER_49_1107 ();
 sg13g2_fill_2 FILLER_49_1119 ();
 sg13g2_fill_2 FILLER_49_1130 ();
 sg13g2_fill_1 FILLER_49_1132 ();
 sg13g2_decap_8 FILLER_49_1193 ();
 sg13g2_decap_4 FILLER_49_1200 ();
 sg13g2_fill_2 FILLER_49_1204 ();
 sg13g2_fill_2 FILLER_49_1219 ();
 sg13g2_fill_2 FILLER_49_1243 ();
 sg13g2_fill_2 FILLER_49_1267 ();
 sg13g2_fill_1 FILLER_49_1309 ();
 sg13g2_fill_2 FILLER_49_1359 ();
 sg13g2_fill_1 FILLER_49_1361 ();
 sg13g2_fill_2 FILLER_49_1407 ();
 sg13g2_fill_1 FILLER_49_1409 ();
 sg13g2_fill_2 FILLER_49_1423 ();
 sg13g2_fill_2 FILLER_49_1438 ();
 sg13g2_fill_1 FILLER_49_1440 ();
 sg13g2_fill_2 FILLER_49_1487 ();
 sg13g2_decap_4 FILLER_49_1524 ();
 sg13g2_fill_1 FILLER_49_1528 ();
 sg13g2_fill_1 FILLER_49_1533 ();
 sg13g2_decap_8 FILLER_49_1547 ();
 sg13g2_decap_8 FILLER_49_1554 ();
 sg13g2_fill_2 FILLER_49_1561 ();
 sg13g2_fill_1 FILLER_49_1563 ();
 sg13g2_decap_8 FILLER_49_1574 ();
 sg13g2_fill_2 FILLER_49_1581 ();
 sg13g2_fill_1 FILLER_49_1595 ();
 sg13g2_decap_4 FILLER_49_1613 ();
 sg13g2_fill_1 FILLER_49_1627 ();
 sg13g2_fill_2 FILLER_49_1668 ();
 sg13g2_fill_1 FILLER_49_1670 ();
 sg13g2_fill_1 FILLER_49_1692 ();
 sg13g2_decap_8 FILLER_49_1703 ();
 sg13g2_fill_1 FILLER_49_1738 ();
 sg13g2_fill_2 FILLER_49_1771 ();
 sg13g2_fill_1 FILLER_49_1773 ();
 sg13g2_fill_2 FILLER_49_1779 ();
 sg13g2_fill_1 FILLER_49_1781 ();
 sg13g2_decap_8 FILLER_49_1822 ();
 sg13g2_fill_2 FILLER_49_1829 ();
 sg13g2_fill_1 FILLER_49_1831 ();
 sg13g2_fill_2 FILLER_49_1902 ();
 sg13g2_fill_2 FILLER_49_2074 ();
 sg13g2_fill_1 FILLER_49_2076 ();
 sg13g2_fill_2 FILLER_49_2120 ();
 sg13g2_fill_1 FILLER_49_2122 ();
 sg13g2_fill_2 FILLER_49_2172 ();
 sg13g2_fill_1 FILLER_49_2174 ();
 sg13g2_fill_1 FILLER_49_2198 ();
 sg13g2_fill_2 FILLER_49_2213 ();
 sg13g2_fill_1 FILLER_49_2233 ();
 sg13g2_fill_2 FILLER_49_2280 ();
 sg13g2_fill_1 FILLER_49_2282 ();
 sg13g2_fill_2 FILLER_49_2323 ();
 sg13g2_fill_1 FILLER_49_2325 ();
 sg13g2_decap_8 FILLER_49_2352 ();
 sg13g2_decap_8 FILLER_49_2359 ();
 sg13g2_decap_8 FILLER_49_2366 ();
 sg13g2_decap_8 FILLER_49_2373 ();
 sg13g2_decap_8 FILLER_49_2380 ();
 sg13g2_decap_8 FILLER_49_2387 ();
 sg13g2_decap_8 FILLER_49_2394 ();
 sg13g2_decap_8 FILLER_49_2401 ();
 sg13g2_decap_8 FILLER_49_2408 ();
 sg13g2_decap_8 FILLER_49_2415 ();
 sg13g2_decap_8 FILLER_49_2422 ();
 sg13g2_decap_8 FILLER_49_2429 ();
 sg13g2_decap_8 FILLER_49_2436 ();
 sg13g2_decap_8 FILLER_49_2443 ();
 sg13g2_decap_8 FILLER_49_2450 ();
 sg13g2_decap_8 FILLER_49_2457 ();
 sg13g2_decap_8 FILLER_49_2464 ();
 sg13g2_decap_8 FILLER_49_2471 ();
 sg13g2_decap_8 FILLER_49_2478 ();
 sg13g2_decap_8 FILLER_49_2485 ();
 sg13g2_decap_8 FILLER_49_2492 ();
 sg13g2_decap_8 FILLER_49_2499 ();
 sg13g2_decap_8 FILLER_49_2506 ();
 sg13g2_decap_8 FILLER_49_2513 ();
 sg13g2_decap_8 FILLER_49_2520 ();
 sg13g2_decap_8 FILLER_49_2527 ();
 sg13g2_decap_8 FILLER_49_2534 ();
 sg13g2_decap_8 FILLER_49_2541 ();
 sg13g2_decap_8 FILLER_49_2548 ();
 sg13g2_decap_8 FILLER_49_2555 ();
 sg13g2_decap_8 FILLER_49_2562 ();
 sg13g2_decap_8 FILLER_49_2569 ();
 sg13g2_decap_8 FILLER_49_2576 ();
 sg13g2_decap_8 FILLER_49_2583 ();
 sg13g2_decap_8 FILLER_49_2590 ();
 sg13g2_decap_8 FILLER_49_2597 ();
 sg13g2_decap_8 FILLER_49_2604 ();
 sg13g2_decap_8 FILLER_49_2611 ();
 sg13g2_decap_8 FILLER_49_2618 ();
 sg13g2_decap_8 FILLER_49_2625 ();
 sg13g2_decap_8 FILLER_49_2632 ();
 sg13g2_decap_8 FILLER_49_2639 ();
 sg13g2_decap_8 FILLER_49_2646 ();
 sg13g2_decap_8 FILLER_49_2653 ();
 sg13g2_decap_8 FILLER_49_2660 ();
 sg13g2_decap_8 FILLER_49_2667 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_decap_8 FILLER_50_147 ();
 sg13g2_decap_8 FILLER_50_154 ();
 sg13g2_decap_8 FILLER_50_161 ();
 sg13g2_decap_8 FILLER_50_168 ();
 sg13g2_decap_8 FILLER_50_175 ();
 sg13g2_decap_8 FILLER_50_182 ();
 sg13g2_decap_8 FILLER_50_189 ();
 sg13g2_decap_8 FILLER_50_196 ();
 sg13g2_decap_8 FILLER_50_203 ();
 sg13g2_decap_8 FILLER_50_210 ();
 sg13g2_decap_8 FILLER_50_217 ();
 sg13g2_decap_8 FILLER_50_224 ();
 sg13g2_decap_8 FILLER_50_231 ();
 sg13g2_decap_8 FILLER_50_238 ();
 sg13g2_decap_8 FILLER_50_245 ();
 sg13g2_decap_8 FILLER_50_252 ();
 sg13g2_decap_8 FILLER_50_259 ();
 sg13g2_decap_8 FILLER_50_266 ();
 sg13g2_decap_8 FILLER_50_273 ();
 sg13g2_decap_8 FILLER_50_280 ();
 sg13g2_decap_8 FILLER_50_287 ();
 sg13g2_decap_8 FILLER_50_294 ();
 sg13g2_decap_8 FILLER_50_301 ();
 sg13g2_decap_8 FILLER_50_308 ();
 sg13g2_decap_8 FILLER_50_315 ();
 sg13g2_decap_8 FILLER_50_322 ();
 sg13g2_decap_8 FILLER_50_329 ();
 sg13g2_decap_8 FILLER_50_336 ();
 sg13g2_decap_8 FILLER_50_343 ();
 sg13g2_decap_8 FILLER_50_350 ();
 sg13g2_decap_8 FILLER_50_357 ();
 sg13g2_decap_8 FILLER_50_364 ();
 sg13g2_decap_8 FILLER_50_371 ();
 sg13g2_decap_8 FILLER_50_378 ();
 sg13g2_decap_8 FILLER_50_385 ();
 sg13g2_decap_8 FILLER_50_392 ();
 sg13g2_decap_8 FILLER_50_399 ();
 sg13g2_decap_8 FILLER_50_406 ();
 sg13g2_decap_8 FILLER_50_413 ();
 sg13g2_decap_8 FILLER_50_420 ();
 sg13g2_decap_8 FILLER_50_427 ();
 sg13g2_decap_8 FILLER_50_434 ();
 sg13g2_decap_8 FILLER_50_441 ();
 sg13g2_decap_8 FILLER_50_448 ();
 sg13g2_fill_2 FILLER_50_486 ();
 sg13g2_fill_1 FILLER_50_506 ();
 sg13g2_decap_4 FILLER_50_517 ();
 sg13g2_fill_2 FILLER_50_556 ();
 sg13g2_fill_2 FILLER_50_584 ();
 sg13g2_fill_1 FILLER_50_586 ();
 sg13g2_fill_1 FILLER_50_622 ();
 sg13g2_fill_1 FILLER_50_644 ();
 sg13g2_fill_1 FILLER_50_666 ();
 sg13g2_fill_1 FILLER_50_688 ();
 sg13g2_fill_1 FILLER_50_706 ();
 sg13g2_fill_2 FILLER_50_716 ();
 sg13g2_fill_1 FILLER_50_718 ();
 sg13g2_fill_2 FILLER_50_736 ();
 sg13g2_fill_2 FILLER_50_766 ();
 sg13g2_fill_2 FILLER_50_800 ();
 sg13g2_fill_1 FILLER_50_824 ();
 sg13g2_fill_1 FILLER_50_864 ();
 sg13g2_fill_1 FILLER_50_890 ();
 sg13g2_fill_2 FILLER_50_900 ();
 sg13g2_fill_2 FILLER_50_928 ();
 sg13g2_fill_1 FILLER_50_930 ();
 sg13g2_fill_1 FILLER_50_941 ();
 sg13g2_fill_2 FILLER_50_947 ();
 sg13g2_decap_4 FILLER_50_959 ();
 sg13g2_fill_2 FILLER_50_963 ();
 sg13g2_fill_2 FILLER_50_969 ();
 sg13g2_decap_8 FILLER_50_989 ();
 sg13g2_fill_1 FILLER_50_996 ();
 sg13g2_decap_8 FILLER_50_1002 ();
 sg13g2_fill_1 FILLER_50_1009 ();
 sg13g2_fill_1 FILLER_50_1063 ();
 sg13g2_fill_1 FILLER_50_1078 ();
 sg13g2_fill_2 FILLER_50_1143 ();
 sg13g2_decap_4 FILLER_50_1189 ();
 sg13g2_fill_2 FILLER_50_1201 ();
 sg13g2_fill_1 FILLER_50_1203 ();
 sg13g2_fill_2 FILLER_50_1217 ();
 sg13g2_fill_1 FILLER_50_1231 ();
 sg13g2_fill_1 FILLER_50_1258 ();
 sg13g2_fill_2 FILLER_50_1269 ();
 sg13g2_fill_1 FILLER_50_1284 ();
 sg13g2_fill_2 FILLER_50_1289 ();
 sg13g2_decap_8 FILLER_50_1334 ();
 sg13g2_fill_2 FILLER_50_1341 ();
 sg13g2_fill_1 FILLER_50_1343 ();
 sg13g2_decap_4 FILLER_50_1348 ();
 sg13g2_fill_2 FILLER_50_1385 ();
 sg13g2_fill_2 FILLER_50_1408 ();
 sg13g2_fill_2 FILLER_50_1451 ();
 sg13g2_fill_1 FILLER_50_1453 ();
 sg13g2_fill_2 FILLER_50_1458 ();
 sg13g2_fill_1 FILLER_50_1460 ();
 sg13g2_fill_1 FILLER_50_1474 ();
 sg13g2_fill_2 FILLER_50_1479 ();
 sg13g2_decap_4 FILLER_50_1489 ();
 sg13g2_fill_2 FILLER_50_1493 ();
 sg13g2_fill_2 FILLER_50_1500 ();
 sg13g2_fill_1 FILLER_50_1502 ();
 sg13g2_fill_2 FILLER_50_1507 ();
 sg13g2_fill_1 FILLER_50_1509 ();
 sg13g2_fill_1 FILLER_50_1518 ();
 sg13g2_fill_1 FILLER_50_1571 ();
 sg13g2_decap_4 FILLER_50_1580 ();
 sg13g2_fill_2 FILLER_50_1584 ();
 sg13g2_fill_2 FILLER_50_1601 ();
 sg13g2_fill_1 FILLER_50_1603 ();
 sg13g2_decap_8 FILLER_50_1608 ();
 sg13g2_decap_8 FILLER_50_1615 ();
 sg13g2_decap_8 FILLER_50_1622 ();
 sg13g2_fill_2 FILLER_50_1629 ();
 sg13g2_decap_4 FILLER_50_1640 ();
 sg13g2_decap_4 FILLER_50_1648 ();
 sg13g2_fill_2 FILLER_50_1696 ();
 sg13g2_fill_2 FILLER_50_1729 ();
 sg13g2_fill_1 FILLER_50_1731 ();
 sg13g2_fill_2 FILLER_50_1776 ();
 sg13g2_fill_1 FILLER_50_1778 ();
 sg13g2_fill_2 FILLER_50_1784 ();
 sg13g2_fill_2 FILLER_50_1791 ();
 sg13g2_fill_2 FILLER_50_1797 ();
 sg13g2_fill_1 FILLER_50_1799 ();
 sg13g2_fill_2 FILLER_50_1815 ();
 sg13g2_fill_1 FILLER_50_1848 ();
 sg13g2_decap_8 FILLER_50_1883 ();
 sg13g2_decap_4 FILLER_50_1890 ();
 sg13g2_fill_1 FILLER_50_1894 ();
 sg13g2_fill_1 FILLER_50_1905 ();
 sg13g2_decap_4 FILLER_50_1910 ();
 sg13g2_decap_4 FILLER_50_1927 ();
 sg13g2_fill_1 FILLER_50_1940 ();
 sg13g2_fill_1 FILLER_50_1954 ();
 sg13g2_fill_2 FILLER_50_1959 ();
 sg13g2_fill_2 FILLER_50_1991 ();
 sg13g2_decap_8 FILLER_50_2002 ();
 sg13g2_fill_1 FILLER_50_2009 ();
 sg13g2_fill_2 FILLER_50_2018 ();
 sg13g2_fill_1 FILLER_50_2020 ();
 sg13g2_fill_2 FILLER_50_2035 ();
 sg13g2_fill_1 FILLER_50_2037 ();
 sg13g2_fill_1 FILLER_50_2061 ();
 sg13g2_decap_8 FILLER_50_2071 ();
 sg13g2_fill_1 FILLER_50_2078 ();
 sg13g2_fill_2 FILLER_50_2084 ();
 sg13g2_fill_1 FILLER_50_2086 ();
 sg13g2_fill_2 FILLER_50_2096 ();
 sg13g2_fill_1 FILLER_50_2098 ();
 sg13g2_fill_1 FILLER_50_2103 ();
 sg13g2_fill_2 FILLER_50_2118 ();
 sg13g2_fill_1 FILLER_50_2120 ();
 sg13g2_decap_4 FILLER_50_2156 ();
 sg13g2_fill_2 FILLER_50_2168 ();
 sg13g2_fill_2 FILLER_50_2201 ();
 sg13g2_fill_1 FILLER_50_2203 ();
 sg13g2_fill_1 FILLER_50_2255 ();
 sg13g2_fill_2 FILLER_50_2312 ();
 sg13g2_fill_1 FILLER_50_2319 ();
 sg13g2_fill_2 FILLER_50_2333 ();
 sg13g2_decap_8 FILLER_50_2348 ();
 sg13g2_decap_8 FILLER_50_2355 ();
 sg13g2_decap_8 FILLER_50_2362 ();
 sg13g2_decap_8 FILLER_50_2369 ();
 sg13g2_decap_8 FILLER_50_2376 ();
 sg13g2_decap_8 FILLER_50_2383 ();
 sg13g2_decap_8 FILLER_50_2390 ();
 sg13g2_decap_8 FILLER_50_2397 ();
 sg13g2_decap_8 FILLER_50_2404 ();
 sg13g2_decap_8 FILLER_50_2411 ();
 sg13g2_decap_8 FILLER_50_2418 ();
 sg13g2_decap_8 FILLER_50_2425 ();
 sg13g2_decap_8 FILLER_50_2432 ();
 sg13g2_decap_8 FILLER_50_2439 ();
 sg13g2_decap_8 FILLER_50_2446 ();
 sg13g2_decap_8 FILLER_50_2453 ();
 sg13g2_decap_8 FILLER_50_2460 ();
 sg13g2_decap_8 FILLER_50_2467 ();
 sg13g2_decap_8 FILLER_50_2474 ();
 sg13g2_decap_8 FILLER_50_2481 ();
 sg13g2_decap_8 FILLER_50_2488 ();
 sg13g2_decap_8 FILLER_50_2495 ();
 sg13g2_decap_8 FILLER_50_2502 ();
 sg13g2_decap_8 FILLER_50_2509 ();
 sg13g2_decap_8 FILLER_50_2516 ();
 sg13g2_decap_8 FILLER_50_2523 ();
 sg13g2_decap_8 FILLER_50_2530 ();
 sg13g2_decap_8 FILLER_50_2537 ();
 sg13g2_decap_8 FILLER_50_2544 ();
 sg13g2_decap_8 FILLER_50_2551 ();
 sg13g2_decap_8 FILLER_50_2558 ();
 sg13g2_decap_8 FILLER_50_2565 ();
 sg13g2_decap_8 FILLER_50_2572 ();
 sg13g2_decap_8 FILLER_50_2579 ();
 sg13g2_decap_8 FILLER_50_2586 ();
 sg13g2_decap_8 FILLER_50_2593 ();
 sg13g2_decap_8 FILLER_50_2600 ();
 sg13g2_decap_8 FILLER_50_2607 ();
 sg13g2_decap_8 FILLER_50_2614 ();
 sg13g2_decap_8 FILLER_50_2621 ();
 sg13g2_decap_8 FILLER_50_2628 ();
 sg13g2_decap_8 FILLER_50_2635 ();
 sg13g2_decap_8 FILLER_50_2642 ();
 sg13g2_decap_8 FILLER_50_2649 ();
 sg13g2_decap_8 FILLER_50_2656 ();
 sg13g2_decap_8 FILLER_50_2663 ();
 sg13g2_decap_4 FILLER_50_2670 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_decap_8 FILLER_51_140 ();
 sg13g2_decap_8 FILLER_51_147 ();
 sg13g2_decap_8 FILLER_51_154 ();
 sg13g2_decap_8 FILLER_51_161 ();
 sg13g2_decap_8 FILLER_51_168 ();
 sg13g2_decap_8 FILLER_51_175 ();
 sg13g2_decap_8 FILLER_51_182 ();
 sg13g2_decap_8 FILLER_51_189 ();
 sg13g2_decap_8 FILLER_51_196 ();
 sg13g2_decap_8 FILLER_51_203 ();
 sg13g2_decap_8 FILLER_51_210 ();
 sg13g2_decap_8 FILLER_51_217 ();
 sg13g2_decap_8 FILLER_51_224 ();
 sg13g2_decap_8 FILLER_51_231 ();
 sg13g2_decap_8 FILLER_51_238 ();
 sg13g2_decap_8 FILLER_51_245 ();
 sg13g2_decap_8 FILLER_51_252 ();
 sg13g2_decap_8 FILLER_51_259 ();
 sg13g2_decap_8 FILLER_51_266 ();
 sg13g2_decap_8 FILLER_51_273 ();
 sg13g2_decap_8 FILLER_51_280 ();
 sg13g2_decap_8 FILLER_51_287 ();
 sg13g2_decap_8 FILLER_51_294 ();
 sg13g2_decap_8 FILLER_51_301 ();
 sg13g2_decap_8 FILLER_51_308 ();
 sg13g2_decap_8 FILLER_51_315 ();
 sg13g2_decap_8 FILLER_51_322 ();
 sg13g2_decap_8 FILLER_51_329 ();
 sg13g2_decap_8 FILLER_51_336 ();
 sg13g2_decap_8 FILLER_51_343 ();
 sg13g2_decap_8 FILLER_51_350 ();
 sg13g2_decap_8 FILLER_51_357 ();
 sg13g2_decap_8 FILLER_51_364 ();
 sg13g2_decap_8 FILLER_51_371 ();
 sg13g2_decap_8 FILLER_51_378 ();
 sg13g2_decap_8 FILLER_51_385 ();
 sg13g2_decap_8 FILLER_51_392 ();
 sg13g2_decap_8 FILLER_51_399 ();
 sg13g2_decap_8 FILLER_51_406 ();
 sg13g2_decap_8 FILLER_51_413 ();
 sg13g2_decap_8 FILLER_51_420 ();
 sg13g2_decap_8 FILLER_51_427 ();
 sg13g2_decap_8 FILLER_51_434 ();
 sg13g2_decap_8 FILLER_51_441 ();
 sg13g2_decap_8 FILLER_51_448 ();
 sg13g2_decap_8 FILLER_51_455 ();
 sg13g2_decap_4 FILLER_51_462 ();
 sg13g2_fill_1 FILLER_51_475 ();
 sg13g2_fill_1 FILLER_51_486 ();
 sg13g2_decap_8 FILLER_51_518 ();
 sg13g2_fill_1 FILLER_51_551 ();
 sg13g2_fill_2 FILLER_51_567 ();
 sg13g2_fill_2 FILLER_51_574 ();
 sg13g2_fill_1 FILLER_51_576 ();
 sg13g2_fill_2 FILLER_51_591 ();
 sg13g2_fill_1 FILLER_51_593 ();
 sg13g2_decap_4 FILLER_51_602 ();
 sg13g2_decap_4 FILLER_51_611 ();
 sg13g2_fill_2 FILLER_51_646 ();
 sg13g2_fill_2 FILLER_51_727 ();
 sg13g2_fill_2 FILLER_51_799 ();
 sg13g2_fill_2 FILLER_51_840 ();
 sg13g2_fill_1 FILLER_51_873 ();
 sg13g2_fill_1 FILLER_51_905 ();
 sg13g2_decap_4 FILLER_51_911 ();
 sg13g2_fill_1 FILLER_51_915 ();
 sg13g2_fill_2 FILLER_51_924 ();
 sg13g2_fill_1 FILLER_51_1057 ();
 sg13g2_fill_2 FILLER_51_1093 ();
 sg13g2_fill_2 FILLER_51_1119 ();
 sg13g2_fill_1 FILLER_51_1121 ();
 sg13g2_fill_2 FILLER_51_1175 ();
 sg13g2_fill_1 FILLER_51_1177 ();
 sg13g2_decap_8 FILLER_51_1194 ();
 sg13g2_fill_2 FILLER_51_1263 ();
 sg13g2_fill_2 FILLER_51_1278 ();
 sg13g2_fill_2 FILLER_51_1290 ();
 sg13g2_fill_1 FILLER_51_1301 ();
 sg13g2_fill_2 FILLER_51_1306 ();
 sg13g2_fill_1 FILLER_51_1321 ();
 sg13g2_fill_2 FILLER_51_1448 ();
 sg13g2_fill_1 FILLER_51_1491 ();
 sg13g2_fill_1 FILLER_51_1518 ();
 sg13g2_fill_1 FILLER_51_1533 ();
 sg13g2_fill_2 FILLER_51_1539 ();
 sg13g2_fill_1 FILLER_51_1541 ();
 sg13g2_fill_2 FILLER_51_1673 ();
 sg13g2_fill_2 FILLER_51_1728 ();
 sg13g2_fill_2 FILLER_51_1788 ();
 sg13g2_fill_2 FILLER_51_1816 ();
 sg13g2_decap_8 FILLER_51_1840 ();
 sg13g2_fill_1 FILLER_51_1847 ();
 sg13g2_fill_2 FILLER_51_1853 ();
 sg13g2_fill_2 FILLER_51_1864 ();
 sg13g2_fill_1 FILLER_51_1866 ();
 sg13g2_fill_1 FILLER_51_1955 ();
 sg13g2_fill_2 FILLER_51_1960 ();
 sg13g2_fill_1 FILLER_51_1962 ();
 sg13g2_fill_1 FILLER_51_2021 ();
 sg13g2_decap_4 FILLER_51_2084 ();
 sg13g2_fill_1 FILLER_51_2114 ();
 sg13g2_decap_4 FILLER_51_2141 ();
 sg13g2_fill_2 FILLER_51_2145 ();
 sg13g2_fill_2 FILLER_51_2152 ();
 sg13g2_fill_1 FILLER_51_2154 ();
 sg13g2_fill_1 FILLER_51_2167 ();
 sg13g2_fill_1 FILLER_51_2177 ();
 sg13g2_fill_2 FILLER_51_2213 ();
 sg13g2_fill_2 FILLER_51_2253 ();
 sg13g2_fill_2 FILLER_51_2263 ();
 sg13g2_fill_1 FILLER_51_2265 ();
 sg13g2_fill_2 FILLER_51_2288 ();
 sg13g2_decap_8 FILLER_51_2342 ();
 sg13g2_decap_8 FILLER_51_2349 ();
 sg13g2_decap_8 FILLER_51_2356 ();
 sg13g2_decap_8 FILLER_51_2363 ();
 sg13g2_decap_8 FILLER_51_2370 ();
 sg13g2_decap_8 FILLER_51_2377 ();
 sg13g2_decap_8 FILLER_51_2384 ();
 sg13g2_decap_8 FILLER_51_2391 ();
 sg13g2_decap_8 FILLER_51_2398 ();
 sg13g2_decap_8 FILLER_51_2405 ();
 sg13g2_decap_8 FILLER_51_2412 ();
 sg13g2_decap_8 FILLER_51_2419 ();
 sg13g2_decap_8 FILLER_51_2426 ();
 sg13g2_decap_8 FILLER_51_2433 ();
 sg13g2_decap_8 FILLER_51_2440 ();
 sg13g2_decap_8 FILLER_51_2447 ();
 sg13g2_decap_8 FILLER_51_2454 ();
 sg13g2_decap_8 FILLER_51_2461 ();
 sg13g2_decap_8 FILLER_51_2468 ();
 sg13g2_decap_8 FILLER_51_2475 ();
 sg13g2_decap_8 FILLER_51_2482 ();
 sg13g2_decap_8 FILLER_51_2489 ();
 sg13g2_decap_8 FILLER_51_2496 ();
 sg13g2_decap_8 FILLER_51_2503 ();
 sg13g2_decap_8 FILLER_51_2510 ();
 sg13g2_decap_8 FILLER_51_2517 ();
 sg13g2_decap_8 FILLER_51_2524 ();
 sg13g2_decap_8 FILLER_51_2531 ();
 sg13g2_decap_8 FILLER_51_2538 ();
 sg13g2_decap_8 FILLER_51_2545 ();
 sg13g2_decap_8 FILLER_51_2552 ();
 sg13g2_decap_8 FILLER_51_2559 ();
 sg13g2_decap_8 FILLER_51_2566 ();
 sg13g2_decap_8 FILLER_51_2573 ();
 sg13g2_decap_8 FILLER_51_2580 ();
 sg13g2_decap_8 FILLER_51_2587 ();
 sg13g2_decap_8 FILLER_51_2594 ();
 sg13g2_decap_8 FILLER_51_2601 ();
 sg13g2_decap_8 FILLER_51_2608 ();
 sg13g2_decap_8 FILLER_51_2615 ();
 sg13g2_decap_8 FILLER_51_2622 ();
 sg13g2_decap_8 FILLER_51_2629 ();
 sg13g2_decap_8 FILLER_51_2636 ();
 sg13g2_decap_8 FILLER_51_2643 ();
 sg13g2_decap_8 FILLER_51_2650 ();
 sg13g2_decap_8 FILLER_51_2657 ();
 sg13g2_decap_8 FILLER_51_2664 ();
 sg13g2_fill_2 FILLER_51_2671 ();
 sg13g2_fill_1 FILLER_51_2673 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_decap_8 FILLER_52_133 ();
 sg13g2_decap_8 FILLER_52_140 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_154 ();
 sg13g2_decap_8 FILLER_52_161 ();
 sg13g2_decap_8 FILLER_52_168 ();
 sg13g2_decap_8 FILLER_52_175 ();
 sg13g2_decap_8 FILLER_52_182 ();
 sg13g2_decap_8 FILLER_52_189 ();
 sg13g2_decap_8 FILLER_52_196 ();
 sg13g2_decap_8 FILLER_52_203 ();
 sg13g2_decap_8 FILLER_52_210 ();
 sg13g2_decap_8 FILLER_52_217 ();
 sg13g2_decap_8 FILLER_52_224 ();
 sg13g2_decap_8 FILLER_52_231 ();
 sg13g2_decap_8 FILLER_52_238 ();
 sg13g2_decap_8 FILLER_52_245 ();
 sg13g2_decap_8 FILLER_52_252 ();
 sg13g2_decap_8 FILLER_52_259 ();
 sg13g2_decap_8 FILLER_52_266 ();
 sg13g2_decap_8 FILLER_52_273 ();
 sg13g2_decap_8 FILLER_52_280 ();
 sg13g2_decap_8 FILLER_52_287 ();
 sg13g2_decap_8 FILLER_52_294 ();
 sg13g2_decap_8 FILLER_52_301 ();
 sg13g2_decap_8 FILLER_52_308 ();
 sg13g2_decap_8 FILLER_52_315 ();
 sg13g2_decap_8 FILLER_52_322 ();
 sg13g2_decap_8 FILLER_52_329 ();
 sg13g2_decap_8 FILLER_52_336 ();
 sg13g2_decap_8 FILLER_52_343 ();
 sg13g2_decap_8 FILLER_52_350 ();
 sg13g2_decap_8 FILLER_52_357 ();
 sg13g2_decap_8 FILLER_52_364 ();
 sg13g2_decap_8 FILLER_52_371 ();
 sg13g2_decap_8 FILLER_52_378 ();
 sg13g2_decap_8 FILLER_52_385 ();
 sg13g2_decap_8 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_decap_8 FILLER_52_406 ();
 sg13g2_decap_8 FILLER_52_413 ();
 sg13g2_decap_8 FILLER_52_420 ();
 sg13g2_decap_8 FILLER_52_427 ();
 sg13g2_decap_8 FILLER_52_434 ();
 sg13g2_decap_8 FILLER_52_441 ();
 sg13g2_fill_1 FILLER_52_448 ();
 sg13g2_fill_2 FILLER_52_475 ();
 sg13g2_fill_1 FILLER_52_576 ();
 sg13g2_fill_2 FILLER_52_582 ();
 sg13g2_fill_1 FILLER_52_584 ();
 sg13g2_decap_4 FILLER_52_637 ();
 sg13g2_fill_1 FILLER_52_641 ();
 sg13g2_fill_2 FILLER_52_651 ();
 sg13g2_fill_1 FILLER_52_700 ();
 sg13g2_fill_1 FILLER_52_727 ();
 sg13g2_fill_2 FILLER_52_744 ();
 sg13g2_fill_2 FILLER_52_751 ();
 sg13g2_fill_1 FILLER_52_753 ();
 sg13g2_fill_2 FILLER_52_846 ();
 sg13g2_fill_1 FILLER_52_848 ();
 sg13g2_decap_4 FILLER_52_872 ();
 sg13g2_fill_2 FILLER_52_885 ();
 sg13g2_fill_1 FILLER_52_887 ();
 sg13g2_fill_2 FILLER_52_944 ();
 sg13g2_fill_1 FILLER_52_950 ();
 sg13g2_decap_4 FILLER_52_955 ();
 sg13g2_fill_2 FILLER_52_959 ();
 sg13g2_decap_4 FILLER_52_979 ();
 sg13g2_fill_2 FILLER_52_983 ();
 sg13g2_fill_2 FILLER_52_998 ();
 sg13g2_fill_1 FILLER_52_1004 ();
 sg13g2_fill_1 FILLER_52_1039 ();
 sg13g2_fill_2 FILLER_52_1054 ();
 sg13g2_fill_2 FILLER_52_1069 ();
 sg13g2_fill_2 FILLER_52_1081 ();
 sg13g2_fill_1 FILLER_52_1088 ();
 sg13g2_fill_2 FILLER_52_1132 ();
 sg13g2_fill_1 FILLER_52_1134 ();
 sg13g2_fill_1 FILLER_52_1140 ();
 sg13g2_fill_2 FILLER_52_1150 ();
 sg13g2_fill_1 FILLER_52_1152 ();
 sg13g2_decap_4 FILLER_52_1193 ();
 sg13g2_fill_2 FILLER_52_1227 ();
 sg13g2_fill_1 FILLER_52_1229 ();
 sg13g2_fill_1 FILLER_52_1234 ();
 sg13g2_fill_2 FILLER_52_1240 ();
 sg13g2_fill_1 FILLER_52_1247 ();
 sg13g2_fill_2 FILLER_52_1253 ();
 sg13g2_fill_1 FILLER_52_1286 ();
 sg13g2_fill_2 FILLER_52_1309 ();
 sg13g2_fill_1 FILLER_52_1311 ();
 sg13g2_fill_1 FILLER_52_1316 ();
 sg13g2_fill_1 FILLER_52_1321 ();
 sg13g2_fill_2 FILLER_52_1330 ();
 sg13g2_fill_1 FILLER_52_1332 ();
 sg13g2_fill_1 FILLER_52_1337 ();
 sg13g2_fill_1 FILLER_52_1416 ();
 sg13g2_fill_1 FILLER_52_1465 ();
 sg13g2_fill_2 FILLER_52_1475 ();
 sg13g2_fill_1 FILLER_52_1487 ();
 sg13g2_fill_2 FILLER_52_1505 ();
 sg13g2_fill_1 FILLER_52_1507 ();
 sg13g2_fill_2 FILLER_52_1512 ();
 sg13g2_fill_2 FILLER_52_1523 ();
 sg13g2_fill_1 FILLER_52_1525 ();
 sg13g2_fill_1 FILLER_52_1556 ();
 sg13g2_fill_2 FILLER_52_1570 ();
 sg13g2_fill_1 FILLER_52_1589 ();
 sg13g2_fill_1 FILLER_52_1608 ();
 sg13g2_fill_1 FILLER_52_1618 ();
 sg13g2_decap_8 FILLER_52_1632 ();
 sg13g2_fill_2 FILLER_52_1639 ();
 sg13g2_fill_1 FILLER_52_1641 ();
 sg13g2_fill_1 FILLER_52_1672 ();
 sg13g2_fill_1 FILLER_52_1686 ();
 sg13g2_fill_2 FILLER_52_1701 ();
 sg13g2_fill_1 FILLER_52_1711 ();
 sg13g2_fill_2 FILLER_52_1732 ();
 sg13g2_fill_2 FILLER_52_1761 ();
 sg13g2_fill_1 FILLER_52_1763 ();
 sg13g2_fill_2 FILLER_52_1768 ();
 sg13g2_fill_1 FILLER_52_1778 ();
 sg13g2_fill_2 FILLER_52_1801 ();
 sg13g2_fill_1 FILLER_52_1812 ();
 sg13g2_fill_2 FILLER_52_1873 ();
 sg13g2_fill_1 FILLER_52_1875 ();
 sg13g2_decap_4 FILLER_52_1902 ();
 sg13g2_fill_2 FILLER_52_1911 ();
 sg13g2_decap_8 FILLER_52_1917 ();
 sg13g2_fill_1 FILLER_52_1924 ();
 sg13g2_fill_2 FILLER_52_1929 ();
 sg13g2_fill_2 FILLER_52_1940 ();
 sg13g2_fill_1 FILLER_52_1942 ();
 sg13g2_fill_1 FILLER_52_1984 ();
 sg13g2_fill_2 FILLER_52_1994 ();
 sg13g2_decap_4 FILLER_52_2013 ();
 sg13g2_fill_1 FILLER_52_2022 ();
 sg13g2_fill_2 FILLER_52_2030 ();
 sg13g2_fill_1 FILLER_52_2040 ();
 sg13g2_fill_2 FILLER_52_2059 ();
 sg13g2_fill_2 FILLER_52_2065 ();
 sg13g2_fill_1 FILLER_52_2072 ();
 sg13g2_fill_2 FILLER_52_2082 ();
 sg13g2_fill_1 FILLER_52_2093 ();
 sg13g2_fill_2 FILLER_52_2098 ();
 sg13g2_decap_8 FILLER_52_2109 ();
 sg13g2_fill_1 FILLER_52_2116 ();
 sg13g2_fill_2 FILLER_52_2134 ();
 sg13g2_fill_1 FILLER_52_2136 ();
 sg13g2_fill_2 FILLER_52_2146 ();
 sg13g2_fill_1 FILLER_52_2148 ();
 sg13g2_fill_2 FILLER_52_2201 ();
 sg13g2_fill_2 FILLER_52_2210 ();
 sg13g2_fill_1 FILLER_52_2212 ();
 sg13g2_fill_1 FILLER_52_2218 ();
 sg13g2_fill_2 FILLER_52_2224 ();
 sg13g2_fill_1 FILLER_52_2226 ();
 sg13g2_fill_2 FILLER_52_2245 ();
 sg13g2_fill_1 FILLER_52_2247 ();
 sg13g2_fill_2 FILLER_52_2261 ();
 sg13g2_fill_2 FILLER_52_2302 ();
 sg13g2_decap_8 FILLER_52_2317 ();
 sg13g2_fill_1 FILLER_52_2324 ();
 sg13g2_fill_2 FILLER_52_2329 ();
 sg13g2_decap_8 FILLER_52_2340 ();
 sg13g2_decap_8 FILLER_52_2347 ();
 sg13g2_decap_8 FILLER_52_2354 ();
 sg13g2_decap_8 FILLER_52_2361 ();
 sg13g2_decap_8 FILLER_52_2368 ();
 sg13g2_decap_8 FILLER_52_2375 ();
 sg13g2_decap_8 FILLER_52_2382 ();
 sg13g2_decap_8 FILLER_52_2389 ();
 sg13g2_decap_8 FILLER_52_2396 ();
 sg13g2_decap_8 FILLER_52_2403 ();
 sg13g2_decap_8 FILLER_52_2410 ();
 sg13g2_decap_8 FILLER_52_2417 ();
 sg13g2_decap_8 FILLER_52_2424 ();
 sg13g2_decap_8 FILLER_52_2431 ();
 sg13g2_decap_8 FILLER_52_2438 ();
 sg13g2_decap_8 FILLER_52_2445 ();
 sg13g2_decap_8 FILLER_52_2452 ();
 sg13g2_decap_8 FILLER_52_2459 ();
 sg13g2_decap_8 FILLER_52_2466 ();
 sg13g2_decap_8 FILLER_52_2473 ();
 sg13g2_decap_8 FILLER_52_2480 ();
 sg13g2_decap_8 FILLER_52_2487 ();
 sg13g2_decap_8 FILLER_52_2494 ();
 sg13g2_decap_8 FILLER_52_2501 ();
 sg13g2_decap_8 FILLER_52_2508 ();
 sg13g2_decap_8 FILLER_52_2515 ();
 sg13g2_decap_8 FILLER_52_2522 ();
 sg13g2_decap_8 FILLER_52_2529 ();
 sg13g2_decap_8 FILLER_52_2536 ();
 sg13g2_decap_8 FILLER_52_2543 ();
 sg13g2_decap_8 FILLER_52_2550 ();
 sg13g2_decap_8 FILLER_52_2557 ();
 sg13g2_decap_8 FILLER_52_2564 ();
 sg13g2_decap_8 FILLER_52_2571 ();
 sg13g2_decap_8 FILLER_52_2578 ();
 sg13g2_decap_8 FILLER_52_2585 ();
 sg13g2_decap_8 FILLER_52_2592 ();
 sg13g2_decap_8 FILLER_52_2599 ();
 sg13g2_decap_8 FILLER_52_2606 ();
 sg13g2_decap_8 FILLER_52_2613 ();
 sg13g2_decap_8 FILLER_52_2620 ();
 sg13g2_decap_8 FILLER_52_2627 ();
 sg13g2_decap_8 FILLER_52_2634 ();
 sg13g2_decap_8 FILLER_52_2641 ();
 sg13g2_decap_8 FILLER_52_2648 ();
 sg13g2_decap_8 FILLER_52_2655 ();
 sg13g2_decap_8 FILLER_52_2662 ();
 sg13g2_decap_4 FILLER_52_2669 ();
 sg13g2_fill_1 FILLER_52_2673 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_133 ();
 sg13g2_decap_8 FILLER_53_140 ();
 sg13g2_decap_8 FILLER_53_147 ();
 sg13g2_decap_8 FILLER_53_154 ();
 sg13g2_decap_8 FILLER_53_161 ();
 sg13g2_decap_8 FILLER_53_168 ();
 sg13g2_decap_8 FILLER_53_175 ();
 sg13g2_decap_8 FILLER_53_182 ();
 sg13g2_decap_8 FILLER_53_189 ();
 sg13g2_decap_8 FILLER_53_196 ();
 sg13g2_decap_8 FILLER_53_203 ();
 sg13g2_decap_8 FILLER_53_210 ();
 sg13g2_decap_8 FILLER_53_217 ();
 sg13g2_decap_8 FILLER_53_224 ();
 sg13g2_decap_8 FILLER_53_231 ();
 sg13g2_decap_8 FILLER_53_238 ();
 sg13g2_decap_8 FILLER_53_245 ();
 sg13g2_decap_8 FILLER_53_252 ();
 sg13g2_decap_8 FILLER_53_259 ();
 sg13g2_decap_8 FILLER_53_266 ();
 sg13g2_decap_8 FILLER_53_273 ();
 sg13g2_decap_8 FILLER_53_280 ();
 sg13g2_decap_8 FILLER_53_287 ();
 sg13g2_decap_8 FILLER_53_294 ();
 sg13g2_decap_8 FILLER_53_301 ();
 sg13g2_decap_8 FILLER_53_308 ();
 sg13g2_decap_8 FILLER_53_315 ();
 sg13g2_decap_8 FILLER_53_322 ();
 sg13g2_decap_8 FILLER_53_329 ();
 sg13g2_decap_8 FILLER_53_336 ();
 sg13g2_decap_8 FILLER_53_343 ();
 sg13g2_decap_8 FILLER_53_350 ();
 sg13g2_decap_8 FILLER_53_357 ();
 sg13g2_decap_8 FILLER_53_364 ();
 sg13g2_decap_8 FILLER_53_371 ();
 sg13g2_decap_8 FILLER_53_378 ();
 sg13g2_decap_8 FILLER_53_385 ();
 sg13g2_decap_8 FILLER_53_392 ();
 sg13g2_decap_8 FILLER_53_399 ();
 sg13g2_decap_8 FILLER_53_406 ();
 sg13g2_decap_8 FILLER_53_413 ();
 sg13g2_decap_8 FILLER_53_420 ();
 sg13g2_decap_8 FILLER_53_427 ();
 sg13g2_decap_8 FILLER_53_434 ();
 sg13g2_decap_8 FILLER_53_441 ();
 sg13g2_decap_8 FILLER_53_448 ();
 sg13g2_fill_2 FILLER_53_499 ();
 sg13g2_fill_1 FILLER_53_524 ();
 sg13g2_fill_2 FILLER_53_534 ();
 sg13g2_fill_2 FILLER_53_605 ();
 sg13g2_fill_1 FILLER_53_607 ();
 sg13g2_fill_2 FILLER_53_618 ();
 sg13g2_fill_1 FILLER_53_620 ();
 sg13g2_decap_4 FILLER_53_636 ();
 sg13g2_fill_2 FILLER_53_650 ();
 sg13g2_fill_1 FILLER_53_661 ();
 sg13g2_fill_2 FILLER_53_670 ();
 sg13g2_fill_1 FILLER_53_672 ();
 sg13g2_fill_2 FILLER_53_704 ();
 sg13g2_fill_1 FILLER_53_706 ();
 sg13g2_fill_2 FILLER_53_767 ();
 sg13g2_fill_2 FILLER_53_804 ();
 sg13g2_fill_2 FILLER_53_901 ();
 sg13g2_fill_2 FILLER_53_907 ();
 sg13g2_fill_1 FILLER_53_913 ();
 sg13g2_decap_4 FILLER_53_923 ();
 sg13g2_fill_2 FILLER_53_927 ();
 sg13g2_decap_8 FILLER_53_933 ();
 sg13g2_fill_2 FILLER_53_940 ();
 sg13g2_fill_1 FILLER_53_942 ();
 sg13g2_fill_1 FILLER_53_1021 ();
 sg13g2_fill_2 FILLER_53_1082 ();
 sg13g2_fill_2 FILLER_53_1089 ();
 sg13g2_fill_2 FILLER_53_1117 ();
 sg13g2_fill_1 FILLER_53_1119 ();
 sg13g2_fill_2 FILLER_53_1137 ();
 sg13g2_fill_1 FILLER_53_1139 ();
 sg13g2_fill_2 FILLER_53_1145 ();
 sg13g2_fill_1 FILLER_53_1147 ();
 sg13g2_decap_4 FILLER_53_1184 ();
 sg13g2_fill_1 FILLER_53_1188 ();
 sg13g2_decap_8 FILLER_53_1194 ();
 sg13g2_fill_1 FILLER_53_1206 ();
 sg13g2_fill_1 FILLER_53_1215 ();
 sg13g2_fill_1 FILLER_53_1225 ();
 sg13g2_decap_4 FILLER_53_1256 ();
 sg13g2_fill_2 FILLER_53_1269 ();
 sg13g2_fill_1 FILLER_53_1271 ();
 sg13g2_fill_1 FILLER_53_1276 ();
 sg13g2_fill_2 FILLER_53_1299 ();
 sg13g2_fill_1 FILLER_53_1332 ();
 sg13g2_decap_8 FILLER_53_1358 ();
 sg13g2_decap_8 FILLER_53_1373 ();
 sg13g2_decap_8 FILLER_53_1380 ();
 sg13g2_fill_1 FILLER_53_1387 ();
 sg13g2_fill_2 FILLER_53_1397 ();
 sg13g2_fill_1 FILLER_53_1399 ();
 sg13g2_decap_8 FILLER_53_1423 ();
 sg13g2_decap_4 FILLER_53_1430 ();
 sg13g2_fill_2 FILLER_53_1434 ();
 sg13g2_fill_2 FILLER_53_1482 ();
 sg13g2_fill_1 FILLER_53_1564 ();
 sg13g2_fill_1 FILLER_53_1570 ();
 sg13g2_decap_8 FILLER_53_1579 ();
 sg13g2_fill_2 FILLER_53_1586 ();
 sg13g2_fill_2 FILLER_53_1670 ();
 sg13g2_fill_1 FILLER_53_1672 ();
 sg13g2_fill_1 FILLER_53_1678 ();
 sg13g2_fill_1 FILLER_53_1717 ();
 sg13g2_fill_2 FILLER_53_1770 ();
 sg13g2_fill_1 FILLER_53_1792 ();
 sg13g2_fill_2 FILLER_53_1832 ();
 sg13g2_fill_1 FILLER_53_1834 ();
 sg13g2_fill_1 FILLER_53_1861 ();
 sg13g2_fill_2 FILLER_53_1871 ();
 sg13g2_fill_1 FILLER_53_1873 ();
 sg13g2_fill_1 FILLER_53_1883 ();
 sg13g2_fill_1 FILLER_53_1908 ();
 sg13g2_fill_1 FILLER_53_1967 ();
 sg13g2_fill_2 FILLER_53_1973 ();
 sg13g2_fill_2 FILLER_53_2013 ();
 sg13g2_fill_1 FILLER_53_2015 ();
 sg13g2_fill_2 FILLER_53_2020 ();
 sg13g2_fill_2 FILLER_53_2041 ();
 sg13g2_fill_2 FILLER_53_2076 ();
 sg13g2_fill_1 FILLER_53_2170 ();
 sg13g2_fill_2 FILLER_53_2291 ();
 sg13g2_decap_8 FILLER_53_2324 ();
 sg13g2_decap_8 FILLER_53_2331 ();
 sg13g2_decap_8 FILLER_53_2338 ();
 sg13g2_decap_8 FILLER_53_2345 ();
 sg13g2_decap_8 FILLER_53_2352 ();
 sg13g2_decap_8 FILLER_53_2359 ();
 sg13g2_decap_8 FILLER_53_2366 ();
 sg13g2_decap_8 FILLER_53_2373 ();
 sg13g2_decap_8 FILLER_53_2380 ();
 sg13g2_decap_8 FILLER_53_2387 ();
 sg13g2_decap_8 FILLER_53_2394 ();
 sg13g2_decap_8 FILLER_53_2401 ();
 sg13g2_decap_8 FILLER_53_2408 ();
 sg13g2_decap_8 FILLER_53_2415 ();
 sg13g2_decap_8 FILLER_53_2422 ();
 sg13g2_decap_8 FILLER_53_2429 ();
 sg13g2_decap_8 FILLER_53_2436 ();
 sg13g2_decap_8 FILLER_53_2443 ();
 sg13g2_decap_8 FILLER_53_2450 ();
 sg13g2_decap_8 FILLER_53_2457 ();
 sg13g2_decap_8 FILLER_53_2464 ();
 sg13g2_decap_8 FILLER_53_2471 ();
 sg13g2_decap_8 FILLER_53_2478 ();
 sg13g2_decap_8 FILLER_53_2485 ();
 sg13g2_decap_8 FILLER_53_2492 ();
 sg13g2_decap_8 FILLER_53_2499 ();
 sg13g2_decap_8 FILLER_53_2506 ();
 sg13g2_decap_8 FILLER_53_2513 ();
 sg13g2_decap_8 FILLER_53_2520 ();
 sg13g2_decap_8 FILLER_53_2527 ();
 sg13g2_decap_8 FILLER_53_2534 ();
 sg13g2_decap_8 FILLER_53_2541 ();
 sg13g2_decap_8 FILLER_53_2548 ();
 sg13g2_decap_8 FILLER_53_2555 ();
 sg13g2_decap_8 FILLER_53_2562 ();
 sg13g2_decap_8 FILLER_53_2569 ();
 sg13g2_decap_8 FILLER_53_2576 ();
 sg13g2_decap_8 FILLER_53_2583 ();
 sg13g2_decap_8 FILLER_53_2590 ();
 sg13g2_decap_8 FILLER_53_2597 ();
 sg13g2_decap_8 FILLER_53_2604 ();
 sg13g2_decap_8 FILLER_53_2611 ();
 sg13g2_decap_8 FILLER_53_2618 ();
 sg13g2_decap_8 FILLER_53_2625 ();
 sg13g2_decap_8 FILLER_53_2632 ();
 sg13g2_decap_8 FILLER_53_2639 ();
 sg13g2_decap_8 FILLER_53_2646 ();
 sg13g2_decap_8 FILLER_53_2653 ();
 sg13g2_decap_8 FILLER_53_2660 ();
 sg13g2_decap_8 FILLER_53_2667 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_decap_8 FILLER_54_133 ();
 sg13g2_decap_8 FILLER_54_140 ();
 sg13g2_decap_8 FILLER_54_147 ();
 sg13g2_decap_8 FILLER_54_154 ();
 sg13g2_decap_8 FILLER_54_161 ();
 sg13g2_decap_8 FILLER_54_168 ();
 sg13g2_decap_8 FILLER_54_175 ();
 sg13g2_decap_8 FILLER_54_182 ();
 sg13g2_decap_8 FILLER_54_189 ();
 sg13g2_decap_8 FILLER_54_196 ();
 sg13g2_decap_8 FILLER_54_203 ();
 sg13g2_decap_8 FILLER_54_210 ();
 sg13g2_decap_8 FILLER_54_217 ();
 sg13g2_decap_8 FILLER_54_224 ();
 sg13g2_decap_8 FILLER_54_231 ();
 sg13g2_decap_8 FILLER_54_238 ();
 sg13g2_decap_8 FILLER_54_245 ();
 sg13g2_decap_8 FILLER_54_252 ();
 sg13g2_decap_8 FILLER_54_259 ();
 sg13g2_decap_8 FILLER_54_266 ();
 sg13g2_decap_8 FILLER_54_273 ();
 sg13g2_decap_8 FILLER_54_280 ();
 sg13g2_decap_8 FILLER_54_287 ();
 sg13g2_decap_8 FILLER_54_294 ();
 sg13g2_decap_8 FILLER_54_301 ();
 sg13g2_decap_8 FILLER_54_308 ();
 sg13g2_decap_8 FILLER_54_315 ();
 sg13g2_decap_8 FILLER_54_322 ();
 sg13g2_decap_8 FILLER_54_329 ();
 sg13g2_decap_8 FILLER_54_336 ();
 sg13g2_decap_8 FILLER_54_343 ();
 sg13g2_decap_8 FILLER_54_350 ();
 sg13g2_decap_8 FILLER_54_357 ();
 sg13g2_decap_8 FILLER_54_364 ();
 sg13g2_decap_8 FILLER_54_371 ();
 sg13g2_decap_8 FILLER_54_378 ();
 sg13g2_decap_8 FILLER_54_385 ();
 sg13g2_decap_8 FILLER_54_392 ();
 sg13g2_decap_8 FILLER_54_399 ();
 sg13g2_decap_8 FILLER_54_406 ();
 sg13g2_decap_8 FILLER_54_413 ();
 sg13g2_decap_8 FILLER_54_420 ();
 sg13g2_decap_8 FILLER_54_427 ();
 sg13g2_decap_8 FILLER_54_434 ();
 sg13g2_decap_8 FILLER_54_441 ();
 sg13g2_decap_8 FILLER_54_448 ();
 sg13g2_decap_4 FILLER_54_455 ();
 sg13g2_fill_2 FILLER_54_459 ();
 sg13g2_fill_1 FILLER_54_532 ();
 sg13g2_fill_1 FILLER_54_541 ();
 sg13g2_decap_4 FILLER_54_547 ();
 sg13g2_fill_1 FILLER_54_575 ();
 sg13g2_decap_4 FILLER_54_636 ();
 sg13g2_fill_2 FILLER_54_640 ();
 sg13g2_decap_8 FILLER_54_678 ();
 sg13g2_decap_4 FILLER_54_714 ();
 sg13g2_fill_2 FILLER_54_718 ();
 sg13g2_decap_8 FILLER_54_728 ();
 sg13g2_decap_4 FILLER_54_746 ();
 sg13g2_fill_1 FILLER_54_763 ();
 sg13g2_fill_2 FILLER_54_777 ();
 sg13g2_fill_1 FILLER_54_779 ();
 sg13g2_fill_2 FILLER_54_789 ();
 sg13g2_fill_1 FILLER_54_791 ();
 sg13g2_fill_2 FILLER_54_824 ();
 sg13g2_fill_1 FILLER_54_826 ();
 sg13g2_fill_1 FILLER_54_879 ();
 sg13g2_decap_8 FILLER_54_927 ();
 sg13g2_fill_2 FILLER_54_947 ();
 sg13g2_fill_1 FILLER_54_954 ();
 sg13g2_fill_2 FILLER_54_964 ();
 sg13g2_fill_1 FILLER_54_966 ();
 sg13g2_fill_1 FILLER_54_1028 ();
 sg13g2_fill_2 FILLER_54_1034 ();
 sg13g2_decap_8 FILLER_54_1044 ();
 sg13g2_fill_2 FILLER_54_1081 ();
 sg13g2_fill_1 FILLER_54_1123 ();
 sg13g2_fill_1 FILLER_54_1168 ();
 sg13g2_decap_8 FILLER_54_1177 ();
 sg13g2_fill_2 FILLER_54_1184 ();
 sg13g2_fill_2 FILLER_54_1226 ();
 sg13g2_fill_1 FILLER_54_1228 ();
 sg13g2_fill_1 FILLER_54_1267 ();
 sg13g2_fill_2 FILLER_54_1277 ();
 sg13g2_fill_1 FILLER_54_1279 ();
 sg13g2_fill_2 FILLER_54_1311 ();
 sg13g2_decap_8 FILLER_54_1357 ();
 sg13g2_decap_4 FILLER_54_1364 ();
 sg13g2_fill_1 FILLER_54_1437 ();
 sg13g2_fill_2 FILLER_54_1457 ();
 sg13g2_fill_2 FILLER_54_1468 ();
 sg13g2_fill_2 FILLER_54_1492 ();
 sg13g2_fill_1 FILLER_54_1494 ();
 sg13g2_fill_1 FILLER_54_1499 ();
 sg13g2_fill_2 FILLER_54_1505 ();
 sg13g2_fill_1 FILLER_54_1507 ();
 sg13g2_fill_2 FILLER_54_1516 ();
 sg13g2_fill_2 FILLER_54_1538 ();
 sg13g2_fill_1 FILLER_54_1540 ();
 sg13g2_decap_4 FILLER_54_1571 ();
 sg13g2_fill_2 FILLER_54_1575 ();
 sg13g2_decap_8 FILLER_54_1587 ();
 sg13g2_decap_8 FILLER_54_1594 ();
 sg13g2_decap_4 FILLER_54_1601 ();
 sg13g2_fill_1 FILLER_54_1605 ();
 sg13g2_fill_1 FILLER_54_1624 ();
 sg13g2_fill_2 FILLER_54_1638 ();
 sg13g2_fill_1 FILLER_54_1640 ();
 sg13g2_decap_4 FILLER_54_1732 ();
 sg13g2_fill_1 FILLER_54_1736 ();
 sg13g2_decap_4 FILLER_54_1772 ();
 sg13g2_fill_2 FILLER_54_1825 ();
 sg13g2_fill_1 FILLER_54_1853 ();
 sg13g2_decap_4 FILLER_54_1900 ();
 sg13g2_fill_2 FILLER_54_1943 ();
 sg13g2_fill_1 FILLER_54_1955 ();
 sg13g2_fill_2 FILLER_54_1971 ();
 sg13g2_fill_1 FILLER_54_1973 ();
 sg13g2_fill_2 FILLER_54_1979 ();
 sg13g2_fill_1 FILLER_54_1981 ();
 sg13g2_fill_2 FILLER_54_1996 ();
 sg13g2_fill_2 FILLER_54_2054 ();
 sg13g2_fill_1 FILLER_54_2056 ();
 sg13g2_fill_1 FILLER_54_2086 ();
 sg13g2_decap_8 FILLER_54_2091 ();
 sg13g2_decap_8 FILLER_54_2098 ();
 sg13g2_decap_8 FILLER_54_2105 ();
 sg13g2_fill_2 FILLER_54_2112 ();
 sg13g2_fill_2 FILLER_54_2118 ();
 sg13g2_fill_1 FILLER_54_2120 ();
 sg13g2_fill_1 FILLER_54_2130 ();
 sg13g2_decap_4 FILLER_54_2145 ();
 sg13g2_fill_2 FILLER_54_2159 ();
 sg13g2_fill_2 FILLER_54_2188 ();
 sg13g2_fill_1 FILLER_54_2190 ();
 sg13g2_fill_2 FILLER_54_2214 ();
 sg13g2_fill_2 FILLER_54_2226 ();
 sg13g2_fill_2 FILLER_54_2237 ();
 sg13g2_fill_2 FILLER_54_2252 ();
 sg13g2_fill_1 FILLER_54_2272 ();
 sg13g2_fill_1 FILLER_54_2278 ();
 sg13g2_fill_2 FILLER_54_2305 ();
 sg13g2_decap_8 FILLER_54_2320 ();
 sg13g2_decap_8 FILLER_54_2327 ();
 sg13g2_decap_8 FILLER_54_2334 ();
 sg13g2_decap_8 FILLER_54_2341 ();
 sg13g2_decap_8 FILLER_54_2348 ();
 sg13g2_decap_8 FILLER_54_2355 ();
 sg13g2_decap_8 FILLER_54_2362 ();
 sg13g2_decap_8 FILLER_54_2369 ();
 sg13g2_decap_8 FILLER_54_2376 ();
 sg13g2_decap_8 FILLER_54_2383 ();
 sg13g2_decap_8 FILLER_54_2390 ();
 sg13g2_decap_8 FILLER_54_2397 ();
 sg13g2_decap_8 FILLER_54_2404 ();
 sg13g2_decap_8 FILLER_54_2411 ();
 sg13g2_decap_8 FILLER_54_2418 ();
 sg13g2_decap_8 FILLER_54_2425 ();
 sg13g2_decap_8 FILLER_54_2432 ();
 sg13g2_decap_8 FILLER_54_2439 ();
 sg13g2_decap_8 FILLER_54_2446 ();
 sg13g2_decap_8 FILLER_54_2453 ();
 sg13g2_decap_8 FILLER_54_2460 ();
 sg13g2_decap_8 FILLER_54_2467 ();
 sg13g2_decap_8 FILLER_54_2474 ();
 sg13g2_decap_8 FILLER_54_2481 ();
 sg13g2_decap_8 FILLER_54_2488 ();
 sg13g2_decap_8 FILLER_54_2495 ();
 sg13g2_decap_8 FILLER_54_2502 ();
 sg13g2_decap_8 FILLER_54_2509 ();
 sg13g2_decap_8 FILLER_54_2516 ();
 sg13g2_decap_8 FILLER_54_2523 ();
 sg13g2_decap_8 FILLER_54_2530 ();
 sg13g2_decap_8 FILLER_54_2537 ();
 sg13g2_decap_8 FILLER_54_2544 ();
 sg13g2_decap_8 FILLER_54_2551 ();
 sg13g2_decap_8 FILLER_54_2558 ();
 sg13g2_decap_8 FILLER_54_2565 ();
 sg13g2_decap_8 FILLER_54_2572 ();
 sg13g2_decap_8 FILLER_54_2579 ();
 sg13g2_decap_8 FILLER_54_2586 ();
 sg13g2_decap_8 FILLER_54_2593 ();
 sg13g2_decap_8 FILLER_54_2600 ();
 sg13g2_decap_8 FILLER_54_2607 ();
 sg13g2_decap_8 FILLER_54_2614 ();
 sg13g2_decap_8 FILLER_54_2621 ();
 sg13g2_decap_8 FILLER_54_2628 ();
 sg13g2_decap_8 FILLER_54_2635 ();
 sg13g2_decap_8 FILLER_54_2642 ();
 sg13g2_decap_8 FILLER_54_2649 ();
 sg13g2_decap_8 FILLER_54_2656 ();
 sg13g2_decap_8 FILLER_54_2663 ();
 sg13g2_decap_4 FILLER_54_2670 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_140 ();
 sg13g2_decap_8 FILLER_55_147 ();
 sg13g2_decap_8 FILLER_55_154 ();
 sg13g2_decap_8 FILLER_55_161 ();
 sg13g2_decap_8 FILLER_55_168 ();
 sg13g2_decap_8 FILLER_55_175 ();
 sg13g2_decap_8 FILLER_55_182 ();
 sg13g2_decap_8 FILLER_55_189 ();
 sg13g2_decap_8 FILLER_55_196 ();
 sg13g2_decap_8 FILLER_55_203 ();
 sg13g2_decap_8 FILLER_55_210 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_decap_8 FILLER_55_224 ();
 sg13g2_decap_8 FILLER_55_231 ();
 sg13g2_decap_8 FILLER_55_238 ();
 sg13g2_decap_8 FILLER_55_245 ();
 sg13g2_decap_8 FILLER_55_252 ();
 sg13g2_decap_8 FILLER_55_259 ();
 sg13g2_decap_8 FILLER_55_266 ();
 sg13g2_decap_8 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_280 ();
 sg13g2_decap_8 FILLER_55_287 ();
 sg13g2_decap_8 FILLER_55_294 ();
 sg13g2_decap_8 FILLER_55_301 ();
 sg13g2_decap_8 FILLER_55_308 ();
 sg13g2_decap_8 FILLER_55_315 ();
 sg13g2_decap_8 FILLER_55_322 ();
 sg13g2_decap_8 FILLER_55_329 ();
 sg13g2_decap_8 FILLER_55_336 ();
 sg13g2_decap_8 FILLER_55_343 ();
 sg13g2_decap_8 FILLER_55_350 ();
 sg13g2_decap_8 FILLER_55_357 ();
 sg13g2_decap_8 FILLER_55_364 ();
 sg13g2_decap_8 FILLER_55_371 ();
 sg13g2_decap_8 FILLER_55_378 ();
 sg13g2_decap_8 FILLER_55_385 ();
 sg13g2_decap_8 FILLER_55_392 ();
 sg13g2_decap_8 FILLER_55_399 ();
 sg13g2_decap_8 FILLER_55_406 ();
 sg13g2_decap_8 FILLER_55_413 ();
 sg13g2_decap_8 FILLER_55_420 ();
 sg13g2_decap_8 FILLER_55_427 ();
 sg13g2_decap_8 FILLER_55_434 ();
 sg13g2_decap_8 FILLER_55_441 ();
 sg13g2_decap_8 FILLER_55_448 ();
 sg13g2_decap_8 FILLER_55_455 ();
 sg13g2_decap_4 FILLER_55_462 ();
 sg13g2_fill_1 FILLER_55_466 ();
 sg13g2_fill_2 FILLER_55_485 ();
 sg13g2_fill_2 FILLER_55_492 ();
 sg13g2_fill_1 FILLER_55_494 ();
 sg13g2_fill_2 FILLER_55_504 ();
 sg13g2_fill_1 FILLER_55_506 ();
 sg13g2_fill_1 FILLER_55_550 ();
 sg13g2_fill_2 FILLER_55_556 ();
 sg13g2_fill_1 FILLER_55_572 ();
 sg13g2_fill_2 FILLER_55_583 ();
 sg13g2_fill_1 FILLER_55_585 ();
 sg13g2_fill_1 FILLER_55_599 ();
 sg13g2_fill_2 FILLER_55_628 ();
 sg13g2_decap_4 FILLER_55_678 ();
 sg13g2_fill_2 FILLER_55_682 ();
 sg13g2_fill_2 FILLER_55_697 ();
 sg13g2_decap_4 FILLER_55_707 ();
 sg13g2_fill_2 FILLER_55_719 ();
 sg13g2_fill_1 FILLER_55_721 ();
 sg13g2_fill_2 FILLER_55_769 ();
 sg13g2_fill_2 FILLER_55_775 ();
 sg13g2_fill_1 FILLER_55_777 ();
 sg13g2_fill_1 FILLER_55_830 ();
 sg13g2_decap_4 FILLER_55_836 ();
 sg13g2_fill_2 FILLER_55_845 ();
 sg13g2_fill_2 FILLER_55_851 ();
 sg13g2_fill_2 FILLER_55_875 ();
 sg13g2_fill_2 FILLER_55_890 ();
 sg13g2_fill_1 FILLER_55_892 ();
 sg13g2_fill_2 FILLER_55_932 ();
 sg13g2_fill_1 FILLER_55_934 ();
 sg13g2_fill_2 FILLER_55_970 ();
 sg13g2_decap_8 FILLER_55_993 ();
 sg13g2_decap_4 FILLER_55_1000 ();
 sg13g2_fill_2 FILLER_55_1004 ();
 sg13g2_decap_8 FILLER_55_1010 ();
 sg13g2_fill_2 FILLER_55_1017 ();
 sg13g2_fill_2 FILLER_55_1054 ();
 sg13g2_fill_1 FILLER_55_1087 ();
 sg13g2_decap_8 FILLER_55_1093 ();
 sg13g2_fill_2 FILLER_55_1100 ();
 sg13g2_fill_1 FILLER_55_1102 ();
 sg13g2_fill_2 FILLER_55_1133 ();
 sg13g2_fill_1 FILLER_55_1135 ();
 sg13g2_fill_1 FILLER_55_1145 ();
 sg13g2_fill_2 FILLER_55_1156 ();
 sg13g2_fill_2 FILLER_55_1206 ();
 sg13g2_fill_1 FILLER_55_1208 ();
 sg13g2_fill_2 FILLER_55_1223 ();
 sg13g2_fill_1 FILLER_55_1225 ();
 sg13g2_fill_1 FILLER_55_1235 ();
 sg13g2_fill_2 FILLER_55_1302 ();
 sg13g2_fill_2 FILLER_55_1337 ();
 sg13g2_fill_1 FILLER_55_1361 ();
 sg13g2_fill_1 FILLER_55_1370 ();
 sg13g2_decap_8 FILLER_55_1379 ();
 sg13g2_fill_1 FILLER_55_1386 ();
 sg13g2_fill_2 FILLER_55_1391 ();
 sg13g2_fill_1 FILLER_55_1393 ();
 sg13g2_fill_1 FILLER_55_1399 ();
 sg13g2_fill_2 FILLER_55_1404 ();
 sg13g2_fill_1 FILLER_55_1406 ();
 sg13g2_decap_8 FILLER_55_1570 ();
 sg13g2_fill_1 FILLER_55_1577 ();
 sg13g2_fill_2 FILLER_55_1642 ();
 sg13g2_fill_1 FILLER_55_1644 ();
 sg13g2_decap_8 FILLER_55_1665 ();
 sg13g2_fill_1 FILLER_55_1672 ();
 sg13g2_fill_2 FILLER_55_1677 ();
 sg13g2_fill_2 FILLER_55_1699 ();
 sg13g2_fill_1 FILLER_55_1701 ();
 sg13g2_decap_4 FILLER_55_1710 ();
 sg13g2_fill_1 FILLER_55_1714 ();
 sg13g2_fill_2 FILLER_55_1724 ();
 sg13g2_fill_1 FILLER_55_1726 ();
 sg13g2_decap_4 FILLER_55_1748 ();
 sg13g2_fill_2 FILLER_55_1752 ();
 sg13g2_fill_1 FILLER_55_1759 ();
 sg13g2_fill_2 FILLER_55_1793 ();
 sg13g2_fill_1 FILLER_55_1857 ();
 sg13g2_fill_2 FILLER_55_1867 ();
 sg13g2_fill_1 FILLER_55_1873 ();
 sg13g2_fill_1 FILLER_55_1878 ();
 sg13g2_fill_2 FILLER_55_1889 ();
 sg13g2_fill_1 FILLER_55_1891 ();
 sg13g2_fill_2 FILLER_55_1923 ();
 sg13g2_decap_8 FILLER_55_1937 ();
 sg13g2_decap_4 FILLER_55_1944 ();
 sg13g2_fill_1 FILLER_55_1948 ();
 sg13g2_fill_2 FILLER_55_1963 ();
 sg13g2_fill_2 FILLER_55_2025 ();
 sg13g2_fill_1 FILLER_55_2070 ();
 sg13g2_fill_2 FILLER_55_2140 ();
 sg13g2_fill_1 FILLER_55_2142 ();
 sg13g2_fill_1 FILLER_55_2197 ();
 sg13g2_fill_2 FILLER_55_2258 ();
 sg13g2_decap_8 FILLER_55_2322 ();
 sg13g2_decap_8 FILLER_55_2329 ();
 sg13g2_decap_8 FILLER_55_2336 ();
 sg13g2_decap_8 FILLER_55_2343 ();
 sg13g2_decap_8 FILLER_55_2350 ();
 sg13g2_decap_8 FILLER_55_2357 ();
 sg13g2_decap_8 FILLER_55_2364 ();
 sg13g2_decap_8 FILLER_55_2371 ();
 sg13g2_decap_8 FILLER_55_2378 ();
 sg13g2_decap_8 FILLER_55_2385 ();
 sg13g2_decap_8 FILLER_55_2392 ();
 sg13g2_decap_8 FILLER_55_2399 ();
 sg13g2_decap_8 FILLER_55_2406 ();
 sg13g2_decap_8 FILLER_55_2413 ();
 sg13g2_decap_8 FILLER_55_2420 ();
 sg13g2_decap_8 FILLER_55_2427 ();
 sg13g2_decap_8 FILLER_55_2434 ();
 sg13g2_decap_8 FILLER_55_2441 ();
 sg13g2_decap_8 FILLER_55_2448 ();
 sg13g2_decap_8 FILLER_55_2455 ();
 sg13g2_decap_8 FILLER_55_2462 ();
 sg13g2_decap_8 FILLER_55_2469 ();
 sg13g2_decap_8 FILLER_55_2476 ();
 sg13g2_decap_8 FILLER_55_2483 ();
 sg13g2_decap_8 FILLER_55_2490 ();
 sg13g2_decap_8 FILLER_55_2497 ();
 sg13g2_decap_8 FILLER_55_2504 ();
 sg13g2_decap_8 FILLER_55_2511 ();
 sg13g2_decap_8 FILLER_55_2518 ();
 sg13g2_decap_8 FILLER_55_2525 ();
 sg13g2_decap_8 FILLER_55_2532 ();
 sg13g2_decap_8 FILLER_55_2539 ();
 sg13g2_decap_8 FILLER_55_2546 ();
 sg13g2_decap_8 FILLER_55_2553 ();
 sg13g2_decap_8 FILLER_55_2560 ();
 sg13g2_decap_8 FILLER_55_2567 ();
 sg13g2_decap_8 FILLER_55_2574 ();
 sg13g2_decap_8 FILLER_55_2581 ();
 sg13g2_decap_8 FILLER_55_2588 ();
 sg13g2_decap_8 FILLER_55_2595 ();
 sg13g2_decap_8 FILLER_55_2602 ();
 sg13g2_decap_8 FILLER_55_2609 ();
 sg13g2_decap_8 FILLER_55_2616 ();
 sg13g2_decap_8 FILLER_55_2623 ();
 sg13g2_decap_8 FILLER_55_2630 ();
 sg13g2_decap_8 FILLER_55_2637 ();
 sg13g2_decap_8 FILLER_55_2644 ();
 sg13g2_decap_8 FILLER_55_2651 ();
 sg13g2_decap_8 FILLER_55_2658 ();
 sg13g2_decap_8 FILLER_55_2665 ();
 sg13g2_fill_2 FILLER_55_2672 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_decap_8 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_154 ();
 sg13g2_decap_8 FILLER_56_161 ();
 sg13g2_decap_8 FILLER_56_168 ();
 sg13g2_decap_8 FILLER_56_175 ();
 sg13g2_decap_8 FILLER_56_182 ();
 sg13g2_decap_8 FILLER_56_189 ();
 sg13g2_decap_8 FILLER_56_196 ();
 sg13g2_decap_8 FILLER_56_203 ();
 sg13g2_decap_8 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_217 ();
 sg13g2_decap_8 FILLER_56_224 ();
 sg13g2_decap_8 FILLER_56_231 ();
 sg13g2_decap_8 FILLER_56_238 ();
 sg13g2_decap_8 FILLER_56_245 ();
 sg13g2_decap_8 FILLER_56_252 ();
 sg13g2_decap_8 FILLER_56_259 ();
 sg13g2_decap_8 FILLER_56_266 ();
 sg13g2_decap_8 FILLER_56_273 ();
 sg13g2_decap_8 FILLER_56_280 ();
 sg13g2_decap_8 FILLER_56_287 ();
 sg13g2_decap_8 FILLER_56_294 ();
 sg13g2_decap_8 FILLER_56_301 ();
 sg13g2_decap_8 FILLER_56_308 ();
 sg13g2_decap_8 FILLER_56_315 ();
 sg13g2_decap_8 FILLER_56_322 ();
 sg13g2_decap_8 FILLER_56_329 ();
 sg13g2_decap_8 FILLER_56_336 ();
 sg13g2_decap_8 FILLER_56_343 ();
 sg13g2_decap_8 FILLER_56_350 ();
 sg13g2_decap_8 FILLER_56_357 ();
 sg13g2_decap_8 FILLER_56_364 ();
 sg13g2_decap_8 FILLER_56_371 ();
 sg13g2_decap_8 FILLER_56_378 ();
 sg13g2_decap_8 FILLER_56_385 ();
 sg13g2_decap_8 FILLER_56_392 ();
 sg13g2_decap_8 FILLER_56_399 ();
 sg13g2_decap_8 FILLER_56_406 ();
 sg13g2_decap_8 FILLER_56_413 ();
 sg13g2_decap_8 FILLER_56_420 ();
 sg13g2_decap_8 FILLER_56_427 ();
 sg13g2_decap_8 FILLER_56_434 ();
 sg13g2_decap_8 FILLER_56_441 ();
 sg13g2_decap_8 FILLER_56_448 ();
 sg13g2_decap_8 FILLER_56_455 ();
 sg13g2_decap_4 FILLER_56_462 ();
 sg13g2_fill_1 FILLER_56_492 ();
 sg13g2_fill_1 FILLER_56_498 ();
 sg13g2_fill_2 FILLER_56_534 ();
 sg13g2_fill_1 FILLER_56_561 ();
 sg13g2_fill_1 FILLER_56_575 ();
 sg13g2_fill_1 FILLER_56_610 ();
 sg13g2_fill_2 FILLER_56_629 ();
 sg13g2_fill_1 FILLER_56_631 ();
 sg13g2_fill_1 FILLER_56_649 ();
 sg13g2_fill_1 FILLER_56_655 ();
 sg13g2_fill_1 FILLER_56_682 ();
 sg13g2_fill_1 FILLER_56_714 ();
 sg13g2_fill_2 FILLER_56_729 ();
 sg13g2_fill_1 FILLER_56_731 ();
 sg13g2_fill_2 FILLER_56_741 ();
 sg13g2_fill_1 FILLER_56_743 ();
 sg13g2_fill_1 FILLER_56_748 ();
 sg13g2_fill_1 FILLER_56_758 ();
 sg13g2_fill_2 FILLER_56_763 ();
 sg13g2_decap_4 FILLER_56_779 ();
 sg13g2_fill_1 FILLER_56_783 ();
 sg13g2_fill_2 FILLER_56_788 ();
 sg13g2_fill_1 FILLER_56_794 ();
 sg13g2_fill_2 FILLER_56_822 ();
 sg13g2_fill_2 FILLER_56_834 ();
 sg13g2_fill_2 FILLER_56_862 ();
 sg13g2_fill_1 FILLER_56_876 ();
 sg13g2_fill_2 FILLER_56_891 ();
 sg13g2_fill_1 FILLER_56_893 ();
 sg13g2_fill_1 FILLER_56_913 ();
 sg13g2_fill_2 FILLER_56_936 ();
 sg13g2_fill_1 FILLER_56_938 ();
 sg13g2_fill_2 FILLER_56_944 ();
 sg13g2_fill_1 FILLER_56_946 ();
 sg13g2_fill_1 FILLER_56_982 ();
 sg13g2_decap_4 FILLER_56_987 ();
 sg13g2_fill_1 FILLER_56_991 ();
 sg13g2_decap_4 FILLER_56_1044 ();
 sg13g2_fill_2 FILLER_56_1058 ();
 sg13g2_fill_1 FILLER_56_1060 ();
 sg13g2_fill_2 FILLER_56_1065 ();
 sg13g2_fill_2 FILLER_56_1100 ();
 sg13g2_fill_1 FILLER_56_1133 ();
 sg13g2_decap_4 FILLER_56_1139 ();
 sg13g2_fill_1 FILLER_56_1199 ();
 sg13g2_fill_2 FILLER_56_1234 ();
 sg13g2_fill_1 FILLER_56_1236 ();
 sg13g2_fill_1 FILLER_56_1261 ();
 sg13g2_fill_2 FILLER_56_1273 ();
 sg13g2_fill_2 FILLER_56_1284 ();
 sg13g2_fill_2 FILLER_56_1358 ();
 sg13g2_fill_1 FILLER_56_1368 ();
 sg13g2_fill_2 FILLER_56_1435 ();
 sg13g2_fill_1 FILLER_56_1437 ();
 sg13g2_fill_1 FILLER_56_1447 ();
 sg13g2_fill_2 FILLER_56_1453 ();
 sg13g2_fill_1 FILLER_56_1455 ();
 sg13g2_fill_2 FILLER_56_1465 ();
 sg13g2_fill_2 FILLER_56_1490 ();
 sg13g2_fill_2 FILLER_56_1514 ();
 sg13g2_fill_2 FILLER_56_1551 ();
 sg13g2_fill_1 FILLER_56_1553 ();
 sg13g2_fill_2 FILLER_56_1580 ();
 sg13g2_decap_8 FILLER_56_1590 ();
 sg13g2_decap_8 FILLER_56_1617 ();
 sg13g2_fill_2 FILLER_56_1684 ();
 sg13g2_fill_2 FILLER_56_1700 ();
 sg13g2_fill_1 FILLER_56_1702 ();
 sg13g2_fill_2 FILLER_56_1760 ();
 sg13g2_fill_1 FILLER_56_1762 ();
 sg13g2_decap_4 FILLER_56_1767 ();
 sg13g2_fill_1 FILLER_56_1776 ();
 sg13g2_fill_1 FILLER_56_1803 ();
 sg13g2_fill_2 FILLER_56_1825 ();
 sg13g2_decap_4 FILLER_56_1878 ();
 sg13g2_fill_2 FILLER_56_1882 ();
 sg13g2_decap_4 FILLER_56_1897 ();
 sg13g2_fill_2 FILLER_56_1901 ();
 sg13g2_decap_4 FILLER_56_1907 ();
 sg13g2_decap_4 FILLER_56_1942 ();
 sg13g2_decap_8 FILLER_56_2025 ();
 sg13g2_fill_2 FILLER_56_2032 ();
 sg13g2_fill_1 FILLER_56_2040 ();
 sg13g2_fill_1 FILLER_56_2046 ();
 sg13g2_fill_1 FILLER_56_2051 ();
 sg13g2_decap_4 FILLER_56_2105 ();
 sg13g2_fill_1 FILLER_56_2109 ();
 sg13g2_fill_2 FILLER_56_2136 ();
 sg13g2_fill_1 FILLER_56_2138 ();
 sg13g2_fill_2 FILLER_56_2180 ();
 sg13g2_fill_1 FILLER_56_2182 ();
 sg13g2_decap_4 FILLER_56_2191 ();
 sg13g2_fill_2 FILLER_56_2195 ();
 sg13g2_fill_1 FILLER_56_2207 ();
 sg13g2_fill_2 FILLER_56_2232 ();
 sg13g2_fill_2 FILLER_56_2247 ();
 sg13g2_fill_2 FILLER_56_2305 ();
 sg13g2_fill_1 FILLER_56_2307 ();
 sg13g2_decap_8 FILLER_56_2317 ();
 sg13g2_decap_8 FILLER_56_2324 ();
 sg13g2_decap_8 FILLER_56_2331 ();
 sg13g2_decap_8 FILLER_56_2338 ();
 sg13g2_decap_8 FILLER_56_2345 ();
 sg13g2_decap_8 FILLER_56_2352 ();
 sg13g2_decap_8 FILLER_56_2359 ();
 sg13g2_decap_8 FILLER_56_2366 ();
 sg13g2_decap_8 FILLER_56_2373 ();
 sg13g2_decap_8 FILLER_56_2380 ();
 sg13g2_decap_8 FILLER_56_2387 ();
 sg13g2_decap_8 FILLER_56_2394 ();
 sg13g2_decap_8 FILLER_56_2401 ();
 sg13g2_decap_8 FILLER_56_2408 ();
 sg13g2_decap_8 FILLER_56_2415 ();
 sg13g2_decap_8 FILLER_56_2422 ();
 sg13g2_decap_8 FILLER_56_2429 ();
 sg13g2_decap_8 FILLER_56_2436 ();
 sg13g2_decap_8 FILLER_56_2443 ();
 sg13g2_decap_8 FILLER_56_2450 ();
 sg13g2_decap_8 FILLER_56_2457 ();
 sg13g2_decap_8 FILLER_56_2464 ();
 sg13g2_decap_8 FILLER_56_2471 ();
 sg13g2_decap_8 FILLER_56_2478 ();
 sg13g2_decap_8 FILLER_56_2485 ();
 sg13g2_decap_8 FILLER_56_2492 ();
 sg13g2_decap_8 FILLER_56_2499 ();
 sg13g2_decap_8 FILLER_56_2506 ();
 sg13g2_decap_8 FILLER_56_2513 ();
 sg13g2_decap_8 FILLER_56_2520 ();
 sg13g2_decap_8 FILLER_56_2527 ();
 sg13g2_decap_8 FILLER_56_2534 ();
 sg13g2_decap_8 FILLER_56_2541 ();
 sg13g2_decap_8 FILLER_56_2548 ();
 sg13g2_decap_8 FILLER_56_2555 ();
 sg13g2_decap_8 FILLER_56_2562 ();
 sg13g2_decap_8 FILLER_56_2569 ();
 sg13g2_decap_8 FILLER_56_2576 ();
 sg13g2_decap_8 FILLER_56_2583 ();
 sg13g2_decap_8 FILLER_56_2590 ();
 sg13g2_decap_8 FILLER_56_2597 ();
 sg13g2_decap_8 FILLER_56_2604 ();
 sg13g2_decap_8 FILLER_56_2611 ();
 sg13g2_decap_8 FILLER_56_2618 ();
 sg13g2_decap_8 FILLER_56_2625 ();
 sg13g2_decap_8 FILLER_56_2632 ();
 sg13g2_decap_8 FILLER_56_2639 ();
 sg13g2_decap_8 FILLER_56_2646 ();
 sg13g2_decap_8 FILLER_56_2653 ();
 sg13g2_decap_8 FILLER_56_2660 ();
 sg13g2_decap_8 FILLER_56_2667 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_8 FILLER_57_168 ();
 sg13g2_decap_8 FILLER_57_175 ();
 sg13g2_decap_8 FILLER_57_182 ();
 sg13g2_decap_8 FILLER_57_189 ();
 sg13g2_decap_8 FILLER_57_196 ();
 sg13g2_decap_8 FILLER_57_203 ();
 sg13g2_decap_8 FILLER_57_210 ();
 sg13g2_decap_8 FILLER_57_217 ();
 sg13g2_decap_8 FILLER_57_224 ();
 sg13g2_decap_8 FILLER_57_231 ();
 sg13g2_decap_8 FILLER_57_238 ();
 sg13g2_decap_8 FILLER_57_245 ();
 sg13g2_decap_8 FILLER_57_252 ();
 sg13g2_decap_8 FILLER_57_259 ();
 sg13g2_decap_8 FILLER_57_266 ();
 sg13g2_decap_8 FILLER_57_273 ();
 sg13g2_decap_8 FILLER_57_280 ();
 sg13g2_decap_8 FILLER_57_287 ();
 sg13g2_decap_8 FILLER_57_294 ();
 sg13g2_decap_8 FILLER_57_301 ();
 sg13g2_decap_8 FILLER_57_308 ();
 sg13g2_decap_8 FILLER_57_315 ();
 sg13g2_decap_8 FILLER_57_322 ();
 sg13g2_decap_8 FILLER_57_329 ();
 sg13g2_decap_8 FILLER_57_336 ();
 sg13g2_decap_8 FILLER_57_343 ();
 sg13g2_decap_8 FILLER_57_350 ();
 sg13g2_decap_8 FILLER_57_357 ();
 sg13g2_decap_8 FILLER_57_364 ();
 sg13g2_decap_8 FILLER_57_371 ();
 sg13g2_decap_8 FILLER_57_378 ();
 sg13g2_decap_8 FILLER_57_385 ();
 sg13g2_decap_8 FILLER_57_392 ();
 sg13g2_decap_8 FILLER_57_399 ();
 sg13g2_decap_8 FILLER_57_406 ();
 sg13g2_decap_8 FILLER_57_413 ();
 sg13g2_decap_8 FILLER_57_420 ();
 sg13g2_decap_8 FILLER_57_427 ();
 sg13g2_decap_8 FILLER_57_434 ();
 sg13g2_decap_8 FILLER_57_441 ();
 sg13g2_decap_8 FILLER_57_448 ();
 sg13g2_decap_8 FILLER_57_455 ();
 sg13g2_fill_2 FILLER_57_462 ();
 sg13g2_fill_1 FILLER_57_464 ();
 sg13g2_fill_2 FILLER_57_491 ();
 sg13g2_fill_1 FILLER_57_493 ();
 sg13g2_fill_2 FILLER_57_521 ();
 sg13g2_fill_1 FILLER_57_631 ();
 sg13g2_fill_1 FILLER_57_637 ();
 sg13g2_decap_4 FILLER_57_651 ();
 sg13g2_fill_1 FILLER_57_655 ();
 sg13g2_decap_4 FILLER_57_687 ();
 sg13g2_fill_2 FILLER_57_691 ();
 sg13g2_decap_8 FILLER_57_706 ();
 sg13g2_fill_1 FILLER_57_713 ();
 sg13g2_fill_1 FILLER_57_717 ();
 sg13g2_fill_2 FILLER_57_749 ();
 sg13g2_fill_1 FILLER_57_756 ();
 sg13g2_decap_4 FILLER_57_766 ();
 sg13g2_fill_1 FILLER_57_770 ();
 sg13g2_decap_4 FILLER_57_786 ();
 sg13g2_fill_1 FILLER_57_790 ();
 sg13g2_fill_2 FILLER_57_817 ();
 sg13g2_fill_1 FILLER_57_819 ();
 sg13g2_decap_4 FILLER_57_842 ();
 sg13g2_fill_1 FILLER_57_846 ();
 sg13g2_fill_1 FILLER_57_856 ();
 sg13g2_fill_1 FILLER_57_902 ();
 sg13g2_decap_8 FILLER_57_947 ();
 sg13g2_decap_4 FILLER_57_954 ();
 sg13g2_fill_2 FILLER_57_985 ();
 sg13g2_fill_1 FILLER_57_987 ();
 sg13g2_fill_2 FILLER_57_996 ();
 sg13g2_fill_1 FILLER_57_998 ();
 sg13g2_fill_1 FILLER_57_1016 ();
 sg13g2_fill_2 FILLER_57_1029 ();
 sg13g2_fill_1 FILLER_57_1031 ();
 sg13g2_fill_2 FILLER_57_1084 ();
 sg13g2_fill_1 FILLER_57_1096 ();
 sg13g2_fill_2 FILLER_57_1102 ();
 sg13g2_fill_1 FILLER_57_1104 ();
 sg13g2_fill_1 FILLER_57_1120 ();
 sg13g2_decap_4 FILLER_57_1130 ();
 sg13g2_fill_1 FILLER_57_1134 ();
 sg13g2_fill_1 FILLER_57_1140 ();
 sg13g2_decap_4 FILLER_57_1151 ();
 sg13g2_fill_2 FILLER_57_1174 ();
 sg13g2_fill_2 FILLER_57_1184 ();
 sg13g2_fill_2 FILLER_57_1204 ();
 sg13g2_fill_2 FILLER_57_1211 ();
 sg13g2_fill_2 FILLER_57_1227 ();
 sg13g2_fill_1 FILLER_57_1229 ();
 sg13g2_fill_2 FILLER_57_1235 ();
 sg13g2_fill_1 FILLER_57_1237 ();
 sg13g2_fill_2 FILLER_57_1309 ();
 sg13g2_fill_1 FILLER_57_1311 ();
 sg13g2_fill_2 FILLER_57_1316 ();
 sg13g2_fill_2 FILLER_57_1327 ();
 sg13g2_fill_1 FILLER_57_1343 ();
 sg13g2_decap_8 FILLER_57_1362 ();
 sg13g2_decap_8 FILLER_57_1369 ();
 sg13g2_fill_1 FILLER_57_1376 ();
 sg13g2_fill_2 FILLER_57_1393 ();
 sg13g2_decap_8 FILLER_57_1399 ();
 sg13g2_fill_2 FILLER_57_1406 ();
 sg13g2_fill_1 FILLER_57_1494 ();
 sg13g2_fill_2 FILLER_57_1539 ();
 sg13g2_fill_2 FILLER_57_1555 ();
 sg13g2_fill_2 FILLER_57_1565 ();
 sg13g2_decap_4 FILLER_57_1584 ();
 sg13g2_fill_2 FILLER_57_1588 ();
 sg13g2_decap_8 FILLER_57_1610 ();
 sg13g2_decap_4 FILLER_57_1617 ();
 sg13g2_fill_2 FILLER_57_1621 ();
 sg13g2_decap_8 FILLER_57_1627 ();
 sg13g2_fill_1 FILLER_57_1634 ();
 sg13g2_fill_2 FILLER_57_1639 ();
 sg13g2_decap_8 FILLER_57_1665 ();
 sg13g2_decap_4 FILLER_57_1708 ();
 sg13g2_fill_1 FILLER_57_1712 ();
 sg13g2_fill_1 FILLER_57_1730 ();
 sg13g2_fill_2 FILLER_57_1749 ();
 sg13g2_fill_1 FILLER_57_1751 ();
 sg13g2_fill_2 FILLER_57_1792 ();
 sg13g2_fill_1 FILLER_57_1895 ();
 sg13g2_decap_4 FILLER_57_1912 ();
 sg13g2_fill_2 FILLER_57_1916 ();
 sg13g2_fill_1 FILLER_57_1927 ();
 sg13g2_decap_8 FILLER_57_1949 ();
 sg13g2_decap_4 FILLER_57_1965 ();
 sg13g2_decap_4 FILLER_57_2000 ();
 sg13g2_decap_4 FILLER_57_2008 ();
 sg13g2_fill_1 FILLER_57_2012 ();
 sg13g2_decap_8 FILLER_57_2023 ();
 sg13g2_decap_4 FILLER_57_2040 ();
 sg13g2_fill_2 FILLER_57_2044 ();
 sg13g2_fill_2 FILLER_57_2050 ();
 sg13g2_decap_4 FILLER_57_2057 ();
 sg13g2_decap_8 FILLER_57_2065 ();
 sg13g2_fill_1 FILLER_57_2072 ();
 sg13g2_fill_1 FILLER_57_2086 ();
 sg13g2_decap_4 FILLER_57_2113 ();
 sg13g2_fill_1 FILLER_57_2117 ();
 sg13g2_fill_2 FILLER_57_2173 ();
 sg13g2_fill_1 FILLER_57_2175 ();
 sg13g2_fill_1 FILLER_57_2185 ();
 sg13g2_fill_2 FILLER_57_2190 ();
 sg13g2_fill_2 FILLER_57_2197 ();
 sg13g2_fill_1 FILLER_57_2199 ();
 sg13g2_fill_2 FILLER_57_2213 ();
 sg13g2_fill_1 FILLER_57_2215 ();
 sg13g2_fill_1 FILLER_57_2234 ();
 sg13g2_fill_2 FILLER_57_2239 ();
 sg13g2_decap_4 FILLER_57_2281 ();
 sg13g2_decap_8 FILLER_57_2320 ();
 sg13g2_decap_8 FILLER_57_2327 ();
 sg13g2_decap_8 FILLER_57_2334 ();
 sg13g2_decap_8 FILLER_57_2341 ();
 sg13g2_decap_8 FILLER_57_2348 ();
 sg13g2_decap_8 FILLER_57_2355 ();
 sg13g2_decap_8 FILLER_57_2362 ();
 sg13g2_decap_8 FILLER_57_2369 ();
 sg13g2_decap_8 FILLER_57_2376 ();
 sg13g2_decap_8 FILLER_57_2383 ();
 sg13g2_decap_8 FILLER_57_2390 ();
 sg13g2_decap_8 FILLER_57_2397 ();
 sg13g2_decap_8 FILLER_57_2404 ();
 sg13g2_decap_8 FILLER_57_2411 ();
 sg13g2_decap_8 FILLER_57_2418 ();
 sg13g2_decap_8 FILLER_57_2425 ();
 sg13g2_decap_8 FILLER_57_2432 ();
 sg13g2_decap_8 FILLER_57_2439 ();
 sg13g2_decap_8 FILLER_57_2446 ();
 sg13g2_decap_8 FILLER_57_2453 ();
 sg13g2_decap_8 FILLER_57_2460 ();
 sg13g2_decap_8 FILLER_57_2467 ();
 sg13g2_decap_8 FILLER_57_2474 ();
 sg13g2_decap_8 FILLER_57_2481 ();
 sg13g2_decap_8 FILLER_57_2488 ();
 sg13g2_decap_8 FILLER_57_2495 ();
 sg13g2_decap_8 FILLER_57_2502 ();
 sg13g2_decap_8 FILLER_57_2509 ();
 sg13g2_decap_8 FILLER_57_2516 ();
 sg13g2_decap_8 FILLER_57_2523 ();
 sg13g2_decap_8 FILLER_57_2530 ();
 sg13g2_decap_8 FILLER_57_2537 ();
 sg13g2_decap_8 FILLER_57_2544 ();
 sg13g2_decap_8 FILLER_57_2551 ();
 sg13g2_decap_8 FILLER_57_2558 ();
 sg13g2_decap_8 FILLER_57_2565 ();
 sg13g2_decap_8 FILLER_57_2572 ();
 sg13g2_decap_8 FILLER_57_2579 ();
 sg13g2_decap_8 FILLER_57_2586 ();
 sg13g2_decap_8 FILLER_57_2593 ();
 sg13g2_decap_8 FILLER_57_2600 ();
 sg13g2_decap_8 FILLER_57_2607 ();
 sg13g2_decap_8 FILLER_57_2614 ();
 sg13g2_decap_8 FILLER_57_2621 ();
 sg13g2_decap_8 FILLER_57_2628 ();
 sg13g2_decap_8 FILLER_57_2635 ();
 sg13g2_decap_8 FILLER_57_2642 ();
 sg13g2_decap_8 FILLER_57_2649 ();
 sg13g2_decap_8 FILLER_57_2656 ();
 sg13g2_decap_8 FILLER_57_2663 ();
 sg13g2_decap_4 FILLER_57_2670 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_140 ();
 sg13g2_decap_8 FILLER_58_147 ();
 sg13g2_decap_8 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_decap_8 FILLER_58_182 ();
 sg13g2_decap_8 FILLER_58_189 ();
 sg13g2_decap_8 FILLER_58_196 ();
 sg13g2_decap_8 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_210 ();
 sg13g2_decap_8 FILLER_58_217 ();
 sg13g2_decap_8 FILLER_58_224 ();
 sg13g2_decap_8 FILLER_58_231 ();
 sg13g2_decap_8 FILLER_58_238 ();
 sg13g2_decap_8 FILLER_58_245 ();
 sg13g2_decap_8 FILLER_58_252 ();
 sg13g2_decap_8 FILLER_58_259 ();
 sg13g2_decap_8 FILLER_58_266 ();
 sg13g2_decap_8 FILLER_58_273 ();
 sg13g2_decap_8 FILLER_58_280 ();
 sg13g2_decap_8 FILLER_58_287 ();
 sg13g2_decap_8 FILLER_58_294 ();
 sg13g2_decap_8 FILLER_58_301 ();
 sg13g2_decap_8 FILLER_58_308 ();
 sg13g2_decap_8 FILLER_58_315 ();
 sg13g2_decap_8 FILLER_58_322 ();
 sg13g2_decap_8 FILLER_58_329 ();
 sg13g2_decap_8 FILLER_58_336 ();
 sg13g2_decap_8 FILLER_58_343 ();
 sg13g2_decap_8 FILLER_58_350 ();
 sg13g2_decap_8 FILLER_58_357 ();
 sg13g2_decap_8 FILLER_58_364 ();
 sg13g2_decap_8 FILLER_58_371 ();
 sg13g2_decap_8 FILLER_58_378 ();
 sg13g2_decap_8 FILLER_58_385 ();
 sg13g2_decap_8 FILLER_58_392 ();
 sg13g2_decap_8 FILLER_58_399 ();
 sg13g2_decap_8 FILLER_58_406 ();
 sg13g2_decap_8 FILLER_58_413 ();
 sg13g2_decap_8 FILLER_58_420 ();
 sg13g2_decap_8 FILLER_58_427 ();
 sg13g2_decap_8 FILLER_58_434 ();
 sg13g2_decap_8 FILLER_58_441 ();
 sg13g2_decap_8 FILLER_58_448 ();
 sg13g2_decap_8 FILLER_58_455 ();
 sg13g2_decap_4 FILLER_58_462 ();
 sg13g2_fill_2 FILLER_58_501 ();
 sg13g2_fill_1 FILLER_58_503 ();
 sg13g2_fill_2 FILLER_58_508 ();
 sg13g2_fill_2 FILLER_58_536 ();
 sg13g2_decap_8 FILLER_58_573 ();
 sg13g2_fill_2 FILLER_58_580 ();
 sg13g2_fill_1 FILLER_58_582 ();
 sg13g2_decap_8 FILLER_58_587 ();
 sg13g2_fill_1 FILLER_58_594 ();
 sg13g2_decap_4 FILLER_58_621 ();
 sg13g2_fill_2 FILLER_58_625 ();
 sg13g2_decap_4 FILLER_58_632 ();
 sg13g2_fill_2 FILLER_58_650 ();
 sg13g2_fill_1 FILLER_58_657 ();
 sg13g2_fill_1 FILLER_58_662 ();
 sg13g2_decap_8 FILLER_58_720 ();
 sg13g2_fill_2 FILLER_58_727 ();
 sg13g2_fill_2 FILLER_58_733 ();
 sg13g2_fill_2 FILLER_58_796 ();
 sg13g2_fill_1 FILLER_58_798 ();
 sg13g2_fill_1 FILLER_58_806 ();
 sg13g2_fill_1 FILLER_58_811 ();
 sg13g2_fill_2 FILLER_58_822 ();
 sg13g2_fill_2 FILLER_58_856 ();
 sg13g2_fill_1 FILLER_58_863 ();
 sg13g2_decap_4 FILLER_58_876 ();
 sg13g2_decap_8 FILLER_58_919 ();
 sg13g2_decap_4 FILLER_58_926 ();
 sg13g2_fill_2 FILLER_58_930 ();
 sg13g2_decap_4 FILLER_58_936 ();
 sg13g2_fill_2 FILLER_58_940 ();
 sg13g2_fill_2 FILLER_58_998 ();
 sg13g2_fill_2 FILLER_58_1075 ();
 sg13g2_fill_1 FILLER_58_1077 ();
 sg13g2_fill_1 FILLER_58_1095 ();
 sg13g2_fill_2 FILLER_58_1101 ();
 sg13g2_fill_1 FILLER_58_1107 ();
 sg13g2_fill_2 FILLER_58_1112 ();
 sg13g2_fill_2 FILLER_58_1148 ();
 sg13g2_fill_1 FILLER_58_1176 ();
 sg13g2_fill_2 FILLER_58_1230 ();
 sg13g2_fill_2 FILLER_58_1241 ();
 sg13g2_fill_1 FILLER_58_1248 ();
 sg13g2_fill_2 FILLER_58_1271 ();
 sg13g2_fill_2 FILLER_58_1301 ();
 sg13g2_fill_1 FILLER_58_1311 ();
 sg13g2_fill_1 FILLER_58_1320 ();
 sg13g2_fill_1 FILLER_58_1382 ();
 sg13g2_fill_2 FILLER_58_1387 ();
 sg13g2_decap_8 FILLER_58_1392 ();
 sg13g2_decap_4 FILLER_58_1399 ();
 sg13g2_fill_1 FILLER_58_1403 ();
 sg13g2_fill_2 FILLER_58_1430 ();
 sg13g2_fill_1 FILLER_58_1432 ();
 sg13g2_fill_2 FILLER_58_1441 ();
 sg13g2_fill_1 FILLER_58_1443 ();
 sg13g2_fill_1 FILLER_58_1449 ();
 sg13g2_fill_1 FILLER_58_1459 ();
 sg13g2_fill_1 FILLER_58_1479 ();
 sg13g2_fill_2 FILLER_58_1494 ();
 sg13g2_fill_2 FILLER_58_1505 ();
 sg13g2_fill_1 FILLER_58_1507 ();
 sg13g2_fill_2 FILLER_58_1525 ();
 sg13g2_fill_1 FILLER_58_1527 ();
 sg13g2_fill_2 FILLER_58_1548 ();
 sg13g2_decap_8 FILLER_58_1614 ();
 sg13g2_decap_4 FILLER_58_1673 ();
 sg13g2_fill_1 FILLER_58_1708 ();
 sg13g2_decap_4 FILLER_58_1735 ();
 sg13g2_fill_2 FILLER_58_1743 ();
 sg13g2_fill_2 FILLER_58_1750 ();
 sg13g2_fill_1 FILLER_58_1752 ();
 sg13g2_fill_1 FILLER_58_1775 ();
 sg13g2_fill_2 FILLER_58_1819 ();
 sg13g2_fill_1 FILLER_58_1821 ();
 sg13g2_fill_2 FILLER_58_1826 ();
 sg13g2_fill_1 FILLER_58_1846 ();
 sg13g2_fill_2 FILLER_58_1857 ();
 sg13g2_decap_4 FILLER_58_1877 ();
 sg13g2_fill_2 FILLER_58_1881 ();
 sg13g2_decap_4 FILLER_58_1934 ();
 sg13g2_fill_2 FILLER_58_1938 ();
 sg13g2_fill_2 FILLER_58_1983 ();
 sg13g2_fill_1 FILLER_58_1985 ();
 sg13g2_fill_2 FILLER_58_2022 ();
 sg13g2_fill_1 FILLER_58_2029 ();
 sg13g2_fill_1 FILLER_58_2034 ();
 sg13g2_fill_2 FILLER_58_2084 ();
 sg13g2_fill_1 FILLER_58_2153 ();
 sg13g2_fill_1 FILLER_58_2262 ();
 sg13g2_decap_4 FILLER_58_2297 ();
 sg13g2_fill_2 FILLER_58_2301 ();
 sg13g2_decap_8 FILLER_58_2316 ();
 sg13g2_decap_8 FILLER_58_2323 ();
 sg13g2_decap_8 FILLER_58_2330 ();
 sg13g2_decap_8 FILLER_58_2337 ();
 sg13g2_decap_8 FILLER_58_2344 ();
 sg13g2_decap_8 FILLER_58_2351 ();
 sg13g2_decap_8 FILLER_58_2358 ();
 sg13g2_decap_8 FILLER_58_2365 ();
 sg13g2_decap_8 FILLER_58_2372 ();
 sg13g2_decap_8 FILLER_58_2379 ();
 sg13g2_decap_8 FILLER_58_2386 ();
 sg13g2_decap_8 FILLER_58_2393 ();
 sg13g2_decap_8 FILLER_58_2400 ();
 sg13g2_decap_8 FILLER_58_2407 ();
 sg13g2_decap_8 FILLER_58_2414 ();
 sg13g2_decap_8 FILLER_58_2421 ();
 sg13g2_decap_8 FILLER_58_2428 ();
 sg13g2_decap_8 FILLER_58_2435 ();
 sg13g2_decap_8 FILLER_58_2442 ();
 sg13g2_decap_8 FILLER_58_2449 ();
 sg13g2_decap_8 FILLER_58_2456 ();
 sg13g2_decap_8 FILLER_58_2463 ();
 sg13g2_decap_8 FILLER_58_2470 ();
 sg13g2_decap_8 FILLER_58_2477 ();
 sg13g2_decap_8 FILLER_58_2484 ();
 sg13g2_decap_8 FILLER_58_2491 ();
 sg13g2_decap_8 FILLER_58_2498 ();
 sg13g2_decap_8 FILLER_58_2505 ();
 sg13g2_decap_8 FILLER_58_2512 ();
 sg13g2_decap_8 FILLER_58_2519 ();
 sg13g2_decap_8 FILLER_58_2526 ();
 sg13g2_decap_8 FILLER_58_2533 ();
 sg13g2_decap_8 FILLER_58_2540 ();
 sg13g2_decap_8 FILLER_58_2547 ();
 sg13g2_decap_8 FILLER_58_2554 ();
 sg13g2_decap_8 FILLER_58_2561 ();
 sg13g2_decap_8 FILLER_58_2568 ();
 sg13g2_decap_8 FILLER_58_2575 ();
 sg13g2_decap_8 FILLER_58_2582 ();
 sg13g2_decap_8 FILLER_58_2589 ();
 sg13g2_decap_8 FILLER_58_2596 ();
 sg13g2_decap_8 FILLER_58_2603 ();
 sg13g2_decap_8 FILLER_58_2610 ();
 sg13g2_decap_8 FILLER_58_2617 ();
 sg13g2_decap_8 FILLER_58_2624 ();
 sg13g2_decap_8 FILLER_58_2631 ();
 sg13g2_decap_8 FILLER_58_2638 ();
 sg13g2_decap_8 FILLER_58_2645 ();
 sg13g2_decap_8 FILLER_58_2652 ();
 sg13g2_decap_8 FILLER_58_2659 ();
 sg13g2_decap_8 FILLER_58_2666 ();
 sg13g2_fill_1 FILLER_58_2673 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_decap_8 FILLER_59_140 ();
 sg13g2_decap_8 FILLER_59_147 ();
 sg13g2_decap_8 FILLER_59_154 ();
 sg13g2_decap_8 FILLER_59_161 ();
 sg13g2_decap_8 FILLER_59_168 ();
 sg13g2_decap_8 FILLER_59_175 ();
 sg13g2_decap_8 FILLER_59_182 ();
 sg13g2_decap_8 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_196 ();
 sg13g2_decap_8 FILLER_59_203 ();
 sg13g2_decap_8 FILLER_59_210 ();
 sg13g2_decap_8 FILLER_59_217 ();
 sg13g2_decap_8 FILLER_59_224 ();
 sg13g2_decap_8 FILLER_59_231 ();
 sg13g2_decap_8 FILLER_59_238 ();
 sg13g2_decap_8 FILLER_59_245 ();
 sg13g2_decap_8 FILLER_59_252 ();
 sg13g2_decap_8 FILLER_59_259 ();
 sg13g2_decap_8 FILLER_59_266 ();
 sg13g2_decap_8 FILLER_59_273 ();
 sg13g2_decap_8 FILLER_59_280 ();
 sg13g2_decap_8 FILLER_59_287 ();
 sg13g2_decap_8 FILLER_59_294 ();
 sg13g2_decap_8 FILLER_59_301 ();
 sg13g2_decap_8 FILLER_59_308 ();
 sg13g2_decap_8 FILLER_59_315 ();
 sg13g2_decap_8 FILLER_59_322 ();
 sg13g2_decap_8 FILLER_59_329 ();
 sg13g2_decap_8 FILLER_59_336 ();
 sg13g2_decap_8 FILLER_59_343 ();
 sg13g2_decap_8 FILLER_59_350 ();
 sg13g2_decap_8 FILLER_59_357 ();
 sg13g2_decap_8 FILLER_59_364 ();
 sg13g2_decap_8 FILLER_59_371 ();
 sg13g2_decap_8 FILLER_59_378 ();
 sg13g2_decap_8 FILLER_59_385 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_decap_8 FILLER_59_399 ();
 sg13g2_decap_8 FILLER_59_406 ();
 sg13g2_decap_8 FILLER_59_413 ();
 sg13g2_decap_8 FILLER_59_420 ();
 sg13g2_decap_8 FILLER_59_427 ();
 sg13g2_decap_8 FILLER_59_434 ();
 sg13g2_decap_8 FILLER_59_441 ();
 sg13g2_decap_8 FILLER_59_448 ();
 sg13g2_fill_2 FILLER_59_455 ();
 sg13g2_fill_2 FILLER_59_528 ();
 sg13g2_fill_1 FILLER_59_539 ();
 sg13g2_fill_2 FILLER_59_549 ();
 sg13g2_fill_1 FILLER_59_551 ();
 sg13g2_fill_2 FILLER_59_597 ();
 sg13g2_fill_2 FILLER_59_604 ();
 sg13g2_fill_2 FILLER_59_610 ();
 sg13g2_fill_1 FILLER_59_620 ();
 sg13g2_decap_8 FILLER_59_634 ();
 sg13g2_fill_1 FILLER_59_641 ();
 sg13g2_decap_8 FILLER_59_652 ();
 sg13g2_fill_2 FILLER_59_659 ();
 sg13g2_fill_1 FILLER_59_661 ();
 sg13g2_fill_1 FILLER_59_671 ();
 sg13g2_decap_4 FILLER_59_676 ();
 sg13g2_fill_1 FILLER_59_680 ();
 sg13g2_decap_8 FILLER_59_684 ();
 sg13g2_fill_2 FILLER_59_691 ();
 sg13g2_fill_1 FILLER_59_693 ();
 sg13g2_fill_1 FILLER_59_753 ();
 sg13g2_fill_2 FILLER_59_786 ();
 sg13g2_fill_2 FILLER_59_793 ();
 sg13g2_fill_2 FILLER_59_800 ();
 sg13g2_decap_4 FILLER_59_826 ();
 sg13g2_fill_1 FILLER_59_830 ();
 sg13g2_decap_4 FILLER_59_840 ();
 sg13g2_fill_2 FILLER_59_844 ();
 sg13g2_decap_4 FILLER_59_863 ();
 sg13g2_fill_2 FILLER_59_867 ();
 sg13g2_fill_1 FILLER_59_887 ();
 sg13g2_decap_4 FILLER_59_958 ();
 sg13g2_decap_8 FILLER_59_966 ();
 sg13g2_fill_1 FILLER_59_973 ();
 sg13g2_fill_1 FILLER_59_994 ();
 sg13g2_decap_8 FILLER_59_1000 ();
 sg13g2_decap_8 FILLER_59_1007 ();
 sg13g2_fill_2 FILLER_59_1014 ();
 sg13g2_fill_1 FILLER_59_1016 ();
 sg13g2_fill_2 FILLER_59_1021 ();
 sg13g2_fill_2 FILLER_59_1060 ();
 sg13g2_fill_1 FILLER_59_1098 ();
 sg13g2_fill_2 FILLER_59_1120 ();
 sg13g2_fill_2 FILLER_59_1143 ();
 sg13g2_fill_1 FILLER_59_1145 ();
 sg13g2_fill_2 FILLER_59_1159 ();
 sg13g2_fill_2 FILLER_59_1222 ();
 sg13g2_fill_1 FILLER_59_1294 ();
 sg13g2_decap_8 FILLER_59_1321 ();
 sg13g2_fill_2 FILLER_59_1328 ();
 sg13g2_fill_1 FILLER_59_1335 ();
 sg13g2_fill_2 FILLER_59_1340 ();
 sg13g2_fill_1 FILLER_59_1372 ();
 sg13g2_fill_1 FILLER_59_1429 ();
 sg13g2_fill_1 FILLER_59_1443 ();
 sg13g2_decap_4 FILLER_59_1497 ();
 sg13g2_fill_1 FILLER_59_1501 ();
 sg13g2_fill_1 FILLER_59_1518 ();
 sg13g2_fill_1 FILLER_59_1550 ();
 sg13g2_fill_1 FILLER_59_1559 ();
 sg13g2_decap_4 FILLER_59_1628 ();
 sg13g2_fill_2 FILLER_59_1636 ();
 sg13g2_fill_2 FILLER_59_1664 ();
 sg13g2_fill_1 FILLER_59_1683 ();
 sg13g2_decap_4 FILLER_59_1719 ();
 sg13g2_fill_1 FILLER_59_1771 ();
 sg13g2_fill_2 FILLER_59_1776 ();
 sg13g2_fill_1 FILLER_59_1778 ();
 sg13g2_fill_1 FILLER_59_1814 ();
 sg13g2_fill_2 FILLER_59_1820 ();
 sg13g2_fill_1 FILLER_59_1822 ();
 sg13g2_fill_1 FILLER_59_1836 ();
 sg13g2_fill_2 FILLER_59_1908 ();
 sg13g2_decap_4 FILLER_59_1945 ();
 sg13g2_fill_1 FILLER_59_1949 ();
 sg13g2_fill_1 FILLER_59_1967 ();
 sg13g2_decap_4 FILLER_59_1972 ();
 sg13g2_fill_1 FILLER_59_1976 ();
 sg13g2_decap_8 FILLER_59_1987 ();
 sg13g2_fill_1 FILLER_59_1998 ();
 sg13g2_decap_8 FILLER_59_2068 ();
 sg13g2_decap_4 FILLER_59_2079 ();
 sg13g2_decap_8 FILLER_59_2113 ();
 sg13g2_fill_2 FILLER_59_2130 ();
 sg13g2_fill_1 FILLER_59_2155 ();
 sg13g2_fill_1 FILLER_59_2174 ();
 sg13g2_decap_4 FILLER_59_2213 ();
 sg13g2_fill_2 FILLER_59_2217 ();
 sg13g2_fill_2 FILLER_59_2251 ();
 sg13g2_fill_1 FILLER_59_2253 ();
 sg13g2_fill_2 FILLER_59_2281 ();
 sg13g2_fill_1 FILLER_59_2283 ();
 sg13g2_decap_8 FILLER_59_2319 ();
 sg13g2_decap_8 FILLER_59_2326 ();
 sg13g2_decap_8 FILLER_59_2333 ();
 sg13g2_decap_8 FILLER_59_2340 ();
 sg13g2_decap_8 FILLER_59_2347 ();
 sg13g2_decap_8 FILLER_59_2354 ();
 sg13g2_decap_8 FILLER_59_2361 ();
 sg13g2_decap_8 FILLER_59_2368 ();
 sg13g2_decap_8 FILLER_59_2375 ();
 sg13g2_decap_8 FILLER_59_2382 ();
 sg13g2_decap_8 FILLER_59_2389 ();
 sg13g2_decap_8 FILLER_59_2396 ();
 sg13g2_decap_8 FILLER_59_2403 ();
 sg13g2_decap_8 FILLER_59_2410 ();
 sg13g2_decap_8 FILLER_59_2417 ();
 sg13g2_decap_8 FILLER_59_2424 ();
 sg13g2_decap_8 FILLER_59_2431 ();
 sg13g2_decap_8 FILLER_59_2438 ();
 sg13g2_decap_8 FILLER_59_2445 ();
 sg13g2_decap_8 FILLER_59_2452 ();
 sg13g2_decap_8 FILLER_59_2459 ();
 sg13g2_decap_8 FILLER_59_2466 ();
 sg13g2_decap_8 FILLER_59_2473 ();
 sg13g2_decap_8 FILLER_59_2480 ();
 sg13g2_decap_8 FILLER_59_2487 ();
 sg13g2_decap_8 FILLER_59_2494 ();
 sg13g2_decap_8 FILLER_59_2501 ();
 sg13g2_decap_8 FILLER_59_2508 ();
 sg13g2_decap_8 FILLER_59_2515 ();
 sg13g2_decap_8 FILLER_59_2522 ();
 sg13g2_decap_8 FILLER_59_2529 ();
 sg13g2_decap_8 FILLER_59_2536 ();
 sg13g2_decap_8 FILLER_59_2543 ();
 sg13g2_decap_8 FILLER_59_2550 ();
 sg13g2_decap_8 FILLER_59_2557 ();
 sg13g2_decap_8 FILLER_59_2564 ();
 sg13g2_decap_8 FILLER_59_2571 ();
 sg13g2_decap_8 FILLER_59_2578 ();
 sg13g2_decap_8 FILLER_59_2585 ();
 sg13g2_decap_8 FILLER_59_2592 ();
 sg13g2_decap_8 FILLER_59_2599 ();
 sg13g2_decap_8 FILLER_59_2606 ();
 sg13g2_decap_8 FILLER_59_2613 ();
 sg13g2_decap_8 FILLER_59_2620 ();
 sg13g2_decap_8 FILLER_59_2627 ();
 sg13g2_decap_8 FILLER_59_2634 ();
 sg13g2_decap_8 FILLER_59_2641 ();
 sg13g2_decap_8 FILLER_59_2648 ();
 sg13g2_decap_8 FILLER_59_2655 ();
 sg13g2_decap_8 FILLER_59_2662 ();
 sg13g2_decap_4 FILLER_59_2669 ();
 sg13g2_fill_1 FILLER_59_2673 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_decap_8 FILLER_60_133 ();
 sg13g2_decap_8 FILLER_60_140 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_decap_8 FILLER_60_154 ();
 sg13g2_decap_8 FILLER_60_161 ();
 sg13g2_decap_8 FILLER_60_168 ();
 sg13g2_decap_8 FILLER_60_175 ();
 sg13g2_decap_8 FILLER_60_182 ();
 sg13g2_decap_8 FILLER_60_189 ();
 sg13g2_decap_8 FILLER_60_196 ();
 sg13g2_decap_8 FILLER_60_203 ();
 sg13g2_decap_8 FILLER_60_210 ();
 sg13g2_decap_8 FILLER_60_217 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_decap_8 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_238 ();
 sg13g2_decap_8 FILLER_60_245 ();
 sg13g2_decap_8 FILLER_60_252 ();
 sg13g2_decap_8 FILLER_60_259 ();
 sg13g2_decap_8 FILLER_60_266 ();
 sg13g2_decap_8 FILLER_60_273 ();
 sg13g2_decap_8 FILLER_60_280 ();
 sg13g2_decap_8 FILLER_60_287 ();
 sg13g2_decap_8 FILLER_60_294 ();
 sg13g2_decap_8 FILLER_60_301 ();
 sg13g2_decap_8 FILLER_60_308 ();
 sg13g2_decap_8 FILLER_60_315 ();
 sg13g2_decap_8 FILLER_60_322 ();
 sg13g2_decap_8 FILLER_60_329 ();
 sg13g2_decap_8 FILLER_60_336 ();
 sg13g2_decap_8 FILLER_60_343 ();
 sg13g2_decap_8 FILLER_60_350 ();
 sg13g2_decap_8 FILLER_60_357 ();
 sg13g2_decap_8 FILLER_60_364 ();
 sg13g2_decap_8 FILLER_60_371 ();
 sg13g2_decap_8 FILLER_60_378 ();
 sg13g2_decap_8 FILLER_60_385 ();
 sg13g2_decap_8 FILLER_60_392 ();
 sg13g2_decap_8 FILLER_60_399 ();
 sg13g2_decap_8 FILLER_60_406 ();
 sg13g2_decap_8 FILLER_60_413 ();
 sg13g2_decap_8 FILLER_60_420 ();
 sg13g2_decap_8 FILLER_60_427 ();
 sg13g2_decap_8 FILLER_60_434 ();
 sg13g2_decap_8 FILLER_60_441 ();
 sg13g2_decap_8 FILLER_60_448 ();
 sg13g2_decap_8 FILLER_60_455 ();
 sg13g2_decap_4 FILLER_60_462 ();
 sg13g2_decap_4 FILLER_60_479 ();
 sg13g2_fill_1 FILLER_60_483 ();
 sg13g2_decap_4 FILLER_60_494 ();
 sg13g2_fill_1 FILLER_60_525 ();
 sg13g2_fill_2 FILLER_60_596 ();
 sg13g2_fill_1 FILLER_60_598 ();
 sg13g2_fill_1 FILLER_60_635 ();
 sg13g2_fill_2 FILLER_60_685 ();
 sg13g2_decap_8 FILLER_60_691 ();
 sg13g2_fill_1 FILLER_60_698 ();
 sg13g2_decap_8 FILLER_60_707 ();
 sg13g2_fill_2 FILLER_60_714 ();
 sg13g2_fill_2 FILLER_60_733 ();
 sg13g2_fill_1 FILLER_60_735 ();
 sg13g2_fill_2 FILLER_60_745 ();
 sg13g2_fill_2 FILLER_60_756 ();
 sg13g2_fill_1 FILLER_60_758 ();
 sg13g2_fill_2 FILLER_60_764 ();
 sg13g2_fill_1 FILLER_60_796 ();
 sg13g2_fill_2 FILLER_60_818 ();
 sg13g2_fill_2 FILLER_60_825 ();
 sg13g2_fill_1 FILLER_60_827 ();
 sg13g2_fill_2 FILLER_60_859 ();
 sg13g2_fill_1 FILLER_60_896 ();
 sg13g2_decap_4 FILLER_60_950 ();
 sg13g2_fill_1 FILLER_60_993 ();
 sg13g2_fill_2 FILLER_60_1002 ();
 sg13g2_fill_1 FILLER_60_1004 ();
 sg13g2_fill_1 FILLER_60_1050 ();
 sg13g2_fill_2 FILLER_60_1060 ();
 sg13g2_fill_1 FILLER_60_1080 ();
 sg13g2_fill_2 FILLER_60_1108 ();
 sg13g2_fill_2 FILLER_60_1171 ();
 sg13g2_fill_2 FILLER_60_1180 ();
 sg13g2_fill_2 FILLER_60_1187 ();
 sg13g2_decap_8 FILLER_60_1195 ();
 sg13g2_decap_4 FILLER_60_1202 ();
 sg13g2_fill_2 FILLER_60_1206 ();
 sg13g2_fill_1 FILLER_60_1234 ();
 sg13g2_decap_8 FILLER_60_1263 ();
 sg13g2_fill_2 FILLER_60_1270 ();
 sg13g2_fill_1 FILLER_60_1272 ();
 sg13g2_fill_2 FILLER_60_1278 ();
 sg13g2_fill_1 FILLER_60_1280 ();
 sg13g2_fill_1 FILLER_60_1295 ();
 sg13g2_fill_2 FILLER_60_1305 ();
 sg13g2_fill_1 FILLER_60_1307 ();
 sg13g2_fill_2 FILLER_60_1382 ();
 sg13g2_fill_2 FILLER_60_1398 ();
 sg13g2_fill_1 FILLER_60_1413 ();
 sg13g2_decap_4 FILLER_60_1419 ();
 sg13g2_decap_8 FILLER_60_1427 ();
 sg13g2_decap_8 FILLER_60_1434 ();
 sg13g2_decap_8 FILLER_60_1441 ();
 sg13g2_decap_8 FILLER_60_1448 ();
 sg13g2_fill_1 FILLER_60_1463 ();
 sg13g2_fill_2 FILLER_60_1490 ();
 sg13g2_fill_2 FILLER_60_1518 ();
 sg13g2_fill_1 FILLER_60_1520 ();
 sg13g2_fill_2 FILLER_60_1535 ();
 sg13g2_fill_1 FILLER_60_1537 ();
 sg13g2_fill_1 FILLER_60_1586 ();
 sg13g2_decap_8 FILLER_60_1685 ();
 sg13g2_fill_1 FILLER_60_1692 ();
 sg13g2_fill_1 FILLER_60_1698 ();
 sg13g2_decap_8 FILLER_60_1707 ();
 sg13g2_fill_2 FILLER_60_1745 ();
 sg13g2_fill_1 FILLER_60_1747 ();
 sg13g2_decap_4 FILLER_60_1752 ();
 sg13g2_fill_1 FILLER_60_1760 ();
 sg13g2_fill_2 FILLER_60_1810 ();
 sg13g2_fill_1 FILLER_60_1846 ();
 sg13g2_decap_8 FILLER_60_1860 ();
 sg13g2_fill_2 FILLER_60_1867 ();
 sg13g2_fill_2 FILLER_60_1878 ();
 sg13g2_fill_2 FILLER_60_1915 ();
 sg13g2_fill_1 FILLER_60_1961 ();
 sg13g2_decap_4 FILLER_60_1988 ();
 sg13g2_fill_1 FILLER_60_1992 ();
 sg13g2_decap_4 FILLER_60_1998 ();
 sg13g2_fill_2 FILLER_60_2006 ();
 sg13g2_fill_2 FILLER_60_2031 ();
 sg13g2_decap_8 FILLER_60_2078 ();
 sg13g2_decap_8 FILLER_60_2085 ();
 sg13g2_fill_2 FILLER_60_2092 ();
 sg13g2_fill_2 FILLER_60_2150 ();
 sg13g2_fill_1 FILLER_60_2152 ();
 sg13g2_fill_2 FILLER_60_2179 ();
 sg13g2_fill_1 FILLER_60_2255 ();
 sg13g2_decap_4 FILLER_60_2291 ();
 sg13g2_fill_1 FILLER_60_2295 ();
 sg13g2_fill_2 FILLER_60_2300 ();
 sg13g2_decap_8 FILLER_60_2315 ();
 sg13g2_decap_8 FILLER_60_2322 ();
 sg13g2_decap_8 FILLER_60_2329 ();
 sg13g2_decap_8 FILLER_60_2336 ();
 sg13g2_decap_8 FILLER_60_2343 ();
 sg13g2_decap_8 FILLER_60_2350 ();
 sg13g2_decap_8 FILLER_60_2357 ();
 sg13g2_decap_8 FILLER_60_2364 ();
 sg13g2_decap_8 FILLER_60_2371 ();
 sg13g2_decap_8 FILLER_60_2378 ();
 sg13g2_decap_8 FILLER_60_2385 ();
 sg13g2_decap_8 FILLER_60_2392 ();
 sg13g2_decap_8 FILLER_60_2399 ();
 sg13g2_decap_8 FILLER_60_2406 ();
 sg13g2_decap_8 FILLER_60_2413 ();
 sg13g2_decap_8 FILLER_60_2420 ();
 sg13g2_decap_8 FILLER_60_2427 ();
 sg13g2_decap_8 FILLER_60_2434 ();
 sg13g2_decap_8 FILLER_60_2441 ();
 sg13g2_decap_8 FILLER_60_2448 ();
 sg13g2_decap_8 FILLER_60_2455 ();
 sg13g2_decap_8 FILLER_60_2462 ();
 sg13g2_decap_8 FILLER_60_2469 ();
 sg13g2_decap_8 FILLER_60_2476 ();
 sg13g2_decap_8 FILLER_60_2483 ();
 sg13g2_decap_8 FILLER_60_2490 ();
 sg13g2_decap_8 FILLER_60_2497 ();
 sg13g2_decap_8 FILLER_60_2504 ();
 sg13g2_decap_8 FILLER_60_2511 ();
 sg13g2_decap_8 FILLER_60_2518 ();
 sg13g2_decap_8 FILLER_60_2525 ();
 sg13g2_decap_8 FILLER_60_2532 ();
 sg13g2_decap_8 FILLER_60_2539 ();
 sg13g2_decap_8 FILLER_60_2546 ();
 sg13g2_decap_8 FILLER_60_2553 ();
 sg13g2_decap_8 FILLER_60_2560 ();
 sg13g2_decap_8 FILLER_60_2567 ();
 sg13g2_decap_8 FILLER_60_2574 ();
 sg13g2_decap_8 FILLER_60_2581 ();
 sg13g2_decap_8 FILLER_60_2588 ();
 sg13g2_decap_8 FILLER_60_2595 ();
 sg13g2_decap_8 FILLER_60_2602 ();
 sg13g2_decap_8 FILLER_60_2609 ();
 sg13g2_decap_8 FILLER_60_2616 ();
 sg13g2_decap_8 FILLER_60_2623 ();
 sg13g2_decap_8 FILLER_60_2630 ();
 sg13g2_decap_8 FILLER_60_2637 ();
 sg13g2_decap_8 FILLER_60_2644 ();
 sg13g2_decap_8 FILLER_60_2651 ();
 sg13g2_decap_8 FILLER_60_2658 ();
 sg13g2_decap_8 FILLER_60_2665 ();
 sg13g2_fill_2 FILLER_60_2672 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_decap_8 FILLER_61_133 ();
 sg13g2_decap_8 FILLER_61_140 ();
 sg13g2_decap_8 FILLER_61_147 ();
 sg13g2_decap_8 FILLER_61_154 ();
 sg13g2_decap_8 FILLER_61_161 ();
 sg13g2_decap_8 FILLER_61_168 ();
 sg13g2_decap_8 FILLER_61_175 ();
 sg13g2_decap_8 FILLER_61_182 ();
 sg13g2_decap_8 FILLER_61_189 ();
 sg13g2_decap_8 FILLER_61_196 ();
 sg13g2_decap_8 FILLER_61_203 ();
 sg13g2_decap_8 FILLER_61_210 ();
 sg13g2_decap_8 FILLER_61_217 ();
 sg13g2_decap_8 FILLER_61_224 ();
 sg13g2_decap_8 FILLER_61_231 ();
 sg13g2_decap_8 FILLER_61_238 ();
 sg13g2_decap_8 FILLER_61_245 ();
 sg13g2_decap_8 FILLER_61_252 ();
 sg13g2_decap_8 FILLER_61_259 ();
 sg13g2_decap_8 FILLER_61_266 ();
 sg13g2_decap_8 FILLER_61_273 ();
 sg13g2_decap_8 FILLER_61_280 ();
 sg13g2_decap_8 FILLER_61_287 ();
 sg13g2_decap_8 FILLER_61_294 ();
 sg13g2_decap_8 FILLER_61_301 ();
 sg13g2_decap_8 FILLER_61_308 ();
 sg13g2_decap_8 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_322 ();
 sg13g2_decap_8 FILLER_61_329 ();
 sg13g2_decap_8 FILLER_61_336 ();
 sg13g2_decap_8 FILLER_61_343 ();
 sg13g2_decap_8 FILLER_61_350 ();
 sg13g2_decap_8 FILLER_61_357 ();
 sg13g2_decap_8 FILLER_61_364 ();
 sg13g2_decap_8 FILLER_61_371 ();
 sg13g2_decap_8 FILLER_61_378 ();
 sg13g2_decap_8 FILLER_61_385 ();
 sg13g2_decap_8 FILLER_61_392 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_decap_8 FILLER_61_406 ();
 sg13g2_decap_8 FILLER_61_413 ();
 sg13g2_decap_8 FILLER_61_420 ();
 sg13g2_decap_8 FILLER_61_427 ();
 sg13g2_decap_8 FILLER_61_434 ();
 sg13g2_decap_8 FILLER_61_441 ();
 sg13g2_decap_8 FILLER_61_448 ();
 sg13g2_decap_4 FILLER_61_455 ();
 sg13g2_fill_1 FILLER_61_459 ();
 sg13g2_fill_1 FILLER_61_486 ();
 sg13g2_fill_1 FILLER_61_553 ();
 sg13g2_fill_1 FILLER_61_570 ();
 sg13g2_fill_1 FILLER_61_580 ();
 sg13g2_decap_8 FILLER_61_591 ();
 sg13g2_fill_2 FILLER_61_598 ();
 sg13g2_fill_1 FILLER_61_600 ();
 sg13g2_fill_2 FILLER_61_614 ();
 sg13g2_fill_2 FILLER_61_656 ();
 sg13g2_decap_4 FILLER_61_662 ();
 sg13g2_fill_1 FILLER_61_679 ();
 sg13g2_fill_2 FILLER_61_711 ();
 sg13g2_fill_1 FILLER_61_713 ();
 sg13g2_fill_2 FILLER_61_719 ();
 sg13g2_fill_2 FILLER_61_729 ();
 sg13g2_fill_2 FILLER_61_766 ();
 sg13g2_fill_2 FILLER_61_777 ();
 sg13g2_fill_2 FILLER_61_789 ();
 sg13g2_decap_4 FILLER_61_832 ();
 sg13g2_fill_2 FILLER_61_836 ();
 sg13g2_decap_8 FILLER_61_842 ();
 sg13g2_fill_2 FILLER_61_849 ();
 sg13g2_decap_4 FILLER_61_860 ();
 sg13g2_fill_1 FILLER_61_864 ();
 sg13g2_fill_2 FILLER_61_879 ();
 sg13g2_fill_1 FILLER_61_881 ();
 sg13g2_fill_1 FILLER_61_906 ();
 sg13g2_fill_1 FILLER_61_911 ();
 sg13g2_fill_2 FILLER_61_926 ();
 sg13g2_fill_1 FILLER_61_928 ();
 sg13g2_decap_4 FILLER_61_964 ();
 sg13g2_fill_2 FILLER_61_968 ();
 sg13g2_decap_8 FILLER_61_974 ();
 sg13g2_decap_4 FILLER_61_981 ();
 sg13g2_fill_1 FILLER_61_985 ();
 sg13g2_decap_4 FILLER_61_991 ();
 sg13g2_decap_4 FILLER_61_1000 ();
 sg13g2_fill_2 FILLER_61_1025 ();
 sg13g2_decap_4 FILLER_61_1077 ();
 sg13g2_fill_2 FILLER_61_1099 ();
 sg13g2_fill_1 FILLER_61_1142 ();
 sg13g2_decap_8 FILLER_61_1148 ();
 sg13g2_fill_1 FILLER_61_1155 ();
 sg13g2_decap_4 FILLER_61_1160 ();
 sg13g2_fill_2 FILLER_61_1164 ();
 sg13g2_decap_4 FILLER_61_1211 ();
 sg13g2_decap_4 FILLER_61_1227 ();
 sg13g2_fill_2 FILLER_61_1231 ();
 sg13g2_decap_4 FILLER_61_1243 ();
 sg13g2_fill_1 FILLER_61_1247 ();
 sg13g2_fill_1 FILLER_61_1258 ();
 sg13g2_decap_8 FILLER_61_1269 ();
 sg13g2_fill_2 FILLER_61_1307 ();
 sg13g2_fill_1 FILLER_61_1309 ();
 sg13g2_decap_4 FILLER_61_1327 ();
 sg13g2_fill_1 FILLER_61_1335 ();
 sg13g2_fill_2 FILLER_61_1340 ();
 sg13g2_decap_8 FILLER_61_1351 ();
 sg13g2_decap_8 FILLER_61_1358 ();
 sg13g2_fill_2 FILLER_61_1365 ();
 sg13g2_fill_1 FILLER_61_1367 ();
 sg13g2_fill_1 FILLER_61_1381 ();
 sg13g2_fill_1 FILLER_61_1387 ();
 sg13g2_fill_1 FILLER_61_1402 ();
 sg13g2_fill_2 FILLER_61_1442 ();
 sg13g2_fill_2 FILLER_61_1453 ();
 sg13g2_fill_1 FILLER_61_1464 ();
 sg13g2_decap_4 FILLER_61_1469 ();
 sg13g2_fill_1 FILLER_61_1489 ();
 sg13g2_fill_2 FILLER_61_1499 ();
 sg13g2_fill_1 FILLER_61_1501 ();
 sg13g2_fill_2 FILLER_61_1528 ();
 sg13g2_fill_1 FILLER_61_1530 ();
 sg13g2_fill_1 FILLER_61_1546 ();
 sg13g2_fill_2 FILLER_61_1556 ();
 sg13g2_fill_2 FILLER_61_1579 ();
 sg13g2_fill_2 FILLER_61_1601 ();
 sg13g2_fill_1 FILLER_61_1612 ();
 sg13g2_fill_2 FILLER_61_1618 ();
 sg13g2_decap_8 FILLER_61_1676 ();
 sg13g2_fill_2 FILLER_61_1699 ();
 sg13g2_fill_2 FILLER_61_1736 ();
 sg13g2_fill_1 FILLER_61_1738 ();
 sg13g2_decap_4 FILLER_61_1769 ();
 sg13g2_fill_1 FILLER_61_1829 ();
 sg13g2_fill_2 FILLER_61_1843 ();
 sg13g2_fill_1 FILLER_61_1845 ();
 sg13g2_fill_1 FILLER_61_1872 ();
 sg13g2_fill_2 FILLER_61_1895 ();
 sg13g2_fill_1 FILLER_61_1897 ();
 sg13g2_fill_1 FILLER_61_1985 ();
 sg13g2_fill_2 FILLER_61_2021 ();
 sg13g2_fill_1 FILLER_61_2023 ();
 sg13g2_decap_8 FILLER_61_2040 ();
 sg13g2_fill_2 FILLER_61_2047 ();
 sg13g2_fill_2 FILLER_61_2053 ();
 sg13g2_fill_2 FILLER_61_2090 ();
 sg13g2_fill_1 FILLER_61_2092 ();
 sg13g2_fill_2 FILLER_61_2132 ();
 sg13g2_decap_8 FILLER_61_2152 ();
 sg13g2_fill_2 FILLER_61_2159 ();
 sg13g2_fill_2 FILLER_61_2173 ();
 sg13g2_fill_2 FILLER_61_2180 ();
 sg13g2_fill_2 FILLER_61_2195 ();
 sg13g2_decap_4 FILLER_61_2206 ();
 sg13g2_fill_1 FILLER_61_2210 ();
 sg13g2_fill_1 FILLER_61_2248 ();
 sg13g2_decap_8 FILLER_61_2311 ();
 sg13g2_decap_8 FILLER_61_2318 ();
 sg13g2_decap_8 FILLER_61_2325 ();
 sg13g2_decap_8 FILLER_61_2332 ();
 sg13g2_decap_8 FILLER_61_2339 ();
 sg13g2_decap_8 FILLER_61_2346 ();
 sg13g2_decap_8 FILLER_61_2353 ();
 sg13g2_decap_8 FILLER_61_2360 ();
 sg13g2_decap_8 FILLER_61_2367 ();
 sg13g2_decap_8 FILLER_61_2374 ();
 sg13g2_decap_8 FILLER_61_2381 ();
 sg13g2_decap_8 FILLER_61_2388 ();
 sg13g2_decap_8 FILLER_61_2395 ();
 sg13g2_decap_8 FILLER_61_2402 ();
 sg13g2_decap_8 FILLER_61_2409 ();
 sg13g2_decap_8 FILLER_61_2416 ();
 sg13g2_decap_8 FILLER_61_2423 ();
 sg13g2_decap_8 FILLER_61_2430 ();
 sg13g2_decap_8 FILLER_61_2437 ();
 sg13g2_decap_8 FILLER_61_2444 ();
 sg13g2_decap_8 FILLER_61_2451 ();
 sg13g2_decap_8 FILLER_61_2458 ();
 sg13g2_decap_8 FILLER_61_2465 ();
 sg13g2_decap_8 FILLER_61_2472 ();
 sg13g2_decap_8 FILLER_61_2479 ();
 sg13g2_decap_8 FILLER_61_2486 ();
 sg13g2_decap_8 FILLER_61_2493 ();
 sg13g2_decap_8 FILLER_61_2500 ();
 sg13g2_decap_8 FILLER_61_2507 ();
 sg13g2_decap_8 FILLER_61_2514 ();
 sg13g2_decap_8 FILLER_61_2521 ();
 sg13g2_decap_8 FILLER_61_2528 ();
 sg13g2_decap_8 FILLER_61_2535 ();
 sg13g2_decap_8 FILLER_61_2542 ();
 sg13g2_decap_8 FILLER_61_2549 ();
 sg13g2_decap_8 FILLER_61_2556 ();
 sg13g2_decap_8 FILLER_61_2563 ();
 sg13g2_decap_8 FILLER_61_2570 ();
 sg13g2_decap_8 FILLER_61_2577 ();
 sg13g2_decap_8 FILLER_61_2584 ();
 sg13g2_decap_8 FILLER_61_2591 ();
 sg13g2_decap_8 FILLER_61_2598 ();
 sg13g2_decap_8 FILLER_61_2605 ();
 sg13g2_decap_8 FILLER_61_2612 ();
 sg13g2_decap_8 FILLER_61_2619 ();
 sg13g2_decap_8 FILLER_61_2626 ();
 sg13g2_decap_8 FILLER_61_2633 ();
 sg13g2_decap_8 FILLER_61_2640 ();
 sg13g2_decap_8 FILLER_61_2647 ();
 sg13g2_decap_8 FILLER_61_2654 ();
 sg13g2_decap_8 FILLER_61_2661 ();
 sg13g2_decap_4 FILLER_61_2668 ();
 sg13g2_fill_2 FILLER_61_2672 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_8 FILLER_62_161 ();
 sg13g2_decap_8 FILLER_62_168 ();
 sg13g2_decap_8 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_182 ();
 sg13g2_decap_8 FILLER_62_189 ();
 sg13g2_decap_8 FILLER_62_196 ();
 sg13g2_decap_8 FILLER_62_203 ();
 sg13g2_decap_8 FILLER_62_210 ();
 sg13g2_decap_8 FILLER_62_217 ();
 sg13g2_decap_8 FILLER_62_224 ();
 sg13g2_decap_8 FILLER_62_231 ();
 sg13g2_decap_8 FILLER_62_238 ();
 sg13g2_decap_8 FILLER_62_245 ();
 sg13g2_decap_8 FILLER_62_252 ();
 sg13g2_decap_8 FILLER_62_259 ();
 sg13g2_decap_8 FILLER_62_266 ();
 sg13g2_decap_8 FILLER_62_273 ();
 sg13g2_decap_8 FILLER_62_280 ();
 sg13g2_decap_8 FILLER_62_287 ();
 sg13g2_decap_8 FILLER_62_294 ();
 sg13g2_decap_8 FILLER_62_301 ();
 sg13g2_decap_8 FILLER_62_308 ();
 sg13g2_decap_8 FILLER_62_315 ();
 sg13g2_decap_8 FILLER_62_322 ();
 sg13g2_decap_8 FILLER_62_329 ();
 sg13g2_decap_8 FILLER_62_336 ();
 sg13g2_decap_8 FILLER_62_343 ();
 sg13g2_decap_8 FILLER_62_350 ();
 sg13g2_decap_8 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_364 ();
 sg13g2_decap_8 FILLER_62_371 ();
 sg13g2_decap_8 FILLER_62_378 ();
 sg13g2_decap_8 FILLER_62_385 ();
 sg13g2_decap_8 FILLER_62_392 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_decap_8 FILLER_62_406 ();
 sg13g2_decap_8 FILLER_62_413 ();
 sg13g2_decap_8 FILLER_62_420 ();
 sg13g2_decap_8 FILLER_62_427 ();
 sg13g2_decap_8 FILLER_62_434 ();
 sg13g2_decap_8 FILLER_62_441 ();
 sg13g2_decap_8 FILLER_62_448 ();
 sg13g2_decap_8 FILLER_62_455 ();
 sg13g2_decap_8 FILLER_62_462 ();
 sg13g2_fill_1 FILLER_62_469 ();
 sg13g2_decap_8 FILLER_62_492 ();
 sg13g2_fill_2 FILLER_62_499 ();
 sg13g2_fill_1 FILLER_62_501 ();
 sg13g2_decap_8 FILLER_62_511 ();
 sg13g2_decap_4 FILLER_62_518 ();
 sg13g2_fill_1 FILLER_62_522 ();
 sg13g2_fill_2 FILLER_62_527 ();
 sg13g2_fill_1 FILLER_62_529 ();
 sg13g2_fill_1 FILLER_62_580 ();
 sg13g2_fill_1 FILLER_62_594 ();
 sg13g2_fill_1 FILLER_62_678 ();
 sg13g2_decap_4 FILLER_62_701 ();
 sg13g2_fill_2 FILLER_62_705 ();
 sg13g2_fill_2 FILLER_62_802 ();
 sg13g2_fill_1 FILLER_62_804 ();
 sg13g2_fill_2 FILLER_62_819 ();
 sg13g2_decap_4 FILLER_62_825 ();
 sg13g2_fill_1 FILLER_62_829 ();
 sg13g2_fill_2 FILLER_62_845 ();
 sg13g2_fill_1 FILLER_62_847 ();
 sg13g2_fill_2 FILLER_62_879 ();
 sg13g2_fill_2 FILLER_62_894 ();
 sg13g2_fill_2 FILLER_62_943 ();
 sg13g2_decap_4 FILLER_62_954 ();
 sg13g2_fill_2 FILLER_62_968 ();
 sg13g2_fill_2 FILLER_62_974 ();
 sg13g2_fill_1 FILLER_62_1050 ();
 sg13g2_fill_2 FILLER_62_1055 ();
 sg13g2_fill_1 FILLER_62_1057 ();
 sg13g2_fill_1 FILLER_62_1071 ();
 sg13g2_decap_4 FILLER_62_1111 ();
 sg13g2_fill_1 FILLER_62_1115 ();
 sg13g2_fill_2 FILLER_62_1160 ();
 sg13g2_decap_4 FILLER_62_1217 ();
 sg13g2_fill_1 FILLER_62_1221 ();
 sg13g2_fill_2 FILLER_62_1305 ();
 sg13g2_decap_4 FILLER_62_1338 ();
 sg13g2_fill_2 FILLER_62_1342 ();
 sg13g2_decap_8 FILLER_62_1352 ();
 sg13g2_fill_2 FILLER_62_1359 ();
 sg13g2_fill_1 FILLER_62_1361 ();
 sg13g2_decap_8 FILLER_62_1366 ();
 sg13g2_fill_1 FILLER_62_1373 ();
 sg13g2_fill_1 FILLER_62_1422 ();
 sg13g2_fill_2 FILLER_62_1510 ();
 sg13g2_fill_2 FILLER_62_1538 ();
 sg13g2_fill_2 FILLER_62_1580 ();
 sg13g2_fill_2 FILLER_62_1594 ();
 sg13g2_fill_1 FILLER_62_1596 ();
 sg13g2_fill_2 FILLER_62_1606 ();
 sg13g2_fill_1 FILLER_62_1608 ();
 sg13g2_fill_1 FILLER_62_1622 ();
 sg13g2_fill_2 FILLER_62_1661 ();
 sg13g2_fill_1 FILLER_62_1663 ();
 sg13g2_fill_2 FILLER_62_1687 ();
 sg13g2_fill_1 FILLER_62_1689 ();
 sg13g2_fill_1 FILLER_62_1703 ();
 sg13g2_fill_2 FILLER_62_1709 ();
 sg13g2_fill_1 FILLER_62_1711 ();
 sg13g2_fill_2 FILLER_62_1720 ();
 sg13g2_fill_1 FILLER_62_1722 ();
 sg13g2_fill_2 FILLER_62_1757 ();
 sg13g2_fill_1 FILLER_62_1759 ();
 sg13g2_fill_2 FILLER_62_1770 ();
 sg13g2_fill_1 FILLER_62_1772 ();
 sg13g2_fill_2 FILLER_62_1799 ();
 sg13g2_fill_1 FILLER_62_1810 ();
 sg13g2_fill_2 FILLER_62_1824 ();
 sg13g2_decap_4 FILLER_62_1851 ();
 sg13g2_fill_1 FILLER_62_1872 ();
 sg13g2_fill_1 FILLER_62_1896 ();
 sg13g2_fill_2 FILLER_62_1914 ();
 sg13g2_fill_2 FILLER_62_1929 ();
 sg13g2_fill_1 FILLER_62_1931 ();
 sg13g2_fill_2 FILLER_62_1941 ();
 sg13g2_fill_1 FILLER_62_1943 ();
 sg13g2_fill_1 FILLER_62_1951 ();
 sg13g2_decap_4 FILLER_62_1992 ();
 sg13g2_fill_1 FILLER_62_1996 ();
 sg13g2_decap_8 FILLER_62_2005 ();
 sg13g2_decap_4 FILLER_62_2016 ();
 sg13g2_fill_1 FILLER_62_2025 ();
 sg13g2_fill_2 FILLER_62_2051 ();
 sg13g2_fill_2 FILLER_62_2058 ();
 sg13g2_fill_2 FILLER_62_2074 ();
 sg13g2_fill_1 FILLER_62_2121 ();
 sg13g2_fill_1 FILLER_62_2135 ();
 sg13g2_fill_2 FILLER_62_2239 ();
 sg13g2_fill_1 FILLER_62_2241 ();
 sg13g2_fill_1 FILLER_62_2258 ();
 sg13g2_decap_4 FILLER_62_2290 ();
 sg13g2_fill_1 FILLER_62_2294 ();
 sg13g2_decap_8 FILLER_62_2304 ();
 sg13g2_decap_8 FILLER_62_2311 ();
 sg13g2_decap_8 FILLER_62_2318 ();
 sg13g2_decap_8 FILLER_62_2325 ();
 sg13g2_decap_8 FILLER_62_2332 ();
 sg13g2_decap_8 FILLER_62_2339 ();
 sg13g2_decap_8 FILLER_62_2346 ();
 sg13g2_decap_8 FILLER_62_2353 ();
 sg13g2_decap_8 FILLER_62_2360 ();
 sg13g2_decap_8 FILLER_62_2367 ();
 sg13g2_decap_8 FILLER_62_2374 ();
 sg13g2_decap_8 FILLER_62_2381 ();
 sg13g2_decap_8 FILLER_62_2388 ();
 sg13g2_decap_8 FILLER_62_2395 ();
 sg13g2_decap_8 FILLER_62_2402 ();
 sg13g2_decap_8 FILLER_62_2409 ();
 sg13g2_decap_8 FILLER_62_2416 ();
 sg13g2_decap_8 FILLER_62_2423 ();
 sg13g2_decap_8 FILLER_62_2430 ();
 sg13g2_decap_8 FILLER_62_2437 ();
 sg13g2_decap_8 FILLER_62_2444 ();
 sg13g2_decap_8 FILLER_62_2451 ();
 sg13g2_decap_8 FILLER_62_2458 ();
 sg13g2_decap_8 FILLER_62_2465 ();
 sg13g2_decap_8 FILLER_62_2472 ();
 sg13g2_decap_8 FILLER_62_2479 ();
 sg13g2_decap_8 FILLER_62_2486 ();
 sg13g2_decap_8 FILLER_62_2493 ();
 sg13g2_decap_8 FILLER_62_2500 ();
 sg13g2_decap_8 FILLER_62_2507 ();
 sg13g2_decap_8 FILLER_62_2514 ();
 sg13g2_decap_8 FILLER_62_2521 ();
 sg13g2_decap_8 FILLER_62_2528 ();
 sg13g2_decap_8 FILLER_62_2535 ();
 sg13g2_decap_8 FILLER_62_2542 ();
 sg13g2_decap_8 FILLER_62_2549 ();
 sg13g2_decap_8 FILLER_62_2556 ();
 sg13g2_decap_8 FILLER_62_2563 ();
 sg13g2_decap_8 FILLER_62_2570 ();
 sg13g2_decap_8 FILLER_62_2577 ();
 sg13g2_decap_8 FILLER_62_2584 ();
 sg13g2_decap_8 FILLER_62_2591 ();
 sg13g2_decap_8 FILLER_62_2598 ();
 sg13g2_decap_8 FILLER_62_2605 ();
 sg13g2_decap_8 FILLER_62_2612 ();
 sg13g2_decap_8 FILLER_62_2619 ();
 sg13g2_decap_8 FILLER_62_2626 ();
 sg13g2_decap_8 FILLER_62_2633 ();
 sg13g2_decap_8 FILLER_62_2640 ();
 sg13g2_decap_8 FILLER_62_2647 ();
 sg13g2_decap_8 FILLER_62_2654 ();
 sg13g2_decap_8 FILLER_62_2661 ();
 sg13g2_decap_4 FILLER_62_2668 ();
 sg13g2_fill_2 FILLER_62_2672 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_8 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_140 ();
 sg13g2_decap_8 FILLER_63_147 ();
 sg13g2_decap_8 FILLER_63_154 ();
 sg13g2_decap_8 FILLER_63_161 ();
 sg13g2_decap_8 FILLER_63_168 ();
 sg13g2_decap_8 FILLER_63_175 ();
 sg13g2_decap_8 FILLER_63_182 ();
 sg13g2_decap_8 FILLER_63_189 ();
 sg13g2_decap_8 FILLER_63_196 ();
 sg13g2_decap_8 FILLER_63_203 ();
 sg13g2_decap_8 FILLER_63_210 ();
 sg13g2_decap_8 FILLER_63_217 ();
 sg13g2_decap_8 FILLER_63_224 ();
 sg13g2_decap_8 FILLER_63_231 ();
 sg13g2_decap_8 FILLER_63_238 ();
 sg13g2_decap_8 FILLER_63_245 ();
 sg13g2_decap_8 FILLER_63_252 ();
 sg13g2_decap_8 FILLER_63_259 ();
 sg13g2_decap_8 FILLER_63_266 ();
 sg13g2_decap_8 FILLER_63_273 ();
 sg13g2_decap_8 FILLER_63_280 ();
 sg13g2_decap_8 FILLER_63_287 ();
 sg13g2_decap_8 FILLER_63_294 ();
 sg13g2_decap_8 FILLER_63_301 ();
 sg13g2_decap_8 FILLER_63_308 ();
 sg13g2_decap_8 FILLER_63_315 ();
 sg13g2_decap_8 FILLER_63_322 ();
 sg13g2_decap_8 FILLER_63_329 ();
 sg13g2_decap_8 FILLER_63_336 ();
 sg13g2_decap_8 FILLER_63_343 ();
 sg13g2_decap_8 FILLER_63_350 ();
 sg13g2_decap_8 FILLER_63_357 ();
 sg13g2_decap_8 FILLER_63_364 ();
 sg13g2_decap_8 FILLER_63_371 ();
 sg13g2_decap_8 FILLER_63_378 ();
 sg13g2_decap_8 FILLER_63_385 ();
 sg13g2_decap_8 FILLER_63_392 ();
 sg13g2_decap_8 FILLER_63_399 ();
 sg13g2_decap_8 FILLER_63_406 ();
 sg13g2_decap_8 FILLER_63_413 ();
 sg13g2_decap_8 FILLER_63_420 ();
 sg13g2_decap_8 FILLER_63_427 ();
 sg13g2_decap_8 FILLER_63_434 ();
 sg13g2_decap_8 FILLER_63_441 ();
 sg13g2_decap_8 FILLER_63_448 ();
 sg13g2_decap_8 FILLER_63_455 ();
 sg13g2_decap_4 FILLER_63_462 ();
 sg13g2_fill_1 FILLER_63_466 ();
 sg13g2_fill_1 FILLER_63_498 ();
 sg13g2_fill_2 FILLER_63_540 ();
 sg13g2_fill_1 FILLER_63_542 ();
 sg13g2_fill_1 FILLER_63_583 ();
 sg13g2_fill_1 FILLER_63_602 ();
 sg13g2_fill_1 FILLER_63_633 ();
 sg13g2_decap_4 FILLER_63_638 ();
 sg13g2_fill_2 FILLER_63_642 ();
 sg13g2_fill_2 FILLER_63_653 ();
 sg13g2_fill_2 FILLER_63_673 ();
 sg13g2_fill_1 FILLER_63_675 ();
 sg13g2_fill_2 FILLER_63_707 ();
 sg13g2_fill_2 FILLER_63_713 ();
 sg13g2_fill_2 FILLER_63_725 ();
 sg13g2_fill_1 FILLER_63_727 ();
 sg13g2_decap_4 FILLER_63_745 ();
 sg13g2_fill_2 FILLER_63_749 ();
 sg13g2_fill_2 FILLER_63_760 ();
 sg13g2_fill_1 FILLER_63_767 ();
 sg13g2_fill_2 FILLER_63_809 ();
 sg13g2_decap_4 FILLER_63_851 ();
 sg13g2_decap_8 FILLER_63_897 ();
 sg13g2_decap_4 FILLER_63_904 ();
 sg13g2_fill_2 FILLER_63_913 ();
 sg13g2_fill_1 FILLER_63_915 ();
 sg13g2_fill_2 FILLER_63_954 ();
 sg13g2_fill_1 FILLER_63_956 ();
 sg13g2_fill_2 FILLER_63_1031 ();
 sg13g2_fill_1 FILLER_63_1064 ();
 sg13g2_fill_2 FILLER_63_1070 ();
 sg13g2_fill_2 FILLER_63_1103 ();
 sg13g2_fill_2 FILLER_63_1131 ();
 sg13g2_decap_4 FILLER_63_1159 ();
 sg13g2_fill_1 FILLER_63_1163 ();
 sg13g2_fill_2 FILLER_63_1215 ();
 sg13g2_fill_2 FILLER_63_1275 ();
 sg13g2_fill_1 FILLER_63_1277 ();
 sg13g2_fill_2 FILLER_63_1286 ();
 sg13g2_decap_4 FILLER_63_1297 ();
 sg13g2_fill_2 FILLER_63_1301 ();
 sg13g2_fill_2 FILLER_63_1322 ();
 sg13g2_fill_1 FILLER_63_1324 ();
 sg13g2_fill_1 FILLER_63_1443 ();
 sg13g2_decap_4 FILLER_63_1477 ();
 sg13g2_fill_1 FILLER_63_1481 ();
 sg13g2_fill_1 FILLER_63_1490 ();
 sg13g2_decap_8 FILLER_63_1496 ();
 sg13g2_decap_4 FILLER_63_1503 ();
 sg13g2_fill_1 FILLER_63_1516 ();
 sg13g2_fill_1 FILLER_63_1534 ();
 sg13g2_fill_2 FILLER_63_1544 ();
 sg13g2_fill_1 FILLER_63_1546 ();
 sg13g2_fill_2 FILLER_63_1556 ();
 sg13g2_fill_1 FILLER_63_1558 ();
 sg13g2_fill_1 FILLER_63_1606 ();
 sg13g2_fill_2 FILLER_63_1642 ();
 sg13g2_fill_2 FILLER_63_1683 ();
 sg13g2_decap_8 FILLER_63_1689 ();
 sg13g2_fill_2 FILLER_63_1696 ();
 sg13g2_fill_1 FILLER_63_1698 ();
 sg13g2_fill_2 FILLER_63_1734 ();
 sg13g2_fill_1 FILLER_63_1736 ();
 sg13g2_fill_1 FILLER_63_1760 ();
 sg13g2_fill_1 FILLER_63_1779 ();
 sg13g2_fill_2 FILLER_63_1790 ();
 sg13g2_fill_1 FILLER_63_1792 ();
 sg13g2_fill_1 FILLER_63_1856 ();
 sg13g2_decap_8 FILLER_63_1888 ();
 sg13g2_decap_4 FILLER_63_1899 ();
 sg13g2_fill_1 FILLER_63_1908 ();
 sg13g2_fill_1 FILLER_63_1913 ();
 sg13g2_fill_2 FILLER_63_1918 ();
 sg13g2_fill_2 FILLER_63_1951 ();
 sg13g2_fill_1 FILLER_63_2106 ();
 sg13g2_decap_8 FILLER_63_2133 ();
 sg13g2_decap_8 FILLER_63_2140 ();
 sg13g2_decap_8 FILLER_63_2151 ();
 sg13g2_decap_8 FILLER_63_2158 ();
 sg13g2_fill_2 FILLER_63_2170 ();
 sg13g2_fill_1 FILLER_63_2175 ();
 sg13g2_fill_2 FILLER_63_2180 ();
 sg13g2_fill_2 FILLER_63_2187 ();
 sg13g2_fill_1 FILLER_63_2189 ();
 sg13g2_decap_8 FILLER_63_2199 ();
 sg13g2_decap_4 FILLER_63_2206 ();
 sg13g2_fill_2 FILLER_63_2210 ();
 sg13g2_decap_8 FILLER_63_2217 ();
 sg13g2_fill_2 FILLER_63_2224 ();
 sg13g2_decap_4 FILLER_63_2231 ();
 sg13g2_fill_1 FILLER_63_2235 ();
 sg13g2_decap_4 FILLER_63_2240 ();
 sg13g2_fill_2 FILLER_63_2244 ();
 sg13g2_decap_8 FILLER_63_2312 ();
 sg13g2_decap_8 FILLER_63_2319 ();
 sg13g2_decap_8 FILLER_63_2326 ();
 sg13g2_decap_8 FILLER_63_2333 ();
 sg13g2_decap_8 FILLER_63_2340 ();
 sg13g2_decap_8 FILLER_63_2347 ();
 sg13g2_decap_8 FILLER_63_2354 ();
 sg13g2_decap_8 FILLER_63_2361 ();
 sg13g2_decap_8 FILLER_63_2368 ();
 sg13g2_decap_8 FILLER_63_2375 ();
 sg13g2_decap_8 FILLER_63_2382 ();
 sg13g2_decap_8 FILLER_63_2389 ();
 sg13g2_decap_8 FILLER_63_2396 ();
 sg13g2_decap_8 FILLER_63_2403 ();
 sg13g2_decap_8 FILLER_63_2410 ();
 sg13g2_decap_8 FILLER_63_2417 ();
 sg13g2_decap_8 FILLER_63_2424 ();
 sg13g2_decap_8 FILLER_63_2431 ();
 sg13g2_decap_8 FILLER_63_2438 ();
 sg13g2_decap_8 FILLER_63_2445 ();
 sg13g2_decap_8 FILLER_63_2452 ();
 sg13g2_decap_8 FILLER_63_2459 ();
 sg13g2_decap_8 FILLER_63_2466 ();
 sg13g2_decap_8 FILLER_63_2473 ();
 sg13g2_decap_8 FILLER_63_2480 ();
 sg13g2_decap_8 FILLER_63_2487 ();
 sg13g2_decap_8 FILLER_63_2494 ();
 sg13g2_decap_8 FILLER_63_2501 ();
 sg13g2_decap_8 FILLER_63_2508 ();
 sg13g2_decap_8 FILLER_63_2515 ();
 sg13g2_decap_8 FILLER_63_2522 ();
 sg13g2_decap_8 FILLER_63_2529 ();
 sg13g2_decap_8 FILLER_63_2536 ();
 sg13g2_decap_8 FILLER_63_2543 ();
 sg13g2_decap_8 FILLER_63_2550 ();
 sg13g2_decap_8 FILLER_63_2557 ();
 sg13g2_decap_8 FILLER_63_2564 ();
 sg13g2_decap_8 FILLER_63_2571 ();
 sg13g2_decap_8 FILLER_63_2578 ();
 sg13g2_decap_8 FILLER_63_2585 ();
 sg13g2_decap_8 FILLER_63_2592 ();
 sg13g2_decap_8 FILLER_63_2599 ();
 sg13g2_decap_8 FILLER_63_2606 ();
 sg13g2_decap_8 FILLER_63_2613 ();
 sg13g2_decap_8 FILLER_63_2620 ();
 sg13g2_decap_8 FILLER_63_2627 ();
 sg13g2_decap_8 FILLER_63_2634 ();
 sg13g2_decap_8 FILLER_63_2641 ();
 sg13g2_decap_8 FILLER_63_2648 ();
 sg13g2_decap_8 FILLER_63_2655 ();
 sg13g2_decap_8 FILLER_63_2662 ();
 sg13g2_decap_4 FILLER_63_2669 ();
 sg13g2_fill_1 FILLER_63_2673 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_decap_8 FILLER_64_154 ();
 sg13g2_decap_8 FILLER_64_161 ();
 sg13g2_decap_8 FILLER_64_168 ();
 sg13g2_decap_8 FILLER_64_175 ();
 sg13g2_decap_8 FILLER_64_182 ();
 sg13g2_decap_8 FILLER_64_189 ();
 sg13g2_decap_8 FILLER_64_196 ();
 sg13g2_decap_8 FILLER_64_203 ();
 sg13g2_decap_8 FILLER_64_210 ();
 sg13g2_decap_8 FILLER_64_217 ();
 sg13g2_decap_8 FILLER_64_224 ();
 sg13g2_decap_8 FILLER_64_231 ();
 sg13g2_decap_8 FILLER_64_238 ();
 sg13g2_decap_8 FILLER_64_245 ();
 sg13g2_decap_8 FILLER_64_252 ();
 sg13g2_decap_8 FILLER_64_259 ();
 sg13g2_decap_8 FILLER_64_266 ();
 sg13g2_decap_8 FILLER_64_273 ();
 sg13g2_decap_8 FILLER_64_280 ();
 sg13g2_decap_8 FILLER_64_287 ();
 sg13g2_decap_8 FILLER_64_294 ();
 sg13g2_decap_8 FILLER_64_301 ();
 sg13g2_decap_8 FILLER_64_308 ();
 sg13g2_decap_8 FILLER_64_315 ();
 sg13g2_decap_8 FILLER_64_322 ();
 sg13g2_decap_8 FILLER_64_329 ();
 sg13g2_decap_8 FILLER_64_336 ();
 sg13g2_decap_8 FILLER_64_343 ();
 sg13g2_decap_8 FILLER_64_350 ();
 sg13g2_decap_8 FILLER_64_357 ();
 sg13g2_decap_8 FILLER_64_364 ();
 sg13g2_decap_8 FILLER_64_371 ();
 sg13g2_decap_8 FILLER_64_378 ();
 sg13g2_decap_8 FILLER_64_385 ();
 sg13g2_decap_8 FILLER_64_392 ();
 sg13g2_decap_8 FILLER_64_399 ();
 sg13g2_decap_8 FILLER_64_406 ();
 sg13g2_decap_8 FILLER_64_413 ();
 sg13g2_decap_8 FILLER_64_420 ();
 sg13g2_decap_8 FILLER_64_427 ();
 sg13g2_decap_8 FILLER_64_434 ();
 sg13g2_decap_8 FILLER_64_441 ();
 sg13g2_decap_8 FILLER_64_448 ();
 sg13g2_decap_8 FILLER_64_455 ();
 sg13g2_decap_8 FILLER_64_462 ();
 sg13g2_fill_2 FILLER_64_469 ();
 sg13g2_fill_1 FILLER_64_471 ();
 sg13g2_fill_2 FILLER_64_490 ();
 sg13g2_fill_2 FILLER_64_501 ();
 sg13g2_fill_2 FILLER_64_507 ();
 sg13g2_fill_1 FILLER_64_517 ();
 sg13g2_decap_4 FILLER_64_527 ();
 sg13g2_fill_1 FILLER_64_540 ();
 sg13g2_fill_2 FILLER_64_545 ();
 sg13g2_fill_2 FILLER_64_556 ();
 sg13g2_fill_1 FILLER_64_558 ();
 sg13g2_fill_1 FILLER_64_611 ();
 sg13g2_decap_4 FILLER_64_644 ();
 sg13g2_fill_1 FILLER_64_648 ();
 sg13g2_fill_2 FILLER_64_653 ();
 sg13g2_fill_1 FILLER_64_655 ();
 sg13g2_fill_2 FILLER_64_687 ();
 sg13g2_fill_2 FILLER_64_724 ();
 sg13g2_fill_2 FILLER_64_770 ();
 sg13g2_fill_1 FILLER_64_772 ();
 sg13g2_fill_2 FILLER_64_816 ();
 sg13g2_fill_1 FILLER_64_831 ();
 sg13g2_fill_1 FILLER_64_874 ();
 sg13g2_fill_1 FILLER_64_922 ();
 sg13g2_fill_1 FILLER_64_928 ();
 sg13g2_fill_2 FILLER_64_943 ();
 sg13g2_fill_1 FILLER_64_945 ();
 sg13g2_fill_2 FILLER_64_954 ();
 sg13g2_fill_2 FILLER_64_961 ();
 sg13g2_decap_4 FILLER_64_986 ();
 sg13g2_fill_1 FILLER_64_1021 ();
 sg13g2_fill_1 FILLER_64_1026 ();
 sg13g2_fill_2 FILLER_64_1041 ();
 sg13g2_fill_1 FILLER_64_1043 ();
 sg13g2_fill_2 FILLER_64_1053 ();
 sg13g2_fill_1 FILLER_64_1060 ();
 sg13g2_fill_2 FILLER_64_1087 ();
 sg13g2_fill_1 FILLER_64_1089 ();
 sg13g2_decap_4 FILLER_64_1124 ();
 sg13g2_fill_1 FILLER_64_1128 ();
 sg13g2_fill_1 FILLER_64_1143 ();
 sg13g2_decap_8 FILLER_64_1148 ();
 sg13g2_fill_2 FILLER_64_1155 ();
 sg13g2_fill_1 FILLER_64_1157 ();
 sg13g2_fill_1 FILLER_64_1184 ();
 sg13g2_fill_2 FILLER_64_1314 ();
 sg13g2_fill_2 FILLER_64_1329 ();
 sg13g2_fill_1 FILLER_64_1339 ();
 sg13g2_decap_8 FILLER_64_1357 ();
 sg13g2_fill_1 FILLER_64_1378 ();
 sg13g2_fill_1 FILLER_64_1462 ();
 sg13g2_fill_1 FILLER_64_1541 ();
 sg13g2_fill_2 FILLER_64_1568 ();
 sg13g2_fill_1 FILLER_64_1570 ();
 sg13g2_fill_1 FILLER_64_1595 ();
 sg13g2_fill_2 FILLER_64_1627 ();
 sg13g2_fill_1 FILLER_64_1665 ();
 sg13g2_fill_2 FILLER_64_1671 ();
 sg13g2_fill_1 FILLER_64_1673 ();
 sg13g2_fill_1 FILLER_64_1700 ();
 sg13g2_fill_2 FILLER_64_1722 ();
 sg13g2_fill_1 FILLER_64_1724 ();
 sg13g2_fill_2 FILLER_64_1740 ();
 sg13g2_fill_1 FILLER_64_1742 ();
 sg13g2_fill_1 FILLER_64_1799 ();
 sg13g2_fill_2 FILLER_64_1870 ();
 sg13g2_fill_1 FILLER_64_1872 ();
 sg13g2_decap_8 FILLER_64_1877 ();
 sg13g2_fill_2 FILLER_64_1989 ();
 sg13g2_fill_1 FILLER_64_1991 ();
 sg13g2_fill_2 FILLER_64_2037 ();
 sg13g2_fill_2 FILLER_64_2048 ();
 sg13g2_fill_2 FILLER_64_2059 ();
 sg13g2_fill_2 FILLER_64_2143 ();
 sg13g2_fill_1 FILLER_64_2145 ();
 sg13g2_decap_8 FILLER_64_2167 ();
 sg13g2_fill_2 FILLER_64_2174 ();
 sg13g2_fill_1 FILLER_64_2189 ();
 sg13g2_decap_4 FILLER_64_2216 ();
 sg13g2_decap_4 FILLER_64_2251 ();
 sg13g2_fill_1 FILLER_64_2295 ();
 sg13g2_decap_8 FILLER_64_2300 ();
 sg13g2_decap_8 FILLER_64_2307 ();
 sg13g2_decap_8 FILLER_64_2314 ();
 sg13g2_decap_8 FILLER_64_2321 ();
 sg13g2_decap_8 FILLER_64_2328 ();
 sg13g2_decap_8 FILLER_64_2335 ();
 sg13g2_decap_8 FILLER_64_2342 ();
 sg13g2_decap_8 FILLER_64_2349 ();
 sg13g2_decap_8 FILLER_64_2356 ();
 sg13g2_decap_8 FILLER_64_2363 ();
 sg13g2_decap_8 FILLER_64_2370 ();
 sg13g2_decap_8 FILLER_64_2377 ();
 sg13g2_decap_8 FILLER_64_2384 ();
 sg13g2_decap_8 FILLER_64_2391 ();
 sg13g2_decap_8 FILLER_64_2398 ();
 sg13g2_decap_8 FILLER_64_2405 ();
 sg13g2_decap_8 FILLER_64_2412 ();
 sg13g2_decap_8 FILLER_64_2419 ();
 sg13g2_decap_8 FILLER_64_2426 ();
 sg13g2_decap_8 FILLER_64_2433 ();
 sg13g2_decap_8 FILLER_64_2440 ();
 sg13g2_decap_8 FILLER_64_2447 ();
 sg13g2_decap_8 FILLER_64_2454 ();
 sg13g2_decap_8 FILLER_64_2461 ();
 sg13g2_decap_8 FILLER_64_2468 ();
 sg13g2_decap_8 FILLER_64_2475 ();
 sg13g2_decap_8 FILLER_64_2482 ();
 sg13g2_decap_8 FILLER_64_2489 ();
 sg13g2_decap_8 FILLER_64_2496 ();
 sg13g2_decap_8 FILLER_64_2503 ();
 sg13g2_decap_8 FILLER_64_2510 ();
 sg13g2_decap_8 FILLER_64_2517 ();
 sg13g2_decap_8 FILLER_64_2524 ();
 sg13g2_decap_8 FILLER_64_2531 ();
 sg13g2_decap_8 FILLER_64_2538 ();
 sg13g2_decap_8 FILLER_64_2545 ();
 sg13g2_decap_8 FILLER_64_2552 ();
 sg13g2_decap_8 FILLER_64_2559 ();
 sg13g2_decap_8 FILLER_64_2566 ();
 sg13g2_decap_8 FILLER_64_2573 ();
 sg13g2_decap_8 FILLER_64_2580 ();
 sg13g2_decap_8 FILLER_64_2587 ();
 sg13g2_decap_8 FILLER_64_2594 ();
 sg13g2_decap_8 FILLER_64_2601 ();
 sg13g2_decap_8 FILLER_64_2608 ();
 sg13g2_decap_8 FILLER_64_2615 ();
 sg13g2_decap_8 FILLER_64_2622 ();
 sg13g2_decap_8 FILLER_64_2629 ();
 sg13g2_decap_8 FILLER_64_2636 ();
 sg13g2_decap_8 FILLER_64_2643 ();
 sg13g2_decap_8 FILLER_64_2650 ();
 sg13g2_decap_8 FILLER_64_2657 ();
 sg13g2_decap_8 FILLER_64_2664 ();
 sg13g2_fill_2 FILLER_64_2671 ();
 sg13g2_fill_1 FILLER_64_2673 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_154 ();
 sg13g2_decap_8 FILLER_65_161 ();
 sg13g2_decap_8 FILLER_65_168 ();
 sg13g2_decap_8 FILLER_65_175 ();
 sg13g2_decap_8 FILLER_65_182 ();
 sg13g2_decap_8 FILLER_65_189 ();
 sg13g2_decap_8 FILLER_65_196 ();
 sg13g2_decap_8 FILLER_65_203 ();
 sg13g2_decap_8 FILLER_65_210 ();
 sg13g2_decap_8 FILLER_65_217 ();
 sg13g2_decap_8 FILLER_65_224 ();
 sg13g2_decap_8 FILLER_65_231 ();
 sg13g2_decap_8 FILLER_65_238 ();
 sg13g2_decap_8 FILLER_65_245 ();
 sg13g2_decap_8 FILLER_65_252 ();
 sg13g2_decap_8 FILLER_65_259 ();
 sg13g2_decap_8 FILLER_65_266 ();
 sg13g2_decap_8 FILLER_65_273 ();
 sg13g2_decap_8 FILLER_65_280 ();
 sg13g2_decap_8 FILLER_65_287 ();
 sg13g2_decap_8 FILLER_65_294 ();
 sg13g2_decap_8 FILLER_65_301 ();
 sg13g2_decap_8 FILLER_65_308 ();
 sg13g2_decap_8 FILLER_65_315 ();
 sg13g2_decap_8 FILLER_65_322 ();
 sg13g2_decap_8 FILLER_65_329 ();
 sg13g2_decap_8 FILLER_65_336 ();
 sg13g2_decap_8 FILLER_65_343 ();
 sg13g2_decap_8 FILLER_65_350 ();
 sg13g2_decap_8 FILLER_65_357 ();
 sg13g2_decap_8 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_371 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_decap_8 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_399 ();
 sg13g2_decap_8 FILLER_65_406 ();
 sg13g2_decap_8 FILLER_65_413 ();
 sg13g2_decap_8 FILLER_65_420 ();
 sg13g2_decap_8 FILLER_65_427 ();
 sg13g2_decap_8 FILLER_65_434 ();
 sg13g2_decap_8 FILLER_65_441 ();
 sg13g2_decap_8 FILLER_65_448 ();
 sg13g2_decap_8 FILLER_65_455 ();
 sg13g2_fill_1 FILLER_65_488 ();
 sg13g2_fill_2 FILLER_65_525 ();
 sg13g2_fill_1 FILLER_65_579 ();
 sg13g2_fill_2 FILLER_65_593 ();
 sg13g2_fill_1 FILLER_65_595 ();
 sg13g2_fill_2 FILLER_65_630 ();
 sg13g2_fill_1 FILLER_65_632 ();
 sg13g2_fill_1 FILLER_65_664 ();
 sg13g2_fill_2 FILLER_65_670 ();
 sg13g2_fill_1 FILLER_65_736 ();
 sg13g2_fill_1 FILLER_65_750 ();
 sg13g2_fill_2 FILLER_65_786 ();
 sg13g2_fill_1 FILLER_65_788 ();
 sg13g2_fill_1 FILLER_65_794 ();
 sg13g2_fill_2 FILLER_65_799 ();
 sg13g2_fill_1 FILLER_65_805 ();
 sg13g2_fill_2 FILLER_65_815 ();
 sg13g2_decap_4 FILLER_65_825 ();
 sg13g2_fill_2 FILLER_65_829 ();
 sg13g2_decap_4 FILLER_65_839 ();
 sg13g2_fill_2 FILLER_65_847 ();
 sg13g2_fill_2 FILLER_65_884 ();
 sg13g2_fill_1 FILLER_65_907 ();
 sg13g2_decap_8 FILLER_65_991 ();
 sg13g2_fill_1 FILLER_65_998 ();
 sg13g2_decap_8 FILLER_65_1065 ();
 sg13g2_fill_1 FILLER_65_1072 ();
 sg13g2_fill_2 FILLER_65_1090 ();
 sg13g2_fill_1 FILLER_65_1092 ();
 sg13g2_fill_2 FILLER_65_1110 ();
 sg13g2_decap_4 FILLER_65_1121 ();
 sg13g2_fill_2 FILLER_65_1125 ();
 sg13g2_fill_2 FILLER_65_1135 ();
 sg13g2_fill_2 FILLER_65_1168 ();
 sg13g2_fill_2 FILLER_65_1189 ();
 sg13g2_fill_1 FILLER_65_1191 ();
 sg13g2_fill_2 FILLER_65_1214 ();
 sg13g2_fill_1 FILLER_65_1241 ();
 sg13g2_fill_2 FILLER_65_1251 ();
 sg13g2_fill_2 FILLER_65_1257 ();
 sg13g2_fill_1 FILLER_65_1259 ();
 sg13g2_fill_1 FILLER_65_1268 ();
 sg13g2_fill_2 FILLER_65_1299 ();
 sg13g2_fill_1 FILLER_65_1301 ();
 sg13g2_decap_8 FILLER_65_1325 ();
 sg13g2_fill_2 FILLER_65_1382 ();
 sg13g2_fill_1 FILLER_65_1384 ();
 sg13g2_decap_4 FILLER_65_1419 ();
 sg13g2_fill_1 FILLER_65_1455 ();
 sg13g2_fill_1 FILLER_65_1487 ();
 sg13g2_fill_2 FILLER_65_1493 ();
 sg13g2_fill_1 FILLER_65_1495 ();
 sg13g2_fill_2 FILLER_65_1505 ();
 sg13g2_decap_4 FILLER_65_1511 ();
 sg13g2_fill_1 FILLER_65_1536 ();
 sg13g2_fill_1 FILLER_65_1558 ();
 sg13g2_fill_2 FILLER_65_1568 ();
 sg13g2_fill_2 FILLER_65_1596 ();
 sg13g2_fill_1 FILLER_65_1598 ();
 sg13g2_fill_2 FILLER_65_1602 ();
 sg13g2_fill_2 FILLER_65_1661 ();
 sg13g2_fill_2 FILLER_65_1685 ();
 sg13g2_fill_1 FILLER_65_1687 ();
 sg13g2_fill_1 FILLER_65_1708 ();
 sg13g2_decap_8 FILLER_65_1764 ();
 sg13g2_decap_4 FILLER_65_1771 ();
 sg13g2_fill_2 FILLER_65_1775 ();
 sg13g2_decap_4 FILLER_65_1785 ();
 sg13g2_fill_2 FILLER_65_1833 ();
 sg13g2_fill_1 FILLER_65_1835 ();
 sg13g2_fill_2 FILLER_65_1841 ();
 sg13g2_fill_1 FILLER_65_1843 ();
 sg13g2_fill_2 FILLER_65_1853 ();
 sg13g2_fill_2 FILLER_65_1881 ();
 sg13g2_fill_1 FILLER_65_1883 ();
 sg13g2_decap_8 FILLER_65_1889 ();
 sg13g2_fill_2 FILLER_65_1896 ();
 sg13g2_fill_2 FILLER_65_1916 ();
 sg13g2_fill_2 FILLER_65_1987 ();
 sg13g2_fill_2 FILLER_65_2053 ();
 sg13g2_fill_1 FILLER_65_2055 ();
 sg13g2_fill_1 FILLER_65_2087 ();
 sg13g2_fill_2 FILLER_65_2097 ();
 sg13g2_fill_1 FILLER_65_2099 ();
 sg13g2_fill_2 FILLER_65_2105 ();
 sg13g2_fill_1 FILLER_65_2107 ();
 sg13g2_fill_2 FILLER_65_2121 ();
 sg13g2_fill_1 FILLER_65_2158 ();
 sg13g2_fill_1 FILLER_65_2164 ();
 sg13g2_fill_2 FILLER_65_2178 ();
 sg13g2_fill_1 FILLER_65_2180 ();
 sg13g2_decap_4 FILLER_65_2190 ();
 sg13g2_fill_2 FILLER_65_2198 ();
 sg13g2_fill_1 FILLER_65_2200 ();
 sg13g2_fill_1 FILLER_65_2205 ();
 sg13g2_decap_4 FILLER_65_2263 ();
 sg13g2_fill_1 FILLER_65_2272 ();
 sg13g2_decap_4 FILLER_65_2277 ();
 sg13g2_decap_8 FILLER_65_2306 ();
 sg13g2_decap_8 FILLER_65_2313 ();
 sg13g2_decap_8 FILLER_65_2320 ();
 sg13g2_decap_8 FILLER_65_2327 ();
 sg13g2_decap_8 FILLER_65_2334 ();
 sg13g2_decap_8 FILLER_65_2341 ();
 sg13g2_decap_8 FILLER_65_2348 ();
 sg13g2_decap_8 FILLER_65_2355 ();
 sg13g2_decap_8 FILLER_65_2362 ();
 sg13g2_decap_8 FILLER_65_2369 ();
 sg13g2_decap_8 FILLER_65_2376 ();
 sg13g2_decap_8 FILLER_65_2383 ();
 sg13g2_decap_8 FILLER_65_2390 ();
 sg13g2_decap_8 FILLER_65_2397 ();
 sg13g2_decap_8 FILLER_65_2404 ();
 sg13g2_decap_8 FILLER_65_2411 ();
 sg13g2_decap_8 FILLER_65_2418 ();
 sg13g2_decap_8 FILLER_65_2425 ();
 sg13g2_decap_8 FILLER_65_2432 ();
 sg13g2_decap_8 FILLER_65_2439 ();
 sg13g2_decap_8 FILLER_65_2446 ();
 sg13g2_decap_8 FILLER_65_2453 ();
 sg13g2_decap_8 FILLER_65_2460 ();
 sg13g2_decap_8 FILLER_65_2467 ();
 sg13g2_decap_8 FILLER_65_2474 ();
 sg13g2_decap_8 FILLER_65_2481 ();
 sg13g2_decap_8 FILLER_65_2488 ();
 sg13g2_decap_8 FILLER_65_2495 ();
 sg13g2_decap_8 FILLER_65_2502 ();
 sg13g2_decap_8 FILLER_65_2509 ();
 sg13g2_decap_8 FILLER_65_2516 ();
 sg13g2_decap_8 FILLER_65_2523 ();
 sg13g2_decap_8 FILLER_65_2530 ();
 sg13g2_decap_8 FILLER_65_2537 ();
 sg13g2_decap_8 FILLER_65_2544 ();
 sg13g2_decap_8 FILLER_65_2551 ();
 sg13g2_decap_8 FILLER_65_2558 ();
 sg13g2_decap_8 FILLER_65_2565 ();
 sg13g2_decap_8 FILLER_65_2572 ();
 sg13g2_decap_8 FILLER_65_2579 ();
 sg13g2_decap_8 FILLER_65_2586 ();
 sg13g2_decap_8 FILLER_65_2593 ();
 sg13g2_decap_8 FILLER_65_2600 ();
 sg13g2_decap_8 FILLER_65_2607 ();
 sg13g2_decap_8 FILLER_65_2614 ();
 sg13g2_decap_8 FILLER_65_2621 ();
 sg13g2_decap_8 FILLER_65_2628 ();
 sg13g2_decap_8 FILLER_65_2635 ();
 sg13g2_decap_8 FILLER_65_2642 ();
 sg13g2_decap_8 FILLER_65_2649 ();
 sg13g2_decap_8 FILLER_65_2656 ();
 sg13g2_decap_8 FILLER_65_2663 ();
 sg13g2_decap_4 FILLER_65_2670 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_decap_8 FILLER_66_147 ();
 sg13g2_decap_8 FILLER_66_154 ();
 sg13g2_decap_8 FILLER_66_161 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_decap_8 FILLER_66_182 ();
 sg13g2_decap_8 FILLER_66_189 ();
 sg13g2_decap_8 FILLER_66_196 ();
 sg13g2_decap_8 FILLER_66_203 ();
 sg13g2_decap_8 FILLER_66_210 ();
 sg13g2_decap_8 FILLER_66_217 ();
 sg13g2_decap_8 FILLER_66_224 ();
 sg13g2_decap_8 FILLER_66_231 ();
 sg13g2_decap_8 FILLER_66_238 ();
 sg13g2_decap_8 FILLER_66_245 ();
 sg13g2_decap_8 FILLER_66_252 ();
 sg13g2_decap_8 FILLER_66_259 ();
 sg13g2_decap_8 FILLER_66_266 ();
 sg13g2_decap_8 FILLER_66_273 ();
 sg13g2_decap_8 FILLER_66_280 ();
 sg13g2_decap_8 FILLER_66_287 ();
 sg13g2_decap_8 FILLER_66_294 ();
 sg13g2_decap_8 FILLER_66_301 ();
 sg13g2_decap_8 FILLER_66_308 ();
 sg13g2_decap_8 FILLER_66_315 ();
 sg13g2_decap_8 FILLER_66_322 ();
 sg13g2_decap_8 FILLER_66_329 ();
 sg13g2_decap_8 FILLER_66_336 ();
 sg13g2_decap_8 FILLER_66_343 ();
 sg13g2_decap_8 FILLER_66_350 ();
 sg13g2_decap_8 FILLER_66_357 ();
 sg13g2_decap_8 FILLER_66_364 ();
 sg13g2_decap_8 FILLER_66_371 ();
 sg13g2_decap_8 FILLER_66_378 ();
 sg13g2_decap_8 FILLER_66_385 ();
 sg13g2_decap_8 FILLER_66_392 ();
 sg13g2_decap_8 FILLER_66_399 ();
 sg13g2_decap_8 FILLER_66_406 ();
 sg13g2_decap_8 FILLER_66_413 ();
 sg13g2_decap_8 FILLER_66_420 ();
 sg13g2_decap_8 FILLER_66_427 ();
 sg13g2_decap_8 FILLER_66_434 ();
 sg13g2_decap_8 FILLER_66_441 ();
 sg13g2_decap_8 FILLER_66_448 ();
 sg13g2_decap_8 FILLER_66_455 ();
 sg13g2_decap_8 FILLER_66_462 ();
 sg13g2_decap_4 FILLER_66_469 ();
 sg13g2_fill_1 FILLER_66_477 ();
 sg13g2_decap_4 FILLER_66_505 ();
 sg13g2_fill_2 FILLER_66_513 ();
 sg13g2_decap_4 FILLER_66_524 ();
 sg13g2_fill_1 FILLER_66_528 ();
 sg13g2_fill_1 FILLER_66_545 ();
 sg13g2_fill_1 FILLER_66_563 ();
 sg13g2_fill_2 FILLER_66_572 ();
 sg13g2_fill_1 FILLER_66_574 ();
 sg13g2_decap_4 FILLER_66_579 ();
 sg13g2_fill_1 FILLER_66_591 ();
 sg13g2_fill_2 FILLER_66_602 ();
 sg13g2_fill_2 FILLER_66_633 ();
 sg13g2_fill_2 FILLER_66_645 ();
 sg13g2_fill_1 FILLER_66_651 ();
 sg13g2_fill_2 FILLER_66_739 ();
 sg13g2_fill_1 FILLER_66_741 ();
 sg13g2_fill_1 FILLER_66_765 ();
 sg13g2_fill_1 FILLER_66_783 ();
 sg13g2_decap_4 FILLER_66_827 ();
 sg13g2_fill_2 FILLER_66_858 ();
 sg13g2_fill_1 FILLER_66_864 ();
 sg13g2_fill_2 FILLER_66_874 ();
 sg13g2_fill_1 FILLER_66_881 ();
 sg13g2_fill_1 FILLER_66_908 ();
 sg13g2_decap_4 FILLER_66_1011 ();
 sg13g2_decap_8 FILLER_66_1019 ();
 sg13g2_decap_8 FILLER_66_1026 ();
 sg13g2_decap_8 FILLER_66_1033 ();
 sg13g2_fill_1 FILLER_66_1040 ();
 sg13g2_fill_2 FILLER_66_1045 ();
 sg13g2_fill_1 FILLER_66_1066 ();
 sg13g2_fill_2 FILLER_66_1129 ();
 sg13g2_fill_1 FILLER_66_1131 ();
 sg13g2_fill_2 FILLER_66_1145 ();
 sg13g2_fill_1 FILLER_66_1151 ();
 sg13g2_fill_2 FILLER_66_1168 ();
 sg13g2_fill_2 FILLER_66_1175 ();
 sg13g2_fill_1 FILLER_66_1212 ();
 sg13g2_fill_1 FILLER_66_1244 ();
 sg13g2_fill_2 FILLER_66_1250 ();
 sg13g2_fill_2 FILLER_66_1256 ();
 sg13g2_decap_8 FILLER_66_1287 ();
 sg13g2_fill_1 FILLER_66_1325 ();
 sg13g2_fill_2 FILLER_66_1361 ();
 sg13g2_fill_1 FILLER_66_1433 ();
 sg13g2_decap_4 FILLER_66_1439 ();
 sg13g2_fill_2 FILLER_66_1443 ();
 sg13g2_fill_2 FILLER_66_1449 ();
 sg13g2_fill_1 FILLER_66_1451 ();
 sg13g2_fill_1 FILLER_66_1462 ();
 sg13g2_fill_1 FILLER_66_1524 ();
 sg13g2_fill_1 FILLER_66_1530 ();
 sg13g2_decap_8 FILLER_66_1588 ();
 sg13g2_fill_2 FILLER_66_1603 ();
 sg13g2_fill_1 FILLER_66_1605 ();
 sg13g2_decap_4 FILLER_66_1616 ();
 sg13g2_fill_1 FILLER_66_1620 ();
 sg13g2_decap_4 FILLER_66_1629 ();
 sg13g2_fill_2 FILLER_66_1637 ();
 sg13g2_fill_1 FILLER_66_1639 ();
 sg13g2_fill_2 FILLER_66_1644 ();
 sg13g2_fill_2 FILLER_66_1687 ();
 sg13g2_fill_1 FILLER_66_1689 ();
 sg13g2_fill_2 FILLER_66_1704 ();
 sg13g2_fill_1 FILLER_66_1711 ();
 sg13g2_fill_1 FILLER_66_1725 ();
 sg13g2_fill_2 FILLER_66_1754 ();
 sg13g2_fill_1 FILLER_66_1756 ();
 sg13g2_fill_2 FILLER_66_1815 ();
 sg13g2_decap_4 FILLER_66_1879 ();
 sg13g2_fill_1 FILLER_66_1909 ();
 sg13g2_fill_2 FILLER_66_1959 ();
 sg13g2_fill_1 FILLER_66_1961 ();
 sg13g2_fill_1 FILLER_66_1969 ();
 sg13g2_fill_2 FILLER_66_2004 ();
 sg13g2_fill_1 FILLER_66_2025 ();
 sg13g2_fill_2 FILLER_66_2048 ();
 sg13g2_fill_2 FILLER_66_2063 ();
 sg13g2_fill_1 FILLER_66_2065 ();
 sg13g2_fill_2 FILLER_66_2089 ();
 sg13g2_fill_2 FILLER_66_2100 ();
 sg13g2_fill_1 FILLER_66_2102 ();
 sg13g2_fill_2 FILLER_66_2162 ();
 sg13g2_fill_1 FILLER_66_2164 ();
 sg13g2_fill_2 FILLER_66_2178 ();
 sg13g2_fill_2 FILLER_66_2210 ();
 sg13g2_fill_1 FILLER_66_2212 ();
 sg13g2_fill_2 FILLER_66_2217 ();
 sg13g2_fill_1 FILLER_66_2228 ();
 sg13g2_fill_2 FILLER_66_2277 ();
 sg13g2_fill_1 FILLER_66_2284 ();
 sg13g2_decap_8 FILLER_66_2320 ();
 sg13g2_decap_8 FILLER_66_2327 ();
 sg13g2_decap_8 FILLER_66_2334 ();
 sg13g2_decap_8 FILLER_66_2341 ();
 sg13g2_decap_8 FILLER_66_2348 ();
 sg13g2_decap_8 FILLER_66_2355 ();
 sg13g2_decap_8 FILLER_66_2362 ();
 sg13g2_decap_8 FILLER_66_2369 ();
 sg13g2_decap_8 FILLER_66_2376 ();
 sg13g2_decap_8 FILLER_66_2383 ();
 sg13g2_decap_8 FILLER_66_2390 ();
 sg13g2_decap_8 FILLER_66_2397 ();
 sg13g2_decap_8 FILLER_66_2404 ();
 sg13g2_decap_8 FILLER_66_2411 ();
 sg13g2_decap_8 FILLER_66_2418 ();
 sg13g2_decap_8 FILLER_66_2425 ();
 sg13g2_decap_8 FILLER_66_2432 ();
 sg13g2_decap_8 FILLER_66_2439 ();
 sg13g2_decap_8 FILLER_66_2446 ();
 sg13g2_decap_8 FILLER_66_2453 ();
 sg13g2_decap_8 FILLER_66_2460 ();
 sg13g2_decap_8 FILLER_66_2467 ();
 sg13g2_decap_8 FILLER_66_2474 ();
 sg13g2_decap_8 FILLER_66_2481 ();
 sg13g2_decap_8 FILLER_66_2488 ();
 sg13g2_decap_8 FILLER_66_2495 ();
 sg13g2_decap_8 FILLER_66_2502 ();
 sg13g2_decap_8 FILLER_66_2509 ();
 sg13g2_decap_8 FILLER_66_2516 ();
 sg13g2_decap_8 FILLER_66_2523 ();
 sg13g2_decap_8 FILLER_66_2530 ();
 sg13g2_decap_8 FILLER_66_2537 ();
 sg13g2_decap_8 FILLER_66_2544 ();
 sg13g2_decap_8 FILLER_66_2551 ();
 sg13g2_decap_8 FILLER_66_2558 ();
 sg13g2_decap_8 FILLER_66_2565 ();
 sg13g2_decap_8 FILLER_66_2572 ();
 sg13g2_decap_8 FILLER_66_2579 ();
 sg13g2_decap_8 FILLER_66_2586 ();
 sg13g2_decap_8 FILLER_66_2593 ();
 sg13g2_decap_8 FILLER_66_2600 ();
 sg13g2_decap_8 FILLER_66_2607 ();
 sg13g2_decap_8 FILLER_66_2614 ();
 sg13g2_decap_8 FILLER_66_2621 ();
 sg13g2_decap_8 FILLER_66_2628 ();
 sg13g2_decap_8 FILLER_66_2635 ();
 sg13g2_decap_8 FILLER_66_2642 ();
 sg13g2_decap_8 FILLER_66_2649 ();
 sg13g2_decap_8 FILLER_66_2656 ();
 sg13g2_decap_8 FILLER_66_2663 ();
 sg13g2_decap_4 FILLER_66_2670 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_decap_8 FILLER_67_161 ();
 sg13g2_decap_8 FILLER_67_168 ();
 sg13g2_decap_8 FILLER_67_175 ();
 sg13g2_decap_8 FILLER_67_182 ();
 sg13g2_decap_8 FILLER_67_189 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_203 ();
 sg13g2_decap_8 FILLER_67_210 ();
 sg13g2_decap_8 FILLER_67_217 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_8 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_238 ();
 sg13g2_decap_8 FILLER_67_245 ();
 sg13g2_decap_8 FILLER_67_252 ();
 sg13g2_decap_8 FILLER_67_259 ();
 sg13g2_decap_8 FILLER_67_266 ();
 sg13g2_decap_8 FILLER_67_273 ();
 sg13g2_decap_8 FILLER_67_280 ();
 sg13g2_decap_8 FILLER_67_287 ();
 sg13g2_decap_8 FILLER_67_294 ();
 sg13g2_decap_8 FILLER_67_301 ();
 sg13g2_decap_8 FILLER_67_308 ();
 sg13g2_decap_8 FILLER_67_315 ();
 sg13g2_decap_8 FILLER_67_322 ();
 sg13g2_decap_8 FILLER_67_329 ();
 sg13g2_decap_8 FILLER_67_336 ();
 sg13g2_decap_8 FILLER_67_343 ();
 sg13g2_decap_8 FILLER_67_350 ();
 sg13g2_decap_8 FILLER_67_357 ();
 sg13g2_decap_8 FILLER_67_364 ();
 sg13g2_decap_8 FILLER_67_371 ();
 sg13g2_decap_8 FILLER_67_378 ();
 sg13g2_decap_8 FILLER_67_385 ();
 sg13g2_decap_8 FILLER_67_392 ();
 sg13g2_decap_8 FILLER_67_399 ();
 sg13g2_decap_8 FILLER_67_406 ();
 sg13g2_decap_8 FILLER_67_413 ();
 sg13g2_decap_8 FILLER_67_420 ();
 sg13g2_decap_8 FILLER_67_427 ();
 sg13g2_decap_8 FILLER_67_434 ();
 sg13g2_decap_8 FILLER_67_441 ();
 sg13g2_decap_8 FILLER_67_448 ();
 sg13g2_decap_8 FILLER_67_455 ();
 sg13g2_decap_8 FILLER_67_462 ();
 sg13g2_decap_8 FILLER_67_469 ();
 sg13g2_fill_1 FILLER_67_476 ();
 sg13g2_fill_2 FILLER_67_486 ();
 sg13g2_decap_4 FILLER_67_541 ();
 sg13g2_fill_1 FILLER_67_545 ();
 sg13g2_fill_1 FILLER_67_551 ();
 sg13g2_decap_4 FILLER_67_592 ();
 sg13g2_fill_2 FILLER_67_622 ();
 sg13g2_fill_1 FILLER_67_624 ();
 sg13g2_fill_1 FILLER_67_687 ();
 sg13g2_fill_1 FILLER_67_700 ();
 sg13g2_fill_2 FILLER_67_709 ();
 sg13g2_fill_1 FILLER_67_729 ();
 sg13g2_fill_1 FILLER_67_761 ();
 sg13g2_fill_2 FILLER_67_798 ();
 sg13g2_fill_1 FILLER_67_800 ();
 sg13g2_fill_2 FILLER_67_858 ();
 sg13g2_fill_2 FILLER_67_903 ();
 sg13g2_fill_2 FILLER_67_938 ();
 sg13g2_fill_1 FILLER_67_940 ();
 sg13g2_fill_2 FILLER_67_967 ();
 sg13g2_fill_1 FILLER_67_969 ();
 sg13g2_decap_4 FILLER_67_995 ();
 sg13g2_decap_8 FILLER_67_1003 ();
 sg13g2_fill_2 FILLER_67_1010 ();
 sg13g2_fill_1 FILLER_67_1012 ();
 sg13g2_fill_1 FILLER_67_1021 ();
 sg13g2_fill_1 FILLER_67_1026 ();
 sg13g2_fill_1 FILLER_67_1053 ();
 sg13g2_fill_2 FILLER_67_1143 ();
 sg13g2_fill_2 FILLER_67_1194 ();
 sg13g2_fill_1 FILLER_67_1226 ();
 sg13g2_decap_8 FILLER_67_1266 ();
 sg13g2_fill_1 FILLER_67_1273 ();
 sg13g2_fill_2 FILLER_67_1305 ();
 sg13g2_fill_1 FILLER_67_1307 ();
 sg13g2_fill_2 FILLER_67_1330 ();
 sg13g2_fill_2 FILLER_67_1366 ();
 sg13g2_fill_1 FILLER_67_1368 ();
 sg13g2_fill_2 FILLER_67_1378 ();
 sg13g2_fill_1 FILLER_67_1380 ();
 sg13g2_fill_2 FILLER_67_1397 ();
 sg13g2_fill_1 FILLER_67_1409 ();
 sg13g2_decap_8 FILLER_67_1471 ();
 sg13g2_fill_2 FILLER_67_1487 ();
 sg13g2_fill_1 FILLER_67_1489 ();
 sg13g2_fill_2 FILLER_67_1508 ();
 sg13g2_fill_1 FILLER_67_1510 ();
 sg13g2_fill_1 FILLER_67_1524 ();
 sg13g2_fill_2 FILLER_67_1551 ();
 sg13g2_fill_2 FILLER_67_1571 ();
 sg13g2_decap_8 FILLER_67_1633 ();
 sg13g2_decap_4 FILLER_67_1640 ();
 sg13g2_fill_2 FILLER_67_1662 ();
 sg13g2_fill_2 FILLER_67_1673 ();
 sg13g2_fill_1 FILLER_67_1675 ();
 sg13g2_fill_2 FILLER_67_1712 ();
 sg13g2_fill_2 FILLER_67_1723 ();
 sg13g2_fill_1 FILLER_67_1725 ();
 sg13g2_decap_4 FILLER_67_1757 ();
 sg13g2_decap_4 FILLER_67_1778 ();
 sg13g2_fill_2 FILLER_67_1791 ();
 sg13g2_decap_4 FILLER_67_1797 ();
 sg13g2_fill_2 FILLER_67_1806 ();
 sg13g2_fill_1 FILLER_67_1808 ();
 sg13g2_decap_4 FILLER_67_1817 ();
 sg13g2_fill_1 FILLER_67_1821 ();
 sg13g2_fill_2 FILLER_67_1836 ();
 sg13g2_fill_1 FILLER_67_1842 ();
 sg13g2_fill_2 FILLER_67_1869 ();
 sg13g2_decap_8 FILLER_67_1899 ();
 sg13g2_decap_4 FILLER_67_1906 ();
 sg13g2_fill_1 FILLER_67_1910 ();
 sg13g2_fill_2 FILLER_67_1943 ();
 sg13g2_fill_2 FILLER_67_1954 ();
 sg13g2_fill_1 FILLER_67_1987 ();
 sg13g2_fill_2 FILLER_67_2006 ();
 sg13g2_fill_1 FILLER_67_2008 ();
 sg13g2_fill_1 FILLER_67_2014 ();
 sg13g2_fill_2 FILLER_67_2054 ();
 sg13g2_fill_1 FILLER_67_2078 ();
 sg13g2_fill_1 FILLER_67_2123 ();
 sg13g2_fill_1 FILLER_67_2137 ();
 sg13g2_fill_2 FILLER_67_2148 ();
 sg13g2_fill_2 FILLER_67_2168 ();
 sg13g2_fill_1 FILLER_67_2170 ();
 sg13g2_fill_2 FILLER_67_2185 ();
 sg13g2_fill_1 FILLER_67_2187 ();
 sg13g2_fill_2 FILLER_67_2267 ();
 sg13g2_decap_8 FILLER_67_2308 ();
 sg13g2_decap_8 FILLER_67_2315 ();
 sg13g2_decap_8 FILLER_67_2322 ();
 sg13g2_decap_8 FILLER_67_2329 ();
 sg13g2_decap_8 FILLER_67_2336 ();
 sg13g2_decap_8 FILLER_67_2343 ();
 sg13g2_decap_8 FILLER_67_2350 ();
 sg13g2_decap_8 FILLER_67_2357 ();
 sg13g2_decap_8 FILLER_67_2364 ();
 sg13g2_decap_8 FILLER_67_2371 ();
 sg13g2_decap_8 FILLER_67_2378 ();
 sg13g2_decap_8 FILLER_67_2385 ();
 sg13g2_decap_8 FILLER_67_2392 ();
 sg13g2_decap_8 FILLER_67_2399 ();
 sg13g2_decap_8 FILLER_67_2406 ();
 sg13g2_decap_8 FILLER_67_2413 ();
 sg13g2_decap_8 FILLER_67_2420 ();
 sg13g2_decap_8 FILLER_67_2427 ();
 sg13g2_decap_8 FILLER_67_2434 ();
 sg13g2_decap_8 FILLER_67_2441 ();
 sg13g2_decap_8 FILLER_67_2448 ();
 sg13g2_decap_8 FILLER_67_2455 ();
 sg13g2_decap_8 FILLER_67_2462 ();
 sg13g2_decap_8 FILLER_67_2469 ();
 sg13g2_decap_8 FILLER_67_2476 ();
 sg13g2_decap_8 FILLER_67_2483 ();
 sg13g2_decap_8 FILLER_67_2490 ();
 sg13g2_decap_8 FILLER_67_2497 ();
 sg13g2_decap_8 FILLER_67_2504 ();
 sg13g2_decap_8 FILLER_67_2511 ();
 sg13g2_decap_8 FILLER_67_2518 ();
 sg13g2_decap_8 FILLER_67_2525 ();
 sg13g2_decap_8 FILLER_67_2532 ();
 sg13g2_decap_8 FILLER_67_2539 ();
 sg13g2_decap_8 FILLER_67_2546 ();
 sg13g2_decap_8 FILLER_67_2553 ();
 sg13g2_decap_8 FILLER_67_2560 ();
 sg13g2_decap_8 FILLER_67_2567 ();
 sg13g2_decap_8 FILLER_67_2574 ();
 sg13g2_decap_8 FILLER_67_2581 ();
 sg13g2_decap_8 FILLER_67_2588 ();
 sg13g2_decap_8 FILLER_67_2595 ();
 sg13g2_decap_8 FILLER_67_2602 ();
 sg13g2_decap_8 FILLER_67_2609 ();
 sg13g2_decap_8 FILLER_67_2616 ();
 sg13g2_decap_8 FILLER_67_2623 ();
 sg13g2_decap_8 FILLER_67_2630 ();
 sg13g2_decap_8 FILLER_67_2637 ();
 sg13g2_decap_8 FILLER_67_2644 ();
 sg13g2_decap_8 FILLER_67_2651 ();
 sg13g2_decap_8 FILLER_67_2658 ();
 sg13g2_decap_8 FILLER_67_2665 ();
 sg13g2_fill_2 FILLER_67_2672 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_decap_8 FILLER_68_154 ();
 sg13g2_decap_8 FILLER_68_161 ();
 sg13g2_decap_8 FILLER_68_168 ();
 sg13g2_decap_8 FILLER_68_175 ();
 sg13g2_decap_8 FILLER_68_182 ();
 sg13g2_decap_8 FILLER_68_189 ();
 sg13g2_decap_8 FILLER_68_196 ();
 sg13g2_decap_8 FILLER_68_203 ();
 sg13g2_decap_8 FILLER_68_210 ();
 sg13g2_decap_8 FILLER_68_217 ();
 sg13g2_decap_8 FILLER_68_224 ();
 sg13g2_decap_8 FILLER_68_231 ();
 sg13g2_decap_8 FILLER_68_238 ();
 sg13g2_decap_8 FILLER_68_245 ();
 sg13g2_decap_8 FILLER_68_252 ();
 sg13g2_decap_8 FILLER_68_259 ();
 sg13g2_decap_8 FILLER_68_266 ();
 sg13g2_decap_8 FILLER_68_273 ();
 sg13g2_decap_8 FILLER_68_280 ();
 sg13g2_decap_8 FILLER_68_287 ();
 sg13g2_decap_8 FILLER_68_294 ();
 sg13g2_decap_8 FILLER_68_301 ();
 sg13g2_decap_8 FILLER_68_308 ();
 sg13g2_decap_8 FILLER_68_315 ();
 sg13g2_decap_8 FILLER_68_322 ();
 sg13g2_decap_8 FILLER_68_329 ();
 sg13g2_decap_8 FILLER_68_336 ();
 sg13g2_decap_8 FILLER_68_343 ();
 sg13g2_decap_8 FILLER_68_350 ();
 sg13g2_decap_8 FILLER_68_357 ();
 sg13g2_decap_8 FILLER_68_364 ();
 sg13g2_decap_8 FILLER_68_371 ();
 sg13g2_decap_8 FILLER_68_378 ();
 sg13g2_decap_8 FILLER_68_385 ();
 sg13g2_decap_8 FILLER_68_392 ();
 sg13g2_decap_8 FILLER_68_399 ();
 sg13g2_decap_8 FILLER_68_406 ();
 sg13g2_decap_8 FILLER_68_413 ();
 sg13g2_decap_8 FILLER_68_420 ();
 sg13g2_decap_8 FILLER_68_427 ();
 sg13g2_decap_8 FILLER_68_434 ();
 sg13g2_decap_8 FILLER_68_441 ();
 sg13g2_decap_8 FILLER_68_448 ();
 sg13g2_decap_8 FILLER_68_455 ();
 sg13g2_fill_1 FILLER_68_462 ();
 sg13g2_fill_1 FILLER_68_498 ();
 sg13g2_fill_1 FILLER_68_517 ();
 sg13g2_fill_1 FILLER_68_561 ();
 sg13g2_fill_1 FILLER_68_601 ();
 sg13g2_decap_4 FILLER_68_611 ();
 sg13g2_fill_1 FILLER_68_615 ();
 sg13g2_fill_1 FILLER_68_638 ();
 sg13g2_fill_1 FILLER_68_647 ();
 sg13g2_fill_1 FILLER_68_661 ();
 sg13g2_fill_2 FILLER_68_675 ();
 sg13g2_fill_1 FILLER_68_686 ();
 sg13g2_fill_2 FILLER_68_718 ();
 sg13g2_fill_1 FILLER_68_720 ();
 sg13g2_fill_1 FILLER_68_738 ();
 sg13g2_fill_2 FILLER_68_743 ();
 sg13g2_fill_1 FILLER_68_749 ();
 sg13g2_decap_4 FILLER_68_759 ();
 sg13g2_decap_4 FILLER_68_780 ();
 sg13g2_decap_4 FILLER_68_819 ();
 sg13g2_fill_1 FILLER_68_828 ();
 sg13g2_fill_1 FILLER_68_883 ();
 sg13g2_fill_2 FILLER_68_889 ();
 sg13g2_decap_8 FILLER_68_904 ();
 sg13g2_fill_1 FILLER_68_911 ();
 sg13g2_decap_8 FILLER_68_920 ();
 sg13g2_decap_4 FILLER_68_932 ();
 sg13g2_fill_2 FILLER_68_936 ();
 sg13g2_fill_2 FILLER_68_968 ();
 sg13g2_fill_1 FILLER_68_1026 ();
 sg13g2_fill_1 FILLER_68_1040 ();
 sg13g2_fill_1 FILLER_68_1050 ();
 sg13g2_fill_1 FILLER_68_1055 ();
 sg13g2_decap_4 FILLER_68_1061 ();
 sg13g2_fill_2 FILLER_68_1065 ();
 sg13g2_fill_2 FILLER_68_1092 ();
 sg13g2_fill_2 FILLER_68_1107 ();
 sg13g2_fill_1 FILLER_68_1126 ();
 sg13g2_decap_4 FILLER_68_1245 ();
 sg13g2_fill_2 FILLER_68_1249 ();
 sg13g2_decap_4 FILLER_68_1259 ();
 sg13g2_fill_2 FILLER_68_1267 ();
 sg13g2_fill_1 FILLER_68_1269 ();
 sg13g2_fill_1 FILLER_68_1274 ();
 sg13g2_fill_2 FILLER_68_1283 ();
 sg13g2_fill_2 FILLER_68_1305 ();
 sg13g2_fill_2 FILLER_68_1323 ();
 sg13g2_fill_1 FILLER_68_1325 ();
 sg13g2_fill_2 FILLER_68_1352 ();
 sg13g2_decap_4 FILLER_68_1359 ();
 sg13g2_fill_2 FILLER_68_1443 ();
 sg13g2_fill_2 FILLER_68_1468 ();
 sg13g2_fill_1 FILLER_68_1496 ();
 sg13g2_fill_1 FILLER_68_1523 ();
 sg13g2_fill_2 FILLER_68_1567 ();
 sg13g2_fill_1 FILLER_68_1569 ();
 sg13g2_fill_2 FILLER_68_1617 ();
 sg13g2_fill_1 FILLER_68_1619 ();
 sg13g2_fill_1 FILLER_68_1660 ();
 sg13g2_fill_2 FILLER_68_1666 ();
 sg13g2_fill_2 FILLER_68_1676 ();
 sg13g2_fill_1 FILLER_68_1692 ();
 sg13g2_decap_8 FILLER_68_1702 ();
 sg13g2_fill_1 FILLER_68_1747 ();
 sg13g2_fill_1 FILLER_68_1753 ();
 sg13g2_decap_4 FILLER_68_1763 ();
 sg13g2_fill_2 FILLER_68_1767 ();
 sg13g2_decap_4 FILLER_68_1830 ();
 sg13g2_fill_1 FILLER_68_1838 ();
 sg13g2_fill_2 FILLER_68_1844 ();
 sg13g2_fill_2 FILLER_68_1851 ();
 sg13g2_fill_1 FILLER_68_1853 ();
 sg13g2_fill_1 FILLER_68_1906 ();
 sg13g2_fill_2 FILLER_68_1933 ();
 sg13g2_fill_2 FILLER_68_1961 ();
 sg13g2_fill_1 FILLER_68_1963 ();
 sg13g2_fill_2 FILLER_68_2056 ();
 sg13g2_fill_2 FILLER_68_2093 ();
 sg13g2_decap_4 FILLER_68_2108 ();
 sg13g2_fill_1 FILLER_68_2117 ();
 sg13g2_fill_2 FILLER_68_2122 ();
 sg13g2_fill_1 FILLER_68_2129 ();
 sg13g2_fill_1 FILLER_68_2231 ();
 sg13g2_fill_2 FILLER_68_2266 ();
 sg13g2_fill_1 FILLER_68_2268 ();
 sg13g2_decap_8 FILLER_68_2295 ();
 sg13g2_decap_8 FILLER_68_2302 ();
 sg13g2_decap_8 FILLER_68_2309 ();
 sg13g2_decap_8 FILLER_68_2316 ();
 sg13g2_decap_8 FILLER_68_2323 ();
 sg13g2_decap_8 FILLER_68_2330 ();
 sg13g2_decap_8 FILLER_68_2337 ();
 sg13g2_decap_8 FILLER_68_2344 ();
 sg13g2_decap_8 FILLER_68_2351 ();
 sg13g2_decap_8 FILLER_68_2358 ();
 sg13g2_decap_8 FILLER_68_2365 ();
 sg13g2_decap_8 FILLER_68_2372 ();
 sg13g2_decap_8 FILLER_68_2379 ();
 sg13g2_decap_8 FILLER_68_2386 ();
 sg13g2_decap_8 FILLER_68_2393 ();
 sg13g2_decap_8 FILLER_68_2400 ();
 sg13g2_decap_8 FILLER_68_2407 ();
 sg13g2_decap_8 FILLER_68_2414 ();
 sg13g2_decap_8 FILLER_68_2421 ();
 sg13g2_decap_8 FILLER_68_2428 ();
 sg13g2_decap_8 FILLER_68_2435 ();
 sg13g2_decap_8 FILLER_68_2442 ();
 sg13g2_decap_8 FILLER_68_2449 ();
 sg13g2_decap_8 FILLER_68_2456 ();
 sg13g2_decap_8 FILLER_68_2463 ();
 sg13g2_decap_8 FILLER_68_2470 ();
 sg13g2_decap_8 FILLER_68_2477 ();
 sg13g2_decap_8 FILLER_68_2484 ();
 sg13g2_decap_8 FILLER_68_2491 ();
 sg13g2_decap_8 FILLER_68_2498 ();
 sg13g2_decap_8 FILLER_68_2505 ();
 sg13g2_decap_8 FILLER_68_2512 ();
 sg13g2_decap_8 FILLER_68_2519 ();
 sg13g2_decap_8 FILLER_68_2526 ();
 sg13g2_decap_8 FILLER_68_2533 ();
 sg13g2_decap_8 FILLER_68_2540 ();
 sg13g2_decap_8 FILLER_68_2547 ();
 sg13g2_decap_8 FILLER_68_2554 ();
 sg13g2_decap_8 FILLER_68_2561 ();
 sg13g2_decap_8 FILLER_68_2568 ();
 sg13g2_decap_8 FILLER_68_2575 ();
 sg13g2_decap_8 FILLER_68_2582 ();
 sg13g2_decap_8 FILLER_68_2589 ();
 sg13g2_decap_8 FILLER_68_2596 ();
 sg13g2_decap_8 FILLER_68_2603 ();
 sg13g2_decap_8 FILLER_68_2610 ();
 sg13g2_decap_8 FILLER_68_2617 ();
 sg13g2_decap_8 FILLER_68_2624 ();
 sg13g2_decap_8 FILLER_68_2631 ();
 sg13g2_decap_8 FILLER_68_2638 ();
 sg13g2_decap_8 FILLER_68_2645 ();
 sg13g2_decap_8 FILLER_68_2652 ();
 sg13g2_decap_8 FILLER_68_2659 ();
 sg13g2_decap_8 FILLER_68_2666 ();
 sg13g2_fill_1 FILLER_68_2673 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_decap_8 FILLER_69_147 ();
 sg13g2_decap_8 FILLER_69_154 ();
 sg13g2_decap_8 FILLER_69_161 ();
 sg13g2_decap_8 FILLER_69_168 ();
 sg13g2_decap_8 FILLER_69_175 ();
 sg13g2_decap_8 FILLER_69_182 ();
 sg13g2_decap_8 FILLER_69_189 ();
 sg13g2_decap_8 FILLER_69_196 ();
 sg13g2_decap_8 FILLER_69_203 ();
 sg13g2_decap_8 FILLER_69_210 ();
 sg13g2_decap_8 FILLER_69_217 ();
 sg13g2_decap_8 FILLER_69_224 ();
 sg13g2_decap_8 FILLER_69_231 ();
 sg13g2_decap_8 FILLER_69_238 ();
 sg13g2_decap_8 FILLER_69_245 ();
 sg13g2_decap_8 FILLER_69_252 ();
 sg13g2_decap_8 FILLER_69_259 ();
 sg13g2_decap_8 FILLER_69_266 ();
 sg13g2_decap_8 FILLER_69_273 ();
 sg13g2_decap_8 FILLER_69_280 ();
 sg13g2_decap_8 FILLER_69_287 ();
 sg13g2_decap_8 FILLER_69_294 ();
 sg13g2_decap_8 FILLER_69_301 ();
 sg13g2_decap_8 FILLER_69_308 ();
 sg13g2_decap_8 FILLER_69_315 ();
 sg13g2_decap_8 FILLER_69_322 ();
 sg13g2_decap_8 FILLER_69_329 ();
 sg13g2_decap_8 FILLER_69_336 ();
 sg13g2_decap_8 FILLER_69_343 ();
 sg13g2_decap_8 FILLER_69_350 ();
 sg13g2_decap_8 FILLER_69_357 ();
 sg13g2_decap_8 FILLER_69_364 ();
 sg13g2_decap_8 FILLER_69_371 ();
 sg13g2_decap_8 FILLER_69_378 ();
 sg13g2_decap_8 FILLER_69_385 ();
 sg13g2_decap_8 FILLER_69_392 ();
 sg13g2_decap_8 FILLER_69_399 ();
 sg13g2_decap_8 FILLER_69_406 ();
 sg13g2_decap_8 FILLER_69_413 ();
 sg13g2_decap_8 FILLER_69_420 ();
 sg13g2_decap_8 FILLER_69_427 ();
 sg13g2_decap_8 FILLER_69_434 ();
 sg13g2_decap_8 FILLER_69_441 ();
 sg13g2_decap_8 FILLER_69_448 ();
 sg13g2_decap_8 FILLER_69_455 ();
 sg13g2_decap_8 FILLER_69_462 ();
 sg13g2_decap_4 FILLER_69_469 ();
 sg13g2_fill_1 FILLER_69_473 ();
 sg13g2_decap_8 FILLER_69_478 ();
 sg13g2_decap_4 FILLER_69_485 ();
 sg13g2_fill_1 FILLER_69_489 ();
 sg13g2_fill_2 FILLER_69_533 ();
 sg13g2_fill_1 FILLER_69_535 ();
 sg13g2_fill_2 FILLER_69_552 ();
 sg13g2_fill_1 FILLER_69_554 ();
 sg13g2_fill_2 FILLER_69_581 ();
 sg13g2_decap_4 FILLER_69_618 ();
 sg13g2_fill_1 FILLER_69_622 ();
 sg13g2_fill_2 FILLER_69_633 ();
 sg13g2_fill_2 FILLER_69_666 ();
 sg13g2_fill_1 FILLER_69_681 ();
 sg13g2_fill_1 FILLER_69_698 ();
 sg13g2_fill_2 FILLER_69_760 ();
 sg13g2_fill_1 FILLER_69_862 ();
 sg13g2_decap_8 FILLER_69_867 ();
 sg13g2_decap_4 FILLER_69_874 ();
 sg13g2_decap_8 FILLER_69_913 ();
 sg13g2_fill_2 FILLER_69_920 ();
 sg13g2_fill_2 FILLER_69_944 ();
 sg13g2_fill_1 FILLER_69_946 ();
 sg13g2_fill_1 FILLER_69_978 ();
 sg13g2_fill_2 FILLER_69_988 ();
 sg13g2_fill_1 FILLER_69_990 ();
 sg13g2_fill_2 FILLER_69_1004 ();
 sg13g2_fill_1 FILLER_69_1006 ();
 sg13g2_decap_4 FILLER_69_1142 ();
 sg13g2_fill_1 FILLER_69_1146 ();
 sg13g2_decap_8 FILLER_69_1151 ();
 sg13g2_fill_1 FILLER_69_1158 ();
 sg13g2_fill_1 FILLER_69_1185 ();
 sg13g2_fill_2 FILLER_69_1200 ();
 sg13g2_fill_1 FILLER_69_1202 ();
 sg13g2_fill_2 FILLER_69_1211 ();
 sg13g2_fill_1 FILLER_69_1234 ();
 sg13g2_fill_1 FILLER_69_1248 ();
 sg13g2_decap_4 FILLER_69_1285 ();
 sg13g2_fill_2 FILLER_69_1329 ();
 sg13g2_decap_4 FILLER_69_1340 ();
 sg13g2_fill_1 FILLER_69_1344 ();
 sg13g2_decap_8 FILLER_69_1358 ();
 sg13g2_fill_1 FILLER_69_1423 ();
 sg13g2_fill_1 FILLER_69_1450 ();
 sg13g2_fill_2 FILLER_69_1477 ();
 sg13g2_fill_1 FILLER_69_1479 ();
 sg13g2_fill_2 FILLER_69_1498 ();
 sg13g2_fill_1 FILLER_69_1500 ();
 sg13g2_fill_1 FILLER_69_1535 ();
 sg13g2_fill_1 FILLER_69_1567 ();
 sg13g2_decap_8 FILLER_69_1591 ();
 sg13g2_fill_2 FILLER_69_1598 ();
 sg13g2_fill_1 FILLER_69_1600 ();
 sg13g2_fill_1 FILLER_69_1623 ();
 sg13g2_fill_2 FILLER_69_1629 ();
 sg13g2_fill_1 FILLER_69_1631 ();
 sg13g2_fill_1 FILLER_69_1640 ();
 sg13g2_fill_2 FILLER_69_1659 ();
 sg13g2_fill_1 FILLER_69_1661 ();
 sg13g2_fill_1 FILLER_69_1697 ();
 sg13g2_decap_8 FILLER_69_1712 ();
 sg13g2_fill_2 FILLER_69_1740 ();
 sg13g2_fill_2 FILLER_69_1785 ();
 sg13g2_fill_1 FILLER_69_1787 ();
 sg13g2_fill_2 FILLER_69_1798 ();
 sg13g2_fill_1 FILLER_69_1800 ();
 sg13g2_fill_2 FILLER_69_1810 ();
 sg13g2_fill_1 FILLER_69_1812 ();
 sg13g2_fill_2 FILLER_69_1844 ();
 sg13g2_fill_1 FILLER_69_1846 ();
 sg13g2_fill_2 FILLER_69_1866 ();
 sg13g2_fill_1 FILLER_69_1868 ();
 sg13g2_fill_2 FILLER_69_1894 ();
 sg13g2_fill_1 FILLER_69_1896 ();
 sg13g2_fill_2 FILLER_69_1906 ();
 sg13g2_fill_1 FILLER_69_1935 ();
 sg13g2_fill_2 FILLER_69_1962 ();
 sg13g2_fill_2 FILLER_69_1969 ();
 sg13g2_fill_1 FILLER_69_1971 ();
 sg13g2_fill_1 FILLER_69_1994 ();
 sg13g2_fill_2 FILLER_69_1999 ();
 sg13g2_fill_2 FILLER_69_2014 ();
 sg13g2_fill_2 FILLER_69_2021 ();
 sg13g2_fill_1 FILLER_69_2023 ();
 sg13g2_fill_2 FILLER_69_2051 ();
 sg13g2_fill_1 FILLER_69_2058 ();
 sg13g2_fill_1 FILLER_69_2069 ();
 sg13g2_fill_1 FILLER_69_2091 ();
 sg13g2_decap_8 FILLER_69_2144 ();
 sg13g2_fill_2 FILLER_69_2163 ();
 sg13g2_decap_8 FILLER_69_2192 ();
 sg13g2_fill_2 FILLER_69_2199 ();
 sg13g2_decap_4 FILLER_69_2209 ();
 sg13g2_fill_2 FILLER_69_2243 ();
 sg13g2_fill_1 FILLER_69_2245 ();
 sg13g2_fill_1 FILLER_69_2256 ();
 sg13g2_fill_2 FILLER_69_2266 ();
 sg13g2_decap_8 FILLER_69_2304 ();
 sg13g2_decap_8 FILLER_69_2311 ();
 sg13g2_decap_8 FILLER_69_2318 ();
 sg13g2_decap_8 FILLER_69_2325 ();
 sg13g2_decap_8 FILLER_69_2332 ();
 sg13g2_decap_8 FILLER_69_2339 ();
 sg13g2_decap_8 FILLER_69_2346 ();
 sg13g2_decap_8 FILLER_69_2353 ();
 sg13g2_decap_8 FILLER_69_2360 ();
 sg13g2_decap_8 FILLER_69_2367 ();
 sg13g2_decap_8 FILLER_69_2374 ();
 sg13g2_decap_8 FILLER_69_2381 ();
 sg13g2_decap_8 FILLER_69_2388 ();
 sg13g2_decap_8 FILLER_69_2395 ();
 sg13g2_decap_8 FILLER_69_2402 ();
 sg13g2_decap_8 FILLER_69_2409 ();
 sg13g2_decap_8 FILLER_69_2416 ();
 sg13g2_decap_8 FILLER_69_2423 ();
 sg13g2_decap_8 FILLER_69_2430 ();
 sg13g2_decap_8 FILLER_69_2437 ();
 sg13g2_decap_8 FILLER_69_2444 ();
 sg13g2_decap_8 FILLER_69_2451 ();
 sg13g2_decap_8 FILLER_69_2458 ();
 sg13g2_decap_8 FILLER_69_2465 ();
 sg13g2_decap_8 FILLER_69_2472 ();
 sg13g2_decap_8 FILLER_69_2479 ();
 sg13g2_decap_8 FILLER_69_2486 ();
 sg13g2_decap_8 FILLER_69_2493 ();
 sg13g2_decap_8 FILLER_69_2500 ();
 sg13g2_decap_8 FILLER_69_2507 ();
 sg13g2_decap_8 FILLER_69_2514 ();
 sg13g2_decap_8 FILLER_69_2521 ();
 sg13g2_decap_8 FILLER_69_2528 ();
 sg13g2_decap_8 FILLER_69_2535 ();
 sg13g2_decap_8 FILLER_69_2542 ();
 sg13g2_decap_8 FILLER_69_2549 ();
 sg13g2_decap_8 FILLER_69_2556 ();
 sg13g2_decap_8 FILLER_69_2563 ();
 sg13g2_decap_8 FILLER_69_2570 ();
 sg13g2_decap_8 FILLER_69_2577 ();
 sg13g2_decap_8 FILLER_69_2584 ();
 sg13g2_decap_8 FILLER_69_2591 ();
 sg13g2_decap_8 FILLER_69_2598 ();
 sg13g2_decap_8 FILLER_69_2605 ();
 sg13g2_decap_8 FILLER_69_2612 ();
 sg13g2_decap_8 FILLER_69_2619 ();
 sg13g2_decap_8 FILLER_69_2626 ();
 sg13g2_decap_8 FILLER_69_2633 ();
 sg13g2_decap_8 FILLER_69_2640 ();
 sg13g2_decap_8 FILLER_69_2647 ();
 sg13g2_decap_8 FILLER_69_2654 ();
 sg13g2_decap_8 FILLER_69_2661 ();
 sg13g2_decap_4 FILLER_69_2668 ();
 sg13g2_fill_2 FILLER_69_2672 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_decap_8 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_182 ();
 sg13g2_decap_8 FILLER_70_189 ();
 sg13g2_decap_8 FILLER_70_196 ();
 sg13g2_decap_8 FILLER_70_203 ();
 sg13g2_decap_8 FILLER_70_210 ();
 sg13g2_decap_8 FILLER_70_217 ();
 sg13g2_decap_8 FILLER_70_224 ();
 sg13g2_decap_8 FILLER_70_231 ();
 sg13g2_decap_8 FILLER_70_238 ();
 sg13g2_decap_8 FILLER_70_245 ();
 sg13g2_decap_8 FILLER_70_252 ();
 sg13g2_decap_8 FILLER_70_259 ();
 sg13g2_decap_8 FILLER_70_266 ();
 sg13g2_decap_8 FILLER_70_273 ();
 sg13g2_decap_8 FILLER_70_280 ();
 sg13g2_decap_8 FILLER_70_287 ();
 sg13g2_decap_8 FILLER_70_294 ();
 sg13g2_decap_8 FILLER_70_301 ();
 sg13g2_decap_8 FILLER_70_308 ();
 sg13g2_decap_8 FILLER_70_315 ();
 sg13g2_decap_8 FILLER_70_322 ();
 sg13g2_decap_8 FILLER_70_329 ();
 sg13g2_decap_8 FILLER_70_336 ();
 sg13g2_decap_8 FILLER_70_343 ();
 sg13g2_decap_8 FILLER_70_350 ();
 sg13g2_decap_8 FILLER_70_357 ();
 sg13g2_decap_8 FILLER_70_364 ();
 sg13g2_decap_8 FILLER_70_371 ();
 sg13g2_decap_8 FILLER_70_378 ();
 sg13g2_decap_8 FILLER_70_385 ();
 sg13g2_decap_8 FILLER_70_392 ();
 sg13g2_decap_8 FILLER_70_399 ();
 sg13g2_decap_8 FILLER_70_406 ();
 sg13g2_decap_8 FILLER_70_413 ();
 sg13g2_decap_8 FILLER_70_420 ();
 sg13g2_decap_8 FILLER_70_427 ();
 sg13g2_decap_8 FILLER_70_434 ();
 sg13g2_decap_8 FILLER_70_441 ();
 sg13g2_decap_8 FILLER_70_448 ();
 sg13g2_decap_8 FILLER_70_455 ();
 sg13g2_decap_8 FILLER_70_462 ();
 sg13g2_decap_8 FILLER_70_469 ();
 sg13g2_decap_4 FILLER_70_476 ();
 sg13g2_fill_2 FILLER_70_480 ();
 sg13g2_fill_2 FILLER_70_522 ();
 sg13g2_fill_2 FILLER_70_550 ();
 sg13g2_decap_4 FILLER_70_561 ();
 sg13g2_fill_1 FILLER_70_609 ();
 sg13g2_fill_2 FILLER_70_645 ();
 sg13g2_fill_1 FILLER_70_647 ();
 sg13g2_fill_1 FILLER_70_657 ();
 sg13g2_fill_1 FILLER_70_692 ();
 sg13g2_decap_8 FILLER_70_702 ();
 sg13g2_decap_8 FILLER_70_709 ();
 sg13g2_decap_4 FILLER_70_716 ();
 sg13g2_fill_2 FILLER_70_725 ();
 sg13g2_fill_2 FILLER_70_732 ();
 sg13g2_fill_1 FILLER_70_734 ();
 sg13g2_decap_4 FILLER_70_749 ();
 sg13g2_fill_2 FILLER_70_753 ();
 sg13g2_fill_2 FILLER_70_764 ();
 sg13g2_fill_1 FILLER_70_797 ();
 sg13g2_fill_1 FILLER_70_825 ();
 sg13g2_fill_1 FILLER_70_882 ();
 sg13g2_fill_2 FILLER_70_892 ();
 sg13g2_fill_2 FILLER_70_934 ();
 sg13g2_fill_2 FILLER_70_971 ();
 sg13g2_fill_2 FILLER_70_1021 ();
 sg13g2_fill_1 FILLER_70_1023 ();
 sg13g2_fill_1 FILLER_70_1042 ();
 sg13g2_fill_2 FILLER_70_1078 ();
 sg13g2_fill_2 FILLER_70_1112 ();
 sg13g2_fill_1 FILLER_70_1114 ();
 sg13g2_decap_4 FILLER_70_1124 ();
 sg13g2_fill_1 FILLER_70_1132 ();
 sg13g2_decap_4 FILLER_70_1148 ();
 sg13g2_fill_1 FILLER_70_1152 ();
 sg13g2_fill_2 FILLER_70_1157 ();
 sg13g2_fill_1 FILLER_70_1159 ();
 sg13g2_fill_1 FILLER_70_1186 ();
 sg13g2_fill_1 FILLER_70_1213 ();
 sg13g2_fill_2 FILLER_70_1235 ();
 sg13g2_fill_2 FILLER_70_1263 ();
 sg13g2_fill_1 FILLER_70_1265 ();
 sg13g2_fill_1 FILLER_70_1284 ();
 sg13g2_fill_2 FILLER_70_1290 ();
 sg13g2_decap_8 FILLER_70_1301 ();
 sg13g2_fill_2 FILLER_70_1334 ();
 sg13g2_fill_1 FILLER_70_1345 ();
 sg13g2_fill_1 FILLER_70_1381 ();
 sg13g2_decap_4 FILLER_70_1387 ();
 sg13g2_fill_2 FILLER_70_1404 ();
 sg13g2_decap_4 FILLER_70_1409 ();
 sg13g2_fill_1 FILLER_70_1413 ();
 sg13g2_decap_4 FILLER_70_1423 ();
 sg13g2_fill_2 FILLER_70_1427 ();
 sg13g2_fill_1 FILLER_70_1433 ();
 sg13g2_fill_2 FILLER_70_1438 ();
 sg13g2_fill_2 FILLER_70_1449 ();
 sg13g2_fill_2 FILLER_70_1503 ();
 sg13g2_fill_1 FILLER_70_1505 ();
 sg13g2_fill_2 FILLER_70_1549 ();
 sg13g2_fill_2 FILLER_70_1561 ();
 sg13g2_fill_2 FILLER_70_1624 ();
 sg13g2_fill_1 FILLER_70_1630 ();
 sg13g2_fill_2 FILLER_70_1636 ();
 sg13g2_fill_1 FILLER_70_1638 ();
 sg13g2_decap_8 FILLER_70_1669 ();
 sg13g2_decap_8 FILLER_70_1676 ();
 sg13g2_fill_2 FILLER_70_1718 ();
 sg13g2_fill_2 FILLER_70_1751 ();
 sg13g2_fill_1 FILLER_70_1787 ();
 sg13g2_fill_2 FILLER_70_1802 ();
 sg13g2_fill_2 FILLER_70_1856 ();
 sg13g2_fill_1 FILLER_70_1872 ();
 sg13g2_fill_2 FILLER_70_1886 ();
 sg13g2_fill_2 FILLER_70_1913 ();
 sg13g2_decap_4 FILLER_70_1920 ();
 sg13g2_fill_2 FILLER_70_1924 ();
 sg13g2_fill_2 FILLER_70_1943 ();
 sg13g2_fill_1 FILLER_70_1945 ();
 sg13g2_fill_1 FILLER_70_1958 ();
 sg13g2_fill_1 FILLER_70_1963 ();
 sg13g2_decap_8 FILLER_70_1990 ();
 sg13g2_fill_2 FILLER_70_1997 ();
 sg13g2_decap_4 FILLER_70_2006 ();
 sg13g2_fill_1 FILLER_70_2010 ();
 sg13g2_fill_1 FILLER_70_2047 ();
 sg13g2_fill_2 FILLER_70_2067 ();
 sg13g2_decap_4 FILLER_70_2095 ();
 sg13g2_fill_2 FILLER_70_2161 ();
 sg13g2_fill_1 FILLER_70_2163 ();
 sg13g2_fill_1 FILLER_70_2211 ();
 sg13g2_fill_1 FILLER_70_2221 ();
 sg13g2_fill_2 FILLER_70_2244 ();
 sg13g2_fill_1 FILLER_70_2246 ();
 sg13g2_fill_2 FILLER_70_2251 ();
 sg13g2_fill_1 FILLER_70_2253 ();
 sg13g2_decap_8 FILLER_70_2311 ();
 sg13g2_decap_8 FILLER_70_2318 ();
 sg13g2_decap_8 FILLER_70_2325 ();
 sg13g2_decap_8 FILLER_70_2332 ();
 sg13g2_decap_8 FILLER_70_2339 ();
 sg13g2_decap_8 FILLER_70_2346 ();
 sg13g2_decap_8 FILLER_70_2353 ();
 sg13g2_decap_8 FILLER_70_2360 ();
 sg13g2_decap_8 FILLER_70_2367 ();
 sg13g2_decap_8 FILLER_70_2374 ();
 sg13g2_decap_8 FILLER_70_2381 ();
 sg13g2_decap_8 FILLER_70_2388 ();
 sg13g2_decap_8 FILLER_70_2395 ();
 sg13g2_decap_8 FILLER_70_2402 ();
 sg13g2_decap_8 FILLER_70_2409 ();
 sg13g2_decap_8 FILLER_70_2416 ();
 sg13g2_decap_8 FILLER_70_2423 ();
 sg13g2_decap_8 FILLER_70_2430 ();
 sg13g2_decap_8 FILLER_70_2437 ();
 sg13g2_decap_8 FILLER_70_2444 ();
 sg13g2_decap_8 FILLER_70_2451 ();
 sg13g2_decap_8 FILLER_70_2458 ();
 sg13g2_decap_8 FILLER_70_2465 ();
 sg13g2_decap_8 FILLER_70_2472 ();
 sg13g2_decap_8 FILLER_70_2479 ();
 sg13g2_decap_8 FILLER_70_2486 ();
 sg13g2_decap_8 FILLER_70_2493 ();
 sg13g2_decap_8 FILLER_70_2500 ();
 sg13g2_decap_8 FILLER_70_2507 ();
 sg13g2_decap_8 FILLER_70_2514 ();
 sg13g2_decap_8 FILLER_70_2521 ();
 sg13g2_decap_8 FILLER_70_2528 ();
 sg13g2_decap_8 FILLER_70_2535 ();
 sg13g2_decap_8 FILLER_70_2542 ();
 sg13g2_decap_8 FILLER_70_2549 ();
 sg13g2_decap_8 FILLER_70_2556 ();
 sg13g2_decap_8 FILLER_70_2563 ();
 sg13g2_decap_8 FILLER_70_2570 ();
 sg13g2_decap_8 FILLER_70_2577 ();
 sg13g2_decap_8 FILLER_70_2584 ();
 sg13g2_decap_8 FILLER_70_2591 ();
 sg13g2_decap_8 FILLER_70_2598 ();
 sg13g2_decap_8 FILLER_70_2605 ();
 sg13g2_decap_8 FILLER_70_2612 ();
 sg13g2_decap_8 FILLER_70_2619 ();
 sg13g2_decap_8 FILLER_70_2626 ();
 sg13g2_decap_8 FILLER_70_2633 ();
 sg13g2_decap_8 FILLER_70_2640 ();
 sg13g2_decap_8 FILLER_70_2647 ();
 sg13g2_decap_8 FILLER_70_2654 ();
 sg13g2_decap_8 FILLER_70_2661 ();
 sg13g2_decap_4 FILLER_70_2668 ();
 sg13g2_fill_2 FILLER_70_2672 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_8 FILLER_71_154 ();
 sg13g2_decap_8 FILLER_71_161 ();
 sg13g2_decap_8 FILLER_71_168 ();
 sg13g2_decap_8 FILLER_71_175 ();
 sg13g2_decap_8 FILLER_71_182 ();
 sg13g2_decap_8 FILLER_71_189 ();
 sg13g2_decap_8 FILLER_71_196 ();
 sg13g2_decap_8 FILLER_71_203 ();
 sg13g2_decap_8 FILLER_71_210 ();
 sg13g2_decap_8 FILLER_71_217 ();
 sg13g2_decap_8 FILLER_71_224 ();
 sg13g2_decap_8 FILLER_71_231 ();
 sg13g2_decap_8 FILLER_71_238 ();
 sg13g2_decap_8 FILLER_71_245 ();
 sg13g2_decap_8 FILLER_71_252 ();
 sg13g2_decap_8 FILLER_71_259 ();
 sg13g2_decap_8 FILLER_71_266 ();
 sg13g2_decap_8 FILLER_71_273 ();
 sg13g2_decap_8 FILLER_71_280 ();
 sg13g2_decap_8 FILLER_71_287 ();
 sg13g2_decap_8 FILLER_71_294 ();
 sg13g2_decap_8 FILLER_71_301 ();
 sg13g2_decap_8 FILLER_71_308 ();
 sg13g2_decap_8 FILLER_71_315 ();
 sg13g2_decap_8 FILLER_71_322 ();
 sg13g2_decap_8 FILLER_71_329 ();
 sg13g2_decap_8 FILLER_71_336 ();
 sg13g2_decap_8 FILLER_71_343 ();
 sg13g2_decap_8 FILLER_71_350 ();
 sg13g2_decap_8 FILLER_71_357 ();
 sg13g2_decap_8 FILLER_71_364 ();
 sg13g2_decap_8 FILLER_71_371 ();
 sg13g2_decap_8 FILLER_71_378 ();
 sg13g2_decap_8 FILLER_71_385 ();
 sg13g2_decap_8 FILLER_71_392 ();
 sg13g2_decap_8 FILLER_71_399 ();
 sg13g2_decap_8 FILLER_71_406 ();
 sg13g2_decap_8 FILLER_71_413 ();
 sg13g2_decap_8 FILLER_71_420 ();
 sg13g2_decap_8 FILLER_71_427 ();
 sg13g2_decap_8 FILLER_71_434 ();
 sg13g2_decap_8 FILLER_71_441 ();
 sg13g2_decap_8 FILLER_71_448 ();
 sg13g2_decap_8 FILLER_71_455 ();
 sg13g2_decap_8 FILLER_71_462 ();
 sg13g2_decap_8 FILLER_71_469 ();
 sg13g2_decap_8 FILLER_71_476 ();
 sg13g2_decap_4 FILLER_71_483 ();
 sg13g2_fill_2 FILLER_71_487 ();
 sg13g2_decap_8 FILLER_71_521 ();
 sg13g2_fill_2 FILLER_71_528 ();
 sg13g2_fill_2 FILLER_71_588 ();
 sg13g2_fill_2 FILLER_71_603 ();
 sg13g2_decap_8 FILLER_71_614 ();
 sg13g2_fill_2 FILLER_71_625 ();
 sg13g2_decap_4 FILLER_71_632 ();
 sg13g2_fill_2 FILLER_71_680 ();
 sg13g2_fill_1 FILLER_71_783 ();
 sg13g2_fill_1 FILLER_71_865 ();
 sg13g2_fill_2 FILLER_71_870 ();
 sg13g2_decap_4 FILLER_71_890 ();
 sg13g2_fill_2 FILLER_71_917 ();
 sg13g2_fill_2 FILLER_71_928 ();
 sg13g2_fill_1 FILLER_71_930 ();
 sg13g2_decap_8 FILLER_71_935 ();
 sg13g2_decap_4 FILLER_71_942 ();
 sg13g2_fill_1 FILLER_71_946 ();
 sg13g2_fill_1 FILLER_71_959 ();
 sg13g2_fill_1 FILLER_71_983 ();
 sg13g2_fill_2 FILLER_71_1002 ();
 sg13g2_fill_1 FILLER_71_1004 ();
 sg13g2_fill_1 FILLER_71_1083 ();
 sg13g2_fill_2 FILLER_71_1197 ();
 sg13g2_fill_1 FILLER_71_1199 ();
 sg13g2_fill_2 FILLER_71_1204 ();
 sg13g2_decap_8 FILLER_71_1232 ();
 sg13g2_fill_1 FILLER_71_1239 ();
 sg13g2_fill_1 FILLER_71_1249 ();
 sg13g2_fill_1 FILLER_71_1280 ();
 sg13g2_fill_2 FILLER_71_1312 ();
 sg13g2_fill_2 FILLER_71_1319 ();
 sg13g2_fill_1 FILLER_71_1400 ();
 sg13g2_fill_2 FILLER_71_1405 ();
 sg13g2_decap_8 FILLER_71_1434 ();
 sg13g2_decap_4 FILLER_71_1441 ();
 sg13g2_fill_2 FILLER_71_1491 ();
 sg13g2_fill_2 FILLER_71_1530 ();
 sg13g2_fill_1 FILLER_71_1532 ();
 sg13g2_fill_1 FILLER_71_1589 ();
 sg13g2_fill_1 FILLER_71_1594 ();
 sg13g2_fill_2 FILLER_71_1613 ();
 sg13g2_fill_1 FILLER_71_1664 ();
 sg13g2_fill_1 FILLER_71_1700 ();
 sg13g2_fill_2 FILLER_71_1718 ();
 sg13g2_decap_4 FILLER_71_1739 ();
 sg13g2_decap_4 FILLER_71_1769 ();
 sg13g2_fill_1 FILLER_71_1799 ();
 sg13g2_fill_2 FILLER_71_1840 ();
 sg13g2_fill_1 FILLER_71_1842 ();
 sg13g2_fill_1 FILLER_71_1869 ();
 sg13g2_fill_2 FILLER_71_1896 ();
 sg13g2_fill_2 FILLER_71_1955 ();
 sg13g2_fill_2 FILLER_71_1970 ();
 sg13g2_fill_1 FILLER_71_1972 ();
 sg13g2_fill_1 FILLER_71_1983 ();
 sg13g2_decap_8 FILLER_71_2013 ();
 sg13g2_fill_2 FILLER_71_2020 ();
 sg13g2_fill_1 FILLER_71_2026 ();
 sg13g2_fill_2 FILLER_71_2032 ();
 sg13g2_fill_1 FILLER_71_2034 ();
 sg13g2_fill_2 FILLER_71_2040 ();
 sg13g2_fill_2 FILLER_71_2047 ();
 sg13g2_decap_4 FILLER_71_2075 ();
 sg13g2_fill_1 FILLER_71_2079 ();
 sg13g2_decap_4 FILLER_71_2085 ();
 sg13g2_decap_4 FILLER_71_2093 ();
 sg13g2_fill_1 FILLER_71_2097 ();
 sg13g2_decap_4 FILLER_71_2112 ();
 sg13g2_fill_2 FILLER_71_2147 ();
 sg13g2_fill_2 FILLER_71_2184 ();
 sg13g2_fill_1 FILLER_71_2186 ();
 sg13g2_fill_2 FILLER_71_2205 ();
 sg13g2_decap_4 FILLER_71_2216 ();
 sg13g2_fill_2 FILLER_71_2225 ();
 sg13g2_fill_2 FILLER_71_2235 ();
 sg13g2_fill_2 FILLER_71_2262 ();
 sg13g2_fill_1 FILLER_71_2264 ();
 sg13g2_fill_1 FILLER_71_2292 ();
 sg13g2_decap_8 FILLER_71_2306 ();
 sg13g2_decap_8 FILLER_71_2313 ();
 sg13g2_decap_8 FILLER_71_2320 ();
 sg13g2_decap_8 FILLER_71_2327 ();
 sg13g2_decap_8 FILLER_71_2334 ();
 sg13g2_decap_8 FILLER_71_2341 ();
 sg13g2_decap_8 FILLER_71_2348 ();
 sg13g2_decap_8 FILLER_71_2355 ();
 sg13g2_decap_8 FILLER_71_2362 ();
 sg13g2_decap_8 FILLER_71_2369 ();
 sg13g2_decap_8 FILLER_71_2376 ();
 sg13g2_decap_8 FILLER_71_2383 ();
 sg13g2_decap_8 FILLER_71_2390 ();
 sg13g2_decap_8 FILLER_71_2397 ();
 sg13g2_decap_8 FILLER_71_2404 ();
 sg13g2_decap_8 FILLER_71_2411 ();
 sg13g2_decap_8 FILLER_71_2418 ();
 sg13g2_decap_8 FILLER_71_2425 ();
 sg13g2_decap_8 FILLER_71_2432 ();
 sg13g2_decap_8 FILLER_71_2439 ();
 sg13g2_decap_8 FILLER_71_2446 ();
 sg13g2_decap_8 FILLER_71_2453 ();
 sg13g2_decap_8 FILLER_71_2460 ();
 sg13g2_decap_8 FILLER_71_2467 ();
 sg13g2_decap_8 FILLER_71_2474 ();
 sg13g2_decap_8 FILLER_71_2481 ();
 sg13g2_decap_8 FILLER_71_2488 ();
 sg13g2_decap_8 FILLER_71_2495 ();
 sg13g2_decap_8 FILLER_71_2502 ();
 sg13g2_decap_8 FILLER_71_2509 ();
 sg13g2_decap_8 FILLER_71_2516 ();
 sg13g2_decap_8 FILLER_71_2523 ();
 sg13g2_decap_8 FILLER_71_2530 ();
 sg13g2_decap_8 FILLER_71_2537 ();
 sg13g2_decap_8 FILLER_71_2544 ();
 sg13g2_decap_8 FILLER_71_2551 ();
 sg13g2_decap_8 FILLER_71_2558 ();
 sg13g2_decap_8 FILLER_71_2565 ();
 sg13g2_decap_8 FILLER_71_2572 ();
 sg13g2_decap_8 FILLER_71_2579 ();
 sg13g2_decap_8 FILLER_71_2586 ();
 sg13g2_decap_8 FILLER_71_2593 ();
 sg13g2_decap_8 FILLER_71_2600 ();
 sg13g2_decap_8 FILLER_71_2607 ();
 sg13g2_decap_8 FILLER_71_2614 ();
 sg13g2_decap_8 FILLER_71_2621 ();
 sg13g2_decap_8 FILLER_71_2628 ();
 sg13g2_decap_8 FILLER_71_2635 ();
 sg13g2_decap_8 FILLER_71_2642 ();
 sg13g2_decap_8 FILLER_71_2649 ();
 sg13g2_decap_8 FILLER_71_2656 ();
 sg13g2_decap_8 FILLER_71_2663 ();
 sg13g2_decap_4 FILLER_71_2670 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_decap_8 FILLER_72_168 ();
 sg13g2_decap_8 FILLER_72_175 ();
 sg13g2_decap_8 FILLER_72_182 ();
 sg13g2_decap_8 FILLER_72_189 ();
 sg13g2_decap_8 FILLER_72_196 ();
 sg13g2_decap_8 FILLER_72_203 ();
 sg13g2_decap_8 FILLER_72_210 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_decap_8 FILLER_72_224 ();
 sg13g2_decap_8 FILLER_72_231 ();
 sg13g2_decap_8 FILLER_72_238 ();
 sg13g2_decap_8 FILLER_72_245 ();
 sg13g2_decap_8 FILLER_72_252 ();
 sg13g2_decap_8 FILLER_72_259 ();
 sg13g2_decap_8 FILLER_72_266 ();
 sg13g2_decap_8 FILLER_72_273 ();
 sg13g2_decap_8 FILLER_72_280 ();
 sg13g2_decap_8 FILLER_72_287 ();
 sg13g2_decap_8 FILLER_72_294 ();
 sg13g2_decap_8 FILLER_72_301 ();
 sg13g2_decap_8 FILLER_72_308 ();
 sg13g2_decap_8 FILLER_72_315 ();
 sg13g2_decap_8 FILLER_72_322 ();
 sg13g2_decap_8 FILLER_72_329 ();
 sg13g2_decap_8 FILLER_72_336 ();
 sg13g2_decap_8 FILLER_72_343 ();
 sg13g2_decap_8 FILLER_72_350 ();
 sg13g2_decap_8 FILLER_72_357 ();
 sg13g2_decap_8 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_371 ();
 sg13g2_decap_8 FILLER_72_378 ();
 sg13g2_decap_8 FILLER_72_385 ();
 sg13g2_decap_8 FILLER_72_392 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_decap_8 FILLER_72_406 ();
 sg13g2_decap_8 FILLER_72_413 ();
 sg13g2_decap_8 FILLER_72_420 ();
 sg13g2_decap_8 FILLER_72_427 ();
 sg13g2_decap_8 FILLER_72_434 ();
 sg13g2_decap_8 FILLER_72_441 ();
 sg13g2_decap_8 FILLER_72_448 ();
 sg13g2_decap_8 FILLER_72_455 ();
 sg13g2_decap_8 FILLER_72_462 ();
 sg13g2_decap_8 FILLER_72_469 ();
 sg13g2_decap_8 FILLER_72_476 ();
 sg13g2_decap_8 FILLER_72_483 ();
 sg13g2_fill_2 FILLER_72_490 ();
 sg13g2_fill_1 FILLER_72_492 ();
 sg13g2_decap_4 FILLER_72_501 ();
 sg13g2_fill_1 FILLER_72_515 ();
 sg13g2_decap_8 FILLER_72_521 ();
 sg13g2_fill_2 FILLER_72_528 ();
 sg13g2_decap_4 FILLER_72_539 ();
 sg13g2_fill_2 FILLER_72_552 ();
 sg13g2_fill_1 FILLER_72_558 ();
 sg13g2_fill_2 FILLER_72_563 ();
 sg13g2_fill_1 FILLER_72_565 ();
 sg13g2_fill_2 FILLER_72_618 ();
 sg13g2_fill_1 FILLER_72_620 ();
 sg13g2_fill_1 FILLER_72_673 ();
 sg13g2_fill_2 FILLER_72_691 ();
 sg13g2_fill_1 FILLER_72_693 ();
 sg13g2_fill_2 FILLER_72_729 ();
 sg13g2_fill_1 FILLER_72_740 ();
 sg13g2_fill_1 FILLER_72_756 ();
 sg13g2_fill_2 FILLER_72_828 ();
 sg13g2_fill_2 FILLER_72_870 ();
 sg13g2_fill_2 FILLER_72_906 ();
 sg13g2_fill_2 FILLER_72_916 ();
 sg13g2_fill_2 FILLER_72_992 ();
 sg13g2_fill_2 FILLER_72_1029 ();
 sg13g2_fill_1 FILLER_72_1031 ();
 sg13g2_fill_2 FILLER_72_1049 ();
 sg13g2_fill_1 FILLER_72_1097 ();
 sg13g2_decap_8 FILLER_72_1103 ();
 sg13g2_fill_2 FILLER_72_1110 ();
 sg13g2_fill_2 FILLER_72_1124 ();
 sg13g2_fill_2 FILLER_72_1140 ();
 sg13g2_fill_1 FILLER_72_1142 ();
 sg13g2_decap_8 FILLER_72_1156 ();
 sg13g2_decap_4 FILLER_72_1163 ();
 sg13g2_fill_1 FILLER_72_1167 ();
 sg13g2_decap_4 FILLER_72_1172 ();
 sg13g2_fill_1 FILLER_72_1176 ();
 sg13g2_fill_1 FILLER_72_1185 ();
 sg13g2_fill_2 FILLER_72_1200 ();
 sg13g2_decap_4 FILLER_72_1216 ();
 sg13g2_fill_2 FILLER_72_1229 ();
 sg13g2_fill_1 FILLER_72_1293 ();
 sg13g2_fill_1 FILLER_72_1303 ();
 sg13g2_fill_2 FILLER_72_1322 ();
 sg13g2_fill_1 FILLER_72_1329 ();
 sg13g2_fill_1 FILLER_72_1339 ();
 sg13g2_decap_8 FILLER_72_1344 ();
 sg13g2_decap_4 FILLER_72_1351 ();
 sg13g2_fill_2 FILLER_72_1355 ();
 sg13g2_fill_1 FILLER_72_1362 ();
 sg13g2_fill_1 FILLER_72_1389 ();
 sg13g2_fill_1 FILLER_72_1416 ();
 sg13g2_fill_2 FILLER_72_1504 ();
 sg13g2_fill_1 FILLER_72_1506 ();
 sg13g2_fill_2 FILLER_72_1546 ();
 sg13g2_fill_2 FILLER_72_1557 ();
 sg13g2_fill_1 FILLER_72_1568 ();
 sg13g2_fill_2 FILLER_72_1578 ();
 sg13g2_fill_1 FILLER_72_1580 ();
 sg13g2_fill_1 FILLER_72_1589 ();
 sg13g2_fill_1 FILLER_72_1599 ();
 sg13g2_fill_2 FILLER_72_1604 ();
 sg13g2_fill_1 FILLER_72_1606 ();
 sg13g2_fill_2 FILLER_72_1611 ();
 sg13g2_fill_1 FILLER_72_1613 ();
 sg13g2_fill_2 FILLER_72_1628 ();
 sg13g2_fill_1 FILLER_72_1630 ();
 sg13g2_fill_1 FILLER_72_1644 ();
 sg13g2_fill_1 FILLER_72_1671 ();
 sg13g2_fill_2 FILLER_72_1677 ();
 sg13g2_fill_1 FILLER_72_1679 ();
 sg13g2_fill_2 FILLER_72_1693 ();
 sg13g2_fill_1 FILLER_72_1695 ();
 sg13g2_fill_2 FILLER_72_1704 ();
 sg13g2_fill_1 FILLER_72_1706 ();
 sg13g2_fill_2 FILLER_72_1755 ();
 sg13g2_fill_1 FILLER_72_1757 ();
 sg13g2_decap_4 FILLER_72_1800 ();
 sg13g2_fill_1 FILLER_72_1804 ();
 sg13g2_fill_1 FILLER_72_1810 ();
 sg13g2_decap_4 FILLER_72_1815 ();
 sg13g2_fill_2 FILLER_72_1819 ();
 sg13g2_decap_4 FILLER_72_1860 ();
 sg13g2_fill_2 FILLER_72_1864 ();
 sg13g2_fill_1 FILLER_72_1897 ();
 sg13g2_fill_1 FILLER_72_1925 ();
 sg13g2_fill_2 FILLER_72_1930 ();
 sg13g2_fill_2 FILLER_72_2007 ();
 sg13g2_fill_1 FILLER_72_2009 ();
 sg13g2_fill_2 FILLER_72_2023 ();
 sg13g2_fill_1 FILLER_72_2051 ();
 sg13g2_fill_1 FILLER_72_2079 ();
 sg13g2_fill_2 FILLER_72_2144 ();
 sg13g2_fill_2 FILLER_72_2172 ();
 sg13g2_fill_1 FILLER_72_2174 ();
 sg13g2_decap_4 FILLER_72_2211 ();
 sg13g2_fill_1 FILLER_72_2246 ();
 sg13g2_decap_8 FILLER_72_2287 ();
 sg13g2_decap_8 FILLER_72_2294 ();
 sg13g2_decap_8 FILLER_72_2301 ();
 sg13g2_decap_8 FILLER_72_2308 ();
 sg13g2_decap_8 FILLER_72_2315 ();
 sg13g2_decap_8 FILLER_72_2322 ();
 sg13g2_decap_8 FILLER_72_2329 ();
 sg13g2_decap_8 FILLER_72_2336 ();
 sg13g2_decap_8 FILLER_72_2343 ();
 sg13g2_decap_8 FILLER_72_2350 ();
 sg13g2_decap_8 FILLER_72_2357 ();
 sg13g2_decap_8 FILLER_72_2364 ();
 sg13g2_decap_8 FILLER_72_2371 ();
 sg13g2_decap_8 FILLER_72_2378 ();
 sg13g2_decap_8 FILLER_72_2385 ();
 sg13g2_decap_8 FILLER_72_2392 ();
 sg13g2_decap_8 FILLER_72_2399 ();
 sg13g2_decap_8 FILLER_72_2406 ();
 sg13g2_decap_8 FILLER_72_2413 ();
 sg13g2_decap_8 FILLER_72_2420 ();
 sg13g2_decap_8 FILLER_72_2427 ();
 sg13g2_decap_8 FILLER_72_2434 ();
 sg13g2_decap_8 FILLER_72_2441 ();
 sg13g2_decap_8 FILLER_72_2448 ();
 sg13g2_decap_8 FILLER_72_2455 ();
 sg13g2_decap_8 FILLER_72_2462 ();
 sg13g2_decap_8 FILLER_72_2469 ();
 sg13g2_decap_8 FILLER_72_2476 ();
 sg13g2_decap_8 FILLER_72_2483 ();
 sg13g2_decap_8 FILLER_72_2490 ();
 sg13g2_decap_8 FILLER_72_2497 ();
 sg13g2_decap_8 FILLER_72_2504 ();
 sg13g2_decap_8 FILLER_72_2511 ();
 sg13g2_decap_8 FILLER_72_2518 ();
 sg13g2_decap_8 FILLER_72_2525 ();
 sg13g2_decap_8 FILLER_72_2532 ();
 sg13g2_decap_8 FILLER_72_2539 ();
 sg13g2_decap_8 FILLER_72_2546 ();
 sg13g2_decap_8 FILLER_72_2553 ();
 sg13g2_decap_8 FILLER_72_2560 ();
 sg13g2_decap_8 FILLER_72_2567 ();
 sg13g2_decap_8 FILLER_72_2574 ();
 sg13g2_decap_8 FILLER_72_2581 ();
 sg13g2_decap_8 FILLER_72_2588 ();
 sg13g2_decap_8 FILLER_72_2595 ();
 sg13g2_decap_8 FILLER_72_2602 ();
 sg13g2_decap_8 FILLER_72_2609 ();
 sg13g2_decap_8 FILLER_72_2616 ();
 sg13g2_decap_8 FILLER_72_2623 ();
 sg13g2_decap_8 FILLER_72_2630 ();
 sg13g2_decap_8 FILLER_72_2637 ();
 sg13g2_decap_8 FILLER_72_2644 ();
 sg13g2_decap_8 FILLER_72_2651 ();
 sg13g2_decap_8 FILLER_72_2658 ();
 sg13g2_decap_8 FILLER_72_2665 ();
 sg13g2_fill_2 FILLER_72_2672 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_decap_8 FILLER_73_175 ();
 sg13g2_decap_8 FILLER_73_182 ();
 sg13g2_decap_8 FILLER_73_189 ();
 sg13g2_decap_8 FILLER_73_196 ();
 sg13g2_decap_8 FILLER_73_203 ();
 sg13g2_decap_8 FILLER_73_210 ();
 sg13g2_decap_8 FILLER_73_217 ();
 sg13g2_decap_8 FILLER_73_224 ();
 sg13g2_decap_8 FILLER_73_231 ();
 sg13g2_decap_8 FILLER_73_238 ();
 sg13g2_decap_8 FILLER_73_245 ();
 sg13g2_decap_8 FILLER_73_252 ();
 sg13g2_decap_8 FILLER_73_259 ();
 sg13g2_decap_8 FILLER_73_266 ();
 sg13g2_decap_8 FILLER_73_273 ();
 sg13g2_decap_8 FILLER_73_280 ();
 sg13g2_decap_8 FILLER_73_287 ();
 sg13g2_decap_8 FILLER_73_294 ();
 sg13g2_decap_8 FILLER_73_301 ();
 sg13g2_decap_8 FILLER_73_308 ();
 sg13g2_decap_8 FILLER_73_315 ();
 sg13g2_decap_8 FILLER_73_322 ();
 sg13g2_decap_8 FILLER_73_329 ();
 sg13g2_decap_8 FILLER_73_336 ();
 sg13g2_decap_8 FILLER_73_343 ();
 sg13g2_decap_8 FILLER_73_350 ();
 sg13g2_decap_8 FILLER_73_357 ();
 sg13g2_decap_8 FILLER_73_364 ();
 sg13g2_decap_8 FILLER_73_371 ();
 sg13g2_decap_8 FILLER_73_378 ();
 sg13g2_decap_8 FILLER_73_385 ();
 sg13g2_decap_8 FILLER_73_392 ();
 sg13g2_decap_8 FILLER_73_399 ();
 sg13g2_decap_8 FILLER_73_406 ();
 sg13g2_decap_8 FILLER_73_413 ();
 sg13g2_decap_8 FILLER_73_420 ();
 sg13g2_decap_8 FILLER_73_427 ();
 sg13g2_decap_8 FILLER_73_434 ();
 sg13g2_decap_8 FILLER_73_441 ();
 sg13g2_decap_8 FILLER_73_448 ();
 sg13g2_decap_8 FILLER_73_455 ();
 sg13g2_decap_8 FILLER_73_462 ();
 sg13g2_decap_8 FILLER_73_469 ();
 sg13g2_decap_8 FILLER_73_476 ();
 sg13g2_fill_2 FILLER_73_483 ();
 sg13g2_fill_1 FILLER_73_485 ();
 sg13g2_fill_2 FILLER_73_512 ();
 sg13g2_fill_1 FILLER_73_545 ();
 sg13g2_fill_2 FILLER_73_554 ();
 sg13g2_fill_1 FILLER_73_561 ();
 sg13g2_fill_2 FILLER_73_567 ();
 sg13g2_fill_1 FILLER_73_569 ();
 sg13g2_fill_2 FILLER_73_595 ();
 sg13g2_fill_2 FILLER_73_659 ();
 sg13g2_fill_2 FILLER_73_675 ();
 sg13g2_fill_2 FILLER_73_696 ();
 sg13g2_fill_1 FILLER_73_698 ();
 sg13g2_decap_4 FILLER_73_759 ();
 sg13g2_decap_4 FILLER_73_768 ();
 sg13g2_fill_2 FILLER_73_772 ();
 sg13g2_fill_2 FILLER_73_798 ();
 sg13g2_fill_1 FILLER_73_809 ();
 sg13g2_decap_4 FILLER_73_870 ();
 sg13g2_fill_2 FILLER_73_874 ();
 sg13g2_fill_2 FILLER_73_901 ();
 sg13g2_fill_2 FILLER_73_930 ();
 sg13g2_decap_8 FILLER_73_950 ();
 sg13g2_fill_1 FILLER_73_957 ();
 sg13g2_fill_2 FILLER_73_988 ();
 sg13g2_fill_2 FILLER_73_1021 ();
 sg13g2_fill_1 FILLER_73_1023 ();
 sg13g2_fill_2 FILLER_73_1028 ();
 sg13g2_fill_2 FILLER_73_1039 ();
 sg13g2_fill_1 FILLER_73_1098 ();
 sg13g2_decap_8 FILLER_73_1168 ();
 sg13g2_fill_1 FILLER_73_1209 ();
 sg13g2_fill_2 FILLER_73_1250 ();
 sg13g2_fill_1 FILLER_73_1252 ();
 sg13g2_fill_2 FILLER_73_1267 ();
 sg13g2_fill_2 FILLER_73_1287 ();
 sg13g2_fill_1 FILLER_73_1289 ();
 sg13g2_fill_2 FILLER_73_1316 ();
 sg13g2_fill_2 FILLER_73_1378 ();
 sg13g2_fill_1 FILLER_73_1380 ();
 sg13g2_fill_2 FILLER_73_1399 ();
 sg13g2_decap_4 FILLER_73_1406 ();
 sg13g2_decap_8 FILLER_73_1415 ();
 sg13g2_decap_4 FILLER_73_1422 ();
 sg13g2_fill_2 FILLER_73_1439 ();
 sg13g2_fill_1 FILLER_73_1441 ();
 sg13g2_fill_2 FILLER_73_1464 ();
 sg13g2_fill_2 FILLER_73_1485 ();
 sg13g2_fill_1 FILLER_73_1487 ();
 sg13g2_fill_1 FILLER_73_1549 ();
 sg13g2_fill_2 FILLER_73_1581 ();
 sg13g2_fill_1 FILLER_73_1583 ();
 sg13g2_fill_1 FILLER_73_1641 ();
 sg13g2_fill_1 FILLER_73_1673 ();
 sg13g2_fill_2 FILLER_73_1683 ();
 sg13g2_fill_1 FILLER_73_1685 ();
 sg13g2_fill_1 FILLER_73_1709 ();
 sg13g2_fill_1 FILLER_73_1727 ();
 sg13g2_fill_1 FILLER_73_1759 ();
 sg13g2_fill_2 FILLER_73_1804 ();
 sg13g2_fill_2 FILLER_73_1819 ();
 sg13g2_fill_1 FILLER_73_1821 ();
 sg13g2_fill_2 FILLER_73_1839 ();
 sg13g2_decap_4 FILLER_73_1850 ();
 sg13g2_fill_1 FILLER_73_1854 ();
 sg13g2_fill_1 FILLER_73_1860 ();
 sg13g2_fill_1 FILLER_73_1865 ();
 sg13g2_fill_1 FILLER_73_1883 ();
 sg13g2_fill_2 FILLER_73_1940 ();
 sg13g2_fill_2 FILLER_73_1946 ();
 sg13g2_fill_1 FILLER_73_1948 ();
 sg13g2_fill_2 FILLER_73_1964 ();
 sg13g2_decap_4 FILLER_73_2027 ();
 sg13g2_fill_1 FILLER_73_2053 ();
 sg13g2_fill_2 FILLER_73_2080 ();
 sg13g2_fill_1 FILLER_73_2082 ();
 sg13g2_fill_2 FILLER_73_2088 ();
 sg13g2_decap_8 FILLER_73_2102 ();
 sg13g2_fill_2 FILLER_73_2113 ();
 sg13g2_fill_1 FILLER_73_2115 ();
 sg13g2_fill_1 FILLER_73_2120 ();
 sg13g2_fill_2 FILLER_73_2130 ();
 sg13g2_fill_2 FILLER_73_2146 ();
 sg13g2_fill_1 FILLER_73_2157 ();
 sg13g2_fill_2 FILLER_73_2180 ();
 sg13g2_fill_1 FILLER_73_2182 ();
 sg13g2_fill_2 FILLER_73_2197 ();
 sg13g2_decap_4 FILLER_73_2212 ();
 sg13g2_decap_8 FILLER_73_2237 ();
 sg13g2_fill_2 FILLER_73_2244 ();
 sg13g2_fill_2 FILLER_73_2250 ();
 sg13g2_decap_8 FILLER_73_2265 ();
 sg13g2_decap_8 FILLER_73_2276 ();
 sg13g2_decap_8 FILLER_73_2283 ();
 sg13g2_decap_8 FILLER_73_2290 ();
 sg13g2_decap_8 FILLER_73_2297 ();
 sg13g2_decap_8 FILLER_73_2304 ();
 sg13g2_decap_8 FILLER_73_2311 ();
 sg13g2_decap_8 FILLER_73_2318 ();
 sg13g2_decap_8 FILLER_73_2325 ();
 sg13g2_decap_8 FILLER_73_2332 ();
 sg13g2_decap_8 FILLER_73_2339 ();
 sg13g2_decap_8 FILLER_73_2346 ();
 sg13g2_decap_8 FILLER_73_2353 ();
 sg13g2_decap_8 FILLER_73_2360 ();
 sg13g2_decap_8 FILLER_73_2367 ();
 sg13g2_decap_8 FILLER_73_2374 ();
 sg13g2_decap_8 FILLER_73_2381 ();
 sg13g2_decap_8 FILLER_73_2388 ();
 sg13g2_decap_8 FILLER_73_2395 ();
 sg13g2_decap_8 FILLER_73_2402 ();
 sg13g2_decap_8 FILLER_73_2409 ();
 sg13g2_decap_8 FILLER_73_2416 ();
 sg13g2_decap_8 FILLER_73_2423 ();
 sg13g2_decap_8 FILLER_73_2430 ();
 sg13g2_decap_8 FILLER_73_2437 ();
 sg13g2_decap_8 FILLER_73_2444 ();
 sg13g2_decap_8 FILLER_73_2451 ();
 sg13g2_decap_8 FILLER_73_2458 ();
 sg13g2_decap_8 FILLER_73_2465 ();
 sg13g2_decap_8 FILLER_73_2472 ();
 sg13g2_decap_8 FILLER_73_2479 ();
 sg13g2_decap_8 FILLER_73_2486 ();
 sg13g2_decap_8 FILLER_73_2493 ();
 sg13g2_decap_8 FILLER_73_2500 ();
 sg13g2_decap_8 FILLER_73_2507 ();
 sg13g2_decap_8 FILLER_73_2514 ();
 sg13g2_decap_8 FILLER_73_2521 ();
 sg13g2_decap_8 FILLER_73_2528 ();
 sg13g2_decap_8 FILLER_73_2535 ();
 sg13g2_decap_8 FILLER_73_2542 ();
 sg13g2_decap_8 FILLER_73_2549 ();
 sg13g2_decap_8 FILLER_73_2556 ();
 sg13g2_decap_8 FILLER_73_2563 ();
 sg13g2_decap_8 FILLER_73_2570 ();
 sg13g2_decap_8 FILLER_73_2577 ();
 sg13g2_decap_8 FILLER_73_2584 ();
 sg13g2_decap_8 FILLER_73_2591 ();
 sg13g2_decap_8 FILLER_73_2598 ();
 sg13g2_decap_8 FILLER_73_2605 ();
 sg13g2_decap_8 FILLER_73_2612 ();
 sg13g2_decap_8 FILLER_73_2619 ();
 sg13g2_decap_8 FILLER_73_2626 ();
 sg13g2_decap_8 FILLER_73_2633 ();
 sg13g2_decap_8 FILLER_73_2640 ();
 sg13g2_decap_8 FILLER_73_2647 ();
 sg13g2_decap_8 FILLER_73_2654 ();
 sg13g2_decap_8 FILLER_73_2661 ();
 sg13g2_decap_4 FILLER_73_2668 ();
 sg13g2_fill_2 FILLER_73_2672 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_decap_8 FILLER_74_175 ();
 sg13g2_decap_8 FILLER_74_182 ();
 sg13g2_decap_8 FILLER_74_189 ();
 sg13g2_decap_8 FILLER_74_196 ();
 sg13g2_decap_8 FILLER_74_203 ();
 sg13g2_decap_8 FILLER_74_210 ();
 sg13g2_decap_8 FILLER_74_217 ();
 sg13g2_decap_8 FILLER_74_224 ();
 sg13g2_decap_8 FILLER_74_231 ();
 sg13g2_decap_8 FILLER_74_238 ();
 sg13g2_decap_8 FILLER_74_245 ();
 sg13g2_decap_8 FILLER_74_252 ();
 sg13g2_decap_8 FILLER_74_259 ();
 sg13g2_decap_8 FILLER_74_266 ();
 sg13g2_decap_8 FILLER_74_273 ();
 sg13g2_decap_8 FILLER_74_280 ();
 sg13g2_decap_8 FILLER_74_287 ();
 sg13g2_decap_8 FILLER_74_294 ();
 sg13g2_decap_8 FILLER_74_301 ();
 sg13g2_decap_8 FILLER_74_308 ();
 sg13g2_decap_8 FILLER_74_315 ();
 sg13g2_decap_8 FILLER_74_322 ();
 sg13g2_decap_8 FILLER_74_329 ();
 sg13g2_decap_8 FILLER_74_336 ();
 sg13g2_decap_8 FILLER_74_343 ();
 sg13g2_decap_8 FILLER_74_350 ();
 sg13g2_decap_8 FILLER_74_357 ();
 sg13g2_decap_8 FILLER_74_364 ();
 sg13g2_decap_8 FILLER_74_371 ();
 sg13g2_decap_8 FILLER_74_378 ();
 sg13g2_decap_8 FILLER_74_385 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_decap_8 FILLER_74_406 ();
 sg13g2_decap_8 FILLER_74_413 ();
 sg13g2_decap_8 FILLER_74_420 ();
 sg13g2_decap_8 FILLER_74_427 ();
 sg13g2_decap_8 FILLER_74_434 ();
 sg13g2_decap_8 FILLER_74_441 ();
 sg13g2_decap_8 FILLER_74_448 ();
 sg13g2_decap_8 FILLER_74_455 ();
 sg13g2_decap_8 FILLER_74_462 ();
 sg13g2_decap_8 FILLER_74_469 ();
 sg13g2_decap_8 FILLER_74_476 ();
 sg13g2_decap_8 FILLER_74_483 ();
 sg13g2_decap_4 FILLER_74_490 ();
 sg13g2_fill_2 FILLER_74_521 ();
 sg13g2_fill_1 FILLER_74_532 ();
 sg13g2_fill_2 FILLER_74_558 ();
 sg13g2_fill_1 FILLER_74_560 ();
 sg13g2_decap_4 FILLER_74_626 ();
 sg13g2_decap_4 FILLER_74_652 ();
 sg13g2_fill_1 FILLER_74_656 ();
 sg13g2_fill_2 FILLER_74_687 ();
 sg13g2_fill_1 FILLER_74_725 ();
 sg13g2_decap_4 FILLER_74_757 ();
 sg13g2_fill_2 FILLER_74_787 ();
 sg13g2_fill_1 FILLER_74_822 ();
 sg13g2_fill_2 FILLER_74_875 ();
 sg13g2_decap_4 FILLER_74_896 ();
 sg13g2_fill_1 FILLER_74_900 ();
 sg13g2_fill_2 FILLER_74_976 ();
 sg13g2_fill_1 FILLER_74_978 ();
 sg13g2_fill_1 FILLER_74_984 ();
 sg13g2_fill_2 FILLER_74_1046 ();
 sg13g2_fill_1 FILLER_74_1048 ();
 sg13g2_fill_2 FILLER_74_1096 ();
 sg13g2_fill_1 FILLER_74_1107 ();
 sg13g2_fill_2 FILLER_74_1113 ();
 sg13g2_fill_2 FILLER_74_1124 ();
 sg13g2_decap_4 FILLER_74_1175 ();
 sg13g2_fill_2 FILLER_74_1192 ();
 sg13g2_fill_1 FILLER_74_1194 ();
 sg13g2_fill_2 FILLER_74_1219 ();
 sg13g2_fill_1 FILLER_74_1221 ();
 sg13g2_fill_1 FILLER_74_1231 ();
 sg13g2_fill_1 FILLER_74_1249 ();
 sg13g2_fill_2 FILLER_74_1297 ();
 sg13g2_fill_2 FILLER_74_1359 ();
 sg13g2_fill_2 FILLER_74_1370 ();
 sg13g2_fill_1 FILLER_74_1372 ();
 sg13g2_fill_1 FILLER_74_1382 ();
 sg13g2_decap_8 FILLER_74_1387 ();
 sg13g2_fill_2 FILLER_74_1394 ();
 sg13g2_fill_1 FILLER_74_1448 ();
 sg13g2_fill_2 FILLER_74_1475 ();
 sg13g2_fill_1 FILLER_74_1477 ();
 sg13g2_fill_1 FILLER_74_1518 ();
 sg13g2_decap_4 FILLER_74_1595 ();
 sg13g2_fill_2 FILLER_74_1599 ();
 sg13g2_fill_1 FILLER_74_1615 ();
 sg13g2_fill_2 FILLER_74_1621 ();
 sg13g2_fill_1 FILLER_74_1654 ();
 sg13g2_fill_1 FILLER_74_1664 ();
 sg13g2_decap_8 FILLER_74_1691 ();
 sg13g2_decap_4 FILLER_74_1703 ();
 sg13g2_fill_1 FILLER_74_1785 ();
 sg13g2_fill_1 FILLER_74_1793 ();
 sg13g2_fill_2 FILLER_74_1813 ();
 sg13g2_fill_1 FILLER_74_1815 ();
 sg13g2_decap_8 FILLER_74_1820 ();
 sg13g2_fill_1 FILLER_74_1827 ();
 sg13g2_fill_1 FILLER_74_1837 ();
 sg13g2_fill_2 FILLER_74_1848 ();
 sg13g2_fill_1 FILLER_74_1885 ();
 sg13g2_fill_1 FILLER_74_1890 ();
 sg13g2_fill_1 FILLER_74_1895 ();
 sg13g2_decap_8 FILLER_74_1900 ();
 sg13g2_fill_2 FILLER_74_1907 ();
 sg13g2_fill_2 FILLER_74_1918 ();
 sg13g2_fill_1 FILLER_74_1920 ();
 sg13g2_decap_8 FILLER_74_1952 ();
 sg13g2_fill_2 FILLER_74_1973 ();
 sg13g2_fill_1 FILLER_74_1975 ();
 sg13g2_fill_2 FILLER_74_1985 ();
 sg13g2_fill_1 FILLER_74_1987 ();
 sg13g2_fill_1 FILLER_74_2002 ();
 sg13g2_decap_8 FILLER_74_2034 ();
 sg13g2_fill_2 FILLER_74_2075 ();
 sg13g2_fill_2 FILLER_74_2082 ();
 sg13g2_fill_1 FILLER_74_2084 ();
 sg13g2_fill_2 FILLER_74_2098 ();
 sg13g2_fill_1 FILLER_74_2100 ();
 sg13g2_fill_2 FILLER_74_2106 ();
 sg13g2_fill_1 FILLER_74_2108 ();
 sg13g2_fill_2 FILLER_74_2160 ();
 sg13g2_fill_1 FILLER_74_2162 ();
 sg13g2_fill_2 FILLER_74_2194 ();
 sg13g2_decap_8 FILLER_74_2279 ();
 sg13g2_decap_8 FILLER_74_2286 ();
 sg13g2_decap_8 FILLER_74_2293 ();
 sg13g2_decap_8 FILLER_74_2300 ();
 sg13g2_decap_8 FILLER_74_2307 ();
 sg13g2_decap_8 FILLER_74_2314 ();
 sg13g2_decap_8 FILLER_74_2321 ();
 sg13g2_decap_8 FILLER_74_2328 ();
 sg13g2_decap_8 FILLER_74_2335 ();
 sg13g2_decap_8 FILLER_74_2342 ();
 sg13g2_decap_8 FILLER_74_2349 ();
 sg13g2_decap_8 FILLER_74_2356 ();
 sg13g2_decap_8 FILLER_74_2363 ();
 sg13g2_decap_8 FILLER_74_2370 ();
 sg13g2_decap_8 FILLER_74_2377 ();
 sg13g2_decap_8 FILLER_74_2384 ();
 sg13g2_decap_8 FILLER_74_2391 ();
 sg13g2_decap_8 FILLER_74_2398 ();
 sg13g2_decap_8 FILLER_74_2405 ();
 sg13g2_decap_8 FILLER_74_2412 ();
 sg13g2_decap_8 FILLER_74_2419 ();
 sg13g2_decap_8 FILLER_74_2426 ();
 sg13g2_decap_8 FILLER_74_2433 ();
 sg13g2_decap_8 FILLER_74_2440 ();
 sg13g2_decap_8 FILLER_74_2447 ();
 sg13g2_decap_8 FILLER_74_2454 ();
 sg13g2_decap_8 FILLER_74_2461 ();
 sg13g2_decap_8 FILLER_74_2468 ();
 sg13g2_decap_8 FILLER_74_2475 ();
 sg13g2_decap_8 FILLER_74_2482 ();
 sg13g2_decap_8 FILLER_74_2489 ();
 sg13g2_decap_8 FILLER_74_2496 ();
 sg13g2_decap_8 FILLER_74_2503 ();
 sg13g2_decap_8 FILLER_74_2510 ();
 sg13g2_decap_8 FILLER_74_2517 ();
 sg13g2_decap_8 FILLER_74_2524 ();
 sg13g2_decap_8 FILLER_74_2531 ();
 sg13g2_decap_8 FILLER_74_2538 ();
 sg13g2_decap_8 FILLER_74_2545 ();
 sg13g2_decap_8 FILLER_74_2552 ();
 sg13g2_decap_8 FILLER_74_2559 ();
 sg13g2_decap_8 FILLER_74_2566 ();
 sg13g2_decap_8 FILLER_74_2573 ();
 sg13g2_decap_8 FILLER_74_2580 ();
 sg13g2_decap_8 FILLER_74_2587 ();
 sg13g2_decap_8 FILLER_74_2594 ();
 sg13g2_decap_8 FILLER_74_2601 ();
 sg13g2_decap_8 FILLER_74_2608 ();
 sg13g2_decap_8 FILLER_74_2615 ();
 sg13g2_decap_8 FILLER_74_2622 ();
 sg13g2_decap_8 FILLER_74_2629 ();
 sg13g2_decap_8 FILLER_74_2636 ();
 sg13g2_decap_8 FILLER_74_2643 ();
 sg13g2_decap_8 FILLER_74_2650 ();
 sg13g2_decap_8 FILLER_74_2657 ();
 sg13g2_decap_8 FILLER_74_2664 ();
 sg13g2_fill_2 FILLER_74_2671 ();
 sg13g2_fill_1 FILLER_74_2673 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_8 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_196 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_224 ();
 sg13g2_decap_8 FILLER_75_231 ();
 sg13g2_decap_8 FILLER_75_238 ();
 sg13g2_decap_8 FILLER_75_245 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_decap_8 FILLER_75_259 ();
 sg13g2_decap_8 FILLER_75_266 ();
 sg13g2_decap_8 FILLER_75_273 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_decap_8 FILLER_75_287 ();
 sg13g2_decap_8 FILLER_75_294 ();
 sg13g2_decap_8 FILLER_75_301 ();
 sg13g2_decap_8 FILLER_75_308 ();
 sg13g2_decap_8 FILLER_75_315 ();
 sg13g2_decap_8 FILLER_75_322 ();
 sg13g2_decap_8 FILLER_75_329 ();
 sg13g2_decap_8 FILLER_75_336 ();
 sg13g2_decap_8 FILLER_75_343 ();
 sg13g2_decap_8 FILLER_75_350 ();
 sg13g2_decap_8 FILLER_75_357 ();
 sg13g2_decap_8 FILLER_75_364 ();
 sg13g2_decap_8 FILLER_75_371 ();
 sg13g2_decap_8 FILLER_75_378 ();
 sg13g2_decap_8 FILLER_75_385 ();
 sg13g2_decap_8 FILLER_75_392 ();
 sg13g2_decap_8 FILLER_75_399 ();
 sg13g2_decap_8 FILLER_75_406 ();
 sg13g2_decap_8 FILLER_75_413 ();
 sg13g2_decap_8 FILLER_75_420 ();
 sg13g2_decap_8 FILLER_75_427 ();
 sg13g2_decap_8 FILLER_75_434 ();
 sg13g2_decap_8 FILLER_75_441 ();
 sg13g2_decap_8 FILLER_75_448 ();
 sg13g2_decap_8 FILLER_75_455 ();
 sg13g2_decap_8 FILLER_75_462 ();
 sg13g2_decap_8 FILLER_75_469 ();
 sg13g2_decap_8 FILLER_75_476 ();
 sg13g2_fill_2 FILLER_75_483 ();
 sg13g2_fill_1 FILLER_75_485 ();
 sg13g2_fill_2 FILLER_75_583 ();
 sg13g2_fill_1 FILLER_75_585 ();
 sg13g2_fill_1 FILLER_75_623 ();
 sg13g2_fill_2 FILLER_75_648 ();
 sg13g2_fill_1 FILLER_75_663 ();
 sg13g2_fill_2 FILLER_75_677 ();
 sg13g2_fill_1 FILLER_75_705 ();
 sg13g2_fill_2 FILLER_75_715 ();
 sg13g2_fill_1 FILLER_75_717 ();
 sg13g2_fill_2 FILLER_75_757 ();
 sg13g2_fill_2 FILLER_75_763 ();
 sg13g2_fill_1 FILLER_75_765 ();
 sg13g2_fill_2 FILLER_75_770 ();
 sg13g2_fill_1 FILLER_75_776 ();
 sg13g2_fill_2 FILLER_75_799 ();
 sg13g2_fill_1 FILLER_75_806 ();
 sg13g2_fill_1 FILLER_75_833 ();
 sg13g2_decap_4 FILLER_75_843 ();
 sg13g2_fill_2 FILLER_75_852 ();
 sg13g2_fill_1 FILLER_75_854 ();
 sg13g2_fill_2 FILLER_75_859 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_fill_1 FILLER_75_927 ();
 sg13g2_fill_1 FILLER_75_954 ();
 sg13g2_fill_1 FILLER_75_986 ();
 sg13g2_fill_2 FILLER_75_992 ();
 sg13g2_fill_1 FILLER_75_994 ();
 sg13g2_fill_2 FILLER_75_1003 ();
 sg13g2_fill_1 FILLER_75_1005 ();
 sg13g2_fill_2 FILLER_75_1024 ();
 sg13g2_fill_1 FILLER_75_1026 ();
 sg13g2_fill_1 FILLER_75_1045 ();
 sg13g2_fill_1 FILLER_75_1055 ();
 sg13g2_fill_1 FILLER_75_1060 ();
 sg13g2_fill_2 FILLER_75_1102 ();
 sg13g2_fill_1 FILLER_75_1104 ();
 sg13g2_fill_2 FILLER_75_1129 ();
 sg13g2_fill_1 FILLER_75_1131 ();
 sg13g2_fill_2 FILLER_75_1220 ();
 sg13g2_fill_1 FILLER_75_1248 ();
 sg13g2_fill_2 FILLER_75_1253 ();
 sg13g2_fill_1 FILLER_75_1255 ();
 sg13g2_fill_2 FILLER_75_1304 ();
 sg13g2_fill_2 FILLER_75_1358 ();
 sg13g2_fill_1 FILLER_75_1360 ();
 sg13g2_fill_2 FILLER_75_1397 ();
 sg13g2_fill_1 FILLER_75_1399 ();
 sg13g2_decap_4 FILLER_75_1426 ();
 sg13g2_fill_2 FILLER_75_1430 ();
 sg13g2_decap_4 FILLER_75_1440 ();
 sg13g2_fill_2 FILLER_75_1452 ();
 sg13g2_fill_1 FILLER_75_1467 ();
 sg13g2_fill_2 FILLER_75_1472 ();
 sg13g2_decap_8 FILLER_75_1482 ();
 sg13g2_fill_2 FILLER_75_1493 ();
 sg13g2_fill_2 FILLER_75_1531 ();
 sg13g2_fill_1 FILLER_75_1533 ();
 sg13g2_fill_2 FILLER_75_1543 ();
 sg13g2_fill_1 FILLER_75_1576 ();
 sg13g2_fill_2 FILLER_75_1603 ();
 sg13g2_fill_2 FILLER_75_1609 ();
 sg13g2_fill_2 FILLER_75_1620 ();
 sg13g2_fill_1 FILLER_75_1626 ();
 sg13g2_fill_2 FILLER_75_1683 ();
 sg13g2_fill_1 FILLER_75_1685 ();
 sg13g2_fill_1 FILLER_75_1708 ();
 sg13g2_fill_1 FILLER_75_1749 ();
 sg13g2_decap_4 FILLER_75_1775 ();
 sg13g2_fill_1 FILLER_75_1779 ();
 sg13g2_fill_1 FILLER_75_1797 ();
 sg13g2_fill_2 FILLER_75_1803 ();
 sg13g2_decap_4 FILLER_75_1822 ();
 sg13g2_fill_1 FILLER_75_1874 ();
 sg13g2_fill_2 FILLER_75_1941 ();
 sg13g2_fill_1 FILLER_75_1943 ();
 sg13g2_fill_1 FILLER_75_2038 ();
 sg13g2_fill_2 FILLER_75_2048 ();
 sg13g2_fill_1 FILLER_75_2050 ();
 sg13g2_fill_1 FILLER_75_2086 ();
 sg13g2_fill_2 FILLER_75_2096 ();
 sg13g2_fill_1 FILLER_75_2154 ();
 sg13g2_decap_4 FILLER_75_2159 ();
 sg13g2_fill_2 FILLER_75_2163 ();
 sg13g2_fill_1 FILLER_75_2169 ();
 sg13g2_fill_2 FILLER_75_2186 ();
 sg13g2_fill_1 FILLER_75_2188 ();
 sg13g2_decap_4 FILLER_75_2223 ();
 sg13g2_fill_1 FILLER_75_2227 ();
 sg13g2_fill_2 FILLER_75_2241 ();
 sg13g2_fill_1 FILLER_75_2260 ();
 sg13g2_fill_1 FILLER_75_2265 ();
 sg13g2_decap_8 FILLER_75_2275 ();
 sg13g2_decap_8 FILLER_75_2282 ();
 sg13g2_decap_8 FILLER_75_2289 ();
 sg13g2_decap_8 FILLER_75_2296 ();
 sg13g2_decap_8 FILLER_75_2303 ();
 sg13g2_decap_8 FILLER_75_2310 ();
 sg13g2_decap_8 FILLER_75_2317 ();
 sg13g2_decap_8 FILLER_75_2324 ();
 sg13g2_decap_8 FILLER_75_2331 ();
 sg13g2_decap_8 FILLER_75_2338 ();
 sg13g2_decap_8 FILLER_75_2345 ();
 sg13g2_decap_8 FILLER_75_2352 ();
 sg13g2_decap_8 FILLER_75_2359 ();
 sg13g2_decap_8 FILLER_75_2366 ();
 sg13g2_decap_8 FILLER_75_2373 ();
 sg13g2_decap_8 FILLER_75_2380 ();
 sg13g2_decap_8 FILLER_75_2387 ();
 sg13g2_decap_8 FILLER_75_2394 ();
 sg13g2_decap_8 FILLER_75_2401 ();
 sg13g2_decap_8 FILLER_75_2408 ();
 sg13g2_decap_8 FILLER_75_2415 ();
 sg13g2_decap_8 FILLER_75_2422 ();
 sg13g2_decap_8 FILLER_75_2429 ();
 sg13g2_decap_8 FILLER_75_2436 ();
 sg13g2_decap_8 FILLER_75_2443 ();
 sg13g2_decap_8 FILLER_75_2450 ();
 sg13g2_decap_8 FILLER_75_2457 ();
 sg13g2_decap_8 FILLER_75_2464 ();
 sg13g2_decap_8 FILLER_75_2471 ();
 sg13g2_decap_8 FILLER_75_2478 ();
 sg13g2_decap_8 FILLER_75_2485 ();
 sg13g2_decap_8 FILLER_75_2492 ();
 sg13g2_decap_8 FILLER_75_2499 ();
 sg13g2_decap_8 FILLER_75_2506 ();
 sg13g2_decap_8 FILLER_75_2513 ();
 sg13g2_decap_8 FILLER_75_2520 ();
 sg13g2_decap_8 FILLER_75_2527 ();
 sg13g2_decap_8 FILLER_75_2534 ();
 sg13g2_decap_8 FILLER_75_2541 ();
 sg13g2_decap_8 FILLER_75_2548 ();
 sg13g2_decap_8 FILLER_75_2555 ();
 sg13g2_decap_8 FILLER_75_2562 ();
 sg13g2_decap_8 FILLER_75_2569 ();
 sg13g2_decap_8 FILLER_75_2576 ();
 sg13g2_decap_8 FILLER_75_2583 ();
 sg13g2_decap_8 FILLER_75_2590 ();
 sg13g2_decap_8 FILLER_75_2597 ();
 sg13g2_decap_8 FILLER_75_2604 ();
 sg13g2_decap_8 FILLER_75_2611 ();
 sg13g2_decap_8 FILLER_75_2618 ();
 sg13g2_decap_8 FILLER_75_2625 ();
 sg13g2_decap_8 FILLER_75_2632 ();
 sg13g2_decap_8 FILLER_75_2639 ();
 sg13g2_decap_8 FILLER_75_2646 ();
 sg13g2_decap_8 FILLER_75_2653 ();
 sg13g2_decap_8 FILLER_75_2660 ();
 sg13g2_decap_8 FILLER_75_2667 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_8 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_decap_8 FILLER_76_273 ();
 sg13g2_decap_8 FILLER_76_280 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_392 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_decap_8 FILLER_76_406 ();
 sg13g2_decap_8 FILLER_76_413 ();
 sg13g2_decap_8 FILLER_76_420 ();
 sg13g2_decap_8 FILLER_76_427 ();
 sg13g2_decap_8 FILLER_76_434 ();
 sg13g2_decap_8 FILLER_76_441 ();
 sg13g2_decap_8 FILLER_76_448 ();
 sg13g2_decap_8 FILLER_76_455 ();
 sg13g2_decap_8 FILLER_76_462 ();
 sg13g2_decap_8 FILLER_76_469 ();
 sg13g2_decap_8 FILLER_76_476 ();
 sg13g2_decap_8 FILLER_76_483 ();
 sg13g2_decap_8 FILLER_76_490 ();
 sg13g2_fill_2 FILLER_76_497 ();
 sg13g2_fill_1 FILLER_76_499 ();
 sg13g2_decap_4 FILLER_76_514 ();
 sg13g2_decap_4 FILLER_76_522 ();
 sg13g2_fill_2 FILLER_76_535 ();
 sg13g2_fill_1 FILLER_76_573 ();
 sg13g2_fill_2 FILLER_76_600 ();
 sg13g2_fill_1 FILLER_76_602 ();
 sg13g2_fill_2 FILLER_76_643 ();
 sg13g2_fill_1 FILLER_76_671 ();
 sg13g2_decap_4 FILLER_76_676 ();
 sg13g2_fill_1 FILLER_76_700 ();
 sg13g2_fill_1 FILLER_76_798 ();
 sg13g2_decap_4 FILLER_76_828 ();
 sg13g2_fill_2 FILLER_76_841 ();
 sg13g2_fill_1 FILLER_76_843 ();
 sg13g2_fill_2 FILLER_76_889 ();
 sg13g2_fill_1 FILLER_76_891 ();
 sg13g2_decap_8 FILLER_76_949 ();
 sg13g2_fill_1 FILLER_76_956 ();
 sg13g2_fill_2 FILLER_76_966 ();
 sg13g2_fill_2 FILLER_76_981 ();
 sg13g2_fill_1 FILLER_76_987 ();
 sg13g2_fill_2 FILLER_76_1000 ();
 sg13g2_fill_1 FILLER_76_1002 ();
 sg13g2_decap_4 FILLER_76_1011 ();
 sg13g2_fill_2 FILLER_76_1041 ();
 sg13g2_fill_2 FILLER_76_1129 ();
 sg13g2_fill_1 FILLER_76_1131 ();
 sg13g2_fill_1 FILLER_76_1142 ();
 sg13g2_fill_2 FILLER_76_1161 ();
 sg13g2_fill_1 FILLER_76_1163 ();
 sg13g2_fill_2 FILLER_76_1177 ();
 sg13g2_fill_2 FILLER_76_1206 ();
 sg13g2_fill_2 FILLER_76_1229 ();
 sg13g2_fill_1 FILLER_76_1240 ();
 sg13g2_fill_2 FILLER_76_1268 ();
 sg13g2_fill_1 FILLER_76_1270 ();
 sg13g2_fill_1 FILLER_76_1306 ();
 sg13g2_fill_2 FILLER_76_1321 ();
 sg13g2_fill_1 FILLER_76_1323 ();
 sg13g2_decap_4 FILLER_76_1337 ();
 sg13g2_fill_2 FILLER_76_1341 ();
 sg13g2_fill_2 FILLER_76_1347 ();
 sg13g2_fill_2 FILLER_76_1354 ();
 sg13g2_fill_1 FILLER_76_1356 ();
 sg13g2_decap_4 FILLER_76_1483 ();
 sg13g2_fill_1 FILLER_76_1505 ();
 sg13g2_fill_2 FILLER_76_1563 ();
 sg13g2_fill_2 FILLER_76_1579 ();
 sg13g2_fill_1 FILLER_76_1581 ();
 sg13g2_fill_2 FILLER_76_1709 ();
 sg13g2_decap_4 FILLER_76_1767 ();
 sg13g2_fill_1 FILLER_76_1802 ();
 sg13g2_fill_2 FILLER_76_1843 ();
 sg13g2_fill_1 FILLER_76_1845 ();
 sg13g2_decap_4 FILLER_76_1894 ();
 sg13g2_fill_2 FILLER_76_1898 ();
 sg13g2_fill_1 FILLER_76_1912 ();
 sg13g2_fill_2 FILLER_76_1918 ();
 sg13g2_fill_1 FILLER_76_1920 ();
 sg13g2_decap_4 FILLER_76_1955 ();
 sg13g2_fill_2 FILLER_76_1959 ();
 sg13g2_fill_2 FILLER_76_2016 ();
 sg13g2_fill_2 FILLER_76_2067 ();
 sg13g2_fill_1 FILLER_76_2114 ();
 sg13g2_fill_2 FILLER_76_2146 ();
 sg13g2_fill_1 FILLER_76_2148 ();
 sg13g2_fill_2 FILLER_76_2158 ();
 sg13g2_fill_1 FILLER_76_2160 ();
 sg13g2_fill_1 FILLER_76_2165 ();
 sg13g2_fill_1 FILLER_76_2179 ();
 sg13g2_fill_1 FILLER_76_2201 ();
 sg13g2_decap_8 FILLER_76_2245 ();
 sg13g2_decap_8 FILLER_76_2252 ();
 sg13g2_decap_8 FILLER_76_2259 ();
 sg13g2_decap_8 FILLER_76_2266 ();
 sg13g2_decap_8 FILLER_76_2273 ();
 sg13g2_decap_8 FILLER_76_2280 ();
 sg13g2_decap_8 FILLER_76_2287 ();
 sg13g2_decap_8 FILLER_76_2294 ();
 sg13g2_decap_8 FILLER_76_2301 ();
 sg13g2_decap_8 FILLER_76_2308 ();
 sg13g2_decap_8 FILLER_76_2315 ();
 sg13g2_decap_8 FILLER_76_2322 ();
 sg13g2_decap_8 FILLER_76_2329 ();
 sg13g2_decap_8 FILLER_76_2336 ();
 sg13g2_decap_8 FILLER_76_2343 ();
 sg13g2_decap_8 FILLER_76_2350 ();
 sg13g2_decap_8 FILLER_76_2357 ();
 sg13g2_decap_8 FILLER_76_2364 ();
 sg13g2_decap_8 FILLER_76_2371 ();
 sg13g2_decap_8 FILLER_76_2378 ();
 sg13g2_decap_8 FILLER_76_2385 ();
 sg13g2_decap_8 FILLER_76_2392 ();
 sg13g2_decap_8 FILLER_76_2399 ();
 sg13g2_decap_8 FILLER_76_2406 ();
 sg13g2_decap_8 FILLER_76_2413 ();
 sg13g2_decap_8 FILLER_76_2420 ();
 sg13g2_decap_8 FILLER_76_2427 ();
 sg13g2_decap_8 FILLER_76_2434 ();
 sg13g2_decap_8 FILLER_76_2441 ();
 sg13g2_decap_8 FILLER_76_2448 ();
 sg13g2_decap_8 FILLER_76_2455 ();
 sg13g2_decap_8 FILLER_76_2462 ();
 sg13g2_decap_8 FILLER_76_2469 ();
 sg13g2_decap_8 FILLER_76_2476 ();
 sg13g2_decap_8 FILLER_76_2483 ();
 sg13g2_decap_8 FILLER_76_2490 ();
 sg13g2_decap_8 FILLER_76_2497 ();
 sg13g2_decap_8 FILLER_76_2504 ();
 sg13g2_decap_8 FILLER_76_2511 ();
 sg13g2_decap_8 FILLER_76_2518 ();
 sg13g2_decap_8 FILLER_76_2525 ();
 sg13g2_decap_8 FILLER_76_2532 ();
 sg13g2_decap_8 FILLER_76_2539 ();
 sg13g2_decap_8 FILLER_76_2546 ();
 sg13g2_decap_8 FILLER_76_2553 ();
 sg13g2_decap_8 FILLER_76_2560 ();
 sg13g2_decap_8 FILLER_76_2567 ();
 sg13g2_decap_8 FILLER_76_2574 ();
 sg13g2_decap_8 FILLER_76_2581 ();
 sg13g2_decap_8 FILLER_76_2588 ();
 sg13g2_decap_8 FILLER_76_2595 ();
 sg13g2_decap_8 FILLER_76_2602 ();
 sg13g2_decap_8 FILLER_76_2609 ();
 sg13g2_decap_8 FILLER_76_2616 ();
 sg13g2_decap_8 FILLER_76_2623 ();
 sg13g2_decap_8 FILLER_76_2630 ();
 sg13g2_decap_8 FILLER_76_2637 ();
 sg13g2_decap_8 FILLER_76_2644 ();
 sg13g2_decap_8 FILLER_76_2651 ();
 sg13g2_decap_8 FILLER_76_2658 ();
 sg13g2_decap_8 FILLER_76_2665 ();
 sg13g2_fill_2 FILLER_76_2672 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_8 FILLER_77_245 ();
 sg13g2_decap_8 FILLER_77_252 ();
 sg13g2_decap_8 FILLER_77_259 ();
 sg13g2_decap_8 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_273 ();
 sg13g2_decap_8 FILLER_77_280 ();
 sg13g2_decap_8 FILLER_77_287 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_decap_8 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_364 ();
 sg13g2_decap_8 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_decap_8 FILLER_77_427 ();
 sg13g2_decap_8 FILLER_77_434 ();
 sg13g2_decap_8 FILLER_77_441 ();
 sg13g2_decap_8 FILLER_77_448 ();
 sg13g2_decap_8 FILLER_77_455 ();
 sg13g2_decap_8 FILLER_77_462 ();
 sg13g2_decap_8 FILLER_77_469 ();
 sg13g2_decap_8 FILLER_77_476 ();
 sg13g2_decap_8 FILLER_77_483 ();
 sg13g2_decap_8 FILLER_77_490 ();
 sg13g2_decap_8 FILLER_77_497 ();
 sg13g2_fill_2 FILLER_77_504 ();
 sg13g2_fill_1 FILLER_77_506 ();
 sg13g2_fill_2 FILLER_77_533 ();
 sg13g2_decap_4 FILLER_77_569 ();
 sg13g2_fill_1 FILLER_77_573 ();
 sg13g2_fill_1 FILLER_77_579 ();
 sg13g2_fill_2 FILLER_77_589 ();
 sg13g2_fill_1 FILLER_77_591 ();
 sg13g2_fill_2 FILLER_77_597 ();
 sg13g2_fill_1 FILLER_77_599 ();
 sg13g2_decap_8 FILLER_77_605 ();
 sg13g2_fill_2 FILLER_77_612 ();
 sg13g2_decap_4 FILLER_77_622 ();
 sg13g2_fill_2 FILLER_77_696 ();
 sg13g2_fill_1 FILLER_77_702 ();
 sg13g2_fill_1 FILLER_77_708 ();
 sg13g2_fill_2 FILLER_77_713 ();
 sg13g2_fill_2 FILLER_77_728 ();
 sg13g2_fill_2 FILLER_77_734 ();
 sg13g2_fill_1 FILLER_77_736 ();
 sg13g2_fill_2 FILLER_77_797 ();
 sg13g2_fill_2 FILLER_77_803 ();
 sg13g2_fill_1 FILLER_77_805 ();
 sg13g2_fill_2 FILLER_77_867 ();
 sg13g2_fill_1 FILLER_77_869 ();
 sg13g2_fill_1 FILLER_77_908 ();
 sg13g2_decap_4 FILLER_77_935 ();
 sg13g2_decap_8 FILLER_77_943 ();
 sg13g2_decap_8 FILLER_77_950 ();
 sg13g2_fill_1 FILLER_77_957 ();
 sg13g2_fill_1 FILLER_77_989 ();
 sg13g2_fill_2 FILLER_77_994 ();
 sg13g2_decap_8 FILLER_77_1005 ();
 sg13g2_fill_1 FILLER_77_1012 ();
 sg13g2_fill_1 FILLER_77_1023 ();
 sg13g2_fill_2 FILLER_77_1050 ();
 sg13g2_fill_2 FILLER_77_1070 ();
 sg13g2_fill_2 FILLER_77_1080 ();
 sg13g2_fill_1 FILLER_77_1099 ();
 sg13g2_fill_1 FILLER_77_1108 ();
 sg13g2_fill_2 FILLER_77_1161 ();
 sg13g2_fill_2 FILLER_77_1215 ();
 sg13g2_fill_1 FILLER_77_1217 ();
 sg13g2_fill_1 FILLER_77_1227 ();
 sg13g2_fill_2 FILLER_77_1280 ();
 sg13g2_fill_1 FILLER_77_1282 ();
 sg13g2_fill_2 FILLER_77_1326 ();
 sg13g2_fill_1 FILLER_77_1328 ();
 sg13g2_fill_2 FILLER_77_1380 ();
 sg13g2_fill_1 FILLER_77_1382 ();
 sg13g2_fill_1 FILLER_77_1396 ();
 sg13g2_fill_2 FILLER_77_1441 ();
 sg13g2_fill_2 FILLER_77_1461 ();
 sg13g2_decap_8 FILLER_77_1512 ();
 sg13g2_fill_2 FILLER_77_1519 ();
 sg13g2_fill_1 FILLER_77_1521 ();
 sg13g2_fill_2 FILLER_77_1531 ();
 sg13g2_fill_2 FILLER_77_1537 ();
 sg13g2_fill_1 FILLER_77_1539 ();
 sg13g2_fill_2 FILLER_77_1549 ();
 sg13g2_fill_1 FILLER_77_1551 ();
 sg13g2_fill_2 FILLER_77_1562 ();
 sg13g2_fill_2 FILLER_77_1599 ();
 sg13g2_fill_1 FILLER_77_1601 ();
 sg13g2_fill_2 FILLER_77_1621 ();
 sg13g2_decap_4 FILLER_77_1706 ();
 sg13g2_fill_1 FILLER_77_1710 ();
 sg13g2_fill_2 FILLER_77_1724 ();
 sg13g2_fill_1 FILLER_77_1726 ();
 sg13g2_fill_2 FILLER_77_1740 ();
 sg13g2_decap_4 FILLER_77_1777 ();
 sg13g2_fill_1 FILLER_77_1781 ();
 sg13g2_decap_8 FILLER_77_1786 ();
 sg13g2_fill_2 FILLER_77_1802 ();
 sg13g2_fill_1 FILLER_77_1804 ();
 sg13g2_decap_8 FILLER_77_1810 ();
 sg13g2_fill_1 FILLER_77_1817 ();
 sg13g2_fill_2 FILLER_77_1910 ();
 sg13g2_fill_1 FILLER_77_1912 ();
 sg13g2_fill_2 FILLER_77_1922 ();
 sg13g2_fill_1 FILLER_77_1924 ();
 sg13g2_fill_2 FILLER_77_2034 ();
 sg13g2_fill_1 FILLER_77_2044 ();
 sg13g2_fill_2 FILLER_77_2050 ();
 sg13g2_decap_4 FILLER_77_2061 ();
 sg13g2_fill_1 FILLER_77_2065 ();
 sg13g2_fill_1 FILLER_77_2080 ();
 sg13g2_fill_2 FILLER_77_2121 ();
 sg13g2_fill_1 FILLER_77_2123 ();
 sg13g2_fill_2 FILLER_77_2176 ();
 sg13g2_fill_1 FILLER_77_2178 ();
 sg13g2_decap_4 FILLER_77_2219 ();
 sg13g2_decap_8 FILLER_77_2240 ();
 sg13g2_decap_8 FILLER_77_2247 ();
 sg13g2_decap_8 FILLER_77_2254 ();
 sg13g2_decap_8 FILLER_77_2261 ();
 sg13g2_decap_8 FILLER_77_2268 ();
 sg13g2_decap_8 FILLER_77_2275 ();
 sg13g2_decap_8 FILLER_77_2282 ();
 sg13g2_decap_8 FILLER_77_2289 ();
 sg13g2_decap_8 FILLER_77_2296 ();
 sg13g2_decap_8 FILLER_77_2303 ();
 sg13g2_decap_8 FILLER_77_2310 ();
 sg13g2_decap_8 FILLER_77_2317 ();
 sg13g2_decap_8 FILLER_77_2324 ();
 sg13g2_decap_8 FILLER_77_2331 ();
 sg13g2_decap_8 FILLER_77_2338 ();
 sg13g2_decap_8 FILLER_77_2345 ();
 sg13g2_decap_8 FILLER_77_2352 ();
 sg13g2_decap_8 FILLER_77_2359 ();
 sg13g2_decap_8 FILLER_77_2366 ();
 sg13g2_decap_8 FILLER_77_2373 ();
 sg13g2_decap_8 FILLER_77_2380 ();
 sg13g2_decap_8 FILLER_77_2387 ();
 sg13g2_decap_8 FILLER_77_2394 ();
 sg13g2_decap_8 FILLER_77_2401 ();
 sg13g2_decap_8 FILLER_77_2408 ();
 sg13g2_decap_8 FILLER_77_2415 ();
 sg13g2_decap_8 FILLER_77_2422 ();
 sg13g2_decap_8 FILLER_77_2429 ();
 sg13g2_decap_8 FILLER_77_2436 ();
 sg13g2_decap_8 FILLER_77_2443 ();
 sg13g2_decap_8 FILLER_77_2450 ();
 sg13g2_decap_8 FILLER_77_2457 ();
 sg13g2_decap_8 FILLER_77_2464 ();
 sg13g2_decap_8 FILLER_77_2471 ();
 sg13g2_decap_8 FILLER_77_2478 ();
 sg13g2_decap_8 FILLER_77_2485 ();
 sg13g2_decap_8 FILLER_77_2492 ();
 sg13g2_decap_8 FILLER_77_2499 ();
 sg13g2_decap_8 FILLER_77_2506 ();
 sg13g2_decap_8 FILLER_77_2513 ();
 sg13g2_decap_8 FILLER_77_2520 ();
 sg13g2_decap_8 FILLER_77_2527 ();
 sg13g2_decap_8 FILLER_77_2534 ();
 sg13g2_decap_8 FILLER_77_2541 ();
 sg13g2_decap_8 FILLER_77_2548 ();
 sg13g2_decap_8 FILLER_77_2555 ();
 sg13g2_decap_8 FILLER_77_2562 ();
 sg13g2_decap_8 FILLER_77_2569 ();
 sg13g2_decap_8 FILLER_77_2576 ();
 sg13g2_decap_8 FILLER_77_2583 ();
 sg13g2_decap_8 FILLER_77_2590 ();
 sg13g2_decap_8 FILLER_77_2597 ();
 sg13g2_decap_8 FILLER_77_2604 ();
 sg13g2_decap_8 FILLER_77_2611 ();
 sg13g2_decap_8 FILLER_77_2618 ();
 sg13g2_decap_8 FILLER_77_2625 ();
 sg13g2_decap_8 FILLER_77_2632 ();
 sg13g2_decap_8 FILLER_77_2639 ();
 sg13g2_decap_8 FILLER_77_2646 ();
 sg13g2_decap_8 FILLER_77_2653 ();
 sg13g2_decap_8 FILLER_77_2660 ();
 sg13g2_decap_8 FILLER_77_2667 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_decap_8 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_259 ();
 sg13g2_decap_8 FILLER_78_266 ();
 sg13g2_decap_8 FILLER_78_273 ();
 sg13g2_decap_8 FILLER_78_280 ();
 sg13g2_decap_8 FILLER_78_287 ();
 sg13g2_decap_8 FILLER_78_294 ();
 sg13g2_decap_8 FILLER_78_301 ();
 sg13g2_decap_8 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_decap_8 FILLER_78_322 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_357 ();
 sg13g2_decap_8 FILLER_78_364 ();
 sg13g2_decap_8 FILLER_78_371 ();
 sg13g2_decap_8 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_decap_8 FILLER_78_406 ();
 sg13g2_decap_8 FILLER_78_413 ();
 sg13g2_decap_8 FILLER_78_420 ();
 sg13g2_decap_8 FILLER_78_427 ();
 sg13g2_decap_8 FILLER_78_434 ();
 sg13g2_decap_8 FILLER_78_441 ();
 sg13g2_decap_8 FILLER_78_448 ();
 sg13g2_decap_8 FILLER_78_455 ();
 sg13g2_decap_8 FILLER_78_462 ();
 sg13g2_decap_8 FILLER_78_469 ();
 sg13g2_decap_8 FILLER_78_476 ();
 sg13g2_decap_8 FILLER_78_483 ();
 sg13g2_decap_8 FILLER_78_490 ();
 sg13g2_decap_8 FILLER_78_497 ();
 sg13g2_decap_8 FILLER_78_504 ();
 sg13g2_decap_8 FILLER_78_511 ();
 sg13g2_decap_4 FILLER_78_518 ();
 sg13g2_fill_1 FILLER_78_522 ();
 sg13g2_fill_2 FILLER_78_540 ();
 sg13g2_fill_1 FILLER_78_542 ();
 sg13g2_fill_2 FILLER_78_567 ();
 sg13g2_fill_2 FILLER_78_582 ();
 sg13g2_fill_1 FILLER_78_584 ();
 sg13g2_decap_4 FILLER_78_594 ();
 sg13g2_fill_2 FILLER_78_598 ();
 sg13g2_fill_2 FILLER_78_639 ();
 sg13g2_fill_1 FILLER_78_641 ();
 sg13g2_fill_1 FILLER_78_646 ();
 sg13g2_decap_8 FILLER_78_656 ();
 sg13g2_fill_2 FILLER_78_675 ();
 sg13g2_fill_2 FILLER_78_686 ();
 sg13g2_fill_2 FILLER_78_695 ();
 sg13g2_fill_1 FILLER_78_697 ();
 sg13g2_decap_4 FILLER_78_715 ();
 sg13g2_fill_2 FILLER_78_759 ();
 sg13g2_fill_1 FILLER_78_761 ();
 sg13g2_fill_2 FILLER_78_792 ();
 sg13g2_fill_2 FILLER_78_815 ();
 sg13g2_fill_2 FILLER_78_839 ();
 sg13g2_fill_1 FILLER_78_841 ();
 sg13g2_fill_2 FILLER_78_873 ();
 sg13g2_fill_1 FILLER_78_875 ();
 sg13g2_fill_1 FILLER_78_903 ();
 sg13g2_decap_8 FILLER_78_935 ();
 sg13g2_decap_8 FILLER_78_942 ();
 sg13g2_decap_8 FILLER_78_949 ();
 sg13g2_decap_4 FILLER_78_956 ();
 sg13g2_fill_2 FILLER_78_991 ();
 sg13g2_fill_2 FILLER_78_1090 ();
 sg13g2_fill_2 FILLER_78_1106 ();
 sg13g2_fill_1 FILLER_78_1108 ();
 sg13g2_fill_2 FILLER_78_1154 ();
 sg13g2_fill_1 FILLER_78_1156 ();
 sg13g2_decap_8 FILLER_78_1161 ();
 sg13g2_decap_8 FILLER_78_1168 ();
 sg13g2_fill_1 FILLER_78_1175 ();
 sg13g2_fill_2 FILLER_78_1198 ();
 sg13g2_decap_4 FILLER_78_1226 ();
 sg13g2_fill_1 FILLER_78_1230 ();
 sg13g2_fill_2 FILLER_78_1262 ();
 sg13g2_fill_2 FILLER_78_1293 ();
 sg13g2_fill_1 FILLER_78_1295 ();
 sg13g2_fill_2 FILLER_78_1322 ();
 sg13g2_fill_1 FILLER_78_1351 ();
 sg13g2_fill_2 FILLER_78_1357 ();
 sg13g2_fill_1 FILLER_78_1359 ();
 sg13g2_fill_2 FILLER_78_1365 ();
 sg13g2_fill_1 FILLER_78_1367 ();
 sg13g2_decap_4 FILLER_78_1402 ();
 sg13g2_fill_2 FILLER_78_1446 ();
 sg13g2_decap_8 FILLER_78_1471 ();
 sg13g2_fill_2 FILLER_78_1478 ();
 sg13g2_fill_1 FILLER_78_1480 ();
 sg13g2_fill_2 FILLER_78_1490 ();
 sg13g2_fill_1 FILLER_78_1492 ();
 sg13g2_fill_2 FILLER_78_1568 ();
 sg13g2_fill_1 FILLER_78_1579 ();
 sg13g2_fill_2 FILLER_78_1594 ();
 sg13g2_fill_1 FILLER_78_1631 ();
 sg13g2_decap_4 FILLER_78_1658 ();
 sg13g2_fill_2 FILLER_78_1662 ();
 sg13g2_fill_2 FILLER_78_1678 ();
 sg13g2_fill_1 FILLER_78_1680 ();
 sg13g2_fill_1 FILLER_78_1736 ();
 sg13g2_decap_4 FILLER_78_1741 ();
 sg13g2_fill_2 FILLER_78_1750 ();
 sg13g2_fill_1 FILLER_78_1752 ();
 sg13g2_fill_2 FILLER_78_1770 ();
 sg13g2_fill_1 FILLER_78_1821 ();
 sg13g2_fill_2 FILLER_78_1834 ();
 sg13g2_fill_2 FILLER_78_1892 ();
 sg13g2_fill_1 FILLER_78_1894 ();
 sg13g2_fill_1 FILLER_78_1899 ();
 sg13g2_fill_1 FILLER_78_1909 ();
 sg13g2_fill_1 FILLER_78_1915 ();
 sg13g2_fill_2 FILLER_78_1951 ();
 sg13g2_fill_1 FILLER_78_1953 ();
 sg13g2_decap_8 FILLER_78_1958 ();
 sg13g2_decap_4 FILLER_78_1965 ();
 sg13g2_fill_1 FILLER_78_1974 ();
 sg13g2_decap_8 FILLER_78_1979 ();
 sg13g2_fill_1 FILLER_78_1986 ();
 sg13g2_fill_2 FILLER_78_2008 ();
 sg13g2_fill_1 FILLER_78_2010 ();
 sg13g2_fill_2 FILLER_78_2016 ();
 sg13g2_fill_1 FILLER_78_2018 ();
 sg13g2_fill_1 FILLER_78_2047 ();
 sg13g2_fill_2 FILLER_78_2117 ();
 sg13g2_fill_2 FILLER_78_2133 ();
 sg13g2_fill_1 FILLER_78_2135 ();
 sg13g2_fill_2 FILLER_78_2145 ();
 sg13g2_fill_2 FILLER_78_2207 ();
 sg13g2_decap_8 FILLER_78_2240 ();
 sg13g2_decap_8 FILLER_78_2247 ();
 sg13g2_decap_8 FILLER_78_2254 ();
 sg13g2_decap_8 FILLER_78_2261 ();
 sg13g2_decap_8 FILLER_78_2268 ();
 sg13g2_decap_8 FILLER_78_2275 ();
 sg13g2_decap_8 FILLER_78_2282 ();
 sg13g2_decap_8 FILLER_78_2289 ();
 sg13g2_decap_8 FILLER_78_2296 ();
 sg13g2_decap_8 FILLER_78_2303 ();
 sg13g2_decap_8 FILLER_78_2310 ();
 sg13g2_decap_8 FILLER_78_2317 ();
 sg13g2_decap_8 FILLER_78_2324 ();
 sg13g2_decap_8 FILLER_78_2331 ();
 sg13g2_decap_8 FILLER_78_2338 ();
 sg13g2_decap_8 FILLER_78_2345 ();
 sg13g2_decap_8 FILLER_78_2352 ();
 sg13g2_decap_8 FILLER_78_2359 ();
 sg13g2_decap_8 FILLER_78_2366 ();
 sg13g2_decap_8 FILLER_78_2373 ();
 sg13g2_decap_8 FILLER_78_2380 ();
 sg13g2_decap_8 FILLER_78_2387 ();
 sg13g2_decap_8 FILLER_78_2394 ();
 sg13g2_decap_8 FILLER_78_2401 ();
 sg13g2_decap_8 FILLER_78_2408 ();
 sg13g2_decap_8 FILLER_78_2415 ();
 sg13g2_decap_8 FILLER_78_2422 ();
 sg13g2_decap_8 FILLER_78_2429 ();
 sg13g2_decap_8 FILLER_78_2436 ();
 sg13g2_decap_8 FILLER_78_2443 ();
 sg13g2_decap_8 FILLER_78_2450 ();
 sg13g2_decap_8 FILLER_78_2457 ();
 sg13g2_decap_8 FILLER_78_2464 ();
 sg13g2_decap_8 FILLER_78_2471 ();
 sg13g2_decap_8 FILLER_78_2478 ();
 sg13g2_decap_8 FILLER_78_2485 ();
 sg13g2_decap_8 FILLER_78_2492 ();
 sg13g2_decap_8 FILLER_78_2499 ();
 sg13g2_decap_8 FILLER_78_2506 ();
 sg13g2_decap_8 FILLER_78_2513 ();
 sg13g2_decap_8 FILLER_78_2520 ();
 sg13g2_decap_8 FILLER_78_2527 ();
 sg13g2_decap_8 FILLER_78_2534 ();
 sg13g2_decap_8 FILLER_78_2541 ();
 sg13g2_decap_8 FILLER_78_2548 ();
 sg13g2_decap_8 FILLER_78_2555 ();
 sg13g2_decap_8 FILLER_78_2562 ();
 sg13g2_decap_8 FILLER_78_2569 ();
 sg13g2_decap_8 FILLER_78_2576 ();
 sg13g2_decap_8 FILLER_78_2583 ();
 sg13g2_decap_8 FILLER_78_2590 ();
 sg13g2_decap_8 FILLER_78_2597 ();
 sg13g2_decap_8 FILLER_78_2604 ();
 sg13g2_decap_8 FILLER_78_2611 ();
 sg13g2_decap_8 FILLER_78_2618 ();
 sg13g2_decap_8 FILLER_78_2625 ();
 sg13g2_decap_8 FILLER_78_2632 ();
 sg13g2_decap_8 FILLER_78_2639 ();
 sg13g2_decap_8 FILLER_78_2646 ();
 sg13g2_decap_8 FILLER_78_2653 ();
 sg13g2_decap_8 FILLER_78_2660 ();
 sg13g2_decap_8 FILLER_78_2667 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_decap_8 FILLER_79_245 ();
 sg13g2_decap_8 FILLER_79_252 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_decap_8 FILLER_79_266 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_decap_8 FILLER_79_280 ();
 sg13g2_decap_8 FILLER_79_287 ();
 sg13g2_decap_8 FILLER_79_294 ();
 sg13g2_decap_8 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_decap_8 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_79_329 ();
 sg13g2_decap_8 FILLER_79_336 ();
 sg13g2_decap_8 FILLER_79_343 ();
 sg13g2_decap_8 FILLER_79_350 ();
 sg13g2_decap_8 FILLER_79_357 ();
 sg13g2_decap_8 FILLER_79_364 ();
 sg13g2_decap_8 FILLER_79_371 ();
 sg13g2_decap_8 FILLER_79_378 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_decap_8 FILLER_79_406 ();
 sg13g2_decap_8 FILLER_79_413 ();
 sg13g2_decap_8 FILLER_79_420 ();
 sg13g2_decap_8 FILLER_79_427 ();
 sg13g2_decap_8 FILLER_79_434 ();
 sg13g2_decap_8 FILLER_79_441 ();
 sg13g2_decap_8 FILLER_79_448 ();
 sg13g2_decap_8 FILLER_79_455 ();
 sg13g2_decap_8 FILLER_79_462 ();
 sg13g2_decap_8 FILLER_79_469 ();
 sg13g2_decap_8 FILLER_79_476 ();
 sg13g2_decap_8 FILLER_79_483 ();
 sg13g2_decap_8 FILLER_79_490 ();
 sg13g2_decap_8 FILLER_79_497 ();
 sg13g2_decap_8 FILLER_79_504 ();
 sg13g2_decap_8 FILLER_79_511 ();
 sg13g2_decap_8 FILLER_79_518 ();
 sg13g2_fill_2 FILLER_79_525 ();
 sg13g2_fill_1 FILLER_79_527 ();
 sg13g2_fill_2 FILLER_79_615 ();
 sg13g2_fill_1 FILLER_79_617 ();
 sg13g2_decap_8 FILLER_79_649 ();
 sg13g2_decap_8 FILLER_79_656 ();
 sg13g2_decap_8 FILLER_79_663 ();
 sg13g2_decap_8 FILLER_79_670 ();
 sg13g2_decap_8 FILLER_79_677 ();
 sg13g2_decap_8 FILLER_79_684 ();
 sg13g2_fill_2 FILLER_79_691 ();
 sg13g2_fill_1 FILLER_79_728 ();
 sg13g2_fill_1 FILLER_79_746 ();
 sg13g2_fill_2 FILLER_79_761 ();
 sg13g2_fill_2 FILLER_79_833 ();
 sg13g2_fill_2 FILLER_79_840 ();
 sg13g2_fill_1 FILLER_79_842 ();
 sg13g2_fill_2 FILLER_79_856 ();
 sg13g2_fill_2 FILLER_79_862 ();
 sg13g2_fill_1 FILLER_79_864 ();
 sg13g2_decap_4 FILLER_79_896 ();
 sg13g2_decap_4 FILLER_79_904 ();
 sg13g2_decap_4 FILLER_79_912 ();
 sg13g2_fill_2 FILLER_79_916 ();
 sg13g2_decap_8 FILLER_79_931 ();
 sg13g2_decap_8 FILLER_79_938 ();
 sg13g2_decap_8 FILLER_79_945 ();
 sg13g2_decap_8 FILLER_79_952 ();
 sg13g2_decap_4 FILLER_79_959 ();
 sg13g2_fill_2 FILLER_79_963 ();
 sg13g2_fill_1 FILLER_79_991 ();
 sg13g2_fill_1 FILLER_79_1024 ();
 sg13g2_decap_4 FILLER_79_1042 ();
 sg13g2_fill_2 FILLER_79_1050 ();
 sg13g2_decap_8 FILLER_79_1056 ();
 sg13g2_decap_8 FILLER_79_1063 ();
 sg13g2_fill_2 FILLER_79_1101 ();
 sg13g2_fill_1 FILLER_79_1103 ();
 sg13g2_fill_2 FILLER_79_1117 ();
 sg13g2_decap_4 FILLER_79_1123 ();
 sg13g2_fill_2 FILLER_79_1140 ();
 sg13g2_decap_8 FILLER_79_1155 ();
 sg13g2_decap_8 FILLER_79_1162 ();
 sg13g2_decap_8 FILLER_79_1169 ();
 sg13g2_decap_8 FILLER_79_1176 ();
 sg13g2_fill_2 FILLER_79_1183 ();
 sg13g2_fill_1 FILLER_79_1185 ();
 sg13g2_decap_8 FILLER_79_1238 ();
 sg13g2_fill_1 FILLER_79_1245 ();
 sg13g2_fill_2 FILLER_79_1298 ();
 sg13g2_fill_1 FILLER_79_1300 ();
 sg13g2_fill_2 FILLER_79_1306 ();
 sg13g2_fill_1 FILLER_79_1308 ();
 sg13g2_fill_1 FILLER_79_1371 ();
 sg13g2_fill_2 FILLER_79_1399 ();
 sg13g2_fill_1 FILLER_79_1401 ();
 sg13g2_fill_1 FILLER_79_1411 ();
 sg13g2_fill_1 FILLER_79_1448 ();
 sg13g2_decap_4 FILLER_79_1475 ();
 sg13g2_decap_8 FILLER_79_1505 ();
 sg13g2_fill_2 FILLER_79_1512 ();
 sg13g2_fill_1 FILLER_79_1518 ();
 sg13g2_decap_8 FILLER_79_1528 ();
 sg13g2_fill_2 FILLER_79_1535 ();
 sg13g2_fill_1 FILLER_79_1537 ();
 sg13g2_fill_2 FILLER_79_1542 ();
 sg13g2_fill_1 FILLER_79_1544 ();
 sg13g2_fill_2 FILLER_79_1646 ();
 sg13g2_fill_1 FILLER_79_1648 ();
 sg13g2_decap_4 FILLER_79_1661 ();
 sg13g2_fill_2 FILLER_79_1725 ();
 sg13g2_fill_2 FILLER_79_1741 ();
 sg13g2_fill_1 FILLER_79_1743 ();
 sg13g2_decap_4 FILLER_79_1789 ();
 sg13g2_fill_1 FILLER_79_1793 ();
 sg13g2_decap_8 FILLER_79_1846 ();
 sg13g2_fill_2 FILLER_79_1862 ();
 sg13g2_fill_1 FILLER_79_1864 ();
 sg13g2_fill_1 FILLER_79_1869 ();
 sg13g2_fill_2 FILLER_79_1901 ();
 sg13g2_fill_2 FILLER_79_1908 ();
 sg13g2_fill_1 FILLER_79_1910 ();
 sg13g2_decap_4 FILLER_79_1945 ();
 sg13g2_decap_4 FILLER_79_2053 ();
 sg13g2_fill_2 FILLER_79_2057 ();
 sg13g2_decap_8 FILLER_79_2063 ();
 sg13g2_decap_8 FILLER_79_2070 ();
 sg13g2_decap_8 FILLER_79_2086 ();
 sg13g2_fill_2 FILLER_79_2093 ();
 sg13g2_fill_2 FILLER_79_2112 ();
 sg13g2_fill_1 FILLER_79_2171 ();
 sg13g2_decap_8 FILLER_79_2229 ();
 sg13g2_decap_8 FILLER_79_2236 ();
 sg13g2_decap_8 FILLER_79_2243 ();
 sg13g2_decap_8 FILLER_79_2250 ();
 sg13g2_decap_8 FILLER_79_2257 ();
 sg13g2_decap_8 FILLER_79_2264 ();
 sg13g2_decap_8 FILLER_79_2271 ();
 sg13g2_decap_8 FILLER_79_2278 ();
 sg13g2_decap_8 FILLER_79_2285 ();
 sg13g2_decap_8 FILLER_79_2292 ();
 sg13g2_decap_8 FILLER_79_2299 ();
 sg13g2_decap_8 FILLER_79_2306 ();
 sg13g2_decap_8 FILLER_79_2313 ();
 sg13g2_decap_8 FILLER_79_2320 ();
 sg13g2_decap_8 FILLER_79_2327 ();
 sg13g2_decap_8 FILLER_79_2334 ();
 sg13g2_decap_8 FILLER_79_2341 ();
 sg13g2_decap_8 FILLER_79_2348 ();
 sg13g2_decap_8 FILLER_79_2355 ();
 sg13g2_decap_8 FILLER_79_2362 ();
 sg13g2_decap_8 FILLER_79_2369 ();
 sg13g2_decap_8 FILLER_79_2376 ();
 sg13g2_decap_8 FILLER_79_2383 ();
 sg13g2_decap_8 FILLER_79_2390 ();
 sg13g2_decap_8 FILLER_79_2397 ();
 sg13g2_decap_8 FILLER_79_2404 ();
 sg13g2_decap_8 FILLER_79_2411 ();
 sg13g2_decap_8 FILLER_79_2418 ();
 sg13g2_decap_8 FILLER_79_2425 ();
 sg13g2_decap_8 FILLER_79_2432 ();
 sg13g2_decap_8 FILLER_79_2439 ();
 sg13g2_decap_8 FILLER_79_2446 ();
 sg13g2_decap_8 FILLER_79_2453 ();
 sg13g2_decap_8 FILLER_79_2460 ();
 sg13g2_decap_8 FILLER_79_2467 ();
 sg13g2_decap_8 FILLER_79_2474 ();
 sg13g2_decap_8 FILLER_79_2481 ();
 sg13g2_decap_8 FILLER_79_2488 ();
 sg13g2_decap_8 FILLER_79_2495 ();
 sg13g2_decap_8 FILLER_79_2502 ();
 sg13g2_decap_8 FILLER_79_2509 ();
 sg13g2_decap_8 FILLER_79_2516 ();
 sg13g2_decap_8 FILLER_79_2523 ();
 sg13g2_decap_8 FILLER_79_2530 ();
 sg13g2_decap_8 FILLER_79_2537 ();
 sg13g2_decap_8 FILLER_79_2544 ();
 sg13g2_decap_8 FILLER_79_2551 ();
 sg13g2_decap_8 FILLER_79_2558 ();
 sg13g2_decap_8 FILLER_79_2565 ();
 sg13g2_decap_8 FILLER_79_2572 ();
 sg13g2_decap_8 FILLER_79_2579 ();
 sg13g2_decap_8 FILLER_79_2586 ();
 sg13g2_decap_8 FILLER_79_2593 ();
 sg13g2_decap_8 FILLER_79_2600 ();
 sg13g2_decap_8 FILLER_79_2607 ();
 sg13g2_decap_8 FILLER_79_2614 ();
 sg13g2_decap_8 FILLER_79_2621 ();
 sg13g2_decap_8 FILLER_79_2628 ();
 sg13g2_decap_8 FILLER_79_2635 ();
 sg13g2_decap_8 FILLER_79_2642 ();
 sg13g2_decap_8 FILLER_79_2649 ();
 sg13g2_decap_8 FILLER_79_2656 ();
 sg13g2_decap_8 FILLER_79_2663 ();
 sg13g2_decap_4 FILLER_79_2670 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_8 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_147 ();
 sg13g2_fill_1 FILLER_80_151 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_8 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_171 ();
 sg13g2_fill_1 FILLER_80_175 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_8 FILLER_80_229 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_decap_8 FILLER_80_243 ();
 sg13g2_decap_8 FILLER_80_250 ();
 sg13g2_decap_8 FILLER_80_257 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_fill_2 FILLER_80_278 ();
 sg13g2_decap_8 FILLER_80_288 ();
 sg13g2_decap_8 FILLER_80_295 ();
 sg13g2_fill_2 FILLER_80_302 ();
 sg13g2_decap_8 FILLER_80_384 ();
 sg13g2_decap_8 FILLER_80_391 ();
 sg13g2_decap_8 FILLER_80_398 ();
 sg13g2_decap_8 FILLER_80_405 ();
 sg13g2_decap_8 FILLER_80_412 ();
 sg13g2_decap_8 FILLER_80_419 ();
 sg13g2_decap_8 FILLER_80_426 ();
 sg13g2_decap_8 FILLER_80_433 ();
 sg13g2_decap_8 FILLER_80_440 ();
 sg13g2_decap_8 FILLER_80_447 ();
 sg13g2_decap_8 FILLER_80_454 ();
 sg13g2_decap_8 FILLER_80_461 ();
 sg13g2_decap_8 FILLER_80_468 ();
 sg13g2_decap_8 FILLER_80_475 ();
 sg13g2_decap_8 FILLER_80_482 ();
 sg13g2_decap_8 FILLER_80_489 ();
 sg13g2_decap_8 FILLER_80_496 ();
 sg13g2_decap_8 FILLER_80_503 ();
 sg13g2_decap_8 FILLER_80_510 ();
 sg13g2_decap_8 FILLER_80_517 ();
 sg13g2_decap_8 FILLER_80_524 ();
 sg13g2_decap_4 FILLER_80_531 ();
 sg13g2_fill_2 FILLER_80_543 ();
 sg13g2_fill_1 FILLER_80_545 ();
 sg13g2_fill_2 FILLER_80_551 ();
 sg13g2_decap_8 FILLER_80_566 ();
 sg13g2_decap_8 FILLER_80_573 ();
 sg13g2_decap_8 FILLER_80_580 ();
 sg13g2_decap_4 FILLER_80_587 ();
 sg13g2_decap_8 FILLER_80_595 ();
 sg13g2_decap_8 FILLER_80_602 ();
 sg13g2_fill_2 FILLER_80_609 ();
 sg13g2_decap_8 FILLER_80_615 ();
 sg13g2_decap_8 FILLER_80_622 ();
 sg13g2_decap_4 FILLER_80_629 ();
 sg13g2_fill_1 FILLER_80_633 ();
 sg13g2_fill_1 FILLER_80_638 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_669 ();
 sg13g2_decap_8 FILLER_80_676 ();
 sg13g2_decap_8 FILLER_80_683 ();
 sg13g2_decap_4 FILLER_80_690 ();
 sg13g2_fill_1 FILLER_80_720 ();
 sg13g2_fill_1 FILLER_80_747 ();
 sg13g2_decap_8 FILLER_80_801 ();
 sg13g2_fill_1 FILLER_80_808 ();
 sg13g2_decap_8 FILLER_80_813 ();
 sg13g2_decap_4 FILLER_80_820 ();
 sg13g2_fill_2 FILLER_80_829 ();
 sg13g2_fill_2 FILLER_80_880 ();
 sg13g2_fill_1 FILLER_80_882 ();
 sg13g2_decap_8 FILLER_80_900 ();
 sg13g2_decap_8 FILLER_80_907 ();
 sg13g2_decap_8 FILLER_80_914 ();
 sg13g2_decap_8 FILLER_80_921 ();
 sg13g2_decap_8 FILLER_80_928 ();
 sg13g2_decap_8 FILLER_80_935 ();
 sg13g2_decap_8 FILLER_80_942 ();
 sg13g2_decap_8 FILLER_80_949 ();
 sg13g2_decap_8 FILLER_80_956 ();
 sg13g2_decap_8 FILLER_80_963 ();
 sg13g2_decap_8 FILLER_80_970 ();
 sg13g2_fill_1 FILLER_80_977 ();
 sg13g2_fill_1 FILLER_80_1004 ();
 sg13g2_decap_8 FILLER_80_1070 ();
 sg13g2_decap_4 FILLER_80_1077 ();
 sg13g2_fill_1 FILLER_80_1081 ();
 sg13g2_fill_2 FILLER_80_1134 ();
 sg13g2_fill_1 FILLER_80_1136 ();
 sg13g2_decap_8 FILLER_80_1145 ();
 sg13g2_decap_8 FILLER_80_1152 ();
 sg13g2_decap_8 FILLER_80_1159 ();
 sg13g2_decap_8 FILLER_80_1166 ();
 sg13g2_decap_8 FILLER_80_1173 ();
 sg13g2_decap_8 FILLER_80_1180 ();
 sg13g2_decap_8 FILLER_80_1187 ();
 sg13g2_fill_1 FILLER_80_1198 ();
 sg13g2_fill_1 FILLER_80_1203 ();
 sg13g2_fill_2 FILLER_80_1213 ();
 sg13g2_fill_1 FILLER_80_1215 ();
 sg13g2_decap_8 FILLER_80_1233 ();
 sg13g2_decap_8 FILLER_80_1240 ();
 sg13g2_decap_8 FILLER_80_1247 ();
 sg13g2_decap_8 FILLER_80_1271 ();
 sg13g2_fill_2 FILLER_80_1278 ();
 sg13g2_fill_2 FILLER_80_1288 ();
 sg13g2_fill_1 FILLER_80_1290 ();
 sg13g2_fill_2 FILLER_80_1304 ();
 sg13g2_fill_1 FILLER_80_1306 ();
 sg13g2_fill_1 FILLER_80_1320 ();
 sg13g2_fill_1 FILLER_80_1330 ();
 sg13g2_fill_1 FILLER_80_1339 ();
 sg13g2_fill_2 FILLER_80_1356 ();
 sg13g2_fill_1 FILLER_80_1358 ();
 sg13g2_fill_2 FILLER_80_1420 ();
 sg13g2_fill_2 FILLER_80_1426 ();
 sg13g2_fill_2 FILLER_80_1458 ();
 sg13g2_fill_1 FILLER_80_1460 ();
 sg13g2_decap_8 FILLER_80_1478 ();
 sg13g2_decap_4 FILLER_80_1485 ();
 sg13g2_fill_1 FILLER_80_1489 ();
 sg13g2_fill_2 FILLER_80_1498 ();
 sg13g2_decap_8 FILLER_80_1509 ();
 sg13g2_decap_8 FILLER_80_1516 ();
 sg13g2_decap_8 FILLER_80_1523 ();
 sg13g2_decap_8 FILLER_80_1530 ();
 sg13g2_decap_4 FILLER_80_1537 ();
 sg13g2_decap_4 FILLER_80_1571 ();
 sg13g2_fill_2 FILLER_80_1587 ();
 sg13g2_fill_1 FILLER_80_1589 ();
 sg13g2_fill_1 FILLER_80_1602 ();
 sg13g2_fill_1 FILLER_80_1612 ();
 sg13g2_decap_8 FILLER_80_1652 ();
 sg13g2_decap_8 FILLER_80_1659 ();
 sg13g2_decap_4 FILLER_80_1666 ();
 sg13g2_fill_2 FILLER_80_1670 ();
 sg13g2_decap_4 FILLER_80_1693 ();
 sg13g2_fill_2 FILLER_80_1697 ();
 sg13g2_fill_2 FILLER_80_1707 ();
 sg13g2_decap_8 FILLER_80_1718 ();
 sg13g2_fill_1 FILLER_80_1725 ();
 sg13g2_fill_1 FILLER_80_1761 ();
 sg13g2_decap_8 FILLER_80_1774 ();
 sg13g2_decap_8 FILLER_80_1781 ();
 sg13g2_decap_8 FILLER_80_1788 ();
 sg13g2_decap_8 FILLER_80_1795 ();
 sg13g2_fill_2 FILLER_80_1802 ();
 sg13g2_fill_1 FILLER_80_1804 ();
 sg13g2_decap_8 FILLER_80_1835 ();
 sg13g2_decap_4 FILLER_80_1842 ();
 sg13g2_fill_2 FILLER_80_1846 ();
 sg13g2_fill_2 FILLER_80_1874 ();
 sg13g2_fill_1 FILLER_80_1876 ();
 sg13g2_decap_8 FILLER_80_1934 ();
 sg13g2_decap_8 FILLER_80_1941 ();
 sg13g2_decap_8 FILLER_80_1948 ();
 sg13g2_fill_2 FILLER_80_1955 ();
 sg13g2_fill_1 FILLER_80_1957 ();
 sg13g2_fill_1 FILLER_80_1971 ();
 sg13g2_decap_4 FILLER_80_1976 ();
 sg13g2_fill_1 FILLER_80_1980 ();
 sg13g2_fill_1 FILLER_80_1985 ();
 sg13g2_fill_2 FILLER_80_2018 ();
 sg13g2_fill_1 FILLER_80_2037 ();
 sg13g2_decap_8 FILLER_80_2051 ();
 sg13g2_decap_8 FILLER_80_2058 ();
 sg13g2_decap_8 FILLER_80_2065 ();
 sg13g2_decap_8 FILLER_80_2072 ();
 sg13g2_decap_4 FILLER_80_2079 ();
 sg13g2_fill_1 FILLER_80_2083 ();
 sg13g2_fill_1 FILLER_80_2131 ();
 sg13g2_fill_1 FILLER_80_2141 ();
 sg13g2_decap_8 FILLER_80_2171 ();
 sg13g2_fill_1 FILLER_80_2204 ();
 sg13g2_fill_2 FILLER_80_2209 ();
 sg13g2_decap_8 FILLER_80_2224 ();
 sg13g2_decap_8 FILLER_80_2231 ();
 sg13g2_decap_8 FILLER_80_2238 ();
 sg13g2_decap_8 FILLER_80_2245 ();
 sg13g2_decap_8 FILLER_80_2252 ();
 sg13g2_decap_8 FILLER_80_2259 ();
 sg13g2_decap_8 FILLER_80_2266 ();
 sg13g2_decap_8 FILLER_80_2273 ();
 sg13g2_decap_8 FILLER_80_2280 ();
 sg13g2_decap_8 FILLER_80_2287 ();
 sg13g2_decap_8 FILLER_80_2294 ();
 sg13g2_decap_8 FILLER_80_2301 ();
 sg13g2_decap_8 FILLER_80_2308 ();
 sg13g2_decap_8 FILLER_80_2315 ();
 sg13g2_decap_8 FILLER_80_2322 ();
 sg13g2_decap_8 FILLER_80_2329 ();
 sg13g2_decap_8 FILLER_80_2336 ();
 sg13g2_decap_8 FILLER_80_2343 ();
 sg13g2_decap_8 FILLER_80_2350 ();
 sg13g2_decap_8 FILLER_80_2357 ();
 sg13g2_decap_8 FILLER_80_2364 ();
 sg13g2_decap_8 FILLER_80_2371 ();
 sg13g2_decap_8 FILLER_80_2378 ();
 sg13g2_decap_8 FILLER_80_2385 ();
 sg13g2_decap_8 FILLER_80_2392 ();
 sg13g2_decap_8 FILLER_80_2399 ();
 sg13g2_decap_8 FILLER_80_2406 ();
 sg13g2_decap_8 FILLER_80_2413 ();
 sg13g2_decap_8 FILLER_80_2420 ();
 sg13g2_decap_8 FILLER_80_2427 ();
 sg13g2_decap_8 FILLER_80_2434 ();
 sg13g2_decap_8 FILLER_80_2441 ();
 sg13g2_decap_8 FILLER_80_2448 ();
 sg13g2_decap_8 FILLER_80_2455 ();
 sg13g2_decap_8 FILLER_80_2462 ();
 sg13g2_decap_8 FILLER_80_2469 ();
 sg13g2_decap_8 FILLER_80_2476 ();
 sg13g2_decap_8 FILLER_80_2483 ();
 sg13g2_decap_8 FILLER_80_2490 ();
 sg13g2_decap_8 FILLER_80_2497 ();
 sg13g2_decap_8 FILLER_80_2504 ();
 sg13g2_decap_8 FILLER_80_2511 ();
 sg13g2_decap_8 FILLER_80_2518 ();
 sg13g2_decap_8 FILLER_80_2525 ();
 sg13g2_decap_8 FILLER_80_2532 ();
 sg13g2_decap_8 FILLER_80_2539 ();
 sg13g2_decap_8 FILLER_80_2546 ();
 sg13g2_decap_8 FILLER_80_2553 ();
 sg13g2_decap_8 FILLER_80_2560 ();
 sg13g2_decap_8 FILLER_80_2567 ();
 sg13g2_decap_8 FILLER_80_2574 ();
 sg13g2_decap_8 FILLER_80_2581 ();
 sg13g2_decap_8 FILLER_80_2588 ();
 sg13g2_decap_8 FILLER_80_2595 ();
 sg13g2_decap_8 FILLER_80_2602 ();
 sg13g2_decap_8 FILLER_80_2609 ();
 sg13g2_decap_8 FILLER_80_2616 ();
 sg13g2_decap_8 FILLER_80_2623 ();
 sg13g2_decap_8 FILLER_80_2630 ();
 sg13g2_decap_8 FILLER_80_2637 ();
 sg13g2_decap_8 FILLER_80_2644 ();
 sg13g2_decap_8 FILLER_80_2651 ();
 sg13g2_decap_8 FILLER_80_2658 ();
 sg13g2_decap_8 FILLER_80_2665 ();
 sg13g2_fill_2 FILLER_80_2672 ();
 assign uio_oe[0] = net12;
 assign uio_oe[1] = net2130;
 assign uio_oe[2] = net13;
 assign uio_oe[3] = net14;
 assign uio_oe[4] = net2131;
 assign uio_oe[5] = net15;
 assign uio_oe[6] = net16;
 assign uio_oe[7] = net17;
 assign uio_out[0] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
 assign uio_out[7] = net23;
endmodule

module tt_um_hpdl1414_uart_atudoroi (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire \pmod_1414.GPout[0] ;
 wire \pmod_1414.GPout[1] ;
 wire \pmod_1414.GPout[2] ;
 wire \pmod_1414.GPout[3] ;
 wire \pmod_1414.GPout[4] ;
 wire \pmod_1414.GPout[5] ;
 wire \pmod_1414.GPout[6] ;
 wire \pmod_1414.GPout[7] ;
 wire \pmod_1414.HPDL_A0 ;
 wire \pmod_1414.HPDL_A1 ;
 wire \pmod_1414.HPDL_D0 ;
 wire \pmod_1414.HPDL_D1 ;
 wire \pmod_1414.HPDL_D2 ;
 wire \pmod_1414.HPDL_D3 ;
 wire \pmod_1414.HPDL_D4 ;
 wire \pmod_1414.HPDL_D5 ;
 wire \pmod_1414.HPDL_D6 ;
 wire \pmod_1414.HPDL_WR1 ;
 wire \pmod_1414.HPDL_WR2 ;
 wire \pmod_1414.HPDL_WR3 ;
 wire \pmod_1414.HPDL_WR4 ;
 wire \pmod_1414.RX.Filter_cnt[0] ;
 wire \pmod_1414.RX.Filter_cnt[1] ;
 wire \pmod_1414.RX.OversamplingCnt[0] ;
 wire \pmod_1414.RX.OversamplingCnt[1] ;
 wire \pmod_1414.RX.OversamplingCnt[2] ;
 wire \pmod_1414.RX.OversamplingCnt[3] ;
 wire \pmod_1414.RX.OversamplingTick ;
 wire \pmod_1414.RX.RxD_bit ;
 wire \pmod_1414.RX.RxD_data[0] ;
 wire \pmod_1414.RX.RxD_data[1] ;
 wire \pmod_1414.RX.RxD_data[2] ;
 wire \pmod_1414.RX.RxD_data[3] ;
 wire \pmod_1414.RX.RxD_data[4] ;
 wire \pmod_1414.RX.RxD_data[5] ;
 wire \pmod_1414.RX.RxD_data[6] ;
 wire \pmod_1414.RX.RxD_data[7] ;
 wire \pmod_1414.RX.RxD_data_ready ;
 wire \pmod_1414.RX.RxD_state[0] ;
 wire \pmod_1414.RX.RxD_state[1] ;
 wire \pmod_1414.RX.RxD_state[2] ;
 wire \pmod_1414.RX.RxD_state[3] ;
 wire \pmod_1414.RX.RxD_sync[0] ;
 wire \pmod_1414.RX.RxD_sync[1] ;
 wire \pmod_1414.RX.tickgen.Acc[0] ;
 wire \pmod_1414.RX.tickgen.Acc[10] ;
 wire \pmod_1414.RX.tickgen.Acc[11] ;
 wire \pmod_1414.RX.tickgen.Acc[12] ;
 wire \pmod_1414.RX.tickgen.Acc[13] ;
 wire \pmod_1414.RX.tickgen.Acc[14] ;
 wire \pmod_1414.RX.tickgen.Acc[1] ;
 wire \pmod_1414.RX.tickgen.Acc[2] ;
 wire \pmod_1414.RX.tickgen.Acc[3] ;
 wire \pmod_1414.RX.tickgen.Acc[4] ;
 wire \pmod_1414.RX.tickgen.Acc[5] ;
 wire \pmod_1414.RX.tickgen.Acc[6] ;
 wire \pmod_1414.RX.tickgen.Acc[7] ;
 wire \pmod_1414.RX.tickgen.Acc[8] ;
 wire \pmod_1414.RX.tickgen.Acc[9] ;
 wire \pmod_1414.mem_strorage.i_w_caret_strobe ;
 wire \pmod_1414.mem_strorage.mem[0][0] ;
 wire \pmod_1414.mem_strorage.mem[0][1] ;
 wire \pmod_1414.mem_strorage.mem[0][2] ;
 wire \pmod_1414.mem_strorage.mem[0][3] ;
 wire \pmod_1414.mem_strorage.mem[0][4] ;
 wire \pmod_1414.mem_strorage.mem[0][5] ;
 wire \pmod_1414.mem_strorage.mem[0][6] ;
 wire \pmod_1414.mem_strorage.mem[10][0] ;
 wire \pmod_1414.mem_strorage.mem[10][1] ;
 wire \pmod_1414.mem_strorage.mem[10][2] ;
 wire \pmod_1414.mem_strorage.mem[10][3] ;
 wire \pmod_1414.mem_strorage.mem[10][4] ;
 wire \pmod_1414.mem_strorage.mem[10][5] ;
 wire \pmod_1414.mem_strorage.mem[10][6] ;
 wire \pmod_1414.mem_strorage.mem[11][0] ;
 wire \pmod_1414.mem_strorage.mem[11][1] ;
 wire \pmod_1414.mem_strorage.mem[11][2] ;
 wire \pmod_1414.mem_strorage.mem[11][3] ;
 wire \pmod_1414.mem_strorage.mem[11][4] ;
 wire \pmod_1414.mem_strorage.mem[11][5] ;
 wire \pmod_1414.mem_strorage.mem[11][6] ;
 wire \pmod_1414.mem_strorage.mem[12][0] ;
 wire \pmod_1414.mem_strorage.mem[12][1] ;
 wire \pmod_1414.mem_strorage.mem[12][2] ;
 wire \pmod_1414.mem_strorage.mem[12][3] ;
 wire \pmod_1414.mem_strorage.mem[12][4] ;
 wire \pmod_1414.mem_strorage.mem[12][5] ;
 wire \pmod_1414.mem_strorage.mem[12][6] ;
 wire \pmod_1414.mem_strorage.mem[13][0] ;
 wire \pmod_1414.mem_strorage.mem[13][1] ;
 wire \pmod_1414.mem_strorage.mem[13][2] ;
 wire \pmod_1414.mem_strorage.mem[13][3] ;
 wire \pmod_1414.mem_strorage.mem[13][4] ;
 wire \pmod_1414.mem_strorage.mem[13][5] ;
 wire \pmod_1414.mem_strorage.mem[13][6] ;
 wire \pmod_1414.mem_strorage.mem[14][0] ;
 wire \pmod_1414.mem_strorage.mem[14][1] ;
 wire \pmod_1414.mem_strorage.mem[14][2] ;
 wire \pmod_1414.mem_strorage.mem[14][3] ;
 wire \pmod_1414.mem_strorage.mem[14][4] ;
 wire \pmod_1414.mem_strorage.mem[14][5] ;
 wire \pmod_1414.mem_strorage.mem[14][6] ;
 wire \pmod_1414.mem_strorage.mem[15][0] ;
 wire \pmod_1414.mem_strorage.mem[15][1] ;
 wire \pmod_1414.mem_strorage.mem[15][2] ;
 wire \pmod_1414.mem_strorage.mem[15][3] ;
 wire \pmod_1414.mem_strorage.mem[15][4] ;
 wire \pmod_1414.mem_strorage.mem[15][5] ;
 wire \pmod_1414.mem_strorage.mem[15][6] ;
 wire \pmod_1414.mem_strorage.mem[1][0] ;
 wire \pmod_1414.mem_strorage.mem[1][1] ;
 wire \pmod_1414.mem_strorage.mem[1][2] ;
 wire \pmod_1414.mem_strorage.mem[1][3] ;
 wire \pmod_1414.mem_strorage.mem[1][4] ;
 wire \pmod_1414.mem_strorage.mem[1][5] ;
 wire \pmod_1414.mem_strorage.mem[1][6] ;
 wire \pmod_1414.mem_strorage.mem[2][0] ;
 wire \pmod_1414.mem_strorage.mem[2][1] ;
 wire \pmod_1414.mem_strorage.mem[2][2] ;
 wire \pmod_1414.mem_strorage.mem[2][3] ;
 wire \pmod_1414.mem_strorage.mem[2][4] ;
 wire \pmod_1414.mem_strorage.mem[2][5] ;
 wire \pmod_1414.mem_strorage.mem[2][6] ;
 wire \pmod_1414.mem_strorage.mem[3][0] ;
 wire \pmod_1414.mem_strorage.mem[3][1] ;
 wire \pmod_1414.mem_strorage.mem[3][2] ;
 wire \pmod_1414.mem_strorage.mem[3][3] ;
 wire \pmod_1414.mem_strorage.mem[3][4] ;
 wire \pmod_1414.mem_strorage.mem[3][5] ;
 wire \pmod_1414.mem_strorage.mem[3][6] ;
 wire \pmod_1414.mem_strorage.mem[4][0] ;
 wire \pmod_1414.mem_strorage.mem[4][1] ;
 wire \pmod_1414.mem_strorage.mem[4][2] ;
 wire \pmod_1414.mem_strorage.mem[4][3] ;
 wire \pmod_1414.mem_strorage.mem[4][4] ;
 wire \pmod_1414.mem_strorage.mem[4][5] ;
 wire \pmod_1414.mem_strorage.mem[4][6] ;
 wire \pmod_1414.mem_strorage.mem[5][0] ;
 wire \pmod_1414.mem_strorage.mem[5][1] ;
 wire \pmod_1414.mem_strorage.mem[5][2] ;
 wire \pmod_1414.mem_strorage.mem[5][3] ;
 wire \pmod_1414.mem_strorage.mem[5][4] ;
 wire \pmod_1414.mem_strorage.mem[5][5] ;
 wire \pmod_1414.mem_strorage.mem[5][6] ;
 wire \pmod_1414.mem_strorage.mem[6][0] ;
 wire \pmod_1414.mem_strorage.mem[6][1] ;
 wire \pmod_1414.mem_strorage.mem[6][2] ;
 wire \pmod_1414.mem_strorage.mem[6][3] ;
 wire \pmod_1414.mem_strorage.mem[6][4] ;
 wire \pmod_1414.mem_strorage.mem[6][5] ;
 wire \pmod_1414.mem_strorage.mem[6][6] ;
 wire \pmod_1414.mem_strorage.mem[7][0] ;
 wire \pmod_1414.mem_strorage.mem[7][1] ;
 wire \pmod_1414.mem_strorage.mem[7][2] ;
 wire \pmod_1414.mem_strorage.mem[7][3] ;
 wire \pmod_1414.mem_strorage.mem[7][4] ;
 wire \pmod_1414.mem_strorage.mem[7][5] ;
 wire \pmod_1414.mem_strorage.mem[7][6] ;
 wire \pmod_1414.mem_strorage.mem[8][0] ;
 wire \pmod_1414.mem_strorage.mem[8][1] ;
 wire \pmod_1414.mem_strorage.mem[8][2] ;
 wire \pmod_1414.mem_strorage.mem[8][3] ;
 wire \pmod_1414.mem_strorage.mem[8][4] ;
 wire \pmod_1414.mem_strorage.mem[8][5] ;
 wire \pmod_1414.mem_strorage.mem[8][6] ;
 wire \pmod_1414.mem_strorage.mem[9][0] ;
 wire \pmod_1414.mem_strorage.mem[9][1] ;
 wire \pmod_1414.mem_strorage.mem[9][2] ;
 wire \pmod_1414.mem_strorage.mem[9][3] ;
 wire \pmod_1414.mem_strorage.mem[9][4] ;
 wire \pmod_1414.mem_strorage.mem[9][5] ;
 wire \pmod_1414.mem_strorage.mem[9][6] ;
 wire \pmod_1414.mem_strorage.r_shift_enable ;
 wire \pmod_1414.r_address_counter[0] ;
 wire \pmod_1414.r_address_counter[1] ;
 wire \pmod_1414.r_address_counter[2] ;
 wire \pmod_1414.r_address_counter[3] ;
 wire \pmod_1414.r_counter[0] ;
 wire \pmod_1414.r_counter[10] ;
 wire \pmod_1414.r_counter[11] ;
 wire \pmod_1414.r_counter[12] ;
 wire \pmod_1414.r_counter[13] ;
 wire \pmod_1414.r_counter[14] ;
 wire \pmod_1414.r_counter[15] ;
 wire \pmod_1414.r_counter[16] ;
 wire \pmod_1414.r_counter[17] ;
 wire \pmod_1414.r_counter[18] ;
 wire \pmod_1414.r_counter[19] ;
 wire \pmod_1414.r_counter[1] ;
 wire \pmod_1414.r_counter[20] ;
 wire \pmod_1414.r_counter[21] ;
 wire \pmod_1414.r_counter[2] ;
 wire \pmod_1414.r_counter[3] ;
 wire \pmod_1414.r_counter[4] ;
 wire \pmod_1414.r_counter[5] ;
 wire \pmod_1414.r_counter[6] ;
 wire \pmod_1414.r_counter[7] ;
 wire \pmod_1414.r_counter[8] ;
 wire \pmod_1414.r_counter[9] ;
 wire \pmod_1414.r_uart_rx_counter[0] ;
 wire \pmod_1414.r_uart_rx_counter[1] ;
 wire \pmod_1414.r_uart_rx_counter[2] ;
 wire \pmod_1414.r_uart_rx_counter[3] ;
 wire net4;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire clknet_0_clk;
 wire net5;
 wire net6;
 wire net7;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;

 sg13g2_inv_1 _1025_ (.Y(_0219_),
    .A(\pmod_1414.r_uart_rx_counter[3] ));
 sg13g2_inv_1 _1026_ (.Y(_0220_),
    .A(\pmod_1414.r_uart_rx_counter[2] ));
 sg13g2_inv_2 _1027_ (.Y(_0221_),
    .A(net231));
 sg13g2_inv_1 _1028_ (.Y(_0222_),
    .A(net226));
 sg13g2_inv_1 _1029_ (.Y(_0223_),
    .A(net502));
 sg13g2_inv_1 _1030_ (.Y(_0224_),
    .A(net536));
 sg13g2_inv_1 _1031_ (.Y(_0225_),
    .A(net508));
 sg13g2_inv_1 _1032_ (.Y(_0226_),
    .A(\pmod_1414.RX.RxD_state[3] ));
 sg13g2_inv_1 _1033_ (.Y(_0227_),
    .A(net302));
 sg13g2_inv_1 _1034_ (.Y(_0228_),
    .A(net413));
 sg13g2_inv_1 _1035_ (.Y(_0229_),
    .A(net481));
 sg13g2_inv_1 _1036_ (.Y(_0230_),
    .A(\pmod_1414.mem_strorage.mem[13][3] ));
 sg13g2_inv_1 _1037_ (.Y(_0231_),
    .A(net459));
 sg13g2_inv_1 _1038_ (.Y(_0232_),
    .A(net390));
 sg13g2_inv_1 _1039_ (.Y(_0233_),
    .A(net471));
 sg13g2_inv_1 _1040_ (.Y(_0234_),
    .A(net431));
 sg13g2_inv_1 _1041_ (.Y(_0235_),
    .A(\pmod_1414.mem_strorage.mem[14][5] ));
 sg13g2_inv_1 _1042_ (.Y(_0236_),
    .A(\pmod_1414.mem_strorage.mem[15][0] ));
 sg13g2_inv_1 _1043_ (.Y(_0237_),
    .A(net475));
 sg13g2_inv_1 _1044_ (.Y(_0238_),
    .A(net511));
 sg13g2_inv_1 _1045_ (.Y(_0239_),
    .A(\pmod_1414.mem_strorage.mem[15][4] ));
 sg13g2_inv_1 _1046_ (.Y(_0240_),
    .A(\pmod_1414.mem_strorage.mem[15][5] ));
 sg13g2_inv_1 _1047_ (.Y(_0241_),
    .A(net204));
 sg13g2_inv_1 _1048_ (.Y(_0242_),
    .A(net322));
 sg13g2_inv_1 _1049_ (.Y(_0243_),
    .A(net549));
 sg13g2_inv_1 _1050_ (.Y(_0244_),
    .A(net300));
 sg13g2_inv_1 _1051_ (.Y(_0245_),
    .A(net521));
 sg13g2_inv_1 _1052_ (.Y(_0246_),
    .A(net524));
 sg13g2_inv_1 _1053_ (.Y(_0247_),
    .A(net529));
 sg13g2_inv_1 _1054_ (.Y(_0248_),
    .A(net296));
 sg13g2_nand2_2 _1055_ (.Y(_0249_),
    .A(\pmod_1414.r_uart_rx_counter[1] ),
    .B(\pmod_1414.r_uart_rx_counter[0] ));
 sg13g2_nand4_1 _1056_ (.B(\pmod_1414.r_uart_rx_counter[2] ),
    .C(net231),
    .A(\pmod_1414.r_uart_rx_counter[3] ),
    .Y(_0250_),
    .D(net232));
 sg13g2_inv_1 _1057_ (.Y(_0251_),
    .A(_0250_));
 sg13g2_nor4_2 _1058_ (.A(net218),
    .B(net221),
    .C(\pmod_1414.GPout[7] ),
    .Y(_0252_),
    .D(net216));
 sg13g2_nor2_1 _1059_ (.A(net228),
    .B(net224),
    .Y(_0253_));
 sg13g2_nand4_1 _1060_ (.B(net222),
    .C(_0252_),
    .A(_0222_),
    .Y(_0254_),
    .D(_0253_));
 sg13g2_nand2_1 _1061_ (.Y(_0255_),
    .A(_0250_),
    .B(net202));
 sg13g2_xor2_1 _1062_ (.B(_0255_),
    .A(_0010_),
    .X(_0256_));
 sg13g2_nor2_1 _1063_ (.A(net231),
    .B(net232),
    .Y(_0257_));
 sg13g2_o21ai_1 _1064_ (.B1(_0249_),
    .Y(_0258_),
    .A1(_0254_),
    .A2(_0257_));
 sg13g2_nand2b_1 _1065_ (.Y(_0259_),
    .B(_0258_),
    .A_N(_0256_));
 sg13g2_nor2_1 _1066_ (.A(\pmod_1414.r_uart_rx_counter[3] ),
    .B(\pmod_1414.r_uart_rx_counter[2] ),
    .Y(_0260_));
 sg13g2_a21oi_1 _1067_ (.A1(_0257_),
    .A2(_0260_),
    .Y(_0261_),
    .B1(_0254_));
 sg13g2_nand2_1 _1068_ (.Y(_0262_),
    .A(_0010_),
    .B(_0261_));
 sg13g2_mux2_1 _1069_ (.A0(_0255_),
    .A1(_0262_),
    .S(_0259_),
    .X(_0263_));
 sg13g2_xnor2_1 _1070_ (.Y(_0169_),
    .A(\pmod_1414.r_uart_rx_counter[3] ),
    .B(_0263_));
 sg13g2_nand2b_1 _1071_ (.Y(_0264_),
    .B(_0255_),
    .A_N(_0261_));
 sg13g2_nand2b_1 _1072_ (.Y(_0265_),
    .B(_0256_),
    .A_N(_0258_));
 sg13g2_nand3_1 _1073_ (.B(_0264_),
    .C(_0265_),
    .A(_0259_),
    .Y(_0266_));
 sg13g2_o21ai_1 _1074_ (.B1(_0266_),
    .Y(_0168_),
    .A1(_0221_),
    .A2(_0264_));
 sg13g2_nand2_1 _1075_ (.Y(_0267_),
    .A(_0054_),
    .B(_0264_));
 sg13g2_mux2_1 _1076_ (.A0(net202),
    .A1(_0255_),
    .S(net231),
    .X(_0268_));
 sg13g2_xnor2_1 _1077_ (.Y(_0167_),
    .A(_0267_),
    .B(_0268_));
 sg13g2_o21ai_1 _1078_ (.B1(_0267_),
    .Y(_0166_),
    .A1(_0221_),
    .A2(_0264_));
 sg13g2_nand3_1 _1079_ (.B(net543),
    .C(\pmod_1414.RX.OversamplingCnt[0] ),
    .A(net234),
    .Y(_0269_));
 sg13g2_or2_1 _1080_ (.X(_0270_),
    .B(_0269_),
    .A(_0227_));
 sg13g2_or2_1 _1081_ (.X(_0271_),
    .B(_0270_),
    .A(net308));
 sg13g2_nor2_1 _1082_ (.A(\pmod_1414.RX.RxD_state[3] ),
    .B(\pmod_1414.RX.RxD_state[2] ),
    .Y(_0272_));
 sg13g2_nand4_1 _1083_ (.B(net508),
    .C(\pmod_1414.RX.RxD_bit ),
    .A(_0224_),
    .Y(_0273_),
    .D(_0272_));
 sg13g2_nor2_1 _1084_ (.A(_0271_),
    .B(net509),
    .Y(_0000_));
 sg13g2_nor2b_2 _1085_ (.A(\pmod_1414.r_address_counter[2] ),
    .B_N(\pmod_1414.r_address_counter[3] ),
    .Y(_0274_));
 sg13g2_mux4_1 _1086_ (.S0(net210),
    .A0(\pmod_1414.mem_strorage.mem[8][0] ),
    .A1(\pmod_1414.mem_strorage.mem[9][0] ),
    .A2(\pmod_1414.mem_strorage.mem[10][0] ),
    .A3(\pmod_1414.mem_strorage.mem[11][0] ),
    .S1(net205),
    .X(_0275_));
 sg13g2_nand2b_1 _1087_ (.Y(_0276_),
    .B(\pmod_1414.r_uart_rx_counter[2] ),
    .A_N(\pmod_1414.r_address_counter[2] ));
 sg13g2_a22oi_1 _1088_ (.Y(_0277_),
    .B1(_0241_),
    .B2(net231),
    .A2(\pmod_1414.r_address_counter[2] ),
    .A1(_0220_));
 sg13g2_xnor2_1 _1089_ (.Y(_0278_),
    .A(net232),
    .B(net209));
 sg13g2_o21ai_1 _1090_ (.B1(_0009_),
    .Y(_0279_),
    .A1(_0219_),
    .A2(\pmod_1414.r_address_counter[3] ));
 sg13g2_a221oi_1 _1091_ (.B2(_0219_),
    .C1(_0279_),
    .B1(\pmod_1414.r_address_counter[3] ),
    .A1(_0221_),
    .Y(_0280_),
    .A2(net204));
 sg13g2_and4_2 _1092_ (.A(_0276_),
    .B(_0277_),
    .C(_0278_),
    .D(_0280_),
    .X(_0281_));
 sg13g2_a21oi_1 _1093_ (.A1(_0274_),
    .A2(_0275_),
    .Y(_0282_),
    .B1(_0281_));
 sg13g2_and2_2 _1094_ (.A(\pmod_1414.r_address_counter[2] ),
    .B(\pmod_1414.r_address_counter[3] ),
    .X(_0283_));
 sg13g2_mux4_1 _1095_ (.S0(net208),
    .A0(\pmod_1414.mem_strorage.mem[12][0] ),
    .A1(\pmod_1414.mem_strorage.mem[13][0] ),
    .A2(\pmod_1414.mem_strorage.mem[14][0] ),
    .A3(\pmod_1414.mem_strorage.mem[15][0] ),
    .S1(net203),
    .X(_0284_));
 sg13g2_nor2_2 _1096_ (.A(\pmod_1414.r_address_counter[2] ),
    .B(\pmod_1414.r_address_counter[3] ),
    .Y(_0285_));
 sg13g2_mux4_1 _1097_ (.S0(net213),
    .A0(\pmod_1414.mem_strorage.mem[0][0] ),
    .A1(\pmod_1414.mem_strorage.mem[1][0] ),
    .A2(\pmod_1414.mem_strorage.mem[2][0] ),
    .A3(\pmod_1414.mem_strorage.mem[3][0] ),
    .S1(net207),
    .X(_0286_));
 sg13g2_nor2b_1 _1098_ (.A(net211),
    .B_N(\pmod_1414.mem_strorage.mem[6][0] ),
    .Y(_0287_));
 sg13g2_a21oi_1 _1099_ (.A1(net211),
    .A2(\pmod_1414.mem_strorage.mem[7][0] ),
    .Y(_0288_),
    .B1(_0287_));
 sg13g2_nand2b_1 _1100_ (.Y(_0289_),
    .B(\pmod_1414.mem_strorage.mem[4][0] ),
    .A_N(net213));
 sg13g2_a21oi_1 _1101_ (.A1(net211),
    .A2(\pmod_1414.mem_strorage.mem[5][0] ),
    .Y(_0290_),
    .B1(net206));
 sg13g2_nor2b_2 _1102_ (.A(\pmod_1414.r_address_counter[3] ),
    .B_N(\pmod_1414.r_address_counter[2] ),
    .Y(_0291_));
 sg13g2_nand2b_1 _1103_ (.Y(_0292_),
    .B(\pmod_1414.r_address_counter[2] ),
    .A_N(\pmod_1414.r_address_counter[3] ));
 sg13g2_a221oi_1 _1104_ (.B2(_0290_),
    .C1(_0292_),
    .B1(_0289_),
    .A1(net206),
    .Y(_0293_),
    .A2(_0288_));
 sg13g2_a221oi_1 _1105_ (.B2(_0286_),
    .C1(_0293_),
    .B1(_0285_),
    .A1(_0283_),
    .Y(_0294_),
    .A2(_0284_));
 sg13g2_nand2_1 _1106_ (.Y(_0001_),
    .A(_0282_),
    .B(_0294_));
 sg13g2_mux4_1 _1107_ (.S0(net209),
    .A0(\pmod_1414.mem_strorage.mem[12][1] ),
    .A1(\pmod_1414.mem_strorage.mem[13][1] ),
    .A2(\pmod_1414.mem_strorage.mem[14][1] ),
    .A3(\pmod_1414.mem_strorage.mem[15][1] ),
    .S1(net204),
    .X(_0295_));
 sg13g2_a21oi_1 _1108_ (.A1(_0283_),
    .A2(_0295_),
    .Y(_0296_),
    .B1(_0281_));
 sg13g2_mux2_1 _1109_ (.A0(\pmod_1414.mem_strorage.mem[8][1] ),
    .A1(\pmod_1414.mem_strorage.mem[9][1] ),
    .S(net210),
    .X(_0297_));
 sg13g2_nor2b_1 _1110_ (.A(net210),
    .B_N(\pmod_1414.mem_strorage.mem[10][1] ),
    .Y(_0298_));
 sg13g2_a21oi_1 _1111_ (.A1(net210),
    .A2(\pmod_1414.mem_strorage.mem[11][1] ),
    .Y(_0299_),
    .B1(_0298_));
 sg13g2_o21ai_1 _1112_ (.B1(_0274_),
    .Y(_0300_),
    .A1(net205),
    .A2(_0297_));
 sg13g2_a21oi_1 _1113_ (.A1(net204),
    .A2(_0299_),
    .Y(_0301_),
    .B1(_0300_));
 sg13g2_mux4_1 _1114_ (.S0(net214),
    .A0(\pmod_1414.mem_strorage.mem[0][1] ),
    .A1(\pmod_1414.mem_strorage.mem[1][1] ),
    .A2(\pmod_1414.mem_strorage.mem[2][1] ),
    .A3(\pmod_1414.mem_strorage.mem[3][1] ),
    .S1(net207),
    .X(_0302_));
 sg13g2_mux4_1 _1115_ (.S0(net206),
    .A0(\pmod_1414.mem_strorage.mem[4][1] ),
    .A1(\pmod_1414.mem_strorage.mem[6][1] ),
    .A2(\pmod_1414.mem_strorage.mem[5][1] ),
    .A3(\pmod_1414.mem_strorage.mem[7][1] ),
    .S1(net213),
    .X(_0303_));
 sg13g2_a221oi_1 _1116_ (.B2(_0291_),
    .C1(_0301_),
    .B1(_0303_),
    .A1(_0285_),
    .Y(_0304_),
    .A2(_0302_));
 sg13g2_nand2_1 _1117_ (.Y(_0002_),
    .A(_0296_),
    .B(_0304_));
 sg13g2_nand2b_1 _1118_ (.Y(_0305_),
    .B(\pmod_1414.mem_strorage.mem[4][2] ),
    .A_N(net213));
 sg13g2_a21oi_1 _1119_ (.A1(net211),
    .A2(\pmod_1414.mem_strorage.mem[5][2] ),
    .Y(_0306_),
    .B1(net206));
 sg13g2_nor2b_1 _1120_ (.A(net211),
    .B_N(\pmod_1414.mem_strorage.mem[6][2] ),
    .Y(_0307_));
 sg13g2_a21oi_1 _1121_ (.A1(net211),
    .A2(\pmod_1414.mem_strorage.mem[7][2] ),
    .Y(_0308_),
    .B1(_0307_));
 sg13g2_a221oi_1 _1122_ (.B2(net206),
    .C1(_0292_),
    .B1(_0308_),
    .A1(_0305_),
    .Y(_0309_),
    .A2(_0306_));
 sg13g2_mux4_1 _1123_ (.S0(net213),
    .A0(\pmod_1414.mem_strorage.mem[0][2] ),
    .A1(\pmod_1414.mem_strorage.mem[1][2] ),
    .A2(\pmod_1414.mem_strorage.mem[2][2] ),
    .A3(\pmod_1414.mem_strorage.mem[3][2] ),
    .S1(net207),
    .X(_0310_));
 sg13g2_mux4_1 _1124_ (.S0(net208),
    .A0(\pmod_1414.mem_strorage.mem[12][2] ),
    .A1(\pmod_1414.mem_strorage.mem[13][2] ),
    .A2(\pmod_1414.mem_strorage.mem[14][2] ),
    .A3(\pmod_1414.mem_strorage.mem[15][2] ),
    .S1(net203),
    .X(_0311_));
 sg13g2_mux4_1 _1125_ (.S0(net209),
    .A0(\pmod_1414.mem_strorage.mem[8][2] ),
    .A1(\pmod_1414.mem_strorage.mem[9][2] ),
    .A2(\pmod_1414.mem_strorage.mem[10][2] ),
    .A3(\pmod_1414.mem_strorage.mem[11][2] ),
    .S1(net204),
    .X(_0312_));
 sg13g2_a221oi_1 _1126_ (.B2(_0283_),
    .C1(_0309_),
    .B1(_0311_),
    .A1(_0285_),
    .Y(_0313_),
    .A2(_0310_));
 sg13g2_a21oi_1 _1127_ (.A1(_0274_),
    .A2(_0312_),
    .Y(_0314_),
    .B1(_0281_));
 sg13g2_nand2_1 _1128_ (.Y(_0003_),
    .A(_0313_),
    .B(_0314_));
 sg13g2_mux4_1 _1129_ (.S0(net209),
    .A0(\pmod_1414.mem_strorage.mem[8][3] ),
    .A1(\pmod_1414.mem_strorage.mem[9][3] ),
    .A2(\pmod_1414.mem_strorage.mem[10][3] ),
    .A3(\pmod_1414.mem_strorage.mem[11][3] ),
    .S1(net205),
    .X(_0315_));
 sg13g2_a21oi_1 _1130_ (.A1(_0274_),
    .A2(_0315_),
    .Y(_0316_),
    .B1(_0281_));
 sg13g2_nor2b_1 _1131_ (.A(net213),
    .B_N(\pmod_1414.mem_strorage.mem[2][3] ),
    .Y(_0317_));
 sg13g2_a21oi_1 _1132_ (.A1(net214),
    .A2(\pmod_1414.mem_strorage.mem[3][3] ),
    .Y(_0318_),
    .B1(_0317_));
 sg13g2_mux2_1 _1133_ (.A0(\pmod_1414.mem_strorage.mem[0][3] ),
    .A1(\pmod_1414.mem_strorage.mem[1][3] ),
    .S(net214),
    .X(_0319_));
 sg13g2_o21ai_1 _1134_ (.B1(_0285_),
    .Y(_0320_),
    .A1(net207),
    .A2(_0319_));
 sg13g2_a21oi_2 _1135_ (.B1(_0320_),
    .Y(_0321_),
    .A2(_0318_),
    .A1(net207));
 sg13g2_mux4_1 _1136_ (.S0(net208),
    .A0(\pmod_1414.mem_strorage.mem[12][3] ),
    .A1(\pmod_1414.mem_strorage.mem[13][3] ),
    .A2(\pmod_1414.mem_strorage.mem[14][3] ),
    .A3(\pmod_1414.mem_strorage.mem[15][3] ),
    .S1(net203),
    .X(_0322_));
 sg13g2_mux4_1 _1137_ (.S0(net206),
    .A0(\pmod_1414.mem_strorage.mem[4][3] ),
    .A1(\pmod_1414.mem_strorage.mem[6][3] ),
    .A2(\pmod_1414.mem_strorage.mem[5][3] ),
    .A3(\pmod_1414.mem_strorage.mem[7][3] ),
    .S1(net211),
    .X(_0323_));
 sg13g2_a221oi_1 _1138_ (.B2(_0291_),
    .C1(_0321_),
    .B1(_0323_),
    .A1(_0283_),
    .Y(_0324_),
    .A2(_0322_));
 sg13g2_nand2_1 _1139_ (.Y(_0004_),
    .A(_0316_),
    .B(_0324_));
 sg13g2_mux2_1 _1140_ (.A0(\pmod_1414.mem_strorage.mem[4][4] ),
    .A1(net556),
    .S(net213),
    .X(_0325_));
 sg13g2_nor2b_1 _1141_ (.A(net212),
    .B_N(\pmod_1414.mem_strorage.mem[6][4] ),
    .Y(_0326_));
 sg13g2_a21oi_1 _1142_ (.A1(net212),
    .A2(\pmod_1414.mem_strorage.mem[7][4] ),
    .Y(_0327_),
    .B1(_0326_));
 sg13g2_a21oi_1 _1143_ (.A1(net204),
    .A2(_0327_),
    .Y(_0328_),
    .B1(_0292_));
 sg13g2_o21ai_1 _1144_ (.B1(_0328_),
    .Y(_0329_),
    .A1(net204),
    .A2(_0325_));
 sg13g2_mux4_1 _1145_ (.S0(net208),
    .A0(\pmod_1414.mem_strorage.mem[12][4] ),
    .A1(\pmod_1414.mem_strorage.mem[13][4] ),
    .A2(\pmod_1414.mem_strorage.mem[14][4] ),
    .A3(\pmod_1414.mem_strorage.mem[15][4] ),
    .S1(net203),
    .X(_0330_));
 sg13g2_mux4_1 _1146_ (.S0(net208),
    .A0(\pmod_1414.mem_strorage.mem[8][4] ),
    .A1(\pmod_1414.mem_strorage.mem[9][4] ),
    .A2(\pmod_1414.mem_strorage.mem[10][4] ),
    .A3(\pmod_1414.mem_strorage.mem[11][4] ),
    .S1(net203),
    .X(_0331_));
 sg13g2_mux4_1 _1147_ (.S0(net214),
    .A0(\pmod_1414.mem_strorage.mem[0][4] ),
    .A1(\pmod_1414.mem_strorage.mem[1][4] ),
    .A2(\pmod_1414.mem_strorage.mem[2][4] ),
    .A3(\pmod_1414.mem_strorage.mem[3][4] ),
    .S1(net207),
    .X(_0332_));
 sg13g2_a22oi_1 _1148_ (.Y(_0333_),
    .B1(_0331_),
    .B2(_0274_),
    .A2(_0330_),
    .A1(_0283_));
 sg13g2_a21oi_1 _1149_ (.A1(_0285_),
    .A2(_0332_),
    .Y(_0334_),
    .B1(_0281_));
 sg13g2_nand3_1 _1150_ (.B(_0333_),
    .C(_0334_),
    .A(_0329_),
    .Y(_0005_));
 sg13g2_mux4_1 _1151_ (.S0(net209),
    .A0(\pmod_1414.mem_strorage.mem[8][5] ),
    .A1(\pmod_1414.mem_strorage.mem[9][5] ),
    .A2(\pmod_1414.mem_strorage.mem[10][5] ),
    .A3(\pmod_1414.mem_strorage.mem[11][5] ),
    .S1(net205),
    .X(_0335_));
 sg13g2_mux4_1 _1152_ (.S0(net215),
    .A0(\pmod_1414.mem_strorage.mem[0][5] ),
    .A1(\pmod_1414.mem_strorage.mem[1][5] ),
    .A2(\pmod_1414.mem_strorage.mem[2][5] ),
    .A3(\pmod_1414.mem_strorage.mem[3][5] ),
    .S1(net207),
    .X(_0336_));
 sg13g2_a22oi_1 _1153_ (.Y(_0337_),
    .B1(_0336_),
    .B2(_0285_),
    .A2(_0335_),
    .A1(_0274_));
 sg13g2_mux4_1 _1154_ (.S0(net208),
    .A0(\pmod_1414.mem_strorage.mem[12][5] ),
    .A1(\pmod_1414.mem_strorage.mem[13][5] ),
    .A2(\pmod_1414.mem_strorage.mem[14][5] ),
    .A3(\pmod_1414.mem_strorage.mem[15][5] ),
    .S1(net203),
    .X(_0338_));
 sg13g2_mux4_1 _1155_ (.S0(net206),
    .A0(\pmod_1414.mem_strorage.mem[4][5] ),
    .A1(\pmod_1414.mem_strorage.mem[6][5] ),
    .A2(\pmod_1414.mem_strorage.mem[5][5] ),
    .A3(\pmod_1414.mem_strorage.mem[7][5] ),
    .S1(net212),
    .X(_0339_));
 sg13g2_a22oi_1 _1156_ (.Y(_0340_),
    .B1(_0339_),
    .B2(_0291_),
    .A2(_0338_),
    .A1(_0283_));
 sg13g2_a21oi_1 _1157_ (.A1(_0337_),
    .A2(_0340_),
    .Y(_0006_),
    .B1(_0281_));
 sg13g2_mux4_1 _1158_ (.S0(net206),
    .A0(\pmod_1414.mem_strorage.mem[4][6] ),
    .A1(\pmod_1414.mem_strorage.mem[6][6] ),
    .A2(\pmod_1414.mem_strorage.mem[5][6] ),
    .A3(\pmod_1414.mem_strorage.mem[7][6] ),
    .S1(net211),
    .X(_0341_));
 sg13g2_mux4_1 _1159_ (.S0(net209),
    .A0(\pmod_1414.mem_strorage.mem[8][6] ),
    .A1(\pmod_1414.mem_strorage.mem[9][6] ),
    .A2(\pmod_1414.mem_strorage.mem[10][6] ),
    .A3(\pmod_1414.mem_strorage.mem[11][6] ),
    .S1(net203),
    .X(_0342_));
 sg13g2_mux4_1 _1160_ (.S0(net208),
    .A0(\pmod_1414.mem_strorage.mem[12][6] ),
    .A1(\pmod_1414.mem_strorage.mem[13][6] ),
    .A2(\pmod_1414.mem_strorage.mem[14][6] ),
    .A3(\pmod_1414.mem_strorage.mem[15][6] ),
    .S1(net203),
    .X(_0343_));
 sg13g2_a22oi_1 _1161_ (.Y(_0344_),
    .B1(_0343_),
    .B2(_0283_),
    .A2(_0342_),
    .A1(_0274_));
 sg13g2_mux4_1 _1162_ (.S0(net213),
    .A0(\pmod_1414.mem_strorage.mem[0][6] ),
    .A1(\pmod_1414.mem_strorage.mem[1][6] ),
    .A2(\pmod_1414.mem_strorage.mem[2][6] ),
    .A3(\pmod_1414.mem_strorage.mem[3][6] ),
    .S1(\pmod_1414.r_address_counter[1] ),
    .X(_0345_));
 sg13g2_a221oi_1 _1163_ (.B2(_0285_),
    .C1(_0281_),
    .B1(_0345_),
    .A1(_0291_),
    .Y(_0346_),
    .A2(_0341_));
 sg13g2_nand2_1 _1164_ (.Y(_0007_),
    .A(_0344_),
    .B(_0346_));
 sg13g2_nand2b_1 _1165_ (.Y(\pmod_1414.HPDL_WR4 ),
    .B(_0283_),
    .A_N(net233));
 sg13g2_nand2b_1 _1166_ (.Y(\pmod_1414.HPDL_WR3 ),
    .B(_0274_),
    .A_N(net233));
 sg13g2_nand2b_1 _1167_ (.Y(\pmod_1414.HPDL_WR2 ),
    .B(_0291_),
    .A_N(net233));
 sg13g2_nand2b_1 _1168_ (.Y(\pmod_1414.HPDL_WR1 ),
    .B(_0285_),
    .A_N(net233));
 sg13g2_nand2_1 _1169_ (.Y(_0347_),
    .A(net209),
    .B(net204));
 sg13g2_xor2_1 _1170_ (.B(net205),
    .A(net208),
    .X(_0035_));
 sg13g2_xnor2_1 _1171_ (.Y(_0036_),
    .A(\pmod_1414.r_address_counter[2] ),
    .B(_0347_));
 sg13g2_nor2_1 _1172_ (.A(_0008_),
    .B(_0347_),
    .Y(_0348_));
 sg13g2_xor2_1 _1173_ (.B(_0348_),
    .A(\pmod_1414.r_address_counter[3] ),
    .X(_0037_));
 sg13g2_xor2_1 _1174_ (.B(net455),
    .A(\pmod_1414.r_counter[0] ),
    .X(_0023_));
 sg13g2_nand3_1 _1175_ (.B(net455),
    .C(net546),
    .A(\pmod_1414.r_counter[0] ),
    .Y(_0349_));
 sg13g2_a21o_1 _1176_ (.A2(net455),
    .A1(\pmod_1414.r_counter[0] ),
    .B1(net546),
    .X(_0350_));
 sg13g2_and2_1 _1177_ (.A(_0349_),
    .B(net547),
    .X(_0027_));
 sg13g2_nand4_1 _1178_ (.B(net455),
    .C(net546),
    .A(\pmod_1414.r_counter[0] ),
    .Y(_0351_),
    .D(net341));
 sg13g2_xnor2_1 _1179_ (.Y(_0028_),
    .A(net341),
    .B(_0349_));
 sg13g2_xnor2_1 _1180_ (.Y(_0029_),
    .A(net322),
    .B(_0351_));
 sg13g2_nor3_2 _1181_ (.A(_0242_),
    .B(_0243_),
    .C(_0351_),
    .Y(_0352_));
 sg13g2_o21ai_1 _1182_ (.B1(_0243_),
    .Y(_0353_),
    .A1(_0242_),
    .A2(_0351_));
 sg13g2_nor2b_1 _1183_ (.A(_0352_),
    .B_N(net550),
    .Y(_0030_));
 sg13g2_xor2_1 _1184_ (.B(_0352_),
    .A(net400),
    .X(_0031_));
 sg13g2_nand2_1 _1185_ (.Y(_0354_),
    .A(\pmod_1414.r_counter[6] ),
    .B(net287));
 sg13g2_nor4_2 _1186_ (.A(_0242_),
    .B(_0243_),
    .C(_0351_),
    .Y(_0355_),
    .D(_0354_));
 sg13g2_a21oi_1 _1187_ (.A1(\pmod_1414.r_counter[6] ),
    .A2(_0352_),
    .Y(_0356_),
    .B1(net287));
 sg13g2_nor2_1 _1188_ (.A(_0355_),
    .B(net288),
    .Y(_0032_));
 sg13g2_and2_1 _1189_ (.A(net552),
    .B(_0355_),
    .X(_0357_));
 sg13g2_xor2_1 _1190_ (.B(_0355_),
    .A(net379),
    .X(_0033_));
 sg13g2_xor2_1 _1191_ (.B(_0357_),
    .A(net369),
    .X(_0034_));
 sg13g2_nand4_1 _1192_ (.B(net379),
    .C(net369),
    .A(net233),
    .Y(_0358_),
    .D(_0355_));
 sg13g2_a21o_1 _1193_ (.A2(_0357_),
    .A1(net369),
    .B1(net233),
    .X(_0359_));
 sg13g2_and2_1 _1194_ (.A(_0358_),
    .B(_0359_),
    .X(_0013_));
 sg13g2_nor2_1 _1195_ (.A(_0244_),
    .B(_0358_),
    .Y(_0360_));
 sg13g2_xnor2_1 _1196_ (.Y(_0014_),
    .A(net300),
    .B(_0358_));
 sg13g2_xor2_1 _1197_ (.B(_0360_),
    .A(net433),
    .X(_0015_));
 sg13g2_nand2_1 _1198_ (.Y(_0361_),
    .A(net433),
    .B(net278));
 sg13g2_nor3_2 _1199_ (.A(_0244_),
    .B(_0358_),
    .C(_0361_),
    .Y(_0362_));
 sg13g2_a21oi_1 _1200_ (.A1(\pmod_1414.r_counter[12] ),
    .A2(_0360_),
    .Y(_0363_),
    .B1(net278));
 sg13g2_nor2_1 _1201_ (.A(_0362_),
    .B(net279),
    .Y(_0016_));
 sg13g2_xor2_1 _1202_ (.B(_0362_),
    .A(net409),
    .X(_0017_));
 sg13g2_nand2_1 _1203_ (.Y(_0364_),
    .A(net409),
    .B(net281));
 sg13g2_nor4_2 _1204_ (.A(_0244_),
    .B(_0358_),
    .C(_0361_),
    .Y(_0365_),
    .D(_0364_));
 sg13g2_a21oi_1 _1205_ (.A1(\pmod_1414.r_counter[14] ),
    .A2(_0362_),
    .Y(_0366_),
    .B1(net281));
 sg13g2_nor2_1 _1206_ (.A(_0365_),
    .B(net282),
    .Y(_0018_));
 sg13g2_xor2_1 _1207_ (.B(_0365_),
    .A(net445),
    .X(_0019_));
 sg13g2_and3_1 _1208_ (.X(_0367_),
    .A(\pmod_1414.r_counter[16] ),
    .B(net309),
    .C(_0365_));
 sg13g2_a21oi_1 _1209_ (.A1(\pmod_1414.r_counter[16] ),
    .A2(_0365_),
    .Y(_0368_),
    .B1(net309));
 sg13g2_nor2_1 _1210_ (.A(_0367_),
    .B(net310),
    .Y(_0020_));
 sg13g2_xor2_1 _1211_ (.B(_0367_),
    .A(net418),
    .X(_0021_));
 sg13g2_and2_1 _1212_ (.A(\pmod_1414.r_counter[18] ),
    .B(net284),
    .X(_0369_));
 sg13g2_and4_2 _1213_ (.A(\pmod_1414.r_counter[16] ),
    .B(net309),
    .C(_0365_),
    .D(_0369_),
    .X(_0370_));
 sg13g2_a21oi_1 _1214_ (.A1(\pmod_1414.r_counter[18] ),
    .A2(_0367_),
    .Y(_0371_),
    .B1(net284));
 sg13g2_nor2_1 _1215_ (.A(_0370_),
    .B(net285),
    .Y(_0022_));
 sg13g2_xor2_1 _1216_ (.B(_0370_),
    .A(net377),
    .X(_0024_));
 sg13g2_and3_1 _1217_ (.X(_0372_),
    .A(\pmod_1414.r_counter[20] ),
    .B(net275),
    .C(_0370_));
 sg13g2_a21oi_1 _1218_ (.A1(\pmod_1414.r_counter[20] ),
    .A2(_0370_),
    .Y(_0373_),
    .B1(net275));
 sg13g2_nor2_1 _1219_ (.A(_0372_),
    .B(net276),
    .Y(_0025_));
 sg13g2_xor2_1 _1220_ (.B(_0372_),
    .A(net271),
    .X(_0026_));
 sg13g2_xor2_1 _1221_ (.B(net336),
    .A(\pmod_1414.RX.tickgen.Acc[0] ),
    .X(_0044_));
 sg13g2_nand3_1 _1222_ (.B(net336),
    .C(net540),
    .A(\pmod_1414.RX.tickgen.Acc[0] ),
    .Y(_0374_));
 sg13g2_a21o_1 _1223_ (.A2(net336),
    .A1(\pmod_1414.RX.tickgen.Acc[0] ),
    .B1(net540),
    .X(_0375_));
 sg13g2_and2_1 _1224_ (.A(_0374_),
    .B(net541),
    .X(_0045_));
 sg13g2_nand2_1 _1225_ (.Y(_0376_),
    .A(_0245_),
    .B(_0374_));
 sg13g2_xnor2_1 _1226_ (.Y(_0046_),
    .A(_0245_),
    .B(_0374_));
 sg13g2_a21oi_1 _1227_ (.A1(_0245_),
    .A2(_0374_),
    .Y(_0377_),
    .B1(_0246_));
 sg13g2_nand2_1 _1228_ (.Y(_0378_),
    .A(\pmod_1414.RX.tickgen.Acc[4] ),
    .B(_0376_));
 sg13g2_xnor2_1 _1229_ (.Y(_0047_),
    .A(_0246_),
    .B(_0376_));
 sg13g2_xor2_1 _1230_ (.B(_0377_),
    .A(net262),
    .X(_0048_));
 sg13g2_o21ai_1 _1231_ (.B1(net262),
    .Y(_0379_),
    .A1(\pmod_1414.RX.tickgen.Acc[5] ),
    .A2(_0378_));
 sg13g2_nand2_1 _1232_ (.Y(_0380_),
    .A(\pmod_1414.RX.tickgen.Acc[6] ),
    .B(_0379_));
 sg13g2_xor2_1 _1233_ (.B(_0379_),
    .A(net425),
    .X(_0049_));
 sg13g2_xor2_1 _1234_ (.B(_0380_),
    .A(net386),
    .X(_0050_));
 sg13g2_o21ai_1 _1235_ (.B1(\pmod_1414.RX.tickgen.Acc[6] ),
    .Y(_0381_),
    .A1(\pmod_1414.RX.tickgen.Acc[5] ),
    .A2(_0377_));
 sg13g2_nor2b_1 _1236_ (.A(\pmod_1414.RX.tickgen.Acc[7] ),
    .B_N(_0381_),
    .Y(_0382_));
 sg13g2_nand2_1 _1237_ (.Y(_0383_),
    .A(net267),
    .B(_0382_));
 sg13g2_xnor2_1 _1238_ (.Y(_0051_),
    .A(net267),
    .B(_0382_));
 sg13g2_xnor2_1 _1239_ (.Y(_0052_),
    .A(net320),
    .B(_0383_));
 sg13g2_nor2_1 _1240_ (.A(\pmod_1414.RX.tickgen.Acc[8] ),
    .B(net320),
    .Y(_0384_));
 sg13g2_nand3b_1 _1241_ (.B(_0381_),
    .C(_0384_),
    .Y(_0385_),
    .A_N(\pmod_1414.RX.tickgen.Acc[7] ));
 sg13g2_xor2_1 _1242_ (.B(_0385_),
    .A(net357),
    .X(_0039_));
 sg13g2_nand3_1 _1243_ (.B(net531),
    .C(_0385_),
    .A(net357),
    .Y(_0386_));
 sg13g2_a21o_1 _1244_ (.A2(_0385_),
    .A1(net357),
    .B1(net531),
    .X(_0387_));
 sg13g2_and2_1 _1245_ (.A(_0386_),
    .B(_0387_),
    .X(_0040_));
 sg13g2_xnor2_1 _1246_ (.Y(_0041_),
    .A(_0247_),
    .B(_0386_));
 sg13g2_a21oi_2 _1247_ (.B1(_0248_),
    .Y(_0388_),
    .A2(_0386_),
    .A1(_0247_));
 sg13g2_nand3_1 _1248_ (.B(_0248_),
    .C(_0386_),
    .A(_0247_),
    .Y(_0389_));
 sg13g2_nor2b_1 _1249_ (.A(net297),
    .B_N(net530),
    .Y(_0042_));
 sg13g2_and2_1 _1250_ (.A(net269),
    .B(_0388_),
    .X(_0038_));
 sg13g2_xor2_1 _1251_ (.B(net297),
    .A(net269),
    .X(_0043_));
 sg13g2_mux2_1 _1252_ (.A0(net439),
    .A1(net2),
    .S(net234),
    .X(_0056_));
 sg13g2_mux2_1 _1253_ (.A0(net454),
    .A1(net439),
    .S(net234),
    .X(_0057_));
 sg13g2_and2_1 _1254_ (.A(net235),
    .B(net202),
    .X(_0390_));
 sg13g2_nand3_1 _1255_ (.B(net202),
    .C(_0260_),
    .A(net235),
    .Y(_0391_));
 sg13g2_nand2_2 _1256_ (.Y(_0392_),
    .A(_0221_),
    .B(net232));
 sg13g2_nor2_2 _1257_ (.A(_0391_),
    .B(_0392_),
    .Y(_0393_));
 sg13g2_nand4_1 _1258_ (.B(\pmod_1414.r_uart_rx_counter[2] ),
    .C(net235),
    .A(\pmod_1414.r_uart_rx_counter[3] ),
    .Y(_0394_),
    .D(net202));
 sg13g2_nand3_1 _1259_ (.B(_0251_),
    .C(net202),
    .A(net235),
    .Y(_0395_));
 sg13g2_nor2_2 _1260_ (.A(_0223_),
    .B(_0395_),
    .Y(_0396_));
 sg13g2_or2_1 _1261_ (.X(_0397_),
    .B(_0395_),
    .A(_0223_));
 sg13g2_nor2_2 _1262_ (.A(_0393_),
    .B(net197),
    .Y(_0398_));
 sg13g2_nand2_1 _1263_ (.Y(_0399_),
    .A(net332),
    .B(_0398_));
 sg13g2_a22oi_1 _1264_ (.Y(_0400_),
    .B1(net195),
    .B2(\pmod_1414.mem_strorage.mem[2][0] ),
    .A2(_0393_),
    .A1(net230));
 sg13g2_nand2_1 _1265_ (.Y(_0058_),
    .A(_0399_),
    .B(_0400_));
 sg13g2_nand2_1 _1266_ (.Y(_0401_),
    .A(net328),
    .B(_0398_));
 sg13g2_a22oi_1 _1267_ (.Y(_0402_),
    .B1(net197),
    .B2(\pmod_1414.mem_strorage.mem[2][1] ),
    .A2(_0393_),
    .A1(net227));
 sg13g2_nand2_1 _1268_ (.Y(_0059_),
    .A(_0401_),
    .B(_0402_));
 sg13g2_nand2_1 _1269_ (.Y(_0403_),
    .A(net375),
    .B(_0398_));
 sg13g2_a22oi_1 _1270_ (.Y(_0404_),
    .B1(net196),
    .B2(\pmod_1414.mem_strorage.mem[2][2] ),
    .A2(_0393_),
    .A1(\pmod_1414.GPout[2] ));
 sg13g2_nand2_1 _1271_ (.Y(_0060_),
    .A(_0403_),
    .B(_0404_));
 sg13g2_nand2_1 _1272_ (.Y(_0405_),
    .A(net364),
    .B(_0398_));
 sg13g2_a22oi_1 _1273_ (.Y(_0406_),
    .B1(net198),
    .B2(\pmod_1414.mem_strorage.mem[2][3] ),
    .A2(_0393_),
    .A1(net223));
 sg13g2_nand2_1 _1274_ (.Y(_0061_),
    .A(_0405_),
    .B(_0406_));
 sg13g2_nand2_1 _1275_ (.Y(_0407_),
    .A(net404),
    .B(_0398_));
 sg13g2_a22oi_1 _1276_ (.Y(_0408_),
    .B1(net196),
    .B2(net402),
    .A2(_0393_),
    .A1(\pmod_1414.GPout[4] ));
 sg13g2_nand2_1 _1277_ (.Y(_0062_),
    .A(_0407_),
    .B(_0408_));
 sg13g2_nand2_1 _1278_ (.Y(_0409_),
    .A(net388),
    .B(_0398_));
 sg13g2_a22oi_1 _1279_ (.Y(_0410_),
    .B1(net193),
    .B2(\pmod_1414.mem_strorage.mem[2][5] ),
    .A2(_0393_),
    .A1(net218));
 sg13g2_nand2_1 _1280_ (.Y(_0063_),
    .A(_0409_),
    .B(_0410_));
 sg13g2_nand2_1 _1281_ (.Y(_0411_),
    .A(net392),
    .B(_0398_));
 sg13g2_a22oi_1 _1282_ (.Y(_0412_),
    .B1(net193),
    .B2(\pmod_1414.mem_strorage.mem[2][6] ),
    .A2(_0393_),
    .A1(net216));
 sg13g2_nand2_1 _1283_ (.Y(_0064_),
    .A(_0411_),
    .B(_0412_));
 sg13g2_nand2b_2 _1284_ (.Y(_0413_),
    .B(\pmod_1414.r_uart_rx_counter[1] ),
    .A_N(net232));
 sg13g2_nor2_2 _1285_ (.A(_0391_),
    .B(_0413_),
    .Y(_0414_));
 sg13g2_nor2_2 _1286_ (.A(net196),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_nand2_1 _1287_ (.Y(_0416_),
    .A(net430),
    .B(_0415_));
 sg13g2_a22oi_1 _1288_ (.Y(_0417_),
    .B1(_0414_),
    .B2(net230),
    .A2(net195),
    .A1(net338));
 sg13g2_nand2_1 _1289_ (.Y(_0065_),
    .A(_0416_),
    .B(_0417_));
 sg13g2_nand2_1 _1290_ (.Y(_0418_),
    .A(net417),
    .B(_0415_));
 sg13g2_a22oi_1 _1291_ (.Y(_0419_),
    .B1(_0414_),
    .B2(net227),
    .A2(net197),
    .A1(net351));
 sg13g2_nand2_1 _1292_ (.Y(_0066_),
    .A(_0418_),
    .B(_0419_));
 sg13g2_nand2_1 _1293_ (.Y(_0420_),
    .A(net408),
    .B(_0415_));
 sg13g2_a22oi_1 _1294_ (.Y(_0421_),
    .B1(_0414_),
    .B2(\pmod_1414.GPout[2] ),
    .A2(net196),
    .A1(net326));
 sg13g2_nand2_1 _1295_ (.Y(_0067_),
    .A(_0420_),
    .B(_0421_));
 sg13g2_nand2_1 _1296_ (.Y(_0422_),
    .A(net366),
    .B(_0415_));
 sg13g2_a22oi_1 _1297_ (.Y(_0423_),
    .B1(_0414_),
    .B2(net223),
    .A2(net198),
    .A1(net345));
 sg13g2_nand2_1 _1298_ (.Y(_0068_),
    .A(_0422_),
    .B(_0423_));
 sg13g2_nand2_1 _1299_ (.Y(_0424_),
    .A(net402),
    .B(_0415_));
 sg13g2_a22oi_1 _1300_ (.Y(_0425_),
    .B1(_0414_),
    .B2(\pmod_1414.GPout[4] ),
    .A2(net196),
    .A1(net334));
 sg13g2_nand2_1 _1301_ (.Y(_0069_),
    .A(_0424_),
    .B(_0425_));
 sg13g2_nand2_1 _1302_ (.Y(_0426_),
    .A(net427),
    .B(_0415_));
 sg13g2_a22oi_1 _1303_ (.Y(_0427_),
    .B1(_0414_),
    .B2(net218),
    .A2(net193),
    .A1(net362));
 sg13g2_nand2_1 _1304_ (.Y(_0070_),
    .A(_0426_),
    .B(_0427_));
 sg13g2_nand2_1 _1305_ (.Y(_0428_),
    .A(net407),
    .B(_0415_));
 sg13g2_a22oi_1 _1306_ (.Y(_0429_),
    .B1(_0414_),
    .B2(net216),
    .A2(net198),
    .A1(net339));
 sg13g2_nand2_1 _1307_ (.Y(_0071_),
    .A(_0428_),
    .B(_0429_));
 sg13g2_nor2_2 _1308_ (.A(_0249_),
    .B(_0391_),
    .Y(_0430_));
 sg13g2_nor2_2 _1309_ (.A(net194),
    .B(_0430_),
    .Y(_0431_));
 sg13g2_nand2_1 _1310_ (.Y(_0432_),
    .A(net338),
    .B(_0431_));
 sg13g2_a22oi_1 _1311_ (.Y(_0433_),
    .B1(_0430_),
    .B2(net230),
    .A2(net195),
    .A1(net318));
 sg13g2_nand2_1 _1312_ (.Y(_0072_),
    .A(_0432_),
    .B(_0433_));
 sg13g2_nand2_1 _1313_ (.Y(_0434_),
    .A(net351),
    .B(_0431_));
 sg13g2_a22oi_1 _1314_ (.Y(_0435_),
    .B1(_0430_),
    .B2(net227),
    .A2(net195),
    .A1(\pmod_1414.mem_strorage.mem[4][1] ));
 sg13g2_nand2_1 _1315_ (.Y(_0073_),
    .A(_0434_),
    .B(_0435_));
 sg13g2_nand2_1 _1316_ (.Y(_0436_),
    .A(net326),
    .B(_0431_));
 sg13g2_a22oi_1 _1317_ (.Y(_0437_),
    .B1(_0430_),
    .B2(net225),
    .A2(net195),
    .A1(\pmod_1414.mem_strorage.mem[4][2] ));
 sg13g2_nand2_1 _1318_ (.Y(_0074_),
    .A(_0436_),
    .B(_0437_));
 sg13g2_nand2_1 _1319_ (.Y(_0438_),
    .A(net345),
    .B(_0431_));
 sg13g2_a22oi_1 _1320_ (.Y(_0439_),
    .B1(_0430_),
    .B2(net223),
    .A2(net194),
    .A1(\pmod_1414.mem_strorage.mem[4][3] ));
 sg13g2_nand2_1 _1321_ (.Y(_0075_),
    .A(_0438_),
    .B(_0439_));
 sg13g2_nand2_1 _1322_ (.Y(_0440_),
    .A(net334),
    .B(_0431_));
 sg13g2_a22oi_1 _1323_ (.Y(_0441_),
    .B1(_0430_),
    .B2(net221),
    .A2(net195),
    .A1(\pmod_1414.mem_strorage.mem[4][4] ));
 sg13g2_nand2_1 _1324_ (.Y(_0076_),
    .A(_0440_),
    .B(_0441_));
 sg13g2_nand2_1 _1325_ (.Y(_0442_),
    .A(net362),
    .B(_0431_));
 sg13g2_a22oi_1 _1326_ (.Y(_0443_),
    .B1(_0430_),
    .B2(net218),
    .A2(net193),
    .A1(\pmod_1414.mem_strorage.mem[4][5] ));
 sg13g2_nand2_1 _1327_ (.Y(_0077_),
    .A(_0442_),
    .B(_0443_));
 sg13g2_nand2_1 _1328_ (.Y(_0444_),
    .A(net339),
    .B(_0431_));
 sg13g2_a22oi_1 _1329_ (.Y(_0445_),
    .B1(_0430_),
    .B2(net216),
    .A2(net198),
    .A1(\pmod_1414.mem_strorage.mem[4][6] ));
 sg13g2_nand2_1 _1330_ (.Y(_0078_),
    .A(_0444_),
    .B(_0445_));
 sg13g2_nand4_1 _1331_ (.B(\pmod_1414.r_uart_rx_counter[2] ),
    .C(net235),
    .A(_0219_),
    .Y(_0446_),
    .D(net202));
 sg13g2_nor3_2 _1332_ (.A(\pmod_1414.r_uart_rx_counter[1] ),
    .B(\pmod_1414.r_uart_rx_counter[0] ),
    .C(_0446_),
    .Y(_0447_));
 sg13g2_nor2_2 _1333_ (.A(net194),
    .B(_0447_),
    .Y(_0448_));
 sg13g2_nand2_1 _1334_ (.Y(_0449_),
    .A(net318),
    .B(_0448_));
 sg13g2_a22oi_1 _1335_ (.Y(_0450_),
    .B1(_0447_),
    .B2(net230),
    .A2(net194),
    .A1(\pmod_1414.mem_strorage.mem[5][0] ));
 sg13g2_nand2_1 _1336_ (.Y(_0079_),
    .A(_0449_),
    .B(_0450_));
 sg13g2_nand2_1 _1337_ (.Y(_0451_),
    .A(net353),
    .B(_0448_));
 sg13g2_a22oi_1 _1338_ (.Y(_0452_),
    .B1(_0447_),
    .B2(net227),
    .A2(net194),
    .A1(\pmod_1414.mem_strorage.mem[5][1] ));
 sg13g2_nand2_1 _1339_ (.Y(_0080_),
    .A(_0451_),
    .B(_0452_));
 sg13g2_nand2_1 _1340_ (.Y(_0453_),
    .A(net330),
    .B(_0448_));
 sg13g2_a22oi_1 _1341_ (.Y(_0454_),
    .B1(_0447_),
    .B2(net225),
    .A2(net194),
    .A1(\pmod_1414.mem_strorage.mem[5][2] ));
 sg13g2_nand2_1 _1342_ (.Y(_0081_),
    .A(_0453_),
    .B(_0454_));
 sg13g2_nand2_1 _1343_ (.Y(_0455_),
    .A(net405),
    .B(_0448_));
 sg13g2_a22oi_1 _1344_ (.Y(_0456_),
    .B1(_0447_),
    .B2(net223),
    .A2(net194),
    .A1(\pmod_1414.mem_strorage.mem[5][3] ));
 sg13g2_nand2_1 _1345_ (.Y(_0082_),
    .A(_0455_),
    .B(_0456_));
 sg13g2_nand2_1 _1346_ (.Y(_0457_),
    .A(net347),
    .B(_0448_));
 sg13g2_a22oi_1 _1347_ (.Y(_0458_),
    .B1(_0447_),
    .B2(net221),
    .A2(net194),
    .A1(\pmod_1414.mem_strorage.mem[5][4] ));
 sg13g2_nand2_1 _1348_ (.Y(_0083_),
    .A(_0457_),
    .B(_0458_));
 sg13g2_nand2_1 _1349_ (.Y(_0459_),
    .A(net367),
    .B(_0448_));
 sg13g2_a22oi_1 _1350_ (.Y(_0460_),
    .B1(_0447_),
    .B2(net218),
    .A2(net193),
    .A1(\pmod_1414.mem_strorage.mem[5][5] ));
 sg13g2_nand2_1 _1351_ (.Y(_0084_),
    .A(_0459_),
    .B(_0460_));
 sg13g2_nand2_1 _1352_ (.Y(_0461_),
    .A(net343),
    .B(_0448_));
 sg13g2_a22oi_1 _1353_ (.Y(_0462_),
    .B1(_0447_),
    .B2(net216),
    .A2(net193),
    .A1(\pmod_1414.mem_strorage.mem[5][6] ));
 sg13g2_nand2_1 _1354_ (.Y(_0085_),
    .A(_0461_),
    .B(_0462_));
 sg13g2_nor2_2 _1355_ (.A(_0249_),
    .B(_0446_),
    .Y(_0463_));
 sg13g2_nor2_2 _1356_ (.A(net191),
    .B(_0463_),
    .Y(_0464_));
 sg13g2_nand2_1 _1357_ (.Y(_0465_),
    .A(net423),
    .B(_0464_));
 sg13g2_a22oi_1 _1358_ (.Y(_0466_),
    .B1(_0463_),
    .B2(net229),
    .A2(net191),
    .A1(net381));
 sg13g2_nand2_1 _1359_ (.Y(_0086_),
    .A(_0465_),
    .B(_0466_));
 sg13g2_nand2_1 _1360_ (.Y(_0467_),
    .A(net512),
    .B(_0464_));
 sg13g2_a22oi_1 _1361_ (.Y(_0468_),
    .B1(_0463_),
    .B2(net226),
    .A2(net193),
    .A1(net294));
 sg13g2_nand2_1 _1362_ (.Y(_0087_),
    .A(_0467_),
    .B(_0468_));
 sg13g2_nand2_1 _1363_ (.Y(_0469_),
    .A(net447),
    .B(_0464_));
 sg13g2_a22oi_1 _1364_ (.Y(_0470_),
    .B1(_0463_),
    .B2(net225),
    .A2(net191),
    .A1(\pmod_1414.mem_strorage.mem[8][2] ));
 sg13g2_nand2_1 _1365_ (.Y(_0088_),
    .A(_0469_),
    .B(_0470_));
 sg13g2_nand2_1 _1366_ (.Y(_0471_),
    .A(net506),
    .B(_0464_));
 sg13g2_a22oi_1 _1367_ (.Y(_0472_),
    .B1(_0463_),
    .B2(net222),
    .A2(net191),
    .A1(net442));
 sg13g2_nand2_1 _1368_ (.Y(_0089_),
    .A(_0471_),
    .B(_0472_));
 sg13g2_nand2_1 _1369_ (.Y(_0473_),
    .A(net411),
    .B(_0464_));
 sg13g2_a22oi_1 _1370_ (.Y(_0474_),
    .B1(_0463_),
    .B2(net221),
    .A2(net191),
    .A1(\pmod_1414.mem_strorage.mem[8][4] ));
 sg13g2_nand2_1 _1371_ (.Y(_0090_),
    .A(_0473_),
    .B(_0474_));
 sg13g2_nand2_1 _1372_ (.Y(_0475_),
    .A(net434),
    .B(_0464_));
 sg13g2_a22oi_1 _1373_ (.Y(_0476_),
    .B1(_0463_),
    .B2(\pmod_1414.GPout[5] ),
    .A2(net190),
    .A1(\pmod_1414.mem_strorage.mem[8][5] ));
 sg13g2_nand2_1 _1374_ (.Y(_0091_),
    .A(_0475_),
    .B(_0476_));
 sg13g2_nand2_1 _1375_ (.Y(_0477_),
    .A(net476),
    .B(_0464_));
 sg13g2_a22oi_1 _1376_ (.Y(_0478_),
    .B1(_0463_),
    .B2(\pmod_1414.GPout[6] ),
    .A2(net199),
    .A1(\pmod_1414.mem_strorage.mem[8][6] ));
 sg13g2_nand2_1 _1377_ (.Y(_0092_),
    .A(_0477_),
    .B(_0478_));
 sg13g2_nand4_1 _1378_ (.B(_0220_),
    .C(net235),
    .A(\pmod_1414.r_uart_rx_counter[3] ),
    .Y(_0479_),
    .D(net202));
 sg13g2_nor3_2 _1379_ (.A(net231),
    .B(net232),
    .C(_0479_),
    .Y(_0480_));
 sg13g2_nor2_2 _1380_ (.A(net189),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_nand2_1 _1381_ (.Y(_0482_),
    .A(net381),
    .B(_0481_));
 sg13g2_a22oi_1 _1382_ (.Y(_0483_),
    .B1(_0480_),
    .B2(net228),
    .A2(net190),
    .A1(\pmod_1414.mem_strorage.mem[9][0] ));
 sg13g2_nand2_1 _1383_ (.Y(_0093_),
    .A(_0482_),
    .B(_0483_));
 sg13g2_nand2_1 _1384_ (.Y(_0484_),
    .A(net294),
    .B(_0481_));
 sg13g2_a22oi_1 _1385_ (.Y(_0485_),
    .B1(_0480_),
    .B2(net227),
    .A2(net191),
    .A1(\pmod_1414.mem_strorage.mem[9][1] ));
 sg13g2_nand2_1 _1386_ (.Y(_0094_),
    .A(_0484_),
    .B(_0485_));
 sg13g2_nand2_1 _1387_ (.Y(_0486_),
    .A(net498),
    .B(_0481_));
 sg13g2_a22oi_1 _1388_ (.Y(_0487_),
    .B1(_0480_),
    .B2(net224),
    .A2(net190),
    .A1(net451));
 sg13g2_nand2_1 _1389_ (.Y(_0095_),
    .A(_0486_),
    .B(_0487_));
 sg13g2_nand2_1 _1390_ (.Y(_0488_),
    .A(net442),
    .B(_0481_));
 sg13g2_a22oi_1 _1391_ (.Y(_0489_),
    .B1(_0480_),
    .B2(net222),
    .A2(net188),
    .A1(net371));
 sg13g2_nand2_1 _1392_ (.Y(_0096_),
    .A(_0488_),
    .B(_0489_));
 sg13g2_nand2_1 _1393_ (.Y(_0490_),
    .A(net449),
    .B(_0481_));
 sg13g2_a22oi_1 _1394_ (.Y(_0491_),
    .B1(_0480_),
    .B2(net220),
    .A2(net188),
    .A1(net403));
 sg13g2_nand2_1 _1395_ (.Y(_0097_),
    .A(_0490_),
    .B(_0491_));
 sg13g2_nand2_1 _1396_ (.Y(_0492_),
    .A(net484),
    .B(_0481_));
 sg13g2_a22oi_1 _1397_ (.Y(_0493_),
    .B1(_0480_),
    .B2(net219),
    .A2(net187),
    .A1(net396));
 sg13g2_nand2_1 _1398_ (.Y(_0098_),
    .A(_0492_),
    .B(_0493_));
 sg13g2_nand2_1 _1399_ (.Y(_0494_),
    .A(net501),
    .B(_0481_));
 sg13g2_a22oi_1 _1400_ (.Y(_0495_),
    .B1(_0480_),
    .B2(net217),
    .A2(net187),
    .A1(net424));
 sg13g2_nand2_1 _1401_ (.Y(_0099_),
    .A(_0494_),
    .B(_0495_));
 sg13g2_nor3_2 _1402_ (.A(net231),
    .B(net232),
    .C(_0391_),
    .Y(_0496_));
 sg13g2_nor2_2 _1403_ (.A(net196),
    .B(_0496_),
    .Y(_0497_));
 sg13g2_nand2_1 _1404_ (.Y(_0498_),
    .A(net304),
    .B(_0497_));
 sg13g2_a22oi_1 _1405_ (.Y(_0499_),
    .B1(_0496_),
    .B2(net230),
    .A2(net195),
    .A1(\pmod_1414.mem_strorage.mem[1][0] ));
 sg13g2_nand2_1 _1406_ (.Y(_0100_),
    .A(_0498_),
    .B(_0499_));
 sg13g2_nand2_1 _1407_ (.Y(_0500_),
    .A(net312),
    .B(_0497_));
 sg13g2_a22oi_1 _1408_ (.Y(_0501_),
    .B1(_0496_),
    .B2(net227),
    .A2(net197),
    .A1(\pmod_1414.mem_strorage.mem[1][1] ));
 sg13g2_nand2_1 _1409_ (.Y(_0101_),
    .A(_0500_),
    .B(_0501_));
 sg13g2_nand2_1 _1410_ (.Y(_0502_),
    .A(net298),
    .B(_0497_));
 sg13g2_a22oi_1 _1411_ (.Y(_0503_),
    .B1(_0496_),
    .B2(net225),
    .A2(net196),
    .A1(\pmod_1414.mem_strorage.mem[1][2] ));
 sg13g2_nand2_1 _1412_ (.Y(_0102_),
    .A(_0502_),
    .B(_0503_));
 sg13g2_nand2_1 _1413_ (.Y(_0504_),
    .A(net292),
    .B(_0497_));
 sg13g2_a22oi_1 _1414_ (.Y(_0505_),
    .B1(_0496_),
    .B2(net223),
    .A2(net198),
    .A1(\pmod_1414.mem_strorage.mem[1][3] ));
 sg13g2_nand2_1 _1415_ (.Y(_0103_),
    .A(_0504_),
    .B(_0505_));
 sg13g2_nand2_1 _1416_ (.Y(_0506_),
    .A(net290),
    .B(_0497_));
 sg13g2_a22oi_1 _1417_ (.Y(_0507_),
    .B1(_0496_),
    .B2(net221),
    .A2(net196),
    .A1(\pmod_1414.mem_strorage.mem[1][4] ));
 sg13g2_nand2_1 _1418_ (.Y(_0104_),
    .A(_0506_),
    .B(_0507_));
 sg13g2_nand2_1 _1419_ (.Y(_0508_),
    .A(net306),
    .B(_0497_));
 sg13g2_a22oi_1 _1420_ (.Y(_0509_),
    .B1(_0496_),
    .B2(net218),
    .A2(net193),
    .A1(\pmod_1414.mem_strorage.mem[1][5] ));
 sg13g2_nand2_1 _1421_ (.Y(_0105_),
    .A(_0508_),
    .B(_0509_));
 sg13g2_nand2_1 _1422_ (.Y(_0510_),
    .A(net314),
    .B(_0497_));
 sg13g2_a22oi_1 _1423_ (.Y(_0511_),
    .B1(_0496_),
    .B2(net216),
    .A2(net198),
    .A1(\pmod_1414.mem_strorage.mem[1][6] ));
 sg13g2_nand2_1 _1424_ (.Y(_0106_),
    .A(_0510_),
    .B(_0511_));
 sg13g2_or2_2 _1425_ (.X(_0512_),
    .B(_0446_),
    .A(_0392_));
 sg13g2_nand2_2 _1426_ (.Y(_0513_),
    .A(net183),
    .B(_0512_));
 sg13g2_nor2_1 _1427_ (.A(net513),
    .B(_0513_),
    .Y(_0514_));
 sg13g2_nor2_1 _1428_ (.A(net507),
    .B(net182),
    .Y(_0515_));
 sg13g2_nor2_1 _1429_ (.A(net230),
    .B(_0512_),
    .Y(_0516_));
 sg13g2_nor3_1 _1430_ (.A(_0514_),
    .B(_0515_),
    .C(_0516_),
    .Y(_0107_));
 sg13g2_nor2_1 _1431_ (.A(net478),
    .B(_0513_),
    .Y(_0517_));
 sg13g2_nor2_1 _1432_ (.A(net227),
    .B(_0512_),
    .Y(_0518_));
 sg13g2_nor2_1 _1433_ (.A(\pmod_1414.mem_strorage.mem[6][1] ),
    .B(net183),
    .Y(_0519_));
 sg13g2_nor3_1 _1434_ (.A(_0517_),
    .B(_0518_),
    .C(_0519_),
    .Y(_0108_));
 sg13g2_nor2_1 _1435_ (.A(net503),
    .B(_0513_),
    .Y(_0520_));
 sg13g2_nor2_1 _1436_ (.A(\pmod_1414.mem_strorage.mem[6][2] ),
    .B(net183),
    .Y(_0521_));
 sg13g2_nor2_1 _1437_ (.A(net225),
    .B(_0512_),
    .Y(_0522_));
 sg13g2_nor3_1 _1438_ (.A(_0520_),
    .B(_0521_),
    .C(_0522_),
    .Y(_0109_));
 sg13g2_nor2_1 _1439_ (.A(net496),
    .B(_0513_),
    .Y(_0523_));
 sg13g2_nor2_1 _1440_ (.A(\pmod_1414.mem_strorage.mem[6][3] ),
    .B(net182),
    .Y(_0524_));
 sg13g2_nor2_1 _1441_ (.A(\pmod_1414.GPout[3] ),
    .B(_0512_),
    .Y(_0525_));
 sg13g2_nor3_1 _1442_ (.A(_0523_),
    .B(_0524_),
    .C(_0525_),
    .Y(_0110_));
 sg13g2_nor2_1 _1443_ (.A(net517),
    .B(_0513_),
    .Y(_0526_));
 sg13g2_nor2_1 _1444_ (.A(net483),
    .B(net182),
    .Y(_0527_));
 sg13g2_nor2_1 _1445_ (.A(net221),
    .B(_0512_),
    .Y(_0528_));
 sg13g2_nor3_1 _1446_ (.A(_0526_),
    .B(_0527_),
    .C(_0528_),
    .Y(_0111_));
 sg13g2_nor2_1 _1447_ (.A(\pmod_1414.mem_strorage.mem[5][5] ),
    .B(_0513_),
    .Y(_0529_));
 sg13g2_nor2_1 _1448_ (.A(net218),
    .B(_0512_),
    .Y(_0530_));
 sg13g2_nor2_1 _1449_ (.A(net469),
    .B(net183),
    .Y(_0531_));
 sg13g2_nor3_1 _1450_ (.A(_0529_),
    .B(_0530_),
    .C(_0531_),
    .Y(_0112_));
 sg13g2_nor2_1 _1451_ (.A(net473),
    .B(_0513_),
    .Y(_0532_));
 sg13g2_nor2_1 _1452_ (.A(\pmod_1414.mem_strorage.mem[6][6] ),
    .B(net183),
    .Y(_0533_));
 sg13g2_nor2_1 _1453_ (.A(net216),
    .B(_0512_),
    .Y(_0534_));
 sg13g2_nor3_1 _1454_ (.A(_0532_),
    .B(_0533_),
    .C(_0534_),
    .Y(_0113_));
 sg13g2_or2_2 _1455_ (.X(_0535_),
    .B(_0446_),
    .A(_0413_));
 sg13g2_nand2_2 _1456_ (.Y(_0536_),
    .A(net182),
    .B(_0535_));
 sg13g2_nor2_1 _1457_ (.A(net507),
    .B(_0536_),
    .Y(_0537_));
 sg13g2_nor2_1 _1458_ (.A(net229),
    .B(_0535_),
    .Y(_0538_));
 sg13g2_nor2_1 _1459_ (.A(net423),
    .B(net182),
    .Y(_0539_));
 sg13g2_nor3_1 _1460_ (.A(_0537_),
    .B(_0538_),
    .C(_0539_),
    .Y(_0114_));
 sg13g2_nor2_1 _1461_ (.A(net533),
    .B(_0536_),
    .Y(_0540_));
 sg13g2_nor2_1 _1462_ (.A(\pmod_1414.GPout[1] ),
    .B(_0535_),
    .Y(_0541_));
 sg13g2_nor2_1 _1463_ (.A(net512),
    .B(_0397_),
    .Y(_0542_));
 sg13g2_nor3_1 _1464_ (.A(_0540_),
    .B(_0541_),
    .C(_0542_),
    .Y(_0115_));
 sg13g2_nor2_1 _1465_ (.A(net516),
    .B(_0536_),
    .Y(_0543_));
 sg13g2_nor2_1 _1466_ (.A(net447),
    .B(net182),
    .Y(_0544_));
 sg13g2_nor2_1 _1467_ (.A(net225),
    .B(_0535_),
    .Y(_0545_));
 sg13g2_nor3_1 _1468_ (.A(_0543_),
    .B(_0544_),
    .C(_0545_),
    .Y(_0116_));
 sg13g2_nor2_1 _1469_ (.A(net520),
    .B(_0536_),
    .Y(_0546_));
 sg13g2_nor2_1 _1470_ (.A(\pmod_1414.GPout[3] ),
    .B(_0535_),
    .Y(_0547_));
 sg13g2_nor2_1 _1471_ (.A(net506),
    .B(net182),
    .Y(_0548_));
 sg13g2_nor3_1 _1472_ (.A(_0546_),
    .B(_0547_),
    .C(_0548_),
    .Y(_0117_));
 sg13g2_nor2_1 _1473_ (.A(net483),
    .B(_0536_),
    .Y(_0549_));
 sg13g2_nor2_1 _1474_ (.A(net221),
    .B(_0535_),
    .Y(_0550_));
 sg13g2_nor2_1 _1475_ (.A(net411),
    .B(net182),
    .Y(_0551_));
 sg13g2_nor3_1 _1476_ (.A(_0549_),
    .B(_0550_),
    .C(_0551_),
    .Y(_0118_));
 sg13g2_nor2_1 _1477_ (.A(net469),
    .B(_0536_),
    .Y(_0552_));
 sg13g2_nor2_1 _1478_ (.A(net434),
    .B(net183),
    .Y(_0553_));
 sg13g2_nor2_1 _1479_ (.A(net218),
    .B(_0535_),
    .Y(_0554_));
 sg13g2_nor3_1 _1480_ (.A(_0552_),
    .B(_0553_),
    .C(_0554_),
    .Y(_0119_));
 sg13g2_nor2_1 _1481_ (.A(net523),
    .B(_0536_),
    .Y(_0555_));
 sg13g2_nor2_1 _1482_ (.A(net476),
    .B(net183),
    .Y(_0556_));
 sg13g2_nor2_1 _1483_ (.A(net216),
    .B(_0535_),
    .Y(_0557_));
 sg13g2_nor3_1 _1484_ (.A(_0555_),
    .B(_0556_),
    .C(_0557_),
    .Y(_0120_));
 sg13g2_nor2_2 _1485_ (.A(_0413_),
    .B(_0479_),
    .Y(_0558_));
 sg13g2_nor2_2 _1486_ (.A(net187),
    .B(_0558_),
    .Y(_0559_));
 sg13g2_nand2_1 _1487_ (.Y(_0560_),
    .A(net421),
    .B(_0559_));
 sg13g2_a22oi_1 _1488_ (.Y(_0561_),
    .B1(_0558_),
    .B2(net228),
    .A2(net190),
    .A1(\pmod_1414.mem_strorage.mem[11][0] ));
 sg13g2_nand2_1 _1489_ (.Y(_0121_),
    .A(_0560_),
    .B(_0561_));
 sg13g2_nand2_1 _1490_ (.Y(_0562_),
    .A(net316),
    .B(_0559_));
 sg13g2_a22oi_1 _1491_ (.Y(_0563_),
    .B1(_0558_),
    .B2(net226),
    .A2(net190),
    .A1(\pmod_1414.mem_strorage.mem[11][1] ));
 sg13g2_nand2_1 _1492_ (.Y(_0122_),
    .A(_0562_),
    .B(_0563_));
 sg13g2_nand2_1 _1493_ (.Y(_0564_),
    .A(net349),
    .B(_0559_));
 sg13g2_a22oi_1 _1494_ (.Y(_0565_),
    .B1(_0558_),
    .B2(net224),
    .A2(net189),
    .A1(\pmod_1414.mem_strorage.mem[11][2] ));
 sg13g2_nand2_1 _1495_ (.Y(_0123_),
    .A(_0564_),
    .B(_0565_));
 sg13g2_nand2_1 _1496_ (.Y(_0566_),
    .A(net398),
    .B(_0559_));
 sg13g2_a22oi_1 _1497_ (.Y(_0567_),
    .B1(_0558_),
    .B2(net223),
    .A2(net188),
    .A1(\pmod_1414.mem_strorage.mem[11][3] ));
 sg13g2_nand2_1 _1498_ (.Y(_0124_),
    .A(_0566_),
    .B(_0567_));
 sg13g2_nand2_1 _1499_ (.Y(_0568_),
    .A(net383),
    .B(_0559_));
 sg13g2_a22oi_1 _1500_ (.Y(_0569_),
    .B1(_0558_),
    .B2(net220),
    .A2(net188),
    .A1(\pmod_1414.mem_strorage.mem[11][4] ));
 sg13g2_nand2_1 _1501_ (.Y(_0125_),
    .A(_0568_),
    .B(_0569_));
 sg13g2_nand2_1 _1502_ (.Y(_0570_),
    .A(net436),
    .B(_0559_));
 sg13g2_a22oi_1 _1503_ (.Y(_0571_),
    .B1(_0558_),
    .B2(net219),
    .A2(net188),
    .A1(\pmod_1414.mem_strorage.mem[11][5] ));
 sg13g2_nand2_1 _1504_ (.Y(_0126_),
    .A(_0570_),
    .B(_0571_));
 sg13g2_nand2_1 _1505_ (.Y(_0572_),
    .A(net373),
    .B(_0559_));
 sg13g2_a22oi_1 _1506_ (.Y(_0573_),
    .B1(_0558_),
    .B2(net217),
    .A2(net187),
    .A1(\pmod_1414.mem_strorage.mem[11][6] ));
 sg13g2_nand2_1 _1507_ (.Y(_0127_),
    .A(_0572_),
    .B(_0573_));
 sg13g2_nor2_2 _1508_ (.A(_0392_),
    .B(_0394_),
    .Y(_0574_));
 sg13g2_nor2_2 _1509_ (.A(net184),
    .B(_0574_),
    .Y(_0575_));
 sg13g2_nand2_1 _1510_ (.Y(_0576_),
    .A(net413),
    .B(_0575_));
 sg13g2_a22oi_1 _1511_ (.Y(_0577_),
    .B1(_0574_),
    .B2(net228),
    .A2(net186),
    .A1(\pmod_1414.mem_strorage.mem[14][0] ));
 sg13g2_nand2_1 _1512_ (.Y(_0128_),
    .A(_0576_),
    .B(_0577_));
 sg13g2_nand2_1 _1513_ (.Y(_0578_),
    .A(net324),
    .B(_0575_));
 sg13g2_a22oi_1 _1514_ (.Y(_0579_),
    .B1(_0574_),
    .B2(net226),
    .A2(net192),
    .A1(\pmod_1414.mem_strorage.mem[14][1] ));
 sg13g2_nand2_1 _1515_ (.Y(_0129_),
    .A(_0578_),
    .B(_0579_));
 sg13g2_a22oi_1 _1516_ (.Y(_0580_),
    .B1(_0575_),
    .B2(\pmod_1414.mem_strorage.mem[13][2] ),
    .A2(_0574_),
    .A1(net224));
 sg13g2_o21ai_1 _1517_ (.B1(_0580_),
    .Y(_0130_),
    .A1(_0233_),
    .A2(net180));
 sg13g2_a22oi_1 _1518_ (.Y(_0581_),
    .B1(_0575_),
    .B2(net505),
    .A2(_0574_),
    .A1(net222));
 sg13g2_o21ai_1 _1519_ (.B1(_0581_),
    .Y(_0131_),
    .A1(_0234_),
    .A2(net180));
 sg13g2_nand2_1 _1520_ (.Y(_0582_),
    .A(net355),
    .B(_0575_));
 sg13g2_a22oi_1 _1521_ (.Y(_0583_),
    .B1(_0574_),
    .B2(net220),
    .A2(net184),
    .A1(\pmod_1414.mem_strorage.mem[14][4] ));
 sg13g2_nand2_1 _1522_ (.Y(_0132_),
    .A(_0582_),
    .B(_0583_));
 sg13g2_a22oi_1 _1523_ (.Y(_0584_),
    .B1(_0575_),
    .B2(net459),
    .A2(_0574_),
    .A1(net219));
 sg13g2_o21ai_1 _1524_ (.B1(_0584_),
    .Y(_0133_),
    .A1(_0235_),
    .A2(net180));
 sg13g2_nand2_1 _1525_ (.Y(_0585_),
    .A(net390),
    .B(_0575_));
 sg13g2_a22oi_1 _1526_ (.Y(_0586_),
    .B1(_0574_),
    .B2(net217),
    .A2(net184),
    .A1(\pmod_1414.mem_strorage.mem[14][6] ));
 sg13g2_nand2_1 _1527_ (.Y(_0134_),
    .A(_0585_),
    .B(_0586_));
 sg13g2_nor2_2 _1528_ (.A(_0394_),
    .B(_0413_),
    .Y(_0587_));
 sg13g2_nor2_2 _1529_ (.A(net184),
    .B(_0587_),
    .Y(_0588_));
 sg13g2_a22oi_1 _1530_ (.Y(_0589_),
    .B1(_0588_),
    .B2(net499),
    .A2(_0587_),
    .A1(net228));
 sg13g2_o21ai_1 _1531_ (.B1(_0589_),
    .Y(_0135_),
    .A1(_0236_),
    .A2(net181));
 sg13g2_a22oi_1 _1532_ (.Y(_0590_),
    .B1(_0588_),
    .B2(net488),
    .A2(_0587_),
    .A1(net226));
 sg13g2_o21ai_1 _1533_ (.B1(_0590_),
    .Y(_0136_),
    .A1(_0237_),
    .A2(net181));
 sg13g2_a22oi_1 _1534_ (.Y(_0591_),
    .B1(_0588_),
    .B2(net471),
    .A2(_0587_),
    .A1(net224));
 sg13g2_o21ai_1 _1535_ (.B1(_0591_),
    .Y(_0137_),
    .A1(_0238_),
    .A2(net180));
 sg13g2_nand2_1 _1536_ (.Y(_0592_),
    .A(net431),
    .B(_0588_));
 sg13g2_a22oi_1 _1537_ (.Y(_0593_),
    .B1(_0587_),
    .B2(net222),
    .A2(net184),
    .A1(\pmod_1414.mem_strorage.mem[15][3] ));
 sg13g2_nand2_1 _1538_ (.Y(_0138_),
    .A(_0592_),
    .B(_0593_));
 sg13g2_a22oi_1 _1539_ (.Y(_0594_),
    .B1(_0588_),
    .B2(net514),
    .A2(_0587_),
    .A1(net220));
 sg13g2_o21ai_1 _1540_ (.B1(_0594_),
    .Y(_0139_),
    .A1(_0239_),
    .A2(net180));
 sg13g2_a22oi_1 _1541_ (.Y(_0595_),
    .B1(_0588_),
    .B2(net489),
    .A2(_0587_),
    .A1(net219));
 sg13g2_o21ai_1 _1542_ (.B1(_0595_),
    .Y(_0140_),
    .A1(_0240_),
    .A2(net180));
 sg13g2_nand2_1 _1543_ (.Y(_0596_),
    .A(net415),
    .B(_0588_));
 sg13g2_a22oi_1 _1544_ (.Y(_0597_),
    .B1(_0587_),
    .B2(net217),
    .A2(net184),
    .A1(\pmod_1414.mem_strorage.mem[15][6] ));
 sg13g2_nand2_1 _1545_ (.Y(_0141_),
    .A(_0596_),
    .B(_0597_));
 sg13g2_nor2_2 _1546_ (.A(_0249_),
    .B(_0479_),
    .Y(_0598_));
 sg13g2_nor2_2 _1547_ (.A(net184),
    .B(_0598_),
    .Y(_0599_));
 sg13g2_nand2_1 _1548_ (.Y(_0600_),
    .A(net440),
    .B(_0599_));
 sg13g2_a22oi_1 _1549_ (.Y(_0601_),
    .B1(_0598_),
    .B2(net229),
    .A2(net186),
    .A1(\pmod_1414.mem_strorage.mem[12][0] ));
 sg13g2_nand2_1 _1550_ (.Y(_0142_),
    .A(_0600_),
    .B(_0601_));
 sg13g2_nand2_1 _1551_ (.Y(_0602_),
    .A(net450),
    .B(_0599_));
 sg13g2_a22oi_1 _1552_ (.Y(_0603_),
    .B1(_0598_),
    .B2(net226),
    .A2(net192),
    .A1(net359));
 sg13g2_nand2_1 _1553_ (.Y(_0143_),
    .A(_0602_),
    .B(_0603_));
 sg13g2_nand2_1 _1554_ (.Y(_0604_),
    .A(net491),
    .B(_0599_));
 sg13g2_a22oi_1 _1555_ (.Y(_0605_),
    .B1(_0598_),
    .B2(net225),
    .A2(net186),
    .A1(\pmod_1414.mem_strorage.mem[12][2] ));
 sg13g2_nand2_1 _1556_ (.Y(_0144_),
    .A(_0604_),
    .B(_0605_));
 sg13g2_nand2_1 _1557_ (.Y(_0606_),
    .A(net457),
    .B(_0599_));
 sg13g2_a22oi_1 _1558_ (.Y(_0607_),
    .B1(_0598_),
    .B2(net223),
    .A2(net185),
    .A1(\pmod_1414.mem_strorage.mem[12][3] ));
 sg13g2_nand2_1 _1559_ (.Y(_0145_),
    .A(_0606_),
    .B(_0607_));
 sg13g2_nand2_1 _1560_ (.Y(_0608_),
    .A(net446),
    .B(_0599_));
 sg13g2_a22oi_1 _1561_ (.Y(_0609_),
    .B1(_0598_),
    .B2(net220),
    .A2(net185),
    .A1(net385));
 sg13g2_nand2_1 _1562_ (.Y(_0146_),
    .A(_0608_),
    .B(_0609_));
 sg13g2_nand2_1 _1563_ (.Y(_0610_),
    .A(net443),
    .B(_0599_));
 sg13g2_a22oi_1 _1564_ (.Y(_0611_),
    .B1(_0598_),
    .B2(net219),
    .A2(net184),
    .A1(\pmod_1414.mem_strorage.mem[12][5] ));
 sg13g2_nand2_1 _1565_ (.Y(_0147_),
    .A(_0610_),
    .B(_0611_));
 sg13g2_nand2_1 _1566_ (.Y(_0612_),
    .A(net428),
    .B(_0599_));
 sg13g2_a22oi_1 _1567_ (.Y(_0613_),
    .B1(_0598_),
    .B2(net217),
    .A2(net185),
    .A1(\pmod_1414.mem_strorage.mem[12][6] ));
 sg13g2_nand2_1 _1568_ (.Y(_0148_),
    .A(_0612_),
    .B(_0613_));
 sg13g2_nor3_2 _1569_ (.A(net231),
    .B(net232),
    .C(_0394_),
    .Y(_0614_));
 sg13g2_nor2_2 _1570_ (.A(net186),
    .B(_0614_),
    .Y(_0615_));
 sg13g2_a22oi_1 _1571_ (.Y(_0616_),
    .B1(_0615_),
    .B2(net480),
    .A2(_0614_),
    .A1(net228));
 sg13g2_o21ai_1 _1572_ (.B1(_0616_),
    .Y(_0149_),
    .A1(_0228_),
    .A2(net181));
 sg13g2_nand2_1 _1573_ (.Y(_0617_),
    .A(net359),
    .B(_0615_));
 sg13g2_a22oi_1 _1574_ (.Y(_0618_),
    .B1(_0614_),
    .B2(net226),
    .A2(net192),
    .A1(net324));
 sg13g2_nand2_1 _1575_ (.Y(_0150_),
    .A(_0617_),
    .B(_0618_));
 sg13g2_a22oi_1 _1576_ (.Y(_0619_),
    .B1(_0615_),
    .B2(\pmod_1414.mem_strorage.mem[12][2] ),
    .A2(_0614_),
    .A1(net224));
 sg13g2_o21ai_1 _1577_ (.B1(_0619_),
    .Y(_0151_),
    .A1(_0229_),
    .A2(net180));
 sg13g2_a22oi_1 _1578_ (.Y(_0620_),
    .B1(_0615_),
    .B2(net486),
    .A2(_0614_),
    .A1(net222));
 sg13g2_o21ai_1 _1579_ (.B1(_0620_),
    .Y(_0152_),
    .A1(_0230_),
    .A2(net181));
 sg13g2_nand2_1 _1580_ (.Y(_0621_),
    .A(net385),
    .B(_0615_));
 sg13g2_a22oi_1 _1581_ (.Y(_0622_),
    .B1(_0614_),
    .B2(net220),
    .A2(net185),
    .A1(net355));
 sg13g2_nand2_1 _1582_ (.Y(_0153_),
    .A(_0621_),
    .B(_0622_));
 sg13g2_a22oi_1 _1583_ (.Y(_0623_),
    .B1(_0615_),
    .B2(net510),
    .A2(_0614_),
    .A1(net219));
 sg13g2_o21ai_1 _1584_ (.B1(_0623_),
    .Y(_0154_),
    .A1(_0231_),
    .A2(net180));
 sg13g2_a22oi_1 _1585_ (.Y(_0624_),
    .B1(_0615_),
    .B2(net438),
    .A2(_0614_),
    .A1(net217));
 sg13g2_o21ai_1 _1586_ (.B1(_0624_),
    .Y(_0155_),
    .A1(_0232_),
    .A2(net181));
 sg13g2_mux2_1 _1587_ (.A0(net228),
    .A1(net534),
    .S(_0395_),
    .X(_0156_));
 sg13g2_nand2_1 _1588_ (.Y(_0625_),
    .A(net475),
    .B(net201));
 sg13g2_o21ai_1 _1589_ (.B1(_0625_),
    .Y(_0157_),
    .A1(_0222_),
    .A2(net201));
 sg13g2_mux2_1 _1590_ (.A0(net224),
    .A1(net511),
    .S(net201),
    .X(_0158_));
 sg13g2_mux2_1 _1591_ (.A0(net222),
    .A1(net535),
    .S(net201),
    .X(_0159_));
 sg13g2_mux2_1 _1592_ (.A0(net220),
    .A1(net538),
    .S(net201),
    .X(_0160_));
 sg13g2_mux2_1 _1593_ (.A0(net219),
    .A1(net532),
    .S(net201),
    .X(_0161_));
 sg13g2_mux2_1 _1594_ (.A0(net217),
    .A1(net528),
    .S(net201),
    .X(_0162_));
 sg13g2_nor2_1 _1595_ (.A(net493),
    .B(net468),
    .Y(_0626_));
 sg13g2_nand2b_1 _1596_ (.Y(_0627_),
    .B(_0626_),
    .A_N(\pmod_1414.RX.RxD_sync[1] ));
 sg13g2_nand3_1 _1597_ (.B(\pmod_1414.RX.Filter_cnt[1] ),
    .C(\pmod_1414.RX.RxD_sync[1] ),
    .A(\pmod_1414.RX.Filter_cnt[0] ),
    .Y(_0628_));
 sg13g2_nand3_1 _1598_ (.B(_0627_),
    .C(_0628_),
    .A(net234),
    .Y(_0629_));
 sg13g2_mux2_1 _1599_ (.A0(net273),
    .A1(\pmod_1414.RX.Filter_cnt[0] ),
    .S(_0629_),
    .X(_0163_));
 sg13g2_xnor2_1 _1600_ (.Y(_0630_),
    .A(net454),
    .B(net273));
 sg13g2_nor2_1 _1601_ (.A(_0629_),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_xor2_1 _1602_ (.B(_0631_),
    .A(net468),
    .X(_0164_));
 sg13g2_nand3_1 _1603_ (.B(net468),
    .C(\pmod_1414.RX.OversamplingTick ),
    .A(net493),
    .Y(_0632_));
 sg13g2_nand2_1 _1604_ (.Y(_0633_),
    .A(\pmod_1414.RX.OversamplingTick ),
    .B(_0626_));
 sg13g2_nand2_1 _1605_ (.Y(_0634_),
    .A(\pmod_1414.RX.RxD_bit ),
    .B(_0633_));
 sg13g2_nand2_1 _1606_ (.Y(_0165_),
    .A(net494),
    .B(_0634_));
 sg13g2_nor2_1 _1607_ (.A(_0226_),
    .B(_0271_),
    .Y(_0635_));
 sg13g2_mux2_1 _1608_ (.A0(net360),
    .A1(\pmod_1414.RX.RxD_data[1] ),
    .S(_0635_),
    .X(_0170_));
 sg13g2_mux2_1 _1609_ (.A0(net461),
    .A1(net452),
    .S(net200),
    .X(_0171_));
 sg13g2_mux2_1 _1610_ (.A0(net452),
    .A1(\pmod_1414.RX.RxD_data[3] ),
    .S(net200),
    .X(_0172_));
 sg13g2_mux2_1 _1611_ (.A0(net464),
    .A1(\pmod_1414.RX.RxD_data[4] ),
    .S(net200),
    .X(_0173_));
 sg13g2_mux2_1 _1612_ (.A0(net485),
    .A1(net462),
    .S(net200),
    .X(_0174_));
 sg13g2_mux2_1 _1613_ (.A0(net462),
    .A1(\pmod_1414.RX.RxD_data[6] ),
    .S(net200),
    .X(_0175_));
 sg13g2_mux2_1 _1614_ (.A0(net466),
    .A1(\pmod_1414.RX.RxD_data[7] ),
    .S(net200),
    .X(_0176_));
 sg13g2_mux2_1 _1615_ (.A0(net518),
    .A1(\pmod_1414.RX.RxD_bit ),
    .S(net200),
    .X(_0177_));
 sg13g2_nor2_1 _1616_ (.A(\pmod_1414.RX.RxD_state[0] ),
    .B(\pmod_1414.RX.RxD_state[1] ),
    .Y(_0636_));
 sg13g2_nor3_1 _1617_ (.A(net557),
    .B(\pmod_1414.RX.RxD_state[1] ),
    .C(\pmod_1414.RX.RxD_state[2] ),
    .Y(_0637_));
 sg13g2_and2_1 _1618_ (.A(_0226_),
    .B(net558),
    .X(_0638_));
 sg13g2_nand2_1 _1619_ (.Y(_0639_),
    .A(net234),
    .B(_0638_));
 sg13g2_nand2b_1 _1620_ (.Y(_0640_),
    .B(\pmod_1414.RX.OversamplingCnt[0] ),
    .A_N(net234));
 sg13g2_nand2_1 _1621_ (.Y(_0641_),
    .A(net264),
    .B(net234));
 sg13g2_o21ai_1 _1622_ (.B1(_0640_),
    .Y(_0178_),
    .A1(_0638_),
    .A2(net265));
 sg13g2_a21o_1 _1623_ (.A2(\pmod_1414.RX.OversamplingCnt[0] ),
    .A1(net234),
    .B1(net543),
    .X(_0642_));
 sg13g2_and3_1 _1624_ (.X(_0179_),
    .A(_0269_),
    .B(_0639_),
    .C(net544));
 sg13g2_nand2_1 _1625_ (.Y(_0643_),
    .A(_0270_),
    .B(_0639_));
 sg13g2_a21oi_1 _1626_ (.A1(_0227_),
    .A2(_0269_),
    .Y(_0180_),
    .B1(_0643_));
 sg13g2_nand3_1 _1627_ (.B(_0270_),
    .C(_0639_),
    .A(net308),
    .Y(_0644_));
 sg13g2_o21ai_1 _1628_ (.B1(_0644_),
    .Y(_0181_),
    .A1(_0271_),
    .A2(_0638_));
 sg13g2_o21ai_1 _1629_ (.B1(net201),
    .Y(_0182_),
    .A1(_0223_),
    .A2(_0390_));
 sg13g2_nor2_2 _1630_ (.A(_0392_),
    .B(_0479_),
    .Y(_0645_));
 sg13g2_nor2_2 _1631_ (.A(net187),
    .B(_0645_),
    .Y(_0646_));
 sg13g2_nand2_1 _1632_ (.Y(_0647_),
    .A(net394),
    .B(_0646_));
 sg13g2_a22oi_1 _1633_ (.Y(_0648_),
    .B1(_0645_),
    .B2(net228),
    .A2(net190),
    .A1(\pmod_1414.mem_strorage.mem[10][0] ));
 sg13g2_nand2_1 _1634_ (.Y(_0183_),
    .A(_0647_),
    .B(_0648_));
 sg13g2_nand2_1 _1635_ (.Y(_0194_),
    .A(net420),
    .B(_0646_));
 sg13g2_a22oi_1 _1636_ (.Y(_0195_),
    .B1(_0645_),
    .B2(net226),
    .A2(net190),
    .A1(net316));
 sg13g2_nand2_1 _1637_ (.Y(_0184_),
    .A(_0194_),
    .B(_0195_));
 sg13g2_nand2_1 _1638_ (.Y(_0196_),
    .A(net451),
    .B(_0646_));
 sg13g2_a22oi_1 _1639_ (.Y(_0197_),
    .B1(_0645_),
    .B2(net224),
    .A2(net190),
    .A1(net349));
 sg13g2_nand2_1 _1640_ (.Y(_0185_),
    .A(_0196_),
    .B(_0197_));
 sg13g2_nand2_1 _1641_ (.Y(_0198_),
    .A(net371),
    .B(_0646_));
 sg13g2_a22oi_1 _1642_ (.Y(_0199_),
    .B1(_0645_),
    .B2(net222),
    .A2(net187),
    .A1(\pmod_1414.mem_strorage.mem[10][3] ));
 sg13g2_nand2_1 _1643_ (.Y(_0186_),
    .A(_0198_),
    .B(_0199_));
 sg13g2_nand2_1 _1644_ (.Y(_0200_),
    .A(net403),
    .B(_0646_));
 sg13g2_a22oi_1 _1645_ (.Y(_0201_),
    .B1(_0645_),
    .B2(net220),
    .A2(net188),
    .A1(net383));
 sg13g2_nand2_1 _1646_ (.Y(_0187_),
    .A(_0200_),
    .B(_0201_));
 sg13g2_nand2_1 _1647_ (.Y(_0202_),
    .A(net396),
    .B(_0646_));
 sg13g2_a22oi_1 _1648_ (.Y(_0203_),
    .B1(_0645_),
    .B2(net219),
    .A2(net187),
    .A1(\pmod_1414.mem_strorage.mem[10][5] ));
 sg13g2_nand2_1 _1649_ (.Y(_0188_),
    .A(_0202_),
    .B(_0203_));
 sg13g2_nand2_1 _1650_ (.Y(_0204_),
    .A(net424),
    .B(_0646_));
 sg13g2_a22oi_1 _1651_ (.Y(_0205_),
    .B1(_0645_),
    .B2(net217),
    .A2(net187),
    .A1(net373));
 sg13g2_nand2_1 _1652_ (.Y(_0189_),
    .A(_0204_),
    .B(_0205_));
 sg13g2_nor2_1 _1653_ (.A(_0224_),
    .B(_0225_),
    .Y(_0206_));
 sg13g2_nand2_1 _1654_ (.Y(_0207_),
    .A(net536),
    .B(net508));
 sg13g2_nor3_1 _1655_ (.A(\pmod_1414.RX.RxD_state[2] ),
    .B(_0636_),
    .C(_0206_),
    .Y(_0208_));
 sg13g2_o21ai_1 _1656_ (.B1(_0271_),
    .Y(_0209_),
    .A1(\pmod_1414.RX.RxD_state[3] ),
    .A2(_0208_));
 sg13g2_nand2_1 _1657_ (.Y(_0210_),
    .A(net536),
    .B(_0209_));
 sg13g2_nand3_1 _1658_ (.B(_0272_),
    .C(_0636_),
    .A(net553),
    .Y(_0211_));
 sg13g2_nand3_1 _1659_ (.B(_0225_),
    .C(_0209_),
    .A(net536),
    .Y(_0212_));
 sg13g2_nand2_1 _1660_ (.Y(_0213_),
    .A(net526),
    .B(_0209_));
 sg13g2_a21oi_1 _1661_ (.A1(\pmod_1414.RX.RxD_state[3] ),
    .A2(_0207_),
    .Y(_0214_),
    .B1(_0213_));
 sg13g2_a21oi_1 _1662_ (.A1(_0226_),
    .A2(_0212_),
    .Y(_0190_),
    .B1(_0214_));
 sg13g2_a21oi_1 _1663_ (.A1(net200),
    .A2(_0206_),
    .Y(_0215_),
    .B1(net526));
 sg13g2_nor2_1 _1664_ (.A(_0214_),
    .B(_0215_),
    .Y(_0191_));
 sg13g2_o21ai_1 _1665_ (.B1(net539),
    .Y(_0216_),
    .A1(net526),
    .A2(_0207_));
 sg13g2_a22oi_1 _1666_ (.Y(_0192_),
    .B1(_0216_),
    .B2(_0209_),
    .A2(_0210_),
    .A1(_0225_));
 sg13g2_a21o_1 _1667_ (.A2(net539),
    .A1(_0224_),
    .B1(_0637_),
    .X(_0217_));
 sg13g2_nand3_1 _1668_ (.B(net554),
    .C(_0217_),
    .A(_0209_),
    .Y(_0218_));
 sg13g2_o21ai_1 _1669_ (.B1(net555),
    .Y(_0193_),
    .A1(_0224_),
    .A2(_0209_));
 sg13g2_dfrbp_1 _1670_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net113),
    .D(_0056_),
    .Q_N(_0783_),
    .Q(\pmod_1414.RX.RxD_sync[0] ));
 sg13g2_dfrbp_1 _1671_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net40),
    .D(_0057_),
    .Q_N(_0782_),
    .Q(\pmod_1414.RX.RxD_sync[1] ));
 sg13g2_dfrbp_1 _1672_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net39),
    .D(net333),
    .Q_N(_0781_),
    .Q(\pmod_1414.mem_strorage.mem[1][0] ));
 sg13g2_dfrbp_1 _1673_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net38),
    .D(net329),
    .Q_N(_0780_),
    .Q(\pmod_1414.mem_strorage.mem[1][1] ));
 sg13g2_dfrbp_1 _1674_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net37),
    .D(net376),
    .Q_N(_0779_),
    .Q(\pmod_1414.mem_strorage.mem[1][2] ));
 sg13g2_dfrbp_1 _1675_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net36),
    .D(net365),
    .Q_N(_0778_),
    .Q(\pmod_1414.mem_strorage.mem[1][3] ));
 sg13g2_dfrbp_1 _1676_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net35),
    .D(_0062_),
    .Q_N(_0777_),
    .Q(\pmod_1414.mem_strorage.mem[1][4] ));
 sg13g2_dfrbp_1 _1677_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net34),
    .D(net389),
    .Q_N(_0776_),
    .Q(\pmod_1414.mem_strorage.mem[1][5] ));
 sg13g2_dfrbp_1 _1678_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net33),
    .D(net393),
    .Q_N(_0775_),
    .Q(\pmod_1414.mem_strorage.mem[1][6] ));
 sg13g2_dfrbp_1 _1679_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net32),
    .D(_0065_),
    .Q_N(_0774_),
    .Q(\pmod_1414.mem_strorage.mem[2][0] ));
 sg13g2_dfrbp_1 _1680_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net31),
    .D(_0066_),
    .Q_N(_0773_),
    .Q(\pmod_1414.mem_strorage.mem[2][1] ));
 sg13g2_dfrbp_1 _1681_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net30),
    .D(_0067_),
    .Q_N(_0772_),
    .Q(\pmod_1414.mem_strorage.mem[2][2] ));
 sg13g2_dfrbp_1 _1682_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net29),
    .D(_0068_),
    .Q_N(_0771_),
    .Q(\pmod_1414.mem_strorage.mem[2][3] ));
 sg13g2_dfrbp_1 _1683_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net28),
    .D(_0069_),
    .Q_N(_0770_),
    .Q(\pmod_1414.mem_strorage.mem[2][4] ));
 sg13g2_dfrbp_1 _1684_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net27),
    .D(_0070_),
    .Q_N(_0769_),
    .Q(\pmod_1414.mem_strorage.mem[2][5] ));
 sg13g2_dfrbp_1 _1685_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net26),
    .D(_0071_),
    .Q_N(_0768_),
    .Q(\pmod_1414.mem_strorage.mem[2][6] ));
 sg13g2_dfrbp_1 _1686_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net25),
    .D(_0072_),
    .Q_N(_0767_),
    .Q(\pmod_1414.mem_strorage.mem[3][0] ));
 sg13g2_dfrbp_1 _1687_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net24),
    .D(net352),
    .Q_N(_0766_),
    .Q(\pmod_1414.mem_strorage.mem[3][1] ));
 sg13g2_dfrbp_1 _1688_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net23),
    .D(net327),
    .Q_N(_0765_),
    .Q(\pmod_1414.mem_strorage.mem[3][2] ));
 sg13g2_dfrbp_1 _1689_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net22),
    .D(net346),
    .Q_N(_0764_),
    .Q(\pmod_1414.mem_strorage.mem[3][3] ));
 sg13g2_dfrbp_1 _1690_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net21),
    .D(net335),
    .Q_N(_0763_),
    .Q(\pmod_1414.mem_strorage.mem[3][4] ));
 sg13g2_dfrbp_1 _1691_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net20),
    .D(net363),
    .Q_N(_0762_),
    .Q(\pmod_1414.mem_strorage.mem[3][5] ));
 sg13g2_dfrbp_1 _1692_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net19),
    .D(net340),
    .Q_N(_0761_),
    .Q(\pmod_1414.mem_strorage.mem[3][6] ));
 sg13g2_dfrbp_1 _1693_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net18),
    .D(net319),
    .Q_N(_0760_),
    .Q(\pmod_1414.mem_strorage.mem[4][0] ));
 sg13g2_dfrbp_1 _1694_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net17),
    .D(net354),
    .Q_N(_0759_),
    .Q(\pmod_1414.mem_strorage.mem[4][1] ));
 sg13g2_dfrbp_1 _1695_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net16),
    .D(net331),
    .Q_N(_0758_),
    .Q(\pmod_1414.mem_strorage.mem[4][2] ));
 sg13g2_dfrbp_1 _1696_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net15),
    .D(net406),
    .Q_N(_0757_),
    .Q(\pmod_1414.mem_strorage.mem[4][3] ));
 sg13g2_dfrbp_1 _1697_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net14),
    .D(net348),
    .Q_N(_0756_),
    .Q(\pmod_1414.mem_strorage.mem[4][4] ));
 sg13g2_dfrbp_1 _1698_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net13),
    .D(net368),
    .Q_N(_0755_),
    .Q(\pmod_1414.mem_strorage.mem[4][5] ));
 sg13g2_dfrbp_1 _1699_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net12),
    .D(net344),
    .Q_N(_0754_),
    .Q(\pmod_1414.mem_strorage.mem[4][6] ));
 sg13g2_dfrbp_1 _1700_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net11),
    .D(_0086_),
    .Q_N(_0753_),
    .Q(\pmod_1414.mem_strorage.mem[7][0] ));
 sg13g2_dfrbp_1 _1701_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net10),
    .D(_0087_),
    .Q_N(_0752_),
    .Q(\pmod_1414.mem_strorage.mem[7][1] ));
 sg13g2_dfrbp_1 _1702_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net9),
    .D(net448),
    .Q_N(_0751_),
    .Q(\pmod_1414.mem_strorage.mem[7][2] ));
 sg13g2_dfrbp_1 _1703_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net8),
    .D(_0089_),
    .Q_N(_0750_),
    .Q(\pmod_1414.mem_strorage.mem[7][3] ));
 sg13g2_dfrbp_1 _1704_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net7),
    .D(net412),
    .Q_N(_0749_),
    .Q(\pmod_1414.mem_strorage.mem[7][4] ));
 sg13g2_dfrbp_1 _1705_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net252),
    .D(net435),
    .Q_N(_0748_),
    .Q(\pmod_1414.mem_strorage.mem[7][5] ));
 sg13g2_dfrbp_1 _1706_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net251),
    .D(net477),
    .Q_N(_0747_),
    .Q(\pmod_1414.mem_strorage.mem[7][6] ));
 sg13g2_dfrbp_1 _1707_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net250),
    .D(net382),
    .Q_N(_0746_),
    .Q(\pmod_1414.mem_strorage.mem[8][0] ));
 sg13g2_dfrbp_1 _1708_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net249),
    .D(net295),
    .Q_N(_0745_),
    .Q(\pmod_1414.mem_strorage.mem[8][1] ));
 sg13g2_dfrbp_1 _1709_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net168),
    .D(_0095_),
    .Q_N(_0744_),
    .Q(\pmod_1414.mem_strorage.mem[8][2] ));
 sg13g2_dfrbp_1 _1710_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net167),
    .D(_0096_),
    .Q_N(_0743_),
    .Q(\pmod_1414.mem_strorage.mem[8][3] ));
 sg13g2_dfrbp_1 _1711_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net166),
    .D(_0097_),
    .Q_N(_0742_),
    .Q(\pmod_1414.mem_strorage.mem[8][4] ));
 sg13g2_dfrbp_1 _1712_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net165),
    .D(_0098_),
    .Q_N(_0741_),
    .Q(\pmod_1414.mem_strorage.mem[8][5] ));
 sg13g2_dfrbp_1 _1713_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net164),
    .D(_0099_),
    .Q_N(_0740_),
    .Q(\pmod_1414.mem_strorage.mem[8][6] ));
 sg13g2_dfrbp_1 _1714_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net163),
    .D(net305),
    .Q_N(_0739_),
    .Q(\pmod_1414.mem_strorage.mem[0][0] ));
 sg13g2_dfrbp_1 _1715_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net162),
    .D(net313),
    .Q_N(_0738_),
    .Q(\pmod_1414.mem_strorage.mem[0][1] ));
 sg13g2_dfrbp_1 _1716_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net153),
    .D(net299),
    .Q_N(_0737_),
    .Q(\pmod_1414.mem_strorage.mem[0][2] ));
 sg13g2_dfrbp_1 _1717_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net129),
    .D(net293),
    .Q_N(_0736_),
    .Q(\pmod_1414.mem_strorage.mem[0][3] ));
 sg13g2_dfrbp_1 _1718_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net128),
    .D(net291),
    .Q_N(_0735_),
    .Q(\pmod_1414.mem_strorage.mem[0][4] ));
 sg13g2_dfrbp_1 _1719_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net127),
    .D(net307),
    .Q_N(_0734_),
    .Q(\pmod_1414.mem_strorage.mem[0][5] ));
 sg13g2_dfrbp_1 _1720_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net126),
    .D(net315),
    .Q_N(_0733_),
    .Q(\pmod_1414.mem_strorage.mem[0][6] ));
 sg13g2_dfrbp_1 _1721_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net125),
    .D(_0107_),
    .Q_N(_0732_),
    .Q(\pmod_1414.mem_strorage.mem[5][0] ));
 sg13g2_dfrbp_1 _1722_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net124),
    .D(net479),
    .Q_N(_0731_),
    .Q(\pmod_1414.mem_strorage.mem[5][1] ));
 sg13g2_dfrbp_1 _1723_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net123),
    .D(net504),
    .Q_N(_0730_),
    .Q(\pmod_1414.mem_strorage.mem[5][2] ));
 sg13g2_dfrbp_1 _1724_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net122),
    .D(net497),
    .Q_N(_0729_),
    .Q(\pmod_1414.mem_strorage.mem[5][3] ));
 sg13g2_dfrbp_1 _1725_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net121),
    .D(_0111_),
    .Q_N(_0728_),
    .Q(\pmod_1414.mem_strorage.mem[5][4] ));
 sg13g2_dfrbp_1 _1726_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net120),
    .D(net470),
    .Q_N(_0727_),
    .Q(\pmod_1414.mem_strorage.mem[5][5] ));
 sg13g2_dfrbp_1 _1727_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net119),
    .D(net474),
    .Q_N(_0726_),
    .Q(\pmod_1414.mem_strorage.mem[5][6] ));
 sg13g2_dfrbp_1 _1728_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net118),
    .D(_0114_),
    .Q_N(_0725_),
    .Q(\pmod_1414.mem_strorage.mem[6][0] ));
 sg13g2_dfrbp_1 _1729_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net117),
    .D(_0115_),
    .Q_N(_0724_),
    .Q(\pmod_1414.mem_strorage.mem[6][1] ));
 sg13g2_dfrbp_1 _1730_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net116),
    .D(_0116_),
    .Q_N(_0723_),
    .Q(\pmod_1414.mem_strorage.mem[6][2] ));
 sg13g2_dfrbp_1 _1731_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net115),
    .D(_0117_),
    .Q_N(_0722_),
    .Q(\pmod_1414.mem_strorage.mem[6][3] ));
 sg13g2_dfrbp_1 _1732_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net114),
    .D(_0118_),
    .Q_N(_0721_),
    .Q(\pmod_1414.mem_strorage.mem[6][4] ));
 sg13g2_dfrbp_1 _1733_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net112),
    .D(_0119_),
    .Q_N(_0720_),
    .Q(\pmod_1414.mem_strorage.mem[6][5] ));
 sg13g2_dfrbp_1 _1734_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net111),
    .D(_0120_),
    .Q_N(_0719_),
    .Q(\pmod_1414.mem_strorage.mem[6][6] ));
 sg13g2_dfrbp_1 _1735_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net110),
    .D(net422),
    .Q_N(_0718_),
    .Q(\pmod_1414.mem_strorage.mem[10][0] ));
 sg13g2_dfrbp_1 _1736_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net109),
    .D(net317),
    .Q_N(_0717_),
    .Q(\pmod_1414.mem_strorage.mem[10][1] ));
 sg13g2_dfrbp_1 _1737_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net108),
    .D(net350),
    .Q_N(_0716_),
    .Q(\pmod_1414.mem_strorage.mem[10][2] ));
 sg13g2_dfrbp_1 _1738_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net107),
    .D(net399),
    .Q_N(_0715_),
    .Q(\pmod_1414.mem_strorage.mem[10][3] ));
 sg13g2_dfrbp_1 _1739_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net106),
    .D(net384),
    .Q_N(_0714_),
    .Q(\pmod_1414.mem_strorage.mem[10][4] ));
 sg13g2_dfrbp_1 _1740_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net105),
    .D(net437),
    .Q_N(_0713_),
    .Q(\pmod_1414.mem_strorage.mem[10][5] ));
 sg13g2_dfrbp_1 _1741_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net104),
    .D(net374),
    .Q_N(_0712_),
    .Q(\pmod_1414.mem_strorage.mem[10][6] ));
 sg13g2_dfrbp_1 _1742_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net103),
    .D(net414),
    .Q_N(_0711_),
    .Q(\pmod_1414.mem_strorage.mem[13][0] ));
 sg13g2_dfrbp_1 _1743_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net102),
    .D(net325),
    .Q_N(_0710_),
    .Q(\pmod_1414.mem_strorage.mem[13][1] ));
 sg13g2_dfrbp_1 _1744_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net101),
    .D(net472),
    .Q_N(_0709_),
    .Q(\pmod_1414.mem_strorage.mem[13][2] ));
 sg13g2_dfrbp_1 _1745_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net100),
    .D(_0131_),
    .Q_N(_0708_),
    .Q(\pmod_1414.mem_strorage.mem[13][3] ));
 sg13g2_dfrbp_1 _1746_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net99),
    .D(net356),
    .Q_N(_0707_),
    .Q(\pmod_1414.mem_strorage.mem[13][4] ));
 sg13g2_dfrbp_1 _1747_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net98),
    .D(net460),
    .Q_N(_0706_),
    .Q(\pmod_1414.mem_strorage.mem[13][5] ));
 sg13g2_dfrbp_1 _1748_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net97),
    .D(net391),
    .Q_N(_0705_),
    .Q(\pmod_1414.mem_strorage.mem[13][6] ));
 sg13g2_dfrbp_1 _1749_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net96),
    .D(net500),
    .Q_N(_0704_),
    .Q(\pmod_1414.mem_strorage.mem[14][0] ));
 sg13g2_dfrbp_1 _1750_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net95),
    .D(_0136_),
    .Q_N(_0703_),
    .Q(\pmod_1414.mem_strorage.mem[14][1] ));
 sg13g2_dfrbp_1 _1751_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net94),
    .D(_0137_),
    .Q_N(_0702_),
    .Q(\pmod_1414.mem_strorage.mem[14][2] ));
 sg13g2_dfrbp_1 _1752_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net93),
    .D(net432),
    .Q_N(_0701_),
    .Q(\pmod_1414.mem_strorage.mem[14][3] ));
 sg13g2_dfrbp_1 _1753_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net92),
    .D(net515),
    .Q_N(_0700_),
    .Q(\pmod_1414.mem_strorage.mem[14][4] ));
 sg13g2_dfrbp_1 _1754_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net91),
    .D(net490),
    .Q_N(_0699_),
    .Q(\pmod_1414.mem_strorage.mem[14][5] ));
 sg13g2_dfrbp_1 _1755_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net90),
    .D(net416),
    .Q_N(_0698_),
    .Q(\pmod_1414.mem_strorage.mem[14][6] ));
 sg13g2_dfrbp_1 _1756_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net89),
    .D(net441),
    .Q_N(_0697_),
    .Q(\pmod_1414.mem_strorage.mem[11][0] ));
 sg13g2_dfrbp_1 _1757_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net88),
    .D(_0143_),
    .Q_N(_0696_),
    .Q(\pmod_1414.mem_strorage.mem[11][1] ));
 sg13g2_dfrbp_1 _1758_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net87),
    .D(net492),
    .Q_N(_0695_),
    .Q(\pmod_1414.mem_strorage.mem[11][2] ));
 sg13g2_dfrbp_1 _1759_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net86),
    .D(net458),
    .Q_N(_0694_),
    .Q(\pmod_1414.mem_strorage.mem[11][3] ));
 sg13g2_dfrbp_1 _1760_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net85),
    .D(_0146_),
    .Q_N(_0693_),
    .Q(\pmod_1414.mem_strorage.mem[11][4] ));
 sg13g2_dfrbp_1 _1761_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net84),
    .D(net444),
    .Q_N(_0692_),
    .Q(\pmod_1414.mem_strorage.mem[11][5] ));
 sg13g2_dfrbp_1 _1762_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net83),
    .D(net429),
    .Q_N(_0691_),
    .Q(\pmod_1414.mem_strorage.mem[11][6] ));
 sg13g2_dfrbp_1 _1763_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net82),
    .D(_0149_),
    .Q_N(_0690_),
    .Q(\pmod_1414.mem_strorage.mem[12][0] ));
 sg13g2_dfrbp_1 _1764_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net81),
    .D(_0150_),
    .Q_N(_0689_),
    .Q(\pmod_1414.mem_strorage.mem[12][1] ));
 sg13g2_dfrbp_1 _1765_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net80),
    .D(net482),
    .Q_N(_0688_),
    .Q(\pmod_1414.mem_strorage.mem[12][2] ));
 sg13g2_dfrbp_1 _1766_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net79),
    .D(net487),
    .Q_N(_0687_),
    .Q(\pmod_1414.mem_strorage.mem[12][3] ));
 sg13g2_dfrbp_1 _1767_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net78),
    .D(_0153_),
    .Q_N(_0686_),
    .Q(\pmod_1414.mem_strorage.mem[12][4] ));
 sg13g2_dfrbp_1 _1768_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net77),
    .D(_0154_),
    .Q_N(_0685_),
    .Q(\pmod_1414.mem_strorage.mem[12][5] ));
 sg13g2_dfrbp_1 _1769_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net76),
    .D(_0155_),
    .Q_N(_0684_),
    .Q(\pmod_1414.mem_strorage.mem[12][6] ));
 sg13g2_dfrbp_1 _1770_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net75),
    .D(_0156_),
    .Q_N(_0683_),
    .Q(\pmod_1414.mem_strorage.mem[15][0] ));
 sg13g2_dfrbp_1 _1771_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net74),
    .D(_0157_),
    .Q_N(_0682_),
    .Q(\pmod_1414.mem_strorage.mem[15][1] ));
 sg13g2_dfrbp_1 _1772_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net73),
    .D(_0158_),
    .Q_N(_0681_),
    .Q(\pmod_1414.mem_strorage.mem[15][2] ));
 sg13g2_dfrbp_1 _1773_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net72),
    .D(_0159_),
    .Q_N(_0680_),
    .Q(\pmod_1414.mem_strorage.mem[15][3] ));
 sg13g2_dfrbp_1 _1774_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net71),
    .D(_0160_),
    .Q_N(_0679_),
    .Q(\pmod_1414.mem_strorage.mem[15][4] ));
 sg13g2_dfrbp_1 _1775_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net70),
    .D(_0161_),
    .Q_N(_0678_),
    .Q(\pmod_1414.mem_strorage.mem[15][5] ));
 sg13g2_dfrbp_1 _1776_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net69),
    .D(_0162_),
    .Q_N(_0677_),
    .Q(\pmod_1414.mem_strorage.mem[15][6] ));
 sg13g2_dfrbp_1 _1777_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net68),
    .D(net274),
    .Q_N(_0055_),
    .Q(\pmod_1414.RX.Filter_cnt[0] ));
 sg13g2_dfrbp_1 _1778_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net67),
    .D(_0164_),
    .Q_N(_0676_),
    .Q(\pmod_1414.RX.Filter_cnt[1] ));
 sg13g2_dfrbp_1 _1779_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net130),
    .D(net495),
    .Q_N(_0784_),
    .Q(\pmod_1414.RX.RxD_bit ));
 sg13g2_dfrbp_1 _1780_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net66),
    .D(_0000_),
    .Q_N(_0675_),
    .Q(\pmod_1414.RX.RxD_data_ready ));
 sg13g2_dfrbp_1 _1781_ (.CLK(_0675_),
    .RESET_B(net1),
    .D(_0166_),
    .Q_N(_0054_),
    .Q(\pmod_1414.r_uart_rx_counter[0] ));
 sg13g2_dfrbp_1 _1782_ (.CLK(_0675_),
    .RESET_B(net1),
    .D(_0167_),
    .Q_N(_0674_),
    .Q(\pmod_1414.r_uart_rx_counter[1] ));
 sg13g2_dfrbp_1 _1783_ (.CLK(_0675_),
    .RESET_B(net1),
    .D(_0168_),
    .Q_N(_0010_),
    .Q(\pmod_1414.r_uart_rx_counter[2] ));
 sg13g2_dfrbp_1 _1784_ (.CLK(_0675_),
    .RESET_B(net1),
    .D(_0169_),
    .Q_N(_0673_),
    .Q(\pmod_1414.r_uart_rx_counter[3] ));
 sg13g2_dfrbp_1 _1785_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net60),
    .D(net361),
    .Q_N(_0672_),
    .Q(\pmod_1414.RX.RxD_data[0] ));
 sg13g2_dfrbp_1 _1786_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net59),
    .D(_0171_),
    .Q_N(_0671_),
    .Q(\pmod_1414.RX.RxD_data[1] ));
 sg13g2_dfrbp_1 _1787_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net58),
    .D(net453),
    .Q_N(_0670_),
    .Q(\pmod_1414.RX.RxD_data[2] ));
 sg13g2_dfrbp_1 _1788_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net57),
    .D(net465),
    .Q_N(_0669_),
    .Q(\pmod_1414.RX.RxD_data[3] ));
 sg13g2_dfrbp_1 _1789_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net56),
    .D(_0174_),
    .Q_N(_0668_),
    .Q(\pmod_1414.RX.RxD_data[4] ));
 sg13g2_dfrbp_1 _1790_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net55),
    .D(net463),
    .Q_N(_0667_),
    .Q(\pmod_1414.RX.RxD_data[5] ));
 sg13g2_dfrbp_1 _1791_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net54),
    .D(net467),
    .Q_N(_0666_),
    .Q(\pmod_1414.RX.RxD_data[6] ));
 sg13g2_dfrbp_1 _1792_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net53),
    .D(net519),
    .Q_N(_0665_),
    .Q(\pmod_1414.RX.RxD_data[7] ));
 sg13g2_dfrbp_1 _1793_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net52),
    .D(net266),
    .Q_N(_0053_),
    .Q(\pmod_1414.RX.OversamplingCnt[0] ));
 sg13g2_dfrbp_1 _1794_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net50),
    .D(net545),
    .Q_N(_0664_),
    .Q(\pmod_1414.RX.OversamplingCnt[1] ));
 sg13g2_dfrbp_1 _1795_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net48),
    .D(net303),
    .Q_N(_0663_),
    .Q(\pmod_1414.RX.OversamplingCnt[2] ));
 sg13g2_dfrbp_1 _1796_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net131),
    .D(_0181_),
    .Q_N(_0785_),
    .Q(\pmod_1414.RX.OversamplingCnt[3] ));
 sg13g2_dfrbp_1 _1797_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net132),
    .D(net261),
    .Q_N(_0650_),
    .Q(\pmod_1414.RX.tickgen.Acc[0] ));
 sg13g2_dfrbp_1 _1798_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net133),
    .D(net337),
    .Q_N(_0786_),
    .Q(\pmod_1414.RX.tickgen.Acc[1] ));
 sg13g2_dfrbp_1 _1799_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net134),
    .D(net542),
    .Q_N(_0787_),
    .Q(\pmod_1414.RX.tickgen.Acc[2] ));
 sg13g2_dfrbp_1 _1800_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net135),
    .D(net522),
    .Q_N(_0788_),
    .Q(\pmod_1414.RX.tickgen.Acc[3] ));
 sg13g2_dfrbp_1 _1801_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net136),
    .D(net525),
    .Q_N(_0789_),
    .Q(\pmod_1414.RX.tickgen.Acc[4] ));
 sg13g2_dfrbp_1 _1802_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net137),
    .D(net263),
    .Q_N(_0011_),
    .Q(\pmod_1414.RX.tickgen.Acc[5] ));
 sg13g2_dfrbp_1 _1803_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net138),
    .D(net426),
    .Q_N(_0790_),
    .Q(\pmod_1414.RX.tickgen.Acc[6] ));
 sg13g2_dfrbp_1 _1804_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net139),
    .D(net387),
    .Q_N(_0791_),
    .Q(\pmod_1414.RX.tickgen.Acc[7] ));
 sg13g2_dfrbp_1 _1805_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net140),
    .D(net268),
    .Q_N(_0012_),
    .Q(\pmod_1414.RX.tickgen.Acc[8] ));
 sg13g2_dfrbp_1 _1806_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net141),
    .D(net321),
    .Q_N(_0792_),
    .Q(\pmod_1414.RX.tickgen.Acc[9] ));
 sg13g2_dfrbp_1 _1807_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net142),
    .D(net358),
    .Q_N(_0793_),
    .Q(\pmod_1414.RX.tickgen.Acc[10] ));
 sg13g2_dfrbp_1 _1808_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net143),
    .D(_0040_),
    .Q_N(_0794_),
    .Q(\pmod_1414.RX.tickgen.Acc[11] ));
 sg13g2_dfrbp_1 _1809_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net144),
    .D(_0041_),
    .Q_N(_0795_),
    .Q(\pmod_1414.RX.tickgen.Acc[12] ));
 sg13g2_dfrbp_1 _1810_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net145),
    .D(_0042_),
    .Q_N(_0796_),
    .Q(\pmod_1414.RX.tickgen.Acc[13] ));
 sg13g2_dfrbp_1 _1811_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net146),
    .D(_0043_),
    .Q_N(_0797_),
    .Q(\pmod_1414.RX.tickgen.Acc[14] ));
 sg13g2_dfrbp_1 _1812_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net147),
    .D(net270),
    .Q_N(_0798_),
    .Q(\pmod_1414.RX.OversamplingTick ));
 sg13g2_dfrbp_1 _1813_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net148),
    .D(_0001_),
    .Q_N(_0799_),
    .Q(\pmod_1414.HPDL_D0 ));
 sg13g2_dfrbp_1 _1814_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net149),
    .D(_0002_),
    .Q_N(_0800_),
    .Q(\pmod_1414.HPDL_D1 ));
 sg13g2_dfrbp_1 _1815_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net150),
    .D(_0003_),
    .Q_N(_0801_),
    .Q(\pmod_1414.HPDL_D2 ));
 sg13g2_dfrbp_1 _1816_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net151),
    .D(_0004_),
    .Q_N(_0802_),
    .Q(\pmod_1414.HPDL_D3 ));
 sg13g2_dfrbp_1 _1817_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net152),
    .D(_0005_),
    .Q_N(_0803_),
    .Q(\pmod_1414.HPDL_D4 ));
 sg13g2_dfrbp_1 _1818_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net154),
    .D(_0006_),
    .Q_N(_0804_),
    .Q(\pmod_1414.HPDL_D5 ));
 sg13g2_dfrbp_1 _1819_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net46),
    .D(_0007_),
    .Q_N(_0662_),
    .Q(\pmod_1414.HPDL_D6 ));
 sg13g2_dfrbp_1 _1820_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net155),
    .D(_0182_),
    .Q_N(_0805_),
    .Q(\pmod_1414.mem_strorage.r_shift_enable ));
 sg13g2_dfrbp_1 _1821_ (.CLK(net236),
    .RESET_B(net156),
    .D(\pmod_1414.RX.RxD_data[0] ),
    .Q_N(_0806_),
    .Q(\pmod_1414.GPout[0] ));
 sg13g2_dfrbp_1 _1822_ (.CLK(net236),
    .RESET_B(net157),
    .D(\pmod_1414.RX.RxD_data[1] ),
    .Q_N(_0807_),
    .Q(\pmod_1414.GPout[1] ));
 sg13g2_dfrbp_1 _1823_ (.CLK(net236),
    .RESET_B(net158),
    .D(\pmod_1414.RX.RxD_data[2] ),
    .Q_N(_0808_),
    .Q(\pmod_1414.GPout[2] ));
 sg13g2_dfrbp_1 _1824_ (.CLK(net236),
    .RESET_B(net159),
    .D(\pmod_1414.RX.RxD_data[3] ),
    .Q_N(_0809_),
    .Q(\pmod_1414.GPout[3] ));
 sg13g2_dfrbp_1 _1825_ (.CLK(net236),
    .RESET_B(net160),
    .D(\pmod_1414.RX.RxD_data[4] ),
    .Q_N(_0810_),
    .Q(\pmod_1414.GPout[4] ));
 sg13g2_dfrbp_1 _1826_ (.CLK(net236),
    .RESET_B(net161),
    .D(\pmod_1414.RX.RxD_data[5] ),
    .Q_N(_0811_),
    .Q(\pmod_1414.GPout[5] ));
 sg13g2_dfrbp_1 _1827_ (.CLK(net235),
    .RESET_B(net169),
    .D(\pmod_1414.RX.RxD_data[6] ),
    .Q_N(_0812_),
    .Q(\pmod_1414.GPout[6] ));
 sg13g2_dfrbp_1 _1828_ (.CLK(net235),
    .RESET_B(net44),
    .D(\pmod_1414.RX.RxD_data[7] ),
    .Q_N(_0661_),
    .Q(\pmod_1414.GPout[7] ));
 sg13g2_dfrbp_1 _1829_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net42),
    .D(net395),
    .Q_N(_0660_),
    .Q(\pmod_1414.mem_strorage.mem[9][0] ));
 sg13g2_dfrbp_1 _1830_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net41),
    .D(_0184_),
    .Q_N(_0659_),
    .Q(\pmod_1414.mem_strorage.mem[9][1] ));
 sg13g2_dfrbp_1 _1831_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net65),
    .D(_0185_),
    .Q_N(_0658_),
    .Q(\pmod_1414.mem_strorage.mem[9][2] ));
 sg13g2_dfrbp_1 _1832_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net64),
    .D(net372),
    .Q_N(_0657_),
    .Q(\pmod_1414.mem_strorage.mem[9][3] ));
 sg13g2_dfrbp_1 _1833_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net63),
    .D(_0187_),
    .Q_N(_0656_),
    .Q(\pmod_1414.mem_strorage.mem[9][4] ));
 sg13g2_dfrbp_1 _1834_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net62),
    .D(net397),
    .Q_N(_0655_),
    .Q(\pmod_1414.mem_strorage.mem[9][5] ));
 sg13g2_dfrbp_1 _1835_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net170),
    .D(_0189_),
    .Q_N(_0813_),
    .Q(\pmod_1414.mem_strorage.mem[9][6] ));
 sg13g2_dfrbp_1 _1836_ (.CLK(net233),
    .RESET_B(net1),
    .D(\pmod_1414.HPDL_A0 ),
    .Q_N(\pmod_1414.HPDL_A0 ),
    .Q(\pmod_1414.r_address_counter[0] ));
 sg13g2_dfrbp_1 _1837_ (.CLK(net233),
    .RESET_B(net1),
    .D(_0035_),
    .Q_N(\pmod_1414.HPDL_A1 ),
    .Q(\pmod_1414.r_address_counter[1] ));
 sg13g2_dfrbp_1 _1838_ (.CLK(\pmod_1414.r_counter[10] ),
    .RESET_B(net1),
    .D(_0036_),
    .Q_N(_0008_),
    .Q(\pmod_1414.r_address_counter[2] ));
 sg13g2_dfrbp_1 _1839_ (.CLK(\pmod_1414.r_counter[10] ),
    .RESET_B(net1),
    .D(_0037_),
    .Q_N(_0814_),
    .Q(\pmod_1414.r_address_counter[3] ));
 sg13g2_dfrbp_1 _1840_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net171),
    .D(net260),
    .Q_N(_0649_),
    .Q(\pmod_1414.r_counter[0] ));
 sg13g2_dfrbp_1 _1841_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net172),
    .D(net456),
    .Q_N(_0815_),
    .Q(\pmod_1414.r_counter[1] ));
 sg13g2_dfrbp_1 _1842_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net173),
    .D(net548),
    .Q_N(_0816_),
    .Q(\pmod_1414.r_counter[2] ));
 sg13g2_dfrbp_1 _1843_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net174),
    .D(net342),
    .Q_N(_0817_),
    .Q(\pmod_1414.r_counter[3] ));
 sg13g2_dfrbp_1 _1844_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net175),
    .D(net323),
    .Q_N(_0818_),
    .Q(\pmod_1414.r_counter[4] ));
 sg13g2_dfrbp_1 _1845_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net176),
    .D(net551),
    .Q_N(_0819_),
    .Q(\pmod_1414.r_counter[5] ));
 sg13g2_dfrbp_1 _1846_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net177),
    .D(net401),
    .Q_N(_0820_),
    .Q(\pmod_1414.r_counter[6] ));
 sg13g2_dfrbp_1 _1847_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net178),
    .D(net289),
    .Q_N(_0821_),
    .Q(\pmod_1414.r_counter[7] ));
 sg13g2_dfrbp_1 _1848_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net179),
    .D(net380),
    .Q_N(_0822_),
    .Q(\pmod_1414.r_counter[8] ));
 sg13g2_dfrbp_1 _1849_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net237),
    .D(net370),
    .Q_N(_0823_),
    .Q(\pmod_1414.r_counter[9] ));
 sg13g2_dfrbp_1 _1850_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net238),
    .D(_0013_),
    .Q_N(_0824_),
    .Q(\pmod_1414.r_counter[10] ));
 sg13g2_dfrbp_1 _1851_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net239),
    .D(net301),
    .Q_N(_0825_),
    .Q(\pmod_1414.r_counter[11] ));
 sg13g2_dfrbp_1 _1852_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net240),
    .D(_0015_),
    .Q_N(_0826_),
    .Q(\pmod_1414.r_counter[12] ));
 sg13g2_dfrbp_1 _1853_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net241),
    .D(net280),
    .Q_N(_0827_),
    .Q(\pmod_1414.r_counter[13] ));
 sg13g2_dfrbp_1 _1854_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net242),
    .D(net410),
    .Q_N(_0828_),
    .Q(\pmod_1414.r_counter[14] ));
 sg13g2_dfrbp_1 _1855_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net243),
    .D(net283),
    .Q_N(_0829_),
    .Q(\pmod_1414.r_counter[15] ));
 sg13g2_dfrbp_1 _1856_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net244),
    .D(_0019_),
    .Q_N(_0830_),
    .Q(\pmod_1414.r_counter[16] ));
 sg13g2_dfrbp_1 _1857_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net245),
    .D(net311),
    .Q_N(_0831_),
    .Q(\pmod_1414.r_counter[17] ));
 sg13g2_dfrbp_1 _1858_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net246),
    .D(net419),
    .Q_N(_0832_),
    .Q(\pmod_1414.r_counter[18] ));
 sg13g2_dfrbp_1 _1859_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net247),
    .D(net286),
    .Q_N(_0833_),
    .Q(\pmod_1414.r_counter[19] ));
 sg13g2_dfrbp_1 _1860_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net248),
    .D(net378),
    .Q_N(_0834_),
    .Q(\pmod_1414.r_counter[20] ));
 sg13g2_dfrbp_1 _1861_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net49),
    .D(net277),
    .Q_N(_0835_),
    .Q(\pmod_1414.r_counter[21] ));
 sg13g2_dfrbp_1 _1862_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net61),
    .D(net272),
    .Q_N(_0009_),
    .Q(\pmod_1414.mem_strorage.i_w_caret_strobe ));
 sg13g2_dfrbp_1 _1863_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net51),
    .D(net537),
    .Q_N(_0654_),
    .Q(\pmod_1414.RX.RxD_state[3] ));
 sg13g2_dfrbp_1 _1864_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net47),
    .D(net527),
    .Q_N(_0653_),
    .Q(\pmod_1414.RX.RxD_state[2] ));
 sg13g2_dfrbp_1 _1865_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net43),
    .D(_0192_),
    .Q_N(_0652_),
    .Q(\pmod_1414.RX.RxD_state[1] ));
 sg13g2_dfrbp_1 _1866_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net45),
    .D(_0193_),
    .Q_N(_0651_),
    .Q(\pmod_1414.RX.RxD_state[0] ));
 sg13g2_tiehi _1703__8 (.L_HI(net8));
 sg13g2_tiehi _1702__9 (.L_HI(net9));
 sg13g2_tiehi _1701__10 (.L_HI(net10));
 sg13g2_tiehi _1700__11 (.L_HI(net11));
 sg13g2_tiehi _1699__12 (.L_HI(net12));
 sg13g2_tiehi _1698__13 (.L_HI(net13));
 sg13g2_tiehi _1697__14 (.L_HI(net14));
 sg13g2_tiehi _1696__15 (.L_HI(net15));
 sg13g2_tiehi _1695__16 (.L_HI(net16));
 sg13g2_tiehi _1694__17 (.L_HI(net17));
 sg13g2_tiehi _1693__18 (.L_HI(net18));
 sg13g2_tiehi _1692__19 (.L_HI(net19));
 sg13g2_tiehi _1691__20 (.L_HI(net20));
 sg13g2_tiehi _1690__21 (.L_HI(net21));
 sg13g2_tiehi _1689__22 (.L_HI(net22));
 sg13g2_tiehi _1688__23 (.L_HI(net23));
 sg13g2_tiehi _1687__24 (.L_HI(net24));
 sg13g2_tiehi _1686__25 (.L_HI(net25));
 sg13g2_tiehi _1685__26 (.L_HI(net26));
 sg13g2_tiehi _1684__27 (.L_HI(net27));
 sg13g2_tiehi _1683__28 (.L_HI(net28));
 sg13g2_tiehi _1682__29 (.L_HI(net29));
 sg13g2_tiehi _1681__30 (.L_HI(net30));
 sg13g2_tiehi _1680__31 (.L_HI(net31));
 sg13g2_tiehi _1679__32 (.L_HI(net32));
 sg13g2_tiehi _1678__33 (.L_HI(net33));
 sg13g2_tiehi _1677__34 (.L_HI(net34));
 sg13g2_tiehi _1676__35 (.L_HI(net35));
 sg13g2_tiehi _1675__36 (.L_HI(net36));
 sg13g2_tiehi _1674__37 (.L_HI(net37));
 sg13g2_tiehi _1673__38 (.L_HI(net38));
 sg13g2_tiehi _1672__39 (.L_HI(net39));
 sg13g2_tiehi _1671__40 (.L_HI(net40));
 sg13g2_tiehi _1830__41 (.L_HI(net41));
 sg13g2_tiehi _1829__42 (.L_HI(net42));
 sg13g2_tiehi _1865__43 (.L_HI(net43));
 sg13g2_tiehi _1828__44 (.L_HI(net44));
 sg13g2_tiehi _1866__45 (.L_HI(net45));
 sg13g2_tiehi _1819__46 (.L_HI(net46));
 sg13g2_tiehi _1864__47 (.L_HI(net47));
 sg13g2_tiehi _1795__48 (.L_HI(net48));
 sg13g2_tiehi _1861__49 (.L_HI(net49));
 sg13g2_tiehi _1794__50 (.L_HI(net50));
 sg13g2_tiehi _1863__51 (.L_HI(net51));
 sg13g2_tiehi _1793__52 (.L_HI(net52));
 sg13g2_tiehi _1792__53 (.L_HI(net53));
 sg13g2_tiehi _1791__54 (.L_HI(net54));
 sg13g2_tiehi _1790__55 (.L_HI(net55));
 sg13g2_tiehi _1789__56 (.L_HI(net56));
 sg13g2_tiehi _1788__57 (.L_HI(net57));
 sg13g2_tiehi _1787__58 (.L_HI(net58));
 sg13g2_tiehi _1786__59 (.L_HI(net59));
 sg13g2_tiehi _1785__60 (.L_HI(net60));
 sg13g2_tiehi _1862__61 (.L_HI(net61));
 sg13g2_tiehi _1834__62 (.L_HI(net62));
 sg13g2_tiehi _1833__63 (.L_HI(net63));
 sg13g2_tiehi _1832__64 (.L_HI(net64));
 sg13g2_tiehi _1831__65 (.L_HI(net65));
 sg13g2_tiehi _1780__66 (.L_HI(net66));
 sg13g2_tiehi _1778__67 (.L_HI(net67));
 sg13g2_tiehi _1777__68 (.L_HI(net68));
 sg13g2_tiehi _1776__69 (.L_HI(net69));
 sg13g2_tiehi _1775__70 (.L_HI(net70));
 sg13g2_tiehi _1774__71 (.L_HI(net71));
 sg13g2_tiehi _1773__72 (.L_HI(net72));
 sg13g2_tiehi _1772__73 (.L_HI(net73));
 sg13g2_tiehi _1771__74 (.L_HI(net74));
 sg13g2_tiehi _1770__75 (.L_HI(net75));
 sg13g2_tiehi _1769__76 (.L_HI(net76));
 sg13g2_tiehi _1768__77 (.L_HI(net77));
 sg13g2_tiehi _1767__78 (.L_HI(net78));
 sg13g2_tiehi _1766__79 (.L_HI(net79));
 sg13g2_tiehi _1765__80 (.L_HI(net80));
 sg13g2_tiehi _1764__81 (.L_HI(net81));
 sg13g2_tiehi _1763__82 (.L_HI(net82));
 sg13g2_tiehi _1762__83 (.L_HI(net83));
 sg13g2_tiehi _1761__84 (.L_HI(net84));
 sg13g2_tiehi _1760__85 (.L_HI(net85));
 sg13g2_tiehi _1759__86 (.L_HI(net86));
 sg13g2_tiehi _1758__87 (.L_HI(net87));
 sg13g2_tiehi _1757__88 (.L_HI(net88));
 sg13g2_tiehi _1756__89 (.L_HI(net89));
 sg13g2_tiehi _1755__90 (.L_HI(net90));
 sg13g2_tiehi _1754__91 (.L_HI(net91));
 sg13g2_tiehi _1753__92 (.L_HI(net92));
 sg13g2_tiehi _1752__93 (.L_HI(net93));
 sg13g2_tiehi _1751__94 (.L_HI(net94));
 sg13g2_tiehi _1750__95 (.L_HI(net95));
 sg13g2_tiehi _1749__96 (.L_HI(net96));
 sg13g2_tiehi _1748__97 (.L_HI(net97));
 sg13g2_tiehi _1747__98 (.L_HI(net98));
 sg13g2_tiehi _1746__99 (.L_HI(net99));
 sg13g2_tiehi _1745__100 (.L_HI(net100));
 sg13g2_tiehi _1744__101 (.L_HI(net101));
 sg13g2_tiehi _1743__102 (.L_HI(net102));
 sg13g2_tiehi _1742__103 (.L_HI(net103));
 sg13g2_tiehi _1741__104 (.L_HI(net104));
 sg13g2_tiehi _1740__105 (.L_HI(net105));
 sg13g2_tiehi _1739__106 (.L_HI(net106));
 sg13g2_tiehi _1738__107 (.L_HI(net107));
 sg13g2_tiehi _1737__108 (.L_HI(net108));
 sg13g2_tiehi _1736__109 (.L_HI(net109));
 sg13g2_tiehi _1735__110 (.L_HI(net110));
 sg13g2_tiehi _1734__111 (.L_HI(net111));
 sg13g2_tiehi _1733__112 (.L_HI(net112));
 sg13g2_tiehi _1670__113 (.L_HI(net113));
 sg13g2_tiehi _1732__114 (.L_HI(net114));
 sg13g2_tiehi _1731__115 (.L_HI(net115));
 sg13g2_tiehi _1730__116 (.L_HI(net116));
 sg13g2_tiehi _1729__117 (.L_HI(net117));
 sg13g2_tiehi _1728__118 (.L_HI(net118));
 sg13g2_tiehi _1727__119 (.L_HI(net119));
 sg13g2_tiehi _1726__120 (.L_HI(net120));
 sg13g2_tiehi _1725__121 (.L_HI(net121));
 sg13g2_tiehi _1724__122 (.L_HI(net122));
 sg13g2_tiehi _1723__123 (.L_HI(net123));
 sg13g2_tiehi _1722__124 (.L_HI(net124));
 sg13g2_tiehi _1721__125 (.L_HI(net125));
 sg13g2_tiehi _1720__126 (.L_HI(net126));
 sg13g2_tiehi _1719__127 (.L_HI(net127));
 sg13g2_tiehi _1718__128 (.L_HI(net128));
 sg13g2_tiehi _1717__129 (.L_HI(net129));
 sg13g2_tiehi _1779__130 (.L_HI(net130));
 sg13g2_tiehi _1796__131 (.L_HI(net131));
 sg13g2_tiehi _1797__132 (.L_HI(net132));
 sg13g2_tiehi _1798__133 (.L_HI(net133));
 sg13g2_tiehi _1799__134 (.L_HI(net134));
 sg13g2_tiehi _1800__135 (.L_HI(net135));
 sg13g2_tiehi _1801__136 (.L_HI(net136));
 sg13g2_tiehi _1802__137 (.L_HI(net137));
 sg13g2_tiehi _1803__138 (.L_HI(net138));
 sg13g2_tiehi _1804__139 (.L_HI(net139));
 sg13g2_tiehi _1805__140 (.L_HI(net140));
 sg13g2_tiehi _1806__141 (.L_HI(net141));
 sg13g2_tiehi _1807__142 (.L_HI(net142));
 sg13g2_tiehi _1808__143 (.L_HI(net143));
 sg13g2_tiehi _1809__144 (.L_HI(net144));
 sg13g2_tiehi _1810__145 (.L_HI(net145));
 sg13g2_tiehi _1811__146 (.L_HI(net146));
 sg13g2_tiehi _1812__147 (.L_HI(net147));
 sg13g2_tiehi _1813__148 (.L_HI(net148));
 sg13g2_tiehi _1814__149 (.L_HI(net149));
 sg13g2_tiehi _1815__150 (.L_HI(net150));
 sg13g2_tiehi _1816__151 (.L_HI(net151));
 sg13g2_tiehi _1817__152 (.L_HI(net152));
 sg13g2_tiehi _1716__153 (.L_HI(net153));
 sg13g2_tiehi _1818__154 (.L_HI(net154));
 sg13g2_tiehi _1820__155 (.L_HI(net155));
 sg13g2_tiehi _1821__156 (.L_HI(net156));
 sg13g2_tiehi _1822__157 (.L_HI(net157));
 sg13g2_tiehi _1823__158 (.L_HI(net158));
 sg13g2_tiehi _1824__159 (.L_HI(net159));
 sg13g2_tiehi _1825__160 (.L_HI(net160));
 sg13g2_tiehi _1826__161 (.L_HI(net161));
 sg13g2_tiehi _1715__162 (.L_HI(net162));
 sg13g2_tiehi _1714__163 (.L_HI(net163));
 sg13g2_tiehi _1713__164 (.L_HI(net164));
 sg13g2_tiehi _1712__165 (.L_HI(net165));
 sg13g2_tiehi _1711__166 (.L_HI(net166));
 sg13g2_tiehi _1710__167 (.L_HI(net167));
 sg13g2_tiehi _1709__168 (.L_HI(net168));
 sg13g2_tiehi _1827__169 (.L_HI(net169));
 sg13g2_tiehi _1835__170 (.L_HI(net170));
 sg13g2_tiehi _1840__171 (.L_HI(net171));
 sg13g2_tiehi _1841__172 (.L_HI(net172));
 sg13g2_tiehi _1842__173 (.L_HI(net173));
 sg13g2_tiehi _1843__174 (.L_HI(net174));
 sg13g2_tiehi _1844__175 (.L_HI(net175));
 sg13g2_tiehi _1845__176 (.L_HI(net176));
 sg13g2_tiehi _1846__177 (.L_HI(net177));
 sg13g2_tiehi _1847__178 (.L_HI(net178));
 sg13g2_tiehi _1848__179 (.L_HI(net179));
 sg13g2_tiehi _1849__180 (.L_HI(net237));
 sg13g2_tiehi _1850__181 (.L_HI(net238));
 sg13g2_tiehi _1851__182 (.L_HI(net239));
 sg13g2_tiehi _1852__183 (.L_HI(net240));
 sg13g2_tiehi _1853__184 (.L_HI(net241));
 sg13g2_tiehi _1854__185 (.L_HI(net242));
 sg13g2_tiehi _1855__186 (.L_HI(net243));
 sg13g2_tiehi _1856__187 (.L_HI(net244));
 sg13g2_tiehi _1857__188 (.L_HI(net245));
 sg13g2_tiehi _1858__189 (.L_HI(net246));
 sg13g2_tiehi _1859__190 (.L_HI(net247));
 sg13g2_tiehi _1860__191 (.L_HI(net248));
 sg13g2_tiehi _1708__192 (.L_HI(net249));
 sg13g2_tiehi _1707__193 (.L_HI(net250));
 sg13g2_tiehi _1706__194 (.L_HI(net251));
 sg13g2_tiehi _1705__195 (.L_HI(net252));
 sg13g2_tiehi tt_um_hpdl1414_uart_atudoroi_196 (.L_HI(net253));
 sg13g2_tiehi tt_um_hpdl1414_uart_atudoroi_197 (.L_HI(net254));
 sg13g2_tiehi tt_um_hpdl1414_uart_atudoroi_198 (.L_HI(net255));
 sg13g2_tiehi tt_um_hpdl1414_uart_atudoroi_199 (.L_HI(net256));
 sg13g2_tiehi tt_um_hpdl1414_uart_atudoroi_200 (.L_HI(net257));
 sg13g2_tiehi tt_um_hpdl1414_uart_atudoroi_201 (.L_HI(net258));
 sg13g2_tiehi tt_um_hpdl1414_uart_atudoroi_202 (.L_HI(net259));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_hpdl1414_uart_atudoroi_4 (.L_LO(net4));
 sg13g2_tielo tt_um_hpdl1414_uart_atudoroi_5 (.L_LO(net5));
 sg13g2_tielo tt_um_hpdl1414_uart_atudoroi_6 (.L_LO(net6));
 sg13g2_tiehi _1704__7 (.L_HI(net7));
 sg13g2_buf_1 _2067_ (.A(\pmod_1414.HPDL_A0 ),
    .X(uio_out[0]));
 sg13g2_buf_1 _2068_ (.A(\pmod_1414.HPDL_A1 ),
    .X(uio_out[1]));
 sg13g2_buf_1 _2069_ (.A(\pmod_1414.HPDL_WR1 ),
    .X(uio_out[2]));
 sg13g2_buf_1 _2070_ (.A(\pmod_1414.HPDL_WR2 ),
    .X(uio_out[3]));
 sg13g2_buf_1 _2071_ (.A(\pmod_1414.HPDL_WR3 ),
    .X(uio_out[4]));
 sg13g2_buf_1 _2072_ (.A(\pmod_1414.HPDL_WR4 ),
    .X(uio_out[5]));
 sg13g2_buf_1 _2073_ (.A(\pmod_1414.HPDL_D0 ),
    .X(uo_out[0]));
 sg13g2_buf_1 _2074_ (.A(\pmod_1414.HPDL_D1 ),
    .X(uo_out[1]));
 sg13g2_buf_1 _2075_ (.A(\pmod_1414.HPDL_D2 ),
    .X(uo_out[2]));
 sg13g2_buf_1 _2076_ (.A(\pmod_1414.HPDL_D3 ),
    .X(uo_out[3]));
 sg13g2_buf_1 _2077_ (.A(\pmod_1414.HPDL_D4 ),
    .X(uo_out[4]));
 sg13g2_buf_1 _2078_ (.A(\pmod_1414.HPDL_D5 ),
    .X(uo_out[5]));
 sg13g2_buf_1 _2079_ (.A(\pmod_1414.HPDL_D6 ),
    .X(uo_out[6]));
 sg13g2_buf_2 fanout180 (.A(net181),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_0397_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(net183),
    .X(net182));
 sg13g2_buf_4 fanout183 (.X(net183),
    .A(_0397_));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(net186));
 sg13g2_buf_1 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(net189),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(net188),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(net189),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_0396_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(net192),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(net192),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_0396_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(net199),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(net199),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(net199),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(net197),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(net198),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(net199),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_0396_),
    .X(net199));
 sg13g2_buf_4 fanout200 (.X(net200),
    .A(_0635_));
 sg13g2_buf_4 fanout201 (.X(net201),
    .A(_0395_));
 sg13g2_buf_2 fanout202 (.A(_0254_),
    .X(net202));
 sg13g2_buf_4 fanout203 (.X(net203),
    .A(net205));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(net205));
 sg13g2_buf_4 fanout205 (.X(net205),
    .A(\pmod_1414.r_address_counter[1] ));
 sg13g2_buf_4 fanout206 (.X(net206),
    .A(net207));
 sg13g2_buf_4 fanout207 (.X(net207),
    .A(\pmod_1414.r_address_counter[1] ));
 sg13g2_buf_8 fanout208 (.A(net209),
    .X(net208));
 sg13g2_buf_8 fanout209 (.A(\pmod_1414.r_address_counter[0] ),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(\pmod_1414.r_address_counter[0] ),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(net212),
    .X(net211));
 sg13g2_buf_1 fanout212 (.A(net215),
    .X(net212));
 sg13g2_buf_4 fanout213 (.X(net213),
    .A(net215));
 sg13g2_buf_2 fanout214 (.A(net215),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(\pmod_1414.r_address_counter[0] ),
    .X(net215));
 sg13g2_buf_4 fanout216 (.X(net216),
    .A(\pmod_1414.GPout[6] ));
 sg13g2_buf_4 fanout217 (.X(net217),
    .A(\pmod_1414.GPout[6] ));
 sg13g2_buf_4 fanout218 (.X(net218),
    .A(\pmod_1414.GPout[5] ));
 sg13g2_buf_4 fanout219 (.X(net219),
    .A(\pmod_1414.GPout[5] ));
 sg13g2_buf_4 fanout220 (.X(net220),
    .A(net221));
 sg13g2_buf_4 fanout221 (.X(net221),
    .A(\pmod_1414.GPout[4] ));
 sg13g2_buf_4 fanout222 (.X(net222),
    .A(net223));
 sg13g2_buf_4 fanout223 (.X(net223),
    .A(\pmod_1414.GPout[3] ));
 sg13g2_buf_4 fanout224 (.X(net224),
    .A(net225));
 sg13g2_buf_4 fanout225 (.X(net225),
    .A(\pmod_1414.GPout[2] ));
 sg13g2_buf_4 fanout226 (.X(net226),
    .A(net227));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(\pmod_1414.GPout[1] ));
 sg13g2_buf_4 fanout228 (.X(net228),
    .A(net229));
 sg13g2_buf_2 fanout229 (.A(net230),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(\pmod_1414.GPout[0] ),
    .X(net230));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(\pmod_1414.r_uart_rx_counter[1] ));
 sg13g2_buf_4 fanout232 (.X(net232),
    .A(\pmod_1414.r_uart_rx_counter[0] ));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(\pmod_1414.r_counter[10] ));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(\pmod_1414.RX.OversamplingTick ));
 sg13g2_buf_2 fanout235 (.A(net236),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(\pmod_1414.RX.RxD_data_ready ),
    .X(net236));
 sg13g2_buf_8 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(uio_in[3]),
    .X(net2));
 sg13g2_tielo tt_um_hpdl1414_uart_atudoroi_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0649_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0650_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0011_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0048_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0053_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0641_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0178_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0012_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0051_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold10 (.A(\pmod_1414.RX.tickgen.Acc[14] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0038_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold12 (.A(\pmod_1414.mem_strorage.i_w_caret_strobe ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0026_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0055_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0163_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold16 (.A(\pmod_1414.r_counter[21] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0373_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0025_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold19 (.A(\pmod_1414.r_counter[13] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0363_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0016_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold22 (.A(\pmod_1414.r_counter[15] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0366_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0018_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold25 (.A(\pmod_1414.r_counter[19] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0371_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0022_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold28 (.A(\pmod_1414.r_counter[7] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0356_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0032_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold31 (.A(\pmod_1414.mem_strorage.mem[0][4] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0104_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold33 (.A(\pmod_1414.mem_strorage.mem[0][3] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0103_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold35 (.A(\pmod_1414.mem_strorage.mem[8][1] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0094_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold37 (.A(\pmod_1414.RX.tickgen.Acc[13] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0388_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold39 (.A(\pmod_1414.mem_strorage.mem[0][2] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0102_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold41 (.A(\pmod_1414.r_counter[11] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0014_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold43 (.A(\pmod_1414.RX.OversamplingCnt[2] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0180_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold45 (.A(\pmod_1414.mem_strorage.mem[0][0] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0100_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold47 (.A(\pmod_1414.mem_strorage.mem[0][5] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0105_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold49 (.A(\pmod_1414.RX.OversamplingCnt[3] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold50 (.A(\pmod_1414.r_counter[17] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0368_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0020_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold53 (.A(\pmod_1414.mem_strorage.mem[0][1] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0101_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold55 (.A(\pmod_1414.mem_strorage.mem[0][6] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0106_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold57 (.A(\pmod_1414.mem_strorage.mem[10][1] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0122_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold59 (.A(\pmod_1414.mem_strorage.mem[4][0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0079_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold61 (.A(\pmod_1414.RX.tickgen.Acc[9] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0052_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold63 (.A(\pmod_1414.r_counter[4] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0029_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold65 (.A(\pmod_1414.mem_strorage.mem[13][1] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0129_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold67 (.A(\pmod_1414.mem_strorage.mem[3][2] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0074_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold69 (.A(\pmod_1414.mem_strorage.mem[1][1] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0059_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold71 (.A(\pmod_1414.mem_strorage.mem[4][2] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0081_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold73 (.A(\pmod_1414.mem_strorage.mem[1][0] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0058_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold75 (.A(\pmod_1414.mem_strorage.mem[3][4] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0076_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold77 (.A(\pmod_1414.RX.tickgen.Acc[1] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0044_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold79 (.A(\pmod_1414.mem_strorage.mem[3][0] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold80 (.A(\pmod_1414.mem_strorage.mem[3][6] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0078_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold82 (.A(\pmod_1414.r_counter[3] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0028_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold84 (.A(\pmod_1414.mem_strorage.mem[4][6] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0085_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold86 (.A(\pmod_1414.mem_strorage.mem[3][3] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0075_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold88 (.A(\pmod_1414.mem_strorage.mem[4][4] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0083_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold90 (.A(\pmod_1414.mem_strorage.mem[10][2] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0123_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold92 (.A(\pmod_1414.mem_strorage.mem[3][1] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0073_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold94 (.A(\pmod_1414.mem_strorage.mem[4][1] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0080_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold96 (.A(\pmod_1414.mem_strorage.mem[13][4] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0132_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold98 (.A(\pmod_1414.RX.tickgen.Acc[10] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0039_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold100 (.A(\pmod_1414.mem_strorage.mem[12][1] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold101 (.A(\pmod_1414.RX.RxD_data[0] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0170_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold103 (.A(\pmod_1414.mem_strorage.mem[3][5] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0077_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold105 (.A(\pmod_1414.mem_strorage.mem[1][3] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0061_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold107 (.A(\pmod_1414.mem_strorage.mem[2][3] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold108 (.A(\pmod_1414.mem_strorage.mem[4][5] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0084_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold110 (.A(\pmod_1414.r_counter[9] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0034_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold112 (.A(\pmod_1414.mem_strorage.mem[9][3] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0186_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold114 (.A(\pmod_1414.mem_strorage.mem[10][6] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0127_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold116 (.A(\pmod_1414.mem_strorage.mem[1][2] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0060_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold118 (.A(\pmod_1414.r_counter[20] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0024_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold120 (.A(\pmod_1414.r_counter[8] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0033_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold122 (.A(\pmod_1414.mem_strorage.mem[8][0] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0093_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold124 (.A(\pmod_1414.mem_strorage.mem[10][4] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0125_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold126 (.A(\pmod_1414.mem_strorage.mem[12][4] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold127 (.A(\pmod_1414.RX.tickgen.Acc[7] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0050_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold129 (.A(\pmod_1414.mem_strorage.mem[1][5] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0063_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold131 (.A(\pmod_1414.mem_strorage.mem[13][6] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0134_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold133 (.A(\pmod_1414.mem_strorage.mem[1][6] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0064_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold135 (.A(\pmod_1414.mem_strorage.mem[9][0] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0183_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold137 (.A(\pmod_1414.mem_strorage.mem[9][5] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0188_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold139 (.A(\pmod_1414.mem_strorage.mem[10][3] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0124_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold141 (.A(\pmod_1414.r_counter[6] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0031_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold143 (.A(\pmod_1414.mem_strorage.mem[2][4] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold144 (.A(\pmod_1414.mem_strorage.mem[9][4] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold145 (.A(\pmod_1414.mem_strorage.mem[1][4] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold146 (.A(\pmod_1414.mem_strorage.mem[4][3] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0082_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold148 (.A(\pmod_1414.mem_strorage.mem[2][6] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold149 (.A(\pmod_1414.mem_strorage.mem[2][2] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold150 (.A(\pmod_1414.r_counter[14] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0017_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold152 (.A(\pmod_1414.mem_strorage.mem[7][4] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0090_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold154 (.A(\pmod_1414.mem_strorage.mem[13][0] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0128_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold156 (.A(\pmod_1414.mem_strorage.mem[14][6] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0141_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold158 (.A(\pmod_1414.mem_strorage.mem[2][1] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold159 (.A(\pmod_1414.r_counter[18] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0021_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold161 (.A(\pmod_1414.mem_strorage.mem[9][1] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold162 (.A(\pmod_1414.mem_strorage.mem[10][0] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0121_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold164 (.A(\pmod_1414.mem_strorage.mem[7][0] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold165 (.A(\pmod_1414.mem_strorage.mem[9][6] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold166 (.A(\pmod_1414.RX.tickgen.Acc[6] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0049_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold168 (.A(\pmod_1414.mem_strorage.mem[2][5] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold169 (.A(\pmod_1414.mem_strorage.mem[11][6] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0148_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold171 (.A(\pmod_1414.mem_strorage.mem[2][0] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold172 (.A(\pmod_1414.mem_strorage.mem[14][3] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0138_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold174 (.A(\pmod_1414.r_counter[12] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold175 (.A(\pmod_1414.mem_strorage.mem[7][5] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0091_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold177 (.A(\pmod_1414.mem_strorage.mem[10][5] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0126_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold179 (.A(\pmod_1414.mem_strorage.mem[12][6] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold180 (.A(\pmod_1414.RX.RxD_sync[0] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold181 (.A(\pmod_1414.mem_strorage.mem[11][0] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0142_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold183 (.A(\pmod_1414.mem_strorage.mem[8][3] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold184 (.A(\pmod_1414.mem_strorage.mem[11][5] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0147_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold186 (.A(\pmod_1414.r_counter[16] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold187 (.A(\pmod_1414.mem_strorage.mem[11][4] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold188 (.A(\pmod_1414.mem_strorage.mem[7][2] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0088_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold190 (.A(\pmod_1414.mem_strorage.mem[8][4] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold191 (.A(\pmod_1414.mem_strorage.mem[11][1] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold192 (.A(\pmod_1414.mem_strorage.mem[9][2] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold193 (.A(\pmod_1414.RX.RxD_data[2] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0172_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold195 (.A(\pmod_1414.RX.RxD_sync[1] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold196 (.A(\pmod_1414.r_counter[1] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0023_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold198 (.A(\pmod_1414.mem_strorage.mem[11][3] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0145_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold200 (.A(\pmod_1414.mem_strorage.mem[13][5] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0133_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold202 (.A(\pmod_1414.RX.RxD_data[1] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold203 (.A(\pmod_1414.RX.RxD_data[5] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0175_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold205 (.A(\pmod_1414.RX.RxD_data[3] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0173_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold207 (.A(\pmod_1414.RX.RxD_data[6] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0176_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold209 (.A(\pmod_1414.RX.Filter_cnt[1] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold210 (.A(\pmod_1414.mem_strorage.mem[6][5] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0112_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold212 (.A(\pmod_1414.mem_strorage.mem[14][2] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0130_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold214 (.A(\pmod_1414.mem_strorage.mem[5][6] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0113_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold216 (.A(\pmod_1414.mem_strorage.mem[15][1] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold217 (.A(\pmod_1414.mem_strorage.mem[7][6] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0092_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold219 (.A(\pmod_1414.mem_strorage.mem[5][1] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0108_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold221 (.A(\pmod_1414.mem_strorage.mem[12][0] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold222 (.A(\pmod_1414.mem_strorage.mem[13][2] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0151_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold224 (.A(\pmod_1414.mem_strorage.mem[6][4] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold225 (.A(\pmod_1414.mem_strorage.mem[8][5] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold226 (.A(\pmod_1414.RX.RxD_data[4] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold227 (.A(\pmod_1414.mem_strorage.mem[12][3] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0152_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold229 (.A(\pmod_1414.mem_strorage.mem[14][1] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold230 (.A(\pmod_1414.mem_strorage.mem[14][5] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0140_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold232 (.A(\pmod_1414.mem_strorage.mem[11][2] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0144_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold234 (.A(\pmod_1414.RX.Filter_cnt[0] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0632_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0165_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold237 (.A(\pmod_1414.mem_strorage.mem[5][3] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0110_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold239 (.A(\pmod_1414.mem_strorage.mem[8][2] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold240 (.A(\pmod_1414.mem_strorage.mem[14][0] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0135_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold242 (.A(\pmod_1414.mem_strorage.mem[8][6] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold243 (.A(\pmod_1414.mem_strorage.r_shift_enable ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold244 (.A(\pmod_1414.mem_strorage.mem[5][2] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0109_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold246 (.A(\pmod_1414.mem_strorage.mem[13][3] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold247 (.A(\pmod_1414.mem_strorage.mem[7][3] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold248 (.A(\pmod_1414.mem_strorage.mem[6][0] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold249 (.A(\pmod_1414.RX.RxD_state[1] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0273_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold251 (.A(\pmod_1414.mem_strorage.mem[12][5] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold252 (.A(\pmod_1414.mem_strorage.mem[15][2] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold253 (.A(\pmod_1414.mem_strorage.mem[7][1] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold254 (.A(\pmod_1414.mem_strorage.mem[5][0] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold255 (.A(\pmod_1414.mem_strorage.mem[14][4] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0139_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold257 (.A(\pmod_1414.mem_strorage.mem[6][2] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold258 (.A(\pmod_1414.mem_strorage.mem[5][4] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold259 (.A(\pmod_1414.RX.RxD_data[7] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0177_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold261 (.A(\pmod_1414.mem_strorage.mem[6][3] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold262 (.A(\pmod_1414.RX.tickgen.Acc[3] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0046_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold264 (.A(\pmod_1414.mem_strorage.mem[6][6] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold265 (.A(\pmod_1414.RX.tickgen.Acc[4] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0047_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold267 (.A(\pmod_1414.RX.RxD_state[2] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0191_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold269 (.A(\pmod_1414.mem_strorage.mem[15][6] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold270 (.A(\pmod_1414.RX.tickgen.Acc[12] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0389_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold272 (.A(\pmod_1414.RX.tickgen.Acc[11] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold273 (.A(\pmod_1414.mem_strorage.mem[15][5] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold274 (.A(\pmod_1414.mem_strorage.mem[6][1] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold275 (.A(\pmod_1414.mem_strorage.mem[15][0] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold276 (.A(\pmod_1414.mem_strorage.mem[15][3] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold277 (.A(\pmod_1414.RX.RxD_state[0] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0190_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold279 (.A(\pmod_1414.mem_strorage.mem[15][4] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold280 (.A(\pmod_1414.RX.RxD_state[3] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold281 (.A(\pmod_1414.RX.tickgen.Acc[2] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0375_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0045_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold284 (.A(\pmod_1414.RX.OversamplingCnt[1] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0642_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0179_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold287 (.A(\pmod_1414.r_counter[2] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0350_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0027_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold290 (.A(\pmod_1414.r_counter[5] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0353_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0030_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold293 (.A(\pmod_1414.r_counter[8] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold294 (.A(\pmod_1414.RX.RxD_bit ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0211_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0218_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold297 (.A(\pmod_1414.mem_strorage.mem[5][4] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold298 (.A(\pmod_1414.RX.RxD_state[0] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0637_),
    .X(net558));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_fill_2 FILLER_2_399 ();
 sg13g2_decap_4 FILLER_2_404 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_fill_2 FILLER_3_175 ();
 sg13g2_decap_4 FILLER_3_185 ();
 sg13g2_fill_2 FILLER_3_189 ();
 sg13g2_fill_2 FILLER_3_195 ();
 sg13g2_decap_8 FILLER_3_201 ();
 sg13g2_decap_8 FILLER_3_208 ();
 sg13g2_decap_8 FILLER_3_215 ();
 sg13g2_decap_8 FILLER_3_222 ();
 sg13g2_decap_8 FILLER_3_229 ();
 sg13g2_decap_8 FILLER_3_236 ();
 sg13g2_decap_8 FILLER_3_243 ();
 sg13g2_decap_8 FILLER_3_250 ();
 sg13g2_decap_8 FILLER_3_257 ();
 sg13g2_fill_2 FILLER_3_264 ();
 sg13g2_fill_1 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_decap_4 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_285 ();
 sg13g2_decap_8 FILLER_3_292 ();
 sg13g2_decap_8 FILLER_3_299 ();
 sg13g2_fill_2 FILLER_3_323 ();
 sg13g2_fill_1 FILLER_3_325 ();
 sg13g2_decap_8 FILLER_3_330 ();
 sg13g2_decap_8 FILLER_3_337 ();
 sg13g2_decap_8 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_351 ();
 sg13g2_fill_1 FILLER_3_370 ();
 sg13g2_decap_4 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_4 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_4 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_134 ();
 sg13g2_decap_8 FILLER_4_141 ();
 sg13g2_decap_8 FILLER_4_148 ();
 sg13g2_decap_8 FILLER_4_155 ();
 sg13g2_decap_8 FILLER_4_162 ();
 sg13g2_fill_1 FILLER_4_169 ();
 sg13g2_fill_2 FILLER_4_188 ();
 sg13g2_fill_1 FILLER_4_190 ();
 sg13g2_fill_1 FILLER_4_200 ();
 sg13g2_decap_8 FILLER_4_209 ();
 sg13g2_decap_8 FILLER_4_216 ();
 sg13g2_decap_8 FILLER_4_223 ();
 sg13g2_decap_8 FILLER_4_230 ();
 sg13g2_decap_8 FILLER_4_237 ();
 sg13g2_decap_4 FILLER_4_244 ();
 sg13g2_fill_1 FILLER_4_248 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_fill_2 FILLER_4_259 ();
 sg13g2_fill_2 FILLER_4_290 ();
 sg13g2_fill_1 FILLER_4_292 ();
 sg13g2_fill_1 FILLER_4_310 ();
 sg13g2_decap_4 FILLER_4_345 ();
 sg13g2_fill_1 FILLER_4_349 ();
 sg13g2_fill_2 FILLER_4_363 ();
 sg13g2_fill_1 FILLER_4_365 ();
 sg13g2_fill_2 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_4 FILLER_5_21 ();
 sg13g2_fill_1 FILLER_5_25 ();
 sg13g2_fill_1 FILLER_5_30 ();
 sg13g2_fill_2 FILLER_5_44 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_fill_1 FILLER_5_105 ();
 sg13g2_fill_2 FILLER_5_122 ();
 sg13g2_fill_1 FILLER_5_124 ();
 sg13g2_fill_2 FILLER_5_138 ();
 sg13g2_fill_1 FILLER_5_144 ();
 sg13g2_fill_1 FILLER_5_154 ();
 sg13g2_fill_1 FILLER_5_181 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_4 FILLER_5_238 ();
 sg13g2_fill_1 FILLER_5_242 ();
 sg13g2_fill_2 FILLER_5_325 ();
 sg13g2_fill_2 FILLER_5_336 ();
 sg13g2_fill_1 FILLER_5_338 ();
 sg13g2_fill_2 FILLER_5_373 ();
 sg13g2_fill_2 FILLER_5_401 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_20 ();
 sg13g2_fill_1 FILLER_6_54 ();
 sg13g2_decap_8 FILLER_6_81 ();
 sg13g2_decap_8 FILLER_6_88 ();
 sg13g2_fill_2 FILLER_6_95 ();
 sg13g2_fill_1 FILLER_6_97 ();
 sg13g2_fill_2 FILLER_6_163 ();
 sg13g2_fill_1 FILLER_6_165 ();
 sg13g2_fill_1 FILLER_6_312 ();
 sg13g2_fill_2 FILLER_6_328 ();
 sg13g2_fill_1 FILLER_6_330 ();
 sg13g2_fill_1 FILLER_6_374 ();
 sg13g2_fill_2 FILLER_6_398 ();
 sg13g2_fill_2 FILLER_7_52 ();
 sg13g2_fill_2 FILLER_7_88 ();
 sg13g2_fill_1 FILLER_7_90 ();
 sg13g2_fill_1 FILLER_7_95 ();
 sg13g2_fill_2 FILLER_7_114 ();
 sg13g2_fill_2 FILLER_7_148 ();
 sg13g2_fill_1 FILLER_7_150 ();
 sg13g2_fill_2 FILLER_7_177 ();
 sg13g2_fill_1 FILLER_7_179 ();
 sg13g2_fill_1 FILLER_7_223 ();
 sg13g2_fill_1 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_295 ();
 sg13g2_fill_1 FILLER_7_382 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_160 ();
 sg13g2_fill_1 FILLER_8_206 ();
 sg13g2_fill_2 FILLER_8_281 ();
 sg13g2_fill_1 FILLER_8_283 ();
 sg13g2_fill_1 FILLER_8_382 ();
 sg13g2_fill_1 FILLER_9_26 ();
 sg13g2_fill_1 FILLER_9_56 ();
 sg13g2_fill_2 FILLER_9_71 ();
 sg13g2_fill_1 FILLER_9_90 ();
 sg13g2_fill_1 FILLER_9_105 ();
 sg13g2_fill_1 FILLER_9_115 ();
 sg13g2_fill_2 FILLER_9_129 ();
 sg13g2_fill_1 FILLER_9_149 ();
 sg13g2_fill_2 FILLER_9_176 ();
 sg13g2_fill_1 FILLER_9_178 ();
 sg13g2_fill_2 FILLER_9_188 ();
 sg13g2_fill_2 FILLER_9_207 ();
 sg13g2_fill_1 FILLER_9_209 ();
 sg13g2_decap_4 FILLER_9_227 ();
 sg13g2_fill_2 FILLER_9_231 ();
 sg13g2_fill_2 FILLER_9_319 ();
 sg13g2_fill_1 FILLER_9_321 ();
 sg13g2_fill_1 FILLER_9_353 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_218 ();
 sg13g2_fill_1 FILLER_10_225 ();
 sg13g2_fill_2 FILLER_10_252 ();
 sg13g2_fill_1 FILLER_10_254 ();
 sg13g2_fill_2 FILLER_10_273 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_45 ();
 sg13g2_fill_1 FILLER_11_97 ();
 sg13g2_fill_1 FILLER_11_150 ();
 sg13g2_decap_4 FILLER_11_162 ();
 sg13g2_fill_1 FILLER_11_166 ();
 sg13g2_fill_1 FILLER_11_180 ();
 sg13g2_decap_8 FILLER_11_215 ();
 sg13g2_decap_8 FILLER_11_222 ();
 sg13g2_fill_1 FILLER_11_229 ();
 sg13g2_fill_1 FILLER_11_280 ();
 sg13g2_fill_2 FILLER_11_319 ();
 sg13g2_fill_1 FILLER_11_321 ();
 sg13g2_fill_2 FILLER_11_331 ();
 sg13g2_fill_1 FILLER_11_333 ();
 sg13g2_fill_2 FILLER_12_110 ();
 sg13g2_fill_1 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_129 ();
 sg13g2_decap_4 FILLER_12_136 ();
 sg13g2_decap_4 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_213 ();
 sg13g2_fill_2 FILLER_12_220 ();
 sg13g2_fill_1 FILLER_12_222 ();
 sg13g2_fill_1 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_285 ();
 sg13g2_fill_2 FILLER_12_292 ();
 sg13g2_fill_1 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_fill_1 FILLER_13_115 ();
 sg13g2_fill_1 FILLER_13_134 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_fill_1 FILLER_13_163 ();
 sg13g2_fill_2 FILLER_13_196 ();
 sg13g2_fill_2 FILLER_13_203 ();
 sg13g2_fill_2 FILLER_13_231 ();
 sg13g2_fill_2 FILLER_13_269 ();
 sg13g2_fill_1 FILLER_13_271 ();
 sg13g2_fill_2 FILLER_13_308 ();
 sg13g2_fill_1 FILLER_13_310 ();
 sg13g2_fill_1 FILLER_13_337 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_87 ();
 sg13g2_decap_8 FILLER_14_143 ();
 sg13g2_fill_2 FILLER_14_150 ();
 sg13g2_fill_2 FILLER_14_157 ();
 sg13g2_fill_1 FILLER_14_159 ();
 sg13g2_decap_4 FILLER_14_163 ();
 sg13g2_fill_1 FILLER_14_167 ();
 sg13g2_fill_2 FILLER_14_178 ();
 sg13g2_fill_1 FILLER_14_190 ();
 sg13g2_fill_2 FILLER_14_203 ();
 sg13g2_fill_1 FILLER_14_205 ();
 sg13g2_fill_2 FILLER_14_241 ();
 sg13g2_decap_4 FILLER_14_261 ();
 sg13g2_fill_1 FILLER_14_269 ();
 sg13g2_decap_8 FILLER_14_274 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_291 ();
 sg13g2_fill_1 FILLER_14_318 ();
 sg13g2_fill_2 FILLER_14_328 ();
 sg13g2_fill_1 FILLER_14_330 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_4 ();
 sg13g2_fill_1 FILLER_15_39 ();
 sg13g2_fill_1 FILLER_15_83 ();
 sg13g2_fill_1 FILLER_15_115 ();
 sg13g2_fill_2 FILLER_15_164 ();
 sg13g2_fill_1 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_213 ();
 sg13g2_decap_4 FILLER_15_220 ();
 sg13g2_fill_2 FILLER_15_224 ();
 sg13g2_fill_2 FILLER_15_232 ();
 sg13g2_fill_2 FILLER_15_238 ();
 sg13g2_fill_2 FILLER_15_271 ();
 sg13g2_fill_2 FILLER_15_335 ();
 sg13g2_fill_1 FILLER_15_337 ();
 sg13g2_fill_1 FILLER_15_368 ();
 sg13g2_fill_2 FILLER_15_379 ();
 sg13g2_fill_2 FILLER_15_395 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_2 FILLER_16_26 ();
 sg13g2_fill_2 FILLER_16_146 ();
 sg13g2_decap_4 FILLER_16_163 ();
 sg13g2_decap_8 FILLER_16_179 ();
 sg13g2_fill_2 FILLER_16_186 ();
 sg13g2_fill_1 FILLER_16_188 ();
 sg13g2_decap_4 FILLER_16_215 ();
 sg13g2_fill_2 FILLER_16_219 ();
 sg13g2_fill_2 FILLER_16_237 ();
 sg13g2_decap_4 FILLER_16_247 ();
 sg13g2_fill_2 FILLER_16_255 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_decap_4 FILLER_16_278 ();
 sg13g2_fill_2 FILLER_16_282 ();
 sg13g2_fill_1 FILLER_16_288 ();
 sg13g2_fill_2 FILLER_16_301 ();
 sg13g2_fill_2 FILLER_16_357 ();
 sg13g2_fill_1 FILLER_16_398 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_134 ();
 sg13g2_decap_8 FILLER_17_162 ();
 sg13g2_fill_2 FILLER_17_169 ();
 sg13g2_fill_1 FILLER_17_171 ();
 sg13g2_decap_8 FILLER_17_197 ();
 sg13g2_decap_8 FILLER_17_204 ();
 sg13g2_decap_8 FILLER_17_211 ();
 sg13g2_fill_2 FILLER_17_235 ();
 sg13g2_fill_1 FILLER_17_237 ();
 sg13g2_decap_8 FILLER_17_242 ();
 sg13g2_fill_2 FILLER_17_257 ();
 sg13g2_fill_2 FILLER_17_333 ();
 sg13g2_fill_1 FILLER_17_394 ();
 sg13g2_fill_1 FILLER_18_64 ();
 sg13g2_fill_2 FILLER_18_101 ();
 sg13g2_fill_1 FILLER_18_103 ();
 sg13g2_fill_2 FILLER_18_145 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_fill_2 FILLER_18_179 ();
 sg13g2_fill_2 FILLER_18_185 ();
 sg13g2_decap_4 FILLER_18_193 ();
 sg13g2_decap_8 FILLER_18_205 ();
 sg13g2_decap_8 FILLER_18_212 ();
 sg13g2_fill_2 FILLER_18_225 ();
 sg13g2_fill_1 FILLER_18_325 ();
 sg13g2_fill_2 FILLER_18_373 ();
 sg13g2_fill_2 FILLER_19_30 ();
 sg13g2_fill_1 FILLER_19_59 ();
 sg13g2_fill_2 FILLER_19_117 ();
 sg13g2_fill_1 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_153 ();
 sg13g2_fill_2 FILLER_19_170 ();
 sg13g2_decap_8 FILLER_19_209 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_fill_1 FILLER_19_218 ();
 sg13g2_decap_8 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_241 ();
 sg13g2_fill_2 FILLER_19_292 ();
 sg13g2_fill_1 FILLER_19_294 ();
 sg13g2_fill_1 FILLER_19_351 ();
 sg13g2_fill_1 FILLER_19_366 ();
 sg13g2_fill_2 FILLER_19_388 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_69 ();
 sg13g2_decap_8 FILLER_20_75 ();
 sg13g2_fill_1 FILLER_20_82 ();
 sg13g2_fill_2 FILLER_20_120 ();
 sg13g2_fill_2 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_fill_2 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_fill_2 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_209 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_225 ();
 sg13g2_fill_1 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_244 ();
 sg13g2_decap_4 FILLER_20_251 ();
 sg13g2_fill_2 FILLER_20_289 ();
 sg13g2_fill_1 FILLER_20_336 ();
 sg13g2_fill_1 FILLER_20_363 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_11 ();
 sg13g2_fill_1 FILLER_21_62 ();
 sg13g2_fill_1 FILLER_21_72 ();
 sg13g2_fill_2 FILLER_21_120 ();
 sg13g2_fill_2 FILLER_21_151 ();
 sg13g2_fill_1 FILLER_21_153 ();
 sg13g2_fill_2 FILLER_21_158 ();
 sg13g2_fill_1 FILLER_21_160 ();
 sg13g2_decap_4 FILLER_21_179 ();
 sg13g2_fill_1 FILLER_21_183 ();
 sg13g2_decap_4 FILLER_21_190 ();
 sg13g2_fill_2 FILLER_21_236 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_fill_1 FILLER_21_294 ();
 sg13g2_fill_1 FILLER_21_352 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_30 ();
 sg13g2_decap_8 FILLER_22_52 ();
 sg13g2_fill_1 FILLER_22_59 ();
 sg13g2_fill_2 FILLER_22_95 ();
 sg13g2_fill_2 FILLER_22_158 ();
 sg13g2_fill_1 FILLER_22_160 ();
 sg13g2_decap_8 FILLER_22_199 ();
 sg13g2_fill_1 FILLER_22_215 ();
 sg13g2_fill_1 FILLER_22_265 ();
 sg13g2_fill_2 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_302 ();
 sg13g2_fill_2 FILLER_22_309 ();
 sg13g2_fill_1 FILLER_22_311 ();
 sg13g2_fill_2 FILLER_22_317 ();
 sg13g2_fill_1 FILLER_22_319 ();
 sg13g2_fill_2 FILLER_22_329 ();
 sg13g2_fill_2 FILLER_22_377 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_36 ();
 sg13g2_fill_1 FILLER_23_58 ();
 sg13g2_fill_2 FILLER_23_73 ();
 sg13g2_fill_1 FILLER_23_85 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_fill_1 FILLER_23_110 ();
 sg13g2_fill_2 FILLER_23_150 ();
 sg13g2_fill_2 FILLER_23_191 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_250 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_fill_1 FILLER_23_366 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_41 ();
 sg13g2_fill_2 FILLER_24_58 ();
 sg13g2_fill_1 FILLER_24_60 ();
 sg13g2_fill_2 FILLER_24_81 ();
 sg13g2_fill_1 FILLER_24_109 ();
 sg13g2_fill_1 FILLER_24_127 ();
 sg13g2_fill_1 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_237 ();
 sg13g2_fill_2 FILLER_24_309 ();
 sg13g2_fill_1 FILLER_24_311 ();
 sg13g2_fill_2 FILLER_24_380 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_37 ();
 sg13g2_fill_2 FILLER_25_79 ();
 sg13g2_fill_1 FILLER_25_81 ();
 sg13g2_fill_2 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_93 ();
 sg13g2_fill_1 FILLER_25_102 ();
 sg13g2_fill_1 FILLER_25_118 ();
 sg13g2_fill_2 FILLER_25_128 ();
 sg13g2_fill_1 FILLER_25_130 ();
 sg13g2_fill_2 FILLER_25_144 ();
 sg13g2_fill_1 FILLER_25_146 ();
 sg13g2_fill_2 FILLER_25_157 ();
 sg13g2_fill_1 FILLER_25_159 ();
 sg13g2_fill_1 FILLER_25_165 ();
 sg13g2_fill_2 FILLER_25_178 ();
 sg13g2_fill_2 FILLER_25_195 ();
 sg13g2_fill_2 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_fill_1 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_fill_2 FILLER_25_271 ();
 sg13g2_fill_1 FILLER_25_304 ();
 sg13g2_fill_2 FILLER_25_339 ();
 sg13g2_fill_1 FILLER_25_353 ();
 sg13g2_fill_2 FILLER_25_372 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_36 ();
 sg13g2_fill_1 FILLER_26_90 ();
 sg13g2_fill_2 FILLER_26_133 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_fill_1 FILLER_26_305 ();
 sg13g2_fill_1 FILLER_26_319 ();
 sg13g2_fill_1 FILLER_26_329 ();
 sg13g2_fill_1 FILLER_26_336 ();
 sg13g2_fill_2 FILLER_26_351 ();
 sg13g2_fill_1 FILLER_26_353 ();
 sg13g2_fill_1 FILLER_26_360 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_fill_2 FILLER_27_38 ();
 sg13g2_fill_1 FILLER_27_40 ();
 sg13g2_fill_2 FILLER_27_62 ();
 sg13g2_fill_1 FILLER_27_64 ();
 sg13g2_fill_2 FILLER_27_121 ();
 sg13g2_fill_1 FILLER_27_123 ();
 sg13g2_fill_1 FILLER_27_150 ();
 sg13g2_fill_2 FILLER_27_170 ();
 sg13g2_fill_1 FILLER_27_172 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_fill_2 FILLER_27_206 ();
 sg13g2_fill_2 FILLER_27_221 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_fill_2 FILLER_27_266 ();
 sg13g2_fill_1 FILLER_27_313 ();
 sg13g2_fill_1 FILLER_27_323 ();
 sg13g2_fill_1 FILLER_28_59 ();
 sg13g2_fill_2 FILLER_28_88 ();
 sg13g2_fill_1 FILLER_28_99 ();
 sg13g2_fill_2 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_107 ();
 sg13g2_fill_2 FILLER_28_209 ();
 sg13g2_fill_2 FILLER_28_311 ();
 sg13g2_fill_2 FILLER_28_336 ();
 sg13g2_fill_1 FILLER_28_338 ();
 sg13g2_fill_2 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_28_368 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_50 ();
 sg13g2_fill_1 FILLER_29_52 ();
 sg13g2_fill_2 FILLER_29_59 ();
 sg13g2_fill_1 FILLER_29_61 ();
 sg13g2_fill_1 FILLER_29_93 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_130 ();
 sg13g2_fill_1 FILLER_29_132 ();
 sg13g2_fill_2 FILLER_29_147 ();
 sg13g2_fill_1 FILLER_29_149 ();
 sg13g2_fill_2 FILLER_29_158 ();
 sg13g2_fill_1 FILLER_29_160 ();
 sg13g2_fill_1 FILLER_29_166 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_fill_1 FILLER_29_187 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_fill_1 FILLER_29_234 ();
 sg13g2_fill_2 FILLER_29_248 ();
 sg13g2_fill_1 FILLER_29_276 ();
 sg13g2_fill_2 FILLER_29_344 ();
 sg13g2_fill_1 FILLER_29_346 ();
 sg13g2_fill_1 FILLER_29_360 ();
 sg13g2_fill_2 FILLER_29_391 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_1 FILLER_30_59 ();
 sg13g2_fill_2 FILLER_30_64 ();
 sg13g2_fill_1 FILLER_30_66 ();
 sg13g2_fill_2 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_131 ();
 sg13g2_fill_2 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_223 ();
 sg13g2_fill_2 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_fill_2 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_282 ();
 sg13g2_fill_1 FILLER_30_296 ();
 sg13g2_fill_1 FILLER_30_337 ();
 sg13g2_fill_2 FILLER_30_342 ();
 sg13g2_fill_1 FILLER_30_344 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_23 ();
 sg13g2_fill_2 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_92 ();
 sg13g2_fill_1 FILLER_31_107 ();
 sg13g2_fill_2 FILLER_31_152 ();
 sg13g2_fill_2 FILLER_31_163 ();
 sg13g2_fill_1 FILLER_31_165 ();
 sg13g2_fill_2 FILLER_31_174 ();
 sg13g2_fill_2 FILLER_31_193 ();
 sg13g2_fill_1 FILLER_31_195 ();
 sg13g2_fill_2 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_211 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_fill_1 FILLER_31_261 ();
 sg13g2_fill_1 FILLER_31_307 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_fill_2 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_32_65 ();
 sg13g2_fill_1 FILLER_32_81 ();
 sg13g2_fill_2 FILLER_32_87 ();
 sg13g2_fill_2 FILLER_32_121 ();
 sg13g2_fill_1 FILLER_32_137 ();
 sg13g2_fill_1 FILLER_32_144 ();
 sg13g2_fill_1 FILLER_32_173 ();
 sg13g2_fill_2 FILLER_32_191 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_fill_2 FILLER_32_224 ();
 sg13g2_fill_2 FILLER_32_273 ();
 sg13g2_fill_1 FILLER_32_335 ();
 sg13g2_fill_2 FILLER_32_392 ();
 sg13g2_fill_1 FILLER_32_394 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_35 ();
 sg13g2_fill_1 FILLER_33_43 ();
 sg13g2_fill_2 FILLER_33_74 ();
 sg13g2_fill_1 FILLER_33_166 ();
 sg13g2_fill_2 FILLER_33_186 ();
 sg13g2_fill_1 FILLER_33_188 ();
 sg13g2_fill_1 FILLER_33_204 ();
 sg13g2_fill_2 FILLER_33_269 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_fill_1 FILLER_33_294 ();
 sg13g2_fill_2 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_339 ();
 sg13g2_fill_2 FILLER_33_372 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_2 FILLER_34_38 ();
 sg13g2_fill_1 FILLER_34_40 ();
 sg13g2_fill_2 FILLER_34_47 ();
 sg13g2_fill_1 FILLER_34_49 ();
 sg13g2_fill_2 FILLER_34_68 ();
 sg13g2_fill_1 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_108 ();
 sg13g2_fill_2 FILLER_34_119 ();
 sg13g2_fill_1 FILLER_34_193 ();
 sg13g2_fill_2 FILLER_34_206 ();
 sg13g2_fill_2 FILLER_34_242 ();
 sg13g2_fill_1 FILLER_34_305 ();
 sg13g2_fill_1 FILLER_34_321 ();
 sg13g2_fill_2 FILLER_34_346 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_2 FILLER_35_29 ();
 sg13g2_fill_2 FILLER_35_46 ();
 sg13g2_fill_1 FILLER_35_115 ();
 sg13g2_fill_2 FILLER_35_150 ();
 sg13g2_fill_1 FILLER_35_226 ();
 sg13g2_fill_2 FILLER_35_231 ();
 sg13g2_fill_1 FILLER_35_265 ();
 sg13g2_fill_2 FILLER_35_317 ();
 sg13g2_fill_1 FILLER_35_319 ();
 sg13g2_fill_1 FILLER_35_365 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_118 ();
 sg13g2_fill_1 FILLER_36_120 ();
 sg13g2_fill_2 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_211 ();
 sg13g2_fill_2 FILLER_36_220 ();
 sg13g2_fill_1 FILLER_36_288 ();
 sg13g2_fill_2 FILLER_36_302 ();
 sg13g2_fill_2 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_341 ();
 sg13g2_fill_2 FILLER_36_377 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_29 ();
 sg13g2_fill_2 FILLER_37_40 ();
 sg13g2_fill_2 FILLER_37_81 ();
 sg13g2_fill_2 FILLER_37_182 ();
 sg13g2_fill_2 FILLER_37_249 ();
 sg13g2_fill_2 FILLER_37_260 ();
 sg13g2_fill_1 FILLER_37_262 ();
 sg13g2_fill_2 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_296 ();
 sg13g2_fill_1 FILLER_37_298 ();
 sg13g2_fill_2 FILLER_37_374 ();
 sg13g2_fill_1 FILLER_37_399 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_4 ();
 sg13g2_fill_2 FILLER_38_55 ();
 sg13g2_fill_1 FILLER_38_57 ();
 sg13g2_fill_2 FILLER_38_67 ();
 sg13g2_fill_1 FILLER_38_142 ();
 sg13g2_fill_2 FILLER_38_151 ();
 sg13g2_fill_2 FILLER_38_161 ();
 sg13g2_fill_1 FILLER_38_167 ();
 sg13g2_fill_2 FILLER_38_192 ();
 sg13g2_fill_1 FILLER_38_194 ();
 sg13g2_fill_2 FILLER_38_207 ();
 sg13g2_fill_2 FILLER_38_229 ();
 sg13g2_fill_1 FILLER_38_231 ();
 sg13g2_fill_2 FILLER_38_244 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_346 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net253;
 assign uio_oe[2] = net254;
 assign uio_oe[3] = net255;
 assign uio_oe[4] = net256;
 assign uio_oe[5] = net257;
 assign uio_oe[6] = net258;
 assign uio_oe[7] = net259;
 assign uio_out[6] = net4;
 assign uio_out[7] = net5;
 assign uo_out[7] = net6;
endmodule

module tt_um_cdc_test (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \BNC1_out[0] ;
 wire \BNC1_out[1] ;
 wire \BNC1_out[2] ;
 wire \BNC1_out[3] ;
 wire \BNC1_out[4] ;
 wire \BNC1_out[5] ;
 wire \BNC1_out[6] ;
 wire \BNC1_out[7] ;
 wire \BNC2X_out[0] ;
 wire \BNC2X_out[1] ;
 wire \BNC2X_out[4] ;
 wire \BNC2X_out[5] ;
 wire \BNC2Y_out[0] ;
 wire \BNC2Y_out[1] ;
 wire \BNC2Y_out[4] ;
 wire \BNC2Y_out[5] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire \bnc_image_generator.counter[0] ;
 wire \bnc_image_generator.counter[1] ;
 wire \bnc_image_generator.counter[2] ;
 wire \bnc_image_generator.counter[4] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire clknet_0_clk;
 wire \vga_image_generator.character_hold[0] ;
 wire \vga_image_generator.character_hold[10] ;
 wire \vga_image_generator.character_hold[11] ;
 wire \vga_image_generator.character_hold[12] ;
 wire \vga_image_generator.character_hold[13] ;
 wire \vga_image_generator.character_hold[14] ;
 wire \vga_image_generator.character_hold[15] ;
 wire \vga_image_generator.character_hold[16] ;
 wire \vga_image_generator.character_hold[17] ;
 wire \vga_image_generator.character_hold[1] ;
 wire \vga_image_generator.character_hold[2] ;
 wire \vga_image_generator.character_hold[3] ;
 wire \vga_image_generator.character_hold[4] ;
 wire \vga_image_generator.character_hold[5] ;
 wire \vga_image_generator.character_hold[6] ;
 wire \vga_image_generator.character_hold[7] ;
 wire \vga_image_generator.character_hold[8] ;
 wire \vga_image_generator.character_hold[9] ;
 wire \vga_image_generator.counter[0] ;
 wire \vga_image_generator.counter[10] ;
 wire \vga_image_generator.counter[11] ;
 wire \vga_image_generator.counter[12] ;
 wire \vga_image_generator.counter[13] ;
 wire \vga_image_generator.counter[14] ;
 wire \vga_image_generator.counter[15] ;
 wire \vga_image_generator.counter[16] ;
 wire \vga_image_generator.counter[17] ;
 wire \vga_image_generator.counter[18] ;
 wire \vga_image_generator.counter[19] ;
 wire \vga_image_generator.counter[1] ;
 wire \vga_image_generator.counter[20] ;
 wire \vga_image_generator.counter[21] ;
 wire \vga_image_generator.counter[22] ;
 wire \vga_image_generator.counter[23] ;
 wire \vga_image_generator.counter[24] ;
 wire \vga_image_generator.counter[25] ;
 wire \vga_image_generator.counter[26] ;
 wire \vga_image_generator.counter[27] ;
 wire \vga_image_generator.counter[2] ;
 wire \vga_image_generator.counter[3] ;
 wire \vga_image_generator.counter[4] ;
 wire \vga_image_generator.counter[5] ;
 wire \vga_image_generator.counter[6] ;
 wire \vga_image_generator.counter[7] ;
 wire \vga_image_generator.counter[8] ;
 wire \vga_image_generator.counter[9] ;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;

 sg13g2_inv_1 _0855_ (.Y(_0098_),
    .A(\vga_image_generator.character_hold[1] ));
 sg13g2_inv_1 _0856_ (.Y(_0099_),
    .A(\vga_image_generator.character_hold[7] ));
 sg13g2_inv_1 _0857_ (.Y(_0100_),
    .A(\vga_image_generator.character_hold[9] ));
 sg13g2_inv_1 _0858_ (.Y(_0101_),
    .A(\vga_image_generator.character_hold[13] ));
 sg13g2_inv_1 _0859_ (.Y(_0102_),
    .A(net102));
 sg13g2_inv_1 _0860_ (.Y(_0103_),
    .A(net255));
 sg13g2_inv_1 _0861_ (.Y(_0104_),
    .A(net260));
 sg13g2_inv_1 _0862_ (.Y(_0105_),
    .A(net264));
 sg13g2_inv_4 _0863_ (.A(\hvsync_gen.vpos[8] ),
    .Y(_0106_));
 sg13g2_inv_1 _0864_ (.Y(_0107_),
    .A(net254));
 sg13g2_inv_1 _0865_ (.Y(_0108_),
    .A(\hvsync_gen.vpos[0] ));
 sg13g2_inv_2 _0866_ (.Y(_0109_),
    .A(net236));
 sg13g2_inv_2 _0867_ (.Y(_0110_),
    .A(net234));
 sg13g2_inv_1 _0868_ (.Y(_0111_),
    .A(net247));
 sg13g2_inv_1 _0869_ (.Y(_0112_),
    .A(net232));
 sg13g2_inv_2 _0870_ (.Y(_0113_),
    .A(net197));
 sg13g2_inv_2 _0871_ (.Y(_0114_),
    .A(net287));
 sg13g2_inv_2 _0872_ (.Y(_0115_),
    .A(net2));
 sg13g2_inv_1 _0873_ (.Y(_0116_),
    .A(_0018_));
 sg13g2_inv_1 _0874_ (.Y(_0117_),
    .A(\vga_image_generator.counter[22] ));
 sg13g2_inv_1 _0875_ (.Y(_0118_),
    .A(net275));
 sg13g2_inv_1 _0876_ (.Y(_0119_),
    .A(net269));
 sg13g2_inv_1 _0877_ (.Y(_0120_),
    .A(net201));
 sg13g2_inv_1 _0878_ (.Y(_0121_),
    .A(net163));
 sg13g2_inv_1 _0879_ (.Y(_0122_),
    .A(net175));
 sg13g2_inv_1 _0880_ (.Y(_0123_),
    .A(net182));
 sg13g2_inv_1 _0881_ (.Y(_0124_),
    .A(net193));
 sg13g2_inv_1 _0882_ (.Y(_0125_),
    .A(net170));
 sg13g2_inv_2 _0883_ (.Y(_0126_),
    .A(net194));
 sg13g2_inv_1 _0884_ (.Y(_0127_),
    .A(net218));
 sg13g2_inv_1 _0885_ (.Y(_0128_),
    .A(net204));
 sg13g2_inv_1 _0886_ (.Y(_0129_),
    .A(net292));
 sg13g2_nor2b_2 _0887_ (.A(net234),
    .B_N(net237),
    .Y(_0130_));
 sg13g2_nor2_1 _0888_ (.A(net241),
    .B(net245),
    .Y(_0131_));
 sg13g2_nor2_2 _0889_ (.A(net238),
    .B(\hvsync_gen.hpos[6] ),
    .Y(_0132_));
 sg13g2_or2_2 _0890_ (.X(_0133_),
    .B(net242),
    .A(net238));
 sg13g2_nor2_2 _0891_ (.A(net244),
    .B(_0133_),
    .Y(_0134_));
 sg13g2_nand2b_1 _0892_ (.Y(_0135_),
    .B(_0132_),
    .A_N(net244));
 sg13g2_nor2b_2 _0893_ (.A(net246),
    .B_N(net243),
    .Y(_0136_));
 sg13g2_nand2b_2 _0894_ (.Y(_0137_),
    .B(net244),
    .A_N(net246));
 sg13g2_nor2_1 _0895_ (.A(_0133_),
    .B(_0137_),
    .Y(_0138_));
 sg13g2_and2_2 _0896_ (.A(net253),
    .B(\hvsync_gen.hpos[0] ),
    .X(_0139_));
 sg13g2_nand2_2 _0897_ (.Y(_0140_),
    .A(net253),
    .B(\hvsync_gen.hpos[0] ));
 sg13g2_nor2_2 _0898_ (.A(net252),
    .B(net249),
    .Y(_0141_));
 sg13g2_or2_1 _0899_ (.X(_0142_),
    .B(net250),
    .A(net251));
 sg13g2_nor4_1 _0900_ (.A(_0133_),
    .B(_0137_),
    .C(_0139_),
    .D(_0142_),
    .Y(_0143_));
 sg13g2_nor2b_1 _0901_ (.A(\hvsync_gen.hpos[0] ),
    .B_N(\hvsync_gen.hpos[1] ),
    .Y(_0144_));
 sg13g2_nor2_2 _0902_ (.A(net249),
    .B(\hvsync_gen.hpos[4] ),
    .Y(_0145_));
 sg13g2_nor2_1 _0903_ (.A(net248),
    .B(_0137_),
    .Y(_0146_));
 sg13g2_nand2_1 _0904_ (.Y(_0147_),
    .A(net245),
    .B(_0145_));
 sg13g2_nand4_1 _0905_ (.B(_0136_),
    .C(_0141_),
    .A(_0132_),
    .Y(_0148_),
    .D(_0144_));
 sg13g2_o21ai_1 _0906_ (.B1(_0148_),
    .Y(_0149_),
    .A1(_0134_),
    .A2(_0143_));
 sg13g2_nor2_1 _0907_ (.A(net258),
    .B(net256),
    .Y(_0150_));
 sg13g2_nand2_2 _0908_ (.Y(_0151_),
    .A(net259),
    .B(net261));
 sg13g2_or2_1 _0909_ (.X(_0152_),
    .B(net263),
    .A(net262));
 sg13g2_o21ai_1 _0910_ (.B1(net260),
    .Y(_0153_),
    .A1(net262),
    .A2(net264));
 sg13g2_nor3_1 _0911_ (.A(net258),
    .B(net256),
    .C(net260),
    .Y(_0154_));
 sg13g2_and2_1 _0912_ (.A(_0150_),
    .B(_0153_),
    .X(_0155_));
 sg13g2_nand2b_1 _0913_ (.Y(_0156_),
    .B(net259),
    .A_N(net261));
 sg13g2_nand3b_1 _0914_ (.B(_0150_),
    .C(net259),
    .Y(_0157_),
    .A_N(net262));
 sg13g2_nand2b_2 _0915_ (.Y(_0158_),
    .B(net265),
    .A_N(net263));
 sg13g2_nand2_2 _0916_ (.Y(_0159_),
    .A(net266),
    .B(\hvsync_gen.vpos[0] ));
 sg13g2_or3_1 _0917_ (.A(\hvsync_gen.vpos[9] ),
    .B(_0158_),
    .C(_0159_),
    .X(_0160_));
 sg13g2_o21ai_1 _0918_ (.B1(_0155_),
    .Y(_0161_),
    .A1(_0157_),
    .A2(_0160_));
 sg13g2_nor2_1 _0919_ (.A(_0106_),
    .B(net254),
    .Y(_0162_));
 sg13g2_nand2b_2 _0920_ (.Y(_0163_),
    .B(net242),
    .A_N(net238));
 sg13g2_nor2_1 _0921_ (.A(net245),
    .B(net247),
    .Y(_0164_));
 sg13g2_or2_2 _0922_ (.X(_0165_),
    .B(net247),
    .A(net245));
 sg13g2_nor2_2 _0923_ (.A(_0163_),
    .B(_0165_),
    .Y(_0166_));
 sg13g2_a21oi_1 _0924_ (.A1(net242),
    .A2(_0165_),
    .Y(_0167_),
    .B1(net238));
 sg13g2_nor2b_2 _0925_ (.A(net243),
    .B_N(net246),
    .Y(_0168_));
 sg13g2_nand2b_1 _0926_ (.Y(_0169_),
    .B(net247),
    .A_N(net243));
 sg13g2_nor2_2 _0927_ (.A(_0163_),
    .B(_0169_),
    .Y(_0170_));
 sg13g2_and2_2 _0928_ (.A(net252),
    .B(net249),
    .X(_0171_));
 sg13g2_nand2_2 _0929_ (.Y(_0172_),
    .A(net252),
    .B(net250));
 sg13g2_nor2_2 _0930_ (.A(_0140_),
    .B(_0172_),
    .Y(_0173_));
 sg13g2_nand2_1 _0931_ (.Y(_0174_),
    .A(_0139_),
    .B(_0171_));
 sg13g2_a21o_1 _0932_ (.A2(_0174_),
    .A1(_0170_),
    .B1(_0167_),
    .X(_0175_));
 sg13g2_nand4_1 _0933_ (.B(_0149_),
    .C(_0161_),
    .A(\hvsync_gen.vpos[8] ),
    .Y(_0176_),
    .D(_0175_));
 sg13g2_nor2_1 _0934_ (.A(net253),
    .B(net217),
    .Y(_0177_));
 sg13g2_or2_1 _0935_ (.X(_0178_),
    .B(\hvsync_gen.hpos[0] ),
    .A(net253));
 sg13g2_nor2b_2 _0936_ (.A(net248),
    .B_N(net251),
    .Y(_0179_));
 sg13g2_nand2b_2 _0937_ (.Y(_0180_),
    .B(net252),
    .A_N(net249));
 sg13g2_nor2_1 _0938_ (.A(_0178_),
    .B(_0180_),
    .Y(_0181_));
 sg13g2_nor4_2 _0939_ (.A(\hvsync_gen.hpos[7] ),
    .B(net242),
    .C(net244),
    .Y(_0182_),
    .D(net246));
 sg13g2_nor2_1 _0940_ (.A(net236),
    .B(net234),
    .Y(_0183_));
 sg13g2_nand2_2 _0941_ (.Y(_0184_),
    .A(_0109_),
    .B(_0110_));
 sg13g2_a21oi_1 _0942_ (.A1(_0141_),
    .A2(_0182_),
    .Y(_0185_),
    .B1(_0183_));
 sg13g2_a21o_1 _0943_ (.A2(_0182_),
    .A1(_0181_),
    .B1(_0185_),
    .X(_0186_));
 sg13g2_nand2_1 _0944_ (.Y(_0187_),
    .A(net258),
    .B(net255));
 sg13g2_and3_2 _0945_ (.X(_0188_),
    .A(net257),
    .B(net255),
    .C(net259));
 sg13g2_nand3_1 _0946_ (.B(net255),
    .C(net259),
    .A(net257),
    .Y(_0189_));
 sg13g2_nand4_1 _0947_ (.B(net255),
    .C(net259),
    .A(net257),
    .Y(_0190_),
    .D(net261));
 sg13g2_nor2_1 _0948_ (.A(net266),
    .B(\hvsync_gen.vpos[0] ),
    .Y(_0191_));
 sg13g2_or2_1 _0949_ (.X(_0192_),
    .B(\hvsync_gen.vpos[0] ),
    .A(net266));
 sg13g2_nor2_1 _0950_ (.A(\hvsync_gen.vpos[2] ),
    .B(net263),
    .Y(_0193_));
 sg13g2_or2_2 _0951_ (.X(_0194_),
    .B(net263),
    .A(net265));
 sg13g2_a21oi_1 _0952_ (.A1(_0191_),
    .A2(_0193_),
    .Y(_0195_),
    .B1(_0190_));
 sg13g2_a21oi_1 _0953_ (.A1(\hvsync_gen.vpos[2] ),
    .A2(net266),
    .Y(_0196_),
    .B1(_0152_));
 sg13g2_nand2_1 _0954_ (.Y(_0197_),
    .A(_0171_),
    .B(_0178_));
 sg13g2_nand2_1 _0955_ (.Y(_0198_),
    .A(net240),
    .B(net245));
 sg13g2_and2_2 _0956_ (.A(net243),
    .B(net246),
    .X(_0199_));
 sg13g2_nand2_2 _0957_ (.Y(_0200_),
    .A(net243),
    .B(net247));
 sg13g2_nand3_1 _0958_ (.B(net244),
    .C(net246),
    .A(net242),
    .Y(_0201_));
 sg13g2_nor3_1 _0959_ (.A(_0172_),
    .B(_0177_),
    .C(_0201_),
    .Y(_0202_));
 sg13g2_nor3_1 _0960_ (.A(net238),
    .B(\hvsync_gen.vpos[8] ),
    .C(\hvsync_gen.vpos[9] ),
    .Y(_0203_));
 sg13g2_nand2_1 _0961_ (.Y(_0204_),
    .A(_0188_),
    .B(_0203_));
 sg13g2_nor4_1 _0962_ (.A(_0195_),
    .B(_0196_),
    .C(_0202_),
    .D(_0204_),
    .Y(_0205_));
 sg13g2_a21oi_1 _0963_ (.A1(net251),
    .A2(net253),
    .Y(_0206_),
    .B1(net250));
 sg13g2_nor2_1 _0964_ (.A(net240),
    .B(_0200_),
    .Y(_0207_));
 sg13g2_nor3_1 _0965_ (.A(_0133_),
    .B(_0200_),
    .C(_0206_),
    .Y(_0208_));
 sg13g2_o21ai_1 _0966_ (.B1(net249),
    .Y(_0209_),
    .A1(net251),
    .A2(_0139_));
 sg13g2_a21o_1 _0967_ (.A2(_0209_),
    .A1(_0166_),
    .B1(_0208_),
    .X(_0210_));
 sg13g2_nand2b_1 _0968_ (.Y(_0211_),
    .B(_0151_),
    .A_N(net257));
 sg13g2_nand4_1 _0969_ (.B(net259),
    .C(net261),
    .A(net255),
    .Y(_0212_),
    .D(_0194_));
 sg13g2_nand2b_1 _0970_ (.Y(_0213_),
    .B(net255),
    .A_N(net257));
 sg13g2_nor4_1 _0971_ (.A(_0151_),
    .B(_0158_),
    .C(_0192_),
    .D(_0213_),
    .Y(_0214_));
 sg13g2_nand4_1 _0972_ (.B(_0107_),
    .C(_0187_),
    .A(_0106_),
    .Y(_0215_),
    .D(_0212_));
 sg13g2_a22oi_1 _0973_ (.Y(_0216_),
    .B1(_0210_),
    .B2(_0215_),
    .A2(_0205_),
    .A1(_0186_));
 sg13g2_and2_1 _0974_ (.A(net265),
    .B(net263),
    .X(_0217_));
 sg13g2_nand2_1 _0975_ (.Y(_0218_),
    .A(net265),
    .B(net264));
 sg13g2_a21oi_1 _0976_ (.A1(_0192_),
    .A2(_0217_),
    .Y(_0219_),
    .B1(_0157_));
 sg13g2_nor2_1 _0977_ (.A(_0154_),
    .B(_0219_),
    .Y(_0220_));
 sg13g2_a221oi_1 _0978_ (.B2(\hvsync_gen.vpos[8] ),
    .C1(net254),
    .B1(_0220_),
    .A1(_0176_),
    .Y(_0221_),
    .A2(_0216_));
 sg13g2_nand2_1 _0979_ (.Y(_0222_),
    .A(_0170_),
    .B(_0181_));
 sg13g2_a21oi_1 _0980_ (.A1(_0141_),
    .A2(_0170_),
    .Y(_0223_),
    .B1(_0167_));
 sg13g2_a22oi_1 _0981_ (.Y(_0224_),
    .B1(_0184_),
    .B2(_0223_),
    .A2(_0181_),
    .A1(_0170_));
 sg13g2_a21oi_1 _0982_ (.A1(net242),
    .A2(net243),
    .Y(_0225_),
    .B1(net238));
 sg13g2_nor2_1 _0983_ (.A(_0137_),
    .B(_0163_),
    .Y(_0226_));
 sg13g2_nor2b_1 _0984_ (.A(net251),
    .B_N(net249),
    .Y(_0227_));
 sg13g2_o21ai_1 _0985_ (.B1(net249),
    .Y(_0228_),
    .A1(net252),
    .A2(_0178_));
 sg13g2_a21oi_1 _0986_ (.A1(_0226_),
    .A2(_0228_),
    .Y(_0229_),
    .B1(_0225_));
 sg13g2_a21oi_1 _0987_ (.A1(_0138_),
    .A2(_0197_),
    .Y(_0230_),
    .B1(_0134_));
 sg13g2_and2_2 _0988_ (.A(net250),
    .B(net247),
    .X(_0231_));
 sg13g2_o21ai_1 _0989_ (.B1(_0184_),
    .Y(_0232_),
    .A1(_0135_),
    .A2(_0231_));
 sg13g2_nand2_1 _0990_ (.Y(_0233_),
    .A(_0168_),
    .B(net227));
 sg13g2_nand4_1 _0991_ (.B(_0168_),
    .C(_0177_),
    .A(_0132_),
    .Y(_0234_),
    .D(_0227_));
 sg13g2_a21o_1 _0992_ (.A2(_0234_),
    .A1(_0232_),
    .B1(_0230_),
    .X(_0235_));
 sg13g2_o21ai_1 _0993_ (.B1(_0235_),
    .Y(_0236_),
    .A1(_0224_),
    .A2(_0229_));
 sg13g2_nand3_1 _0994_ (.B(net255),
    .C(net261),
    .A(net257),
    .Y(_0237_));
 sg13g2_o21ai_1 _0995_ (.B1(_0189_),
    .Y(_0238_),
    .A1(_0105_),
    .A2(_0237_));
 sg13g2_nor4_1 _0996_ (.A(\hvsync_gen.vpos[8] ),
    .B(net254),
    .C(_0158_),
    .D(_0159_),
    .Y(_0239_));
 sg13g2_nand2b_2 _0997_ (.Y(_0240_),
    .B(net263),
    .A_N(net265));
 sg13g2_nor4_1 _0998_ (.A(\hvsync_gen.vpos[8] ),
    .B(net254),
    .C(_0192_),
    .D(_0240_),
    .Y(_0241_));
 sg13g2_mux2_1 _0999_ (.A0(_0239_),
    .A1(_0241_),
    .S(_0238_),
    .X(_0242_));
 sg13g2_inv_1 _1000_ (.Y(_0243_),
    .A(_0242_));
 sg13g2_nor3_1 _1001_ (.A(net260),
    .B(_0237_),
    .C(_0243_),
    .Y(_0244_));
 sg13g2_a22oi_1 _1002_ (.Y(_0245_),
    .B1(_0173_),
    .B2(_0184_),
    .A2(_0171_),
    .A1(_0144_));
 sg13g2_o21ai_1 _1003_ (.B1(_0245_),
    .Y(_0246_),
    .A1(_0182_),
    .A2(_0183_));
 sg13g2_a21oi_1 _1004_ (.A1(_0140_),
    .A2(_0141_),
    .Y(_0247_),
    .B1(_0201_));
 sg13g2_a21oi_1 _1005_ (.A1(\hvsync_gen.vpos[2] ),
    .A2(_0192_),
    .Y(_0248_),
    .B1(net263));
 sg13g2_nand4_1 _1006_ (.B(_0188_),
    .C(_0203_),
    .A(net262),
    .Y(_0249_),
    .D(_0248_));
 sg13g2_nor2_1 _1007_ (.A(_0247_),
    .B(_0249_),
    .Y(_0250_));
 sg13g2_a221oi_1 _1008_ (.B2(_0250_),
    .C1(_0221_),
    .B1(_0246_),
    .A1(_0236_),
    .Y(_0251_),
    .A2(_0244_));
 sg13g2_nor2b_1 _1009_ (.A(_0251_),
    .B_N(_0130_),
    .Y(_0252_));
 sg13g2_nor2_1 _1010_ (.A(_0172_),
    .B(_0178_),
    .Y(_0253_));
 sg13g2_a22oi_1 _1011_ (.Y(_0254_),
    .B1(_0253_),
    .B2(_0138_),
    .A2(_0230_),
    .A1(_0184_));
 sg13g2_nand2_1 _1012_ (.Y(_0255_),
    .A(_0222_),
    .B(_0223_));
 sg13g2_nand3_1 _1013_ (.B(_0155_),
    .C(_0162_),
    .A(_0130_),
    .Y(_0256_));
 sg13g2_nor4_1 _1014_ (.A(net266),
    .B(_0108_),
    .C(_0157_),
    .D(_0158_),
    .Y(_0257_));
 sg13g2_nor2_2 _1015_ (.A(net239),
    .B(net237),
    .Y(_0258_));
 sg13g2_nor2_1 _1016_ (.A(net254),
    .B(net1),
    .Y(_0259_));
 sg13g2_o21ai_1 _1017_ (.B1(_0259_),
    .Y(_0260_),
    .A1(net233),
    .A2(_0258_));
 sg13g2_o21ai_1 _1018_ (.B1(_0150_),
    .Y(_0261_),
    .A1(_0104_),
    .A2(_0196_));
 sg13g2_o21ai_1 _1019_ (.B1(_0255_),
    .Y(_0262_),
    .A1(_0257_),
    .A2(_0261_));
 sg13g2_or3_1 _1020_ (.A(_0254_),
    .B(_0256_),
    .C(_0262_),
    .X(_0263_));
 sg13g2_o21ai_1 _1021_ (.B1(_0263_),
    .Y(_0264_),
    .A1(_0106_),
    .A2(_0189_));
 sg13g2_nor3_1 _1022_ (.A(net252),
    .B(\hvsync_gen.hpos[1] ),
    .C(\hvsync_gen.hpos[7] ),
    .Y(_0265_));
 sg13g2_a21oi_1 _1023_ (.A1(_0145_),
    .A2(_0265_),
    .Y(_0266_),
    .B1(_0225_));
 sg13g2_nand2_1 _1024_ (.Y(_0267_),
    .A(net236),
    .B(_0266_));
 sg13g2_nand2_1 _1025_ (.Y(_0268_),
    .A(\hvsync_gen.hpos[0] ),
    .B(_0130_));
 sg13g2_nor4_1 _1026_ (.A(net253),
    .B(_0137_),
    .C(_0163_),
    .D(_0268_),
    .Y(_0269_));
 sg13g2_a22oi_1 _1027_ (.Y(_0270_),
    .B1(_0269_),
    .B2(_0141_),
    .A2(_0267_),
    .A1(_0017_));
 sg13g2_nand3_1 _1028_ (.B(_0139_),
    .C(_0227_),
    .A(_0130_),
    .Y(_0271_));
 sg13g2_nand4_1 _1029_ (.B(_0139_),
    .C(_0170_),
    .A(_0130_),
    .Y(_0272_),
    .D(net227));
 sg13g2_nand2_1 _1030_ (.Y(_0273_),
    .A(net236),
    .B(_0133_));
 sg13g2_nand2_1 _1031_ (.Y(_0274_),
    .A(_0110_),
    .B(_0273_));
 sg13g2_nand2_1 _1032_ (.Y(_0275_),
    .A(net246),
    .B(_0171_));
 sg13g2_nor2_1 _1033_ (.A(net244),
    .B(_0163_),
    .Y(_0276_));
 sg13g2_nand3_1 _1034_ (.B(_0275_),
    .C(_0276_),
    .A(_0130_),
    .Y(_0277_));
 sg13g2_nand2_1 _1035_ (.Y(_0278_),
    .A(_0274_),
    .B(_0277_));
 sg13g2_a21oi_1 _1036_ (.A1(_0272_),
    .A2(_0278_),
    .Y(_0279_),
    .B1(_0270_));
 sg13g2_nor3_1 _1037_ (.A(net253),
    .B(_0180_),
    .C(_0268_),
    .Y(_0280_));
 sg13g2_nand2_1 _1038_ (.Y(_0281_),
    .A(_0138_),
    .B(_0280_));
 sg13g2_a21oi_1 _1039_ (.A1(net251),
    .A2(net253),
    .Y(_0282_),
    .B1(_0133_));
 sg13g2_a21oi_1 _1040_ (.A1(_0145_),
    .A2(_0282_),
    .Y(_0283_),
    .B1(_0109_));
 sg13g2_a21o_1 _1041_ (.A2(_0283_),
    .A1(_0135_),
    .B1(_0112_),
    .X(_0284_));
 sg13g2_nor2_2 _1042_ (.A(_0140_),
    .B(_0275_),
    .Y(_0285_));
 sg13g2_o21ai_1 _1043_ (.B1(net236),
    .Y(_0286_),
    .A1(_0135_),
    .A2(_0285_));
 sg13g2_a22oi_1 _1044_ (.Y(_0287_),
    .B1(_0286_),
    .B2(_0110_),
    .A2(_0284_),
    .A1(_0281_));
 sg13g2_nand2_1 _1045_ (.Y(_0288_),
    .A(net266),
    .B(_0108_));
 sg13g2_nor4_1 _1046_ (.A(net260),
    .B(_0194_),
    .C(_0237_),
    .D(_0288_),
    .Y(_0289_));
 sg13g2_a21oi_1 _1047_ (.A1(_0159_),
    .A2(_0193_),
    .Y(_0290_),
    .B1(_0237_));
 sg13g2_or3_1 _1048_ (.A(_0188_),
    .B(_0289_),
    .C(_0290_),
    .X(_0291_));
 sg13g2_o21ai_1 _1049_ (.B1(_0291_),
    .Y(_0292_),
    .A1(_0279_),
    .A2(_0287_));
 sg13g2_a21o_1 _1050_ (.A2(_0206_),
    .A1(_0166_),
    .B1(_0273_),
    .X(_0293_));
 sg13g2_a22oi_1 _1051_ (.Y(_0294_),
    .B1(_0293_),
    .B2(_0017_),
    .A2(_0280_),
    .A1(_0166_));
 sg13g2_a21oi_1 _1052_ (.A1(_0187_),
    .A2(_0212_),
    .Y(_0295_),
    .B1(_0214_));
 sg13g2_nor3_1 _1053_ (.A(_0133_),
    .B(_0200_),
    .C(_0271_),
    .Y(_0296_));
 sg13g2_nor3_1 _1054_ (.A(_0172_),
    .B(_0183_),
    .C(_0200_),
    .Y(_0297_));
 sg13g2_nor3_1 _1055_ (.A(_0274_),
    .B(_0296_),
    .C(_0297_),
    .Y(_0298_));
 sg13g2_nand2b_2 _1056_ (.Y(_0299_),
    .B(_0217_),
    .A_N(_0159_));
 sg13g2_nor3_1 _1057_ (.A(_0156_),
    .B(_0213_),
    .C(_0299_),
    .Y(_0300_));
 sg13g2_a21oi_1 _1058_ (.A1(net256),
    .A2(_0211_),
    .Y(_0301_),
    .B1(_0300_));
 sg13g2_or4_1 _1059_ (.A(_0294_),
    .B(_0295_),
    .C(_0298_),
    .D(_0301_),
    .X(_0302_));
 sg13g2_a21oi_1 _1060_ (.A1(_0292_),
    .A2(_0302_),
    .Y(_0303_),
    .B1(\hvsync_gen.vpos[8] ));
 sg13g2_nor4_2 _1061_ (.A(_0252_),
    .B(_0260_),
    .C(_0264_),
    .Y(_0304_),
    .D(_0303_));
 sg13g2_inv_1 _1062_ (.Y(_0305_),
    .A(_0304_));
 sg13g2_nor2_1 _1063_ (.A(\BNC2Y_out[0] ),
    .B(_0114_),
    .Y(_0306_));
 sg13g2_o21ai_1 _1064_ (.B1(net1),
    .Y(_0307_),
    .A1(\BNC1_out[0] ),
    .A2(net287));
 sg13g2_o21ai_1 _1065_ (.B1(_0305_),
    .Y(uo_out[0]),
    .A1(_0306_),
    .A2(_0307_));
 sg13g2_nor2_1 _1066_ (.A(net237),
    .B(_0163_),
    .Y(_0308_));
 sg13g2_nand2_1 _1067_ (.Y(_0309_),
    .A(net240),
    .B(_0258_));
 sg13g2_nor2_1 _1068_ (.A(_0151_),
    .B(_0194_),
    .Y(_0310_));
 sg13g2_nor4_1 _1069_ (.A(_0021_),
    .B(_0151_),
    .C(_0194_),
    .D(net228),
    .Y(_0311_));
 sg13g2_nor4_2 _1070_ (.A(_0105_),
    .B(_0106_),
    .C(net229),
    .Y(_0312_),
    .D(net228));
 sg13g2_nor2_1 _1071_ (.A(net226),
    .B(_0312_),
    .Y(_0313_));
 sg13g2_a22oi_1 _1072_ (.Y(_0314_),
    .B1(_0168_),
    .B2(_0171_),
    .A2(_0141_),
    .A1(_0136_));
 sg13g2_nor4_2 _1073_ (.A(net264),
    .B(_0106_),
    .C(net229),
    .Y(_0315_),
    .D(net228));
 sg13g2_nor2b_2 _1074_ (.A(net245),
    .B_N(net240),
    .Y(_0316_));
 sg13g2_nand3_1 _1075_ (.B(_0258_),
    .C(_0316_),
    .A(_0231_),
    .Y(_0317_));
 sg13g2_o21ai_1 _1076_ (.B1(_0317_),
    .Y(_0318_),
    .A1(_0147_),
    .A2(_0309_));
 sg13g2_nor3_1 _1077_ (.A(_0021_),
    .B(net229),
    .C(net228),
    .Y(_0319_));
 sg13g2_nor4_2 _1078_ (.A(_0021_),
    .B(net229),
    .C(net228),
    .Y(_0320_),
    .D(_0240_));
 sg13g2_nor3_1 _1079_ (.A(_0112_),
    .B(_0021_),
    .C(net228),
    .Y(_0321_));
 sg13g2_nor4_2 _1080_ (.A(net265),
    .B(_0021_),
    .C(net229),
    .Y(_0322_),
    .D(net228));
 sg13g2_nor4_2 _1081_ (.A(_0021_),
    .B(net229),
    .C(_0194_),
    .Y(_0323_),
    .D(net228));
 sg13g2_a22oi_1 _1082_ (.Y(_0324_),
    .B1(_0323_),
    .B2(_0110_),
    .A2(net226),
    .A1(net232));
 sg13g2_or2_1 _1083_ (.X(_0325_),
    .B(_0323_),
    .A(net226));
 sg13g2_nand3_1 _1084_ (.B(_0308_),
    .C(_0325_),
    .A(_0146_),
    .Y(_0326_));
 sg13g2_nand2_1 _1085_ (.Y(_0327_),
    .A(_0308_),
    .B(_0319_));
 sg13g2_a22oi_1 _1086_ (.Y(_0328_),
    .B1(net227),
    .B2(_0168_),
    .A2(_0179_),
    .A1(_0136_));
 sg13g2_o21ai_1 _1087_ (.B1(_0326_),
    .Y(_0329_),
    .A1(_0327_),
    .A2(_0328_));
 sg13g2_nor2_1 _1088_ (.A(_0112_),
    .B(net2),
    .Y(_0330_));
 sg13g2_nor2b_2 _1089_ (.A(net240),
    .B_N(net239),
    .Y(_0331_));
 sg13g2_nor2_1 _1090_ (.A(_0179_),
    .B(net227),
    .Y(_0332_));
 sg13g2_xor2_1 _1091_ (.B(net248),
    .A(net251),
    .X(_0333_));
 sg13g2_nor2_1 _1092_ (.A(_0200_),
    .B(_0333_),
    .Y(_0334_));
 sg13g2_nand2_1 _1093_ (.Y(_0335_),
    .A(_0315_),
    .B(_0334_));
 sg13g2_nand2_1 _1094_ (.Y(_0336_),
    .A(_0199_),
    .B(_0333_));
 sg13g2_o21ai_1 _1095_ (.B1(_0335_),
    .Y(_0337_),
    .A1(_0313_),
    .A2(_0336_));
 sg13g2_and3_1 _1096_ (.X(_0338_),
    .A(_0116_),
    .B(_0331_),
    .C(_0337_));
 sg13g2_nand2_1 _1097_ (.Y(_0339_),
    .A(net239),
    .B(net235));
 sg13g2_and4_1 _1098_ (.A(net239),
    .B(net235),
    .C(_0207_),
    .D(_0320_),
    .X(_0340_));
 sg13g2_o21ai_1 _1099_ (.B1(\vga_image_generator.character_hold[16] ),
    .Y(_0341_),
    .A1(_0338_),
    .A2(_0340_));
 sg13g2_nor2_1 _1100_ (.A(net235),
    .B(_0133_),
    .Y(_0342_));
 sg13g2_and4_1 _1101_ (.A(_0110_),
    .B(_0146_),
    .C(_0323_),
    .D(_0342_),
    .X(_0343_));
 sg13g2_nor3_1 _1102_ (.A(_0115_),
    .B(net229),
    .C(_0240_),
    .Y(_0344_));
 sg13g2_or2_1 _1103_ (.X(_0345_),
    .B(_0344_),
    .A(_0310_));
 sg13g2_nand2_1 _1104_ (.Y(_0346_),
    .A(_0131_),
    .B(_0231_));
 sg13g2_o21ai_1 _1105_ (.B1(_0346_),
    .Y(_0347_),
    .A1(net240),
    .A2(_0147_));
 sg13g2_and3_1 _1106_ (.X(_0348_),
    .A(_0258_),
    .B(_0345_),
    .C(_0347_));
 sg13g2_nand3_1 _1107_ (.B(_0231_),
    .C(_0258_),
    .A(_0131_),
    .Y(_0349_));
 sg13g2_nor3_1 _1108_ (.A(net229),
    .B(_0194_),
    .C(_0349_),
    .Y(_0350_));
 sg13g2_o21ai_1 _1109_ (.B1(_0321_),
    .Y(_0351_),
    .A1(_0348_),
    .A2(_0350_));
 sg13g2_and3_1 _1110_ (.X(_0352_),
    .A(net232),
    .B(net225),
    .C(_0342_));
 sg13g2_a21oi_1 _1111_ (.A1(net2),
    .A2(_0233_),
    .Y(_0353_),
    .B1(_0328_));
 sg13g2_a21oi_1 _1112_ (.A1(_0352_),
    .A2(_0353_),
    .Y(_0354_),
    .B1(_0343_));
 sg13g2_a21oi_1 _1113_ (.A1(_0351_),
    .A2(_0354_),
    .Y(_0355_),
    .B1(_0098_));
 sg13g2_or2_1 _1114_ (.X(_0356_),
    .B(net225),
    .A(net226));
 sg13g2_and2_1 _1115_ (.A(_0164_),
    .B(net227),
    .X(_0357_));
 sg13g2_nand2_1 _1116_ (.Y(_0358_),
    .A(\vga_image_generator.character_hold[7] ),
    .B(_0357_));
 sg13g2_nor2_1 _1117_ (.A(_0322_),
    .B(_0332_),
    .Y(_0359_));
 sg13g2_nand2_1 _1118_ (.Y(_0360_),
    .A(\vga_image_generator.character_hold[8] ),
    .B(_0136_));
 sg13g2_o21ai_1 _1119_ (.B1(_0358_),
    .Y(_0361_),
    .A1(_0359_),
    .A2(_0360_));
 sg13g2_xnor2_1 _1120_ (.Y(_0362_),
    .A(net248),
    .B(net247));
 sg13g2_nor2_1 _1121_ (.A(net245),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_nor2_1 _1122_ (.A(_0169_),
    .B(_0180_),
    .Y(_0364_));
 sg13g2_a22oi_1 _1123_ (.Y(_0365_),
    .B1(_0364_),
    .B2(_0315_),
    .A2(_0363_),
    .A1(_0322_));
 sg13g2_nand4_1 _1124_ (.B(_0199_),
    .C(net227),
    .A(\vga_image_generator.character_hold[9] ),
    .Y(_0366_),
    .D(net225));
 sg13g2_o21ai_1 _1125_ (.B1(_0366_),
    .Y(_0367_),
    .A1(_0099_),
    .A2(_0365_));
 sg13g2_a21o_1 _1126_ (.A2(_0361_),
    .A1(_0356_),
    .B1(_0367_),
    .X(_0368_));
 sg13g2_nor2b_1 _1127_ (.A(net235),
    .B_N(net239),
    .Y(_0369_));
 sg13g2_nand3_1 _1128_ (.B(_0368_),
    .C(_0369_),
    .A(net240),
    .Y(_0370_));
 sg13g2_nand2_1 _1129_ (.Y(_0371_),
    .A(net232),
    .B(_0320_));
 sg13g2_nand2_1 _1130_ (.Y(_0372_),
    .A(_0324_),
    .B(_0371_));
 sg13g2_a22oi_1 _1131_ (.Y(_0373_),
    .B1(_0315_),
    .B2(_0141_),
    .A2(_0312_),
    .A1(_0171_));
 sg13g2_inv_1 _1132_ (.Y(_0374_),
    .A(_0373_));
 sg13g2_a21oi_1 _1133_ (.A1(net232),
    .A2(_0374_),
    .Y(_0375_),
    .B1(_0372_));
 sg13g2_nand2_1 _1134_ (.Y(_0376_),
    .A(\vga_image_generator.character_hold[0] ),
    .B(_0182_));
 sg13g2_nor3_1 _1135_ (.A(net235),
    .B(_0375_),
    .C(_0376_),
    .Y(_0377_));
 sg13g2_nor2_1 _1136_ (.A(net250),
    .B(_0218_),
    .Y(_0378_));
 sg13g2_nand2b_1 _1137_ (.Y(_0379_),
    .B(net248),
    .A_N(net264));
 sg13g2_nand3_1 _1138_ (.B(_0194_),
    .C(_0379_),
    .A(_0115_),
    .Y(_0380_));
 sg13g2_o21ai_1 _1139_ (.B1(_0172_),
    .Y(_0381_),
    .A1(_0378_),
    .A2(_0380_));
 sg13g2_a22oi_1 _1140_ (.Y(_0382_),
    .B1(_0381_),
    .B2(net225),
    .A2(_0325_),
    .A1(net2));
 sg13g2_nor2_1 _1141_ (.A(_0142_),
    .B(_0200_),
    .Y(_0383_));
 sg13g2_nor4_1 _1142_ (.A(net234),
    .B(_0142_),
    .C(_0200_),
    .D(_0327_),
    .Y(_0384_));
 sg13g2_nand4_1 _1143_ (.B(_0115_),
    .C(net226),
    .A(net241),
    .Y(_0385_),
    .D(_0334_));
 sg13g2_o21ai_1 _1144_ (.B1(_0385_),
    .Y(_0386_),
    .A1(_0201_),
    .A2(_0382_));
 sg13g2_and3_1 _1145_ (.X(_0387_),
    .A(net232),
    .B(_0258_),
    .C(_0386_));
 sg13g2_o21ai_1 _1146_ (.B1(\vga_image_generator.character_hold[4] ),
    .Y(_0388_),
    .A1(_0384_),
    .A2(_0387_));
 sg13g2_nand3_1 _1147_ (.B(_0342_),
    .C(_0372_),
    .A(_0199_),
    .Y(_0389_));
 sg13g2_a21oi_1 _1148_ (.A1(_0352_),
    .A2(_0383_),
    .Y(_0390_),
    .B1(_0115_));
 sg13g2_nor4_1 _1149_ (.A(net234),
    .B(_0142_),
    .C(_0165_),
    .D(_0327_),
    .Y(_0391_));
 sg13g2_nand4_1 _1150_ (.B(_0018_),
    .C(_0166_),
    .A(net233),
    .Y(_0392_),
    .D(_0311_));
 sg13g2_nand2_1 _1151_ (.Y(_0393_),
    .A(_0115_),
    .B(_0392_));
 sg13g2_o21ai_1 _1152_ (.B1(\vga_image_generator.character_hold[2] ),
    .Y(_0394_),
    .A1(_0391_),
    .A2(_0393_));
 sg13g2_a21oi_1 _1153_ (.A1(_0389_),
    .A2(_0390_),
    .Y(_0395_),
    .B1(_0394_));
 sg13g2_nor2_1 _1154_ (.A(net226),
    .B(_0322_),
    .Y(_0396_));
 sg13g2_nand3_1 _1155_ (.B(_0207_),
    .C(_0369_),
    .A(\vga_image_generator.character_hold[6] ),
    .Y(_0397_));
 sg13g2_a21oi_1 _1156_ (.A1(_0373_),
    .A2(_0396_),
    .Y(_0398_),
    .B1(_0397_));
 sg13g2_nor2b_1 _1157_ (.A(_0018_),
    .B_N(\vga_image_generator.character_hold[12] ),
    .Y(_0399_));
 sg13g2_nand2b_1 _1158_ (.Y(_0400_),
    .B(\vga_image_generator.character_hold[12] ),
    .A_N(_0018_));
 sg13g2_nand2_1 _1159_ (.Y(_0401_),
    .A(net225),
    .B(_0332_));
 sg13g2_a22oi_1 _1160_ (.Y(_0402_),
    .B1(_0316_),
    .B2(_0145_),
    .A2(_0207_),
    .A1(net248));
 sg13g2_nand3b_1 _1161_ (.B(net235),
    .C(\vga_image_generator.character_hold[11] ),
    .Y(_0403_),
    .A_N(net239));
 sg13g2_nand3_1 _1162_ (.B(_0134_),
    .C(_0145_),
    .A(net236),
    .Y(_0404_));
 sg13g2_nand4_1 _1163_ (.B(net240),
    .C(_0199_),
    .A(net248),
    .Y(_0405_),
    .D(_0369_));
 sg13g2_a21oi_1 _1164_ (.A1(_0404_),
    .A2(_0405_),
    .Y(_0406_),
    .B1(_0100_));
 sg13g2_and3_1 _1165_ (.X(_0407_),
    .A(\vga_image_generator.character_hold[15] ),
    .B(net239),
    .C(net235));
 sg13g2_and4_1 _1166_ (.A(\vga_image_generator.character_hold[10] ),
    .B(net236),
    .C(_0132_),
    .D(_0168_),
    .X(_0408_));
 sg13g2_a22oi_1 _1167_ (.Y(_0409_),
    .B1(_0330_),
    .B2(_0312_),
    .A2(net225),
    .A1(net2));
 sg13g2_nor2b_1 _1168_ (.A(_0409_),
    .B_N(_0364_),
    .Y(_0410_));
 sg13g2_o21ai_1 _1169_ (.B1(net264),
    .Y(_0411_),
    .A1(net248),
    .A2(_0111_));
 sg13g2_nand4_1 _1170_ (.B(_0330_),
    .C(_0363_),
    .A(_0322_),
    .Y(_0412_),
    .D(_0411_));
 sg13g2_a22oi_1 _1171_ (.Y(_0413_),
    .B1(_0363_),
    .B2(net226),
    .A2(_0357_),
    .A1(net225));
 sg13g2_a21oi_1 _1172_ (.A1(net234),
    .A2(_0115_),
    .Y(_0414_),
    .B1(_0413_));
 sg13g2_nor2_1 _1173_ (.A(_0410_),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_nand3_1 _1174_ (.B(_0109_),
    .C(_0331_),
    .A(\vga_image_generator.character_hold[5] ),
    .Y(_0416_));
 sg13g2_a21oi_1 _1175_ (.A1(_0412_),
    .A2(_0415_),
    .Y(_0417_),
    .B1(_0416_));
 sg13g2_nor4_1 _1176_ (.A(net239),
    .B(_0109_),
    .C(_0198_),
    .D(_0362_),
    .Y(_0418_));
 sg13g2_a22oi_1 _1177_ (.Y(_0419_),
    .B1(net227),
    .B2(_0136_),
    .A2(_0199_),
    .A1(_0179_));
 sg13g2_nor3_1 _1178_ (.A(_0018_),
    .B(_0163_),
    .C(_0419_),
    .Y(_0420_));
 sg13g2_a22oi_1 _1179_ (.Y(_0421_),
    .B1(_0420_),
    .B2(_0356_),
    .A2(_0418_),
    .A1(_0312_));
 sg13g2_nand3_1 _1180_ (.B(\vga_image_generator.counter[22] ),
    .C(_0316_),
    .A(\vga_image_generator.character_hold[17] ),
    .Y(_0422_));
 sg13g2_nor3_1 _1181_ (.A(_0339_),
    .B(_0362_),
    .C(_0422_),
    .Y(_0423_));
 sg13g2_a22oi_1 _1182_ (.Y(_0424_),
    .B1(_0423_),
    .B2(net226),
    .A2(_0408_),
    .A1(_0320_));
 sg13g2_o21ai_1 _1183_ (.B1(_0424_),
    .Y(_0425_),
    .A1(_0101_),
    .A2(_0421_));
 sg13g2_nand4_1 _1184_ (.B(_0116_),
    .C(_0164_),
    .A(\vga_image_generator.character_hold[14] ),
    .Y(_0426_),
    .D(_0331_));
 sg13g2_a21oi_1 _1185_ (.A1(_0396_),
    .A2(_0401_),
    .Y(_0427_),
    .B1(_0426_));
 sg13g2_nand3_1 _1186_ (.B(_0199_),
    .C(net227),
    .A(\vga_image_generator.character_hold[11] ),
    .Y(_0428_));
 sg13g2_nand3_1 _1187_ (.B(_0141_),
    .C(_0168_),
    .A(\vga_image_generator.character_hold[10] ),
    .Y(_0429_));
 sg13g2_nand2_1 _1188_ (.Y(_0430_),
    .A(_0116_),
    .B(_0132_));
 sg13g2_a21oi_1 _1189_ (.A1(_0428_),
    .A2(_0429_),
    .Y(_0431_),
    .B1(_0430_));
 sg13g2_nand3_1 _1190_ (.B(_0116_),
    .C(_0331_),
    .A(\vga_image_generator.character_hold[15] ),
    .Y(_0432_));
 sg13g2_o21ai_1 _1191_ (.B1(_0115_),
    .Y(_0433_),
    .A1(_0317_),
    .A2(_0324_));
 sg13g2_a21o_1 _1192_ (.A2(_0329_),
    .A1(net232),
    .B1(_0433_),
    .X(_0434_));
 sg13g2_or4_1 _1193_ (.A(_0112_),
    .B(_0309_),
    .C(_0313_),
    .D(_0314_),
    .X(_0435_));
 sg13g2_nand3_1 _1194_ (.B(_0136_),
    .C(_0179_),
    .A(net233),
    .Y(_0436_));
 sg13g2_o21ai_1 _1195_ (.B1(_0436_),
    .Y(_0437_),
    .A1(net234),
    .A2(_0233_));
 sg13g2_nand3_1 _1196_ (.B(_0315_),
    .C(_0437_),
    .A(_0308_),
    .Y(_0438_));
 sg13g2_nand2b_1 _1197_ (.Y(_0439_),
    .B(_0318_),
    .A_N(_0371_));
 sg13g2_nand4_1 _1198_ (.B(_0435_),
    .C(_0438_),
    .A(net2),
    .Y(_0440_),
    .D(_0439_));
 sg13g2_or4_1 _1199_ (.A(_0163_),
    .B(_0169_),
    .C(_0333_),
    .D(_0400_),
    .X(_0441_));
 sg13g2_o21ai_1 _1200_ (.B1(_0441_),
    .Y(_0442_),
    .A1(_0328_),
    .A2(_0432_));
 sg13g2_o21ai_1 _1201_ (.B1(net225),
    .Y(_0443_),
    .A1(_0431_),
    .A2(_0442_));
 sg13g2_nand2b_1 _1202_ (.Y(_0444_),
    .B(_0443_),
    .A_N(_0427_));
 sg13g2_a221oi_1 _1203_ (.B2(_0347_),
    .C1(_0408_),
    .B1(_0407_),
    .A1(_0170_),
    .Y(_0445_),
    .A2(_0399_));
 sg13g2_o21ai_1 _1204_ (.B1(_0445_),
    .Y(_0446_),
    .A1(_0402_),
    .A2(_0403_));
 sg13g2_o21ai_1 _1205_ (.B1(_0325_),
    .Y(_0447_),
    .A1(_0406_),
    .A2(_0446_));
 sg13g2_nand3_1 _1206_ (.B(_0434_),
    .C(_0440_),
    .A(\vga_image_generator.character_hold[3] ),
    .Y(_0448_));
 sg13g2_nor3_1 _1207_ (.A(_0398_),
    .B(_0425_),
    .C(_0444_),
    .Y(_0449_));
 sg13g2_and4_1 _1208_ (.A(_0341_),
    .B(_0370_),
    .C(_0447_),
    .D(_0449_),
    .X(_0450_));
 sg13g2_nor4_1 _1209_ (.A(_0355_),
    .B(_0377_),
    .C(_0395_),
    .D(_0417_),
    .Y(_0451_));
 sg13g2_nand4_1 _1210_ (.B(_0448_),
    .C(_0450_),
    .A(_0388_),
    .Y(_0452_),
    .D(_0451_));
 sg13g2_nand2_1 _1211_ (.Y(_0453_),
    .A(_0304_),
    .B(_0452_));
 sg13g2_o21ai_1 _1212_ (.B1(_0304_),
    .Y(_0454_),
    .A1(_0106_),
    .A2(_0452_));
 sg13g2_nor2_1 _1213_ (.A(net287),
    .B(\BNC1_out[1] ),
    .Y(_0455_));
 sg13g2_o21ai_1 _1214_ (.B1(net289),
    .Y(_0456_),
    .A1(_0114_),
    .A2(\BNC2Y_out[1] ));
 sg13g2_o21ai_1 _1215_ (.B1(_0454_),
    .Y(uo_out[1]),
    .A1(_0455_),
    .A2(_0456_));
 sg13g2_nor2_1 _1216_ (.A(net288),
    .B(\BNC1_out[2] ),
    .Y(_0457_));
 sg13g2_o21ai_1 _1217_ (.B1(net289),
    .Y(_0458_),
    .A1(_0114_),
    .A2(\BNC1_out[5] ));
 sg13g2_o21ai_1 _1218_ (.B1(_0453_),
    .Y(uo_out[2]),
    .A1(_0457_),
    .A2(_0458_));
 sg13g2_nand2b_1 _1219_ (.Y(_0459_),
    .B(\hvsync_gen.vsync ),
    .A_N(net289));
 sg13g2_nor2_1 _1220_ (.A(net287),
    .B(\BNC1_out[3] ),
    .Y(_0460_));
 sg13g2_o21ai_1 _1221_ (.B1(net289),
    .Y(_0461_),
    .A1(_0114_),
    .A2(\BNC1_out[4] ));
 sg13g2_o21ai_1 _1222_ (.B1(_0459_),
    .Y(uo_out[3]),
    .A1(_0460_),
    .A2(_0461_));
 sg13g2_nand2_1 _1223_ (.Y(_0462_),
    .A(_0103_),
    .B(_0304_));
 sg13g2_nor2_1 _1224_ (.A(net287),
    .B(\BNC1_out[4] ),
    .Y(_0463_));
 sg13g2_o21ai_1 _1225_ (.B1(net289),
    .Y(_0464_),
    .A1(_0114_),
    .A2(\BNC2Y_out[4] ));
 sg13g2_or2_1 _1226_ (.X(_0465_),
    .B(_0464_),
    .A(_0463_));
 sg13g2_nand3_1 _1227_ (.B(_0462_),
    .C(_0465_),
    .A(_0454_),
    .Y(uo_out[4]));
 sg13g2_nor2_1 _1228_ (.A(net287),
    .B(\BNC1_out[5] ),
    .Y(_0466_));
 sg13g2_o21ai_1 _1229_ (.B1(net289),
    .Y(_0467_),
    .A1(_0114_),
    .A2(\BNC2Y_out[5] ));
 sg13g2_or2_1 _1230_ (.X(_0468_),
    .B(_0467_),
    .A(_0466_));
 sg13g2_nand3_1 _1231_ (.B(_0462_),
    .C(_0468_),
    .A(_0453_),
    .Y(uo_out[5]));
 sg13g2_nor2_1 _1232_ (.A(net287),
    .B(\BNC1_out[6] ),
    .Y(_0469_));
 sg13g2_o21ai_1 _1233_ (.B1(net289),
    .Y(_0470_),
    .A1(_0114_),
    .A2(\BNC1_out[1] ));
 sg13g2_o21ai_1 _1234_ (.B1(_0453_),
    .Y(uo_out[6]),
    .A1(_0469_),
    .A2(_0470_));
 sg13g2_nor2_1 _1235_ (.A(net288),
    .B(\BNC1_out[7] ),
    .Y(_0471_));
 sg13g2_a21oi_1 _1236_ (.A1(_0113_),
    .A2(net287),
    .Y(_0472_),
    .B1(_0471_));
 sg13g2_mux2_1 _1237_ (.A0(hsync),
    .A1(_0472_),
    .S(net289),
    .X(uo_out[7]));
 sg13g2_and2_1 _1238_ (.A(net286),
    .B(\BNC2X_out[0] ),
    .X(uio_out[0]));
 sg13g2_and2_1 _1239_ (.A(net286),
    .B(\BNC2X_out[1] ),
    .X(uio_out[1]));
 sg13g2_and2_1 _1240_ (.A(net286),
    .B(\BNC1_out[7] ),
    .X(uio_out[2]));
 sg13g2_and2_1 _1241_ (.A(net286),
    .B(\BNC1_out[6] ),
    .X(uio_out[3]));
 sg13g2_and2_1 _1242_ (.A(net286),
    .B(\BNC2X_out[4] ),
    .X(uio_out[4]));
 sg13g2_and2_1 _1243_ (.A(net286),
    .B(\BNC2X_out[5] ),
    .X(uio_out[5]));
 sg13g2_and2_1 _1244_ (.A(net286),
    .B(\BNC1_out[3] ),
    .X(uio_out[6]));
 sg13g2_and2_1 _1245_ (.A(net286),
    .B(\BNC1_out[2] ),
    .X(uio_out[7]));
 sg13g2_nand2_1 _1246_ (.Y(_0473_),
    .A(net213),
    .B(_0118_));
 sg13g2_nor2b_1 _1247_ (.A(net278),
    .B_N(net280),
    .Y(_0474_));
 sg13g2_nor2_1 _1248_ (.A(net278),
    .B(_0473_),
    .Y(_0475_));
 sg13g2_nand2_1 _1249_ (.Y(_0476_),
    .A(net208),
    .B(net275));
 sg13g2_nor2b_1 _1250_ (.A(_0475_),
    .B_N(_0476_),
    .Y(_0477_));
 sg13g2_inv_1 _1251_ (.Y(_0478_),
    .A(_0477_));
 sg13g2_nand2_1 _1252_ (.Y(_0479_),
    .A(_0113_),
    .B(_0478_));
 sg13g2_nor2_2 _1253_ (.A(net213),
    .B(net278),
    .Y(_0480_));
 sg13g2_or2_2 _1254_ (.X(_0481_),
    .B(net278),
    .A(net280));
 sg13g2_nor2_1 _1255_ (.A(_0113_),
    .B(_0118_),
    .Y(_0482_));
 sg13g2_nor2_2 _1256_ (.A(_0113_),
    .B(net276),
    .Y(_0483_));
 sg13g2_a21oi_1 _1257_ (.A1(net279),
    .A2(_0483_),
    .Y(_0484_),
    .B1(net267));
 sg13g2_a221oi_1 _1258_ (.B2(net279),
    .C1(net269),
    .B1(_0483_),
    .A1(_0480_),
    .Y(_0485_),
    .A2(_0482_));
 sg13g2_nor2b_2 _1259_ (.A(net280),
    .B_N(net278),
    .Y(_0486_));
 sg13g2_nor2_2 _1260_ (.A(net275),
    .B(_0486_),
    .Y(_0487_));
 sg13g2_nand2_2 _1261_ (.Y(_0488_),
    .A(net279),
    .B(net276));
 sg13g2_o21ai_1 _1262_ (.B1(net195),
    .Y(_0489_),
    .A1(net272),
    .A2(_0488_));
 sg13g2_nor2_1 _1263_ (.A(_0487_),
    .B(_0489_),
    .Y(_0490_));
 sg13g2_a21oi_1 _1264_ (.A1(_0479_),
    .A2(_0485_),
    .Y(_0008_),
    .B1(_0490_));
 sg13g2_and2_2 _1265_ (.A(net280),
    .B(net278),
    .X(_0491_));
 sg13g2_nand2_2 _1266_ (.Y(_0492_),
    .A(net280),
    .B(net278));
 sg13g2_nand3_1 _1267_ (.B(_0481_),
    .C(_0492_),
    .A(net275),
    .Y(_0493_));
 sg13g2_nor2_1 _1268_ (.A(net213),
    .B(net277),
    .Y(_0494_));
 sg13g2_o21ai_1 _1269_ (.B1(net275),
    .Y(_0495_),
    .A1(_0480_),
    .A2(_0491_));
 sg13g2_and2_1 _1270_ (.A(_0473_),
    .B(_0493_),
    .X(_0496_));
 sg13g2_nor2_1 _1271_ (.A(net272),
    .B(_0496_),
    .Y(_0497_));
 sg13g2_nor2_2 _1272_ (.A(net271),
    .B(net275),
    .Y(_0498_));
 sg13g2_nand2b_1 _1273_ (.Y(_0499_),
    .B(_0496_),
    .A_N(_0498_));
 sg13g2_nand2b_1 _1274_ (.Y(_0500_),
    .B(_0488_),
    .A_N(net280));
 sg13g2_a21oi_1 _1275_ (.A1(net272),
    .A2(_0500_),
    .Y(_0501_),
    .B1(_0498_));
 sg13g2_nand2_1 _1276_ (.Y(_0502_),
    .A(net269),
    .B(_0499_));
 sg13g2_o21ai_1 _1277_ (.B1(net231),
    .Y(_0503_),
    .A1(_0491_),
    .A2(_0501_));
 sg13g2_o21ai_1 _1278_ (.B1(_0503_),
    .Y(_0009_),
    .A1(_0497_),
    .A2(_0502_));
 sg13g2_nor2_1 _1279_ (.A(net276),
    .B(_0491_),
    .Y(_0504_));
 sg13g2_nand2_1 _1280_ (.Y(_0505_),
    .A(net275),
    .B(_0026_));
 sg13g2_o21ai_1 _1281_ (.B1(_0505_),
    .Y(_0506_),
    .A1(net277),
    .A2(_0491_));
 sg13g2_nand2_1 _1282_ (.Y(_0507_),
    .A(_0483_),
    .B(_0486_));
 sg13g2_o21ai_1 _1283_ (.B1(_0507_),
    .Y(_0508_),
    .A1(net270),
    .A2(_0506_));
 sg13g2_o21ai_1 _1284_ (.B1(net280),
    .Y(_0509_),
    .A1(net279),
    .A2(net275));
 sg13g2_or2_1 _1285_ (.X(_0510_),
    .B(_0509_),
    .A(net271));
 sg13g2_a22oi_1 _1286_ (.Y(_0010_),
    .B1(_0510_),
    .B2(_0484_),
    .A2(_0508_),
    .A1(net267));
 sg13g2_o21ai_1 _1287_ (.B1(net273),
    .Y(_0511_),
    .A1(net277),
    .A2(_0480_));
 sg13g2_nand2_1 _1288_ (.Y(_0512_),
    .A(_0479_),
    .B(_0511_));
 sg13g2_o21ai_1 _1289_ (.B1(_0113_),
    .Y(_0513_),
    .A1(net156),
    .A2(_0494_));
 sg13g2_nand2_1 _1290_ (.Y(_0514_),
    .A(net272),
    .B(_0492_));
 sg13g2_nand2_1 _1291_ (.Y(_0515_),
    .A(_0513_),
    .B(_0514_));
 sg13g2_and2_1 _1292_ (.A(net230),
    .B(_0511_),
    .X(_0516_));
 sg13g2_a22oi_1 _1293_ (.Y(_0517_),
    .B1(_0515_),
    .B2(_0516_),
    .A2(_0512_),
    .A1(net269));
 sg13g2_inv_1 _1294_ (.Y(_0011_),
    .A(_0517_));
 sg13g2_xnor2_1 _1295_ (.Y(_0518_),
    .A(net280),
    .B(net277));
 sg13g2_a21oi_1 _1296_ (.A1(_0481_),
    .A2(_0518_),
    .Y(_0519_),
    .B1(net270));
 sg13g2_nand2_1 _1297_ (.Y(_0520_),
    .A(_0474_),
    .B(_0483_));
 sg13g2_nand2_1 _1298_ (.Y(_0521_),
    .A(net267),
    .B(_0520_));
 sg13g2_nor2b_1 _1299_ (.A(_0487_),
    .B_N(_0505_),
    .Y(_0522_));
 sg13g2_o21ai_1 _1300_ (.B1(_0520_),
    .Y(_0523_),
    .A1(net270),
    .A2(_0522_));
 sg13g2_nand2_1 _1301_ (.Y(_0524_),
    .A(net230),
    .B(_0523_));
 sg13g2_o21ai_1 _1302_ (.B1(_0524_),
    .Y(_0012_),
    .A1(_0519_),
    .A2(_0521_));
 sg13g2_o21ai_1 _1303_ (.B1(net272),
    .Y(_0525_),
    .A1(net276),
    .A2(_0481_));
 sg13g2_a21oi_1 _1304_ (.A1(net279),
    .A2(net276),
    .Y(_0526_),
    .B1(net273));
 sg13g2_o21ai_1 _1305_ (.B1(_0526_),
    .Y(_0527_),
    .A1(net276),
    .A2(_0491_));
 sg13g2_nand2_1 _1306_ (.Y(_0528_),
    .A(_0525_),
    .B(_0527_));
 sg13g2_o21ai_1 _1307_ (.B1(_0476_),
    .Y(_0529_),
    .A1(net276),
    .A2(_0492_));
 sg13g2_a21oi_1 _1308_ (.A1(_0113_),
    .A2(_0529_),
    .Y(_0530_),
    .B1(net231));
 sg13g2_a22oi_1 _1309_ (.Y(_0013_),
    .B1(_0530_),
    .B2(_0525_),
    .A2(_0528_),
    .A1(net230));
 sg13g2_a21oi_1 _1310_ (.A1(net104),
    .A2(_0488_),
    .Y(_0531_),
    .B1(net269));
 sg13g2_a21oi_1 _1311_ (.A1(net269),
    .A2(_0526_),
    .Y(_0014_),
    .B1(net105));
 sg13g2_a21oi_2 _1312_ (.B1(net270),
    .Y(_0532_),
    .A2(_0481_),
    .A1(_0118_));
 sg13g2_nor3_1 _1313_ (.A(net267),
    .B(_0474_),
    .C(_0487_),
    .Y(_0533_));
 sg13g2_nand2_1 _1314_ (.Y(_0534_),
    .A(net278),
    .B(net267));
 sg13g2_o21ai_1 _1315_ (.B1(net270),
    .Y(_0535_),
    .A1(_0518_),
    .A2(_0534_));
 sg13g2_nor2_1 _1316_ (.A(_0533_),
    .B(_0535_),
    .Y(_0536_));
 sg13g2_a21oi_1 _1317_ (.A1(_0495_),
    .A2(_0532_),
    .Y(_0000_),
    .B1(_0536_));
 sg13g2_a21o_1 _1318_ (.A2(_0514_),
    .A1(_0473_),
    .B1(_0521_),
    .X(_0537_));
 sg13g2_nor2_1 _1319_ (.A(net271),
    .B(_0487_),
    .Y(_0538_));
 sg13g2_nand2_1 _1320_ (.Y(_0539_),
    .A(_0493_),
    .B(_0538_));
 sg13g2_nand2_1 _1321_ (.Y(_0540_),
    .A(net272),
    .B(_0488_));
 sg13g2_o21ai_1 _1322_ (.B1(_0539_),
    .Y(_0541_),
    .A1(_0475_),
    .A2(_0540_));
 sg13g2_o21ai_1 _1323_ (.B1(_0537_),
    .Y(_0001_),
    .A1(net267),
    .A2(_0541_));
 sg13g2_nand2_1 _1324_ (.Y(_0542_),
    .A(net273),
    .B(_0529_));
 sg13g2_xnor2_1 _1325_ (.Y(_0543_),
    .A(net276),
    .B(_0491_));
 sg13g2_nor2_1 _1326_ (.A(net269),
    .B(_0497_),
    .Y(_0544_));
 sg13g2_nor3_1 _1327_ (.A(net181),
    .B(_0480_),
    .C(_0491_),
    .Y(_0545_));
 sg13g2_o21ai_1 _1328_ (.B1(net269),
    .Y(_0546_),
    .A1(net272),
    .A2(_0545_));
 sg13g2_a21oi_1 _1329_ (.A1(net272),
    .A2(_0543_),
    .Y(_0547_),
    .B1(_0546_));
 sg13g2_a21oi_1 _1330_ (.A1(_0542_),
    .A2(_0544_),
    .Y(_0002_),
    .B1(_0547_));
 sg13g2_o21ai_1 _1331_ (.B1(net268),
    .Y(_0548_),
    .A1(_0113_),
    .A2(_0506_));
 sg13g2_a22oi_1 _1332_ (.Y(_0549_),
    .B1(_0509_),
    .B2(net271),
    .A2(_0498_),
    .A1(_0486_));
 sg13g2_nand2_1 _1333_ (.Y(_0550_),
    .A(net230),
    .B(_0549_));
 sg13g2_o21ai_1 _1334_ (.B1(_0550_),
    .Y(_0003_),
    .A1(_0532_),
    .A2(_0548_));
 sg13g2_a22oi_1 _1335_ (.Y(_0551_),
    .B1(_0486_),
    .B2(_0498_),
    .A2(_0478_),
    .A1(net270));
 sg13g2_o21ai_1 _1336_ (.B1(net274),
    .Y(_0552_),
    .A1(net279),
    .A2(_0494_));
 sg13g2_nor2_1 _1337_ (.A(net267),
    .B(_0532_),
    .Y(_0553_));
 sg13g2_a22oi_1 _1338_ (.Y(_0004_),
    .B1(_0552_),
    .B2(_0553_),
    .A2(_0551_),
    .A1(net267));
 sg13g2_nand3_1 _1339_ (.B(_0481_),
    .C(_0518_),
    .A(net270),
    .Y(_0554_));
 sg13g2_mux2_1 _1340_ (.A0(_0475_),
    .A1(_0522_),
    .S(net270),
    .X(_0555_));
 sg13g2_a21oi_1 _1341_ (.A1(_0474_),
    .A2(_0498_),
    .Y(_0556_),
    .B1(net230));
 sg13g2_a22oi_1 _1342_ (.Y(_0005_),
    .B1(_0556_),
    .B2(_0554_),
    .A2(_0555_),
    .A1(net230));
 sg13g2_nand2_1 _1343_ (.Y(_0557_),
    .A(_0480_),
    .B(_0498_));
 sg13g2_o21ai_1 _1344_ (.B1(_0557_),
    .Y(_0558_),
    .A1(_0504_),
    .A2(_0540_));
 sg13g2_a21oi_1 _1345_ (.A1(_0480_),
    .A2(_0498_),
    .Y(_0559_),
    .B1(net231));
 sg13g2_a22oi_1 _1346_ (.Y(_0006_),
    .B1(_0559_),
    .B2(_0542_),
    .A2(_0558_),
    .A1(net231));
 sg13g2_nand2_1 _1347_ (.Y(_0560_),
    .A(net279),
    .B(_0482_));
 sg13g2_nor3_1 _1348_ (.A(net230),
    .B(net104),
    .C(_0488_),
    .Y(_0561_));
 sg13g2_a21oi_1 _1349_ (.A1(net230),
    .A2(_0560_),
    .Y(_0562_),
    .B1(_0561_));
 sg13g2_inv_1 _1350_ (.Y(_0007_),
    .A(_0562_));
 sg13g2_nand4_1 _1351_ (.B(net256),
    .C(net266),
    .A(net258),
    .Y(_0563_),
    .D(_0162_));
 sg13g2_nor3_1 _1352_ (.A(_0156_),
    .B(_0240_),
    .C(net199),
    .Y(_0016_));
 sg13g2_a21oi_1 _1353_ (.A1(_0109_),
    .A2(_0201_),
    .Y(_0564_),
    .B1(net232));
 sg13g2_nor3_1 _1354_ (.A(net241),
    .B(net235),
    .C(_0165_),
    .Y(_0565_));
 sg13g2_nor4_1 _1355_ (.A(_0110_),
    .B(_0258_),
    .C(_0564_),
    .D(_0565_),
    .Y(_0015_));
 sg13g2_and2_1 _1356_ (.A(net101),
    .B(net292),
    .X(_0027_));
 sg13g2_nor3_1 _1357_ (.A(net281),
    .B(_0480_),
    .C(_0491_),
    .Y(_0028_));
 sg13g2_nor2_1 _1358_ (.A(net281),
    .B(_0543_),
    .Y(_0029_));
 sg13g2_nor2_1 _1359_ (.A(net181),
    .B(_0492_),
    .Y(_0566_));
 sg13g2_o21ai_1 _1360_ (.B1(net292),
    .Y(_0567_),
    .A1(net273),
    .A2(_0566_));
 sg13g2_a21oi_1 _1361_ (.A1(net273),
    .A2(_0566_),
    .Y(_0030_),
    .B1(_0567_));
 sg13g2_nor3_1 _1362_ (.A(_0113_),
    .B(_0118_),
    .C(_0492_),
    .Y(_0568_));
 sg13g2_o21ai_1 _1363_ (.B1(net292),
    .Y(_0569_),
    .A1(net268),
    .A2(_0568_));
 sg13g2_a21oi_1 _1364_ (.A1(net268),
    .A2(_0568_),
    .Y(_0031_),
    .B1(_0569_));
 sg13g2_nand4_1 _1365_ (.B(net234),
    .C(_0134_),
    .A(net236),
    .Y(_0570_),
    .D(_0285_));
 sg13g2_and2_1 _1366_ (.A(net294),
    .B(_0570_),
    .X(_0571_));
 sg13g2_nand2_2 _1367_ (.Y(_0572_),
    .A(net294),
    .B(_0570_));
 sg13g2_nand2_1 _1368_ (.Y(_0573_),
    .A(\hvsync_gen.vpos[0] ),
    .B(_0571_));
 sg13g2_nor3_1 _1369_ (.A(net261),
    .B(_0107_),
    .C(_0218_),
    .Y(_0574_));
 sg13g2_nand4_1 _1370_ (.B(_0154_),
    .C(_0191_),
    .A(_0106_),
    .Y(_0575_),
    .D(_0574_));
 sg13g2_nand2_1 _1371_ (.Y(_0576_),
    .A(net293),
    .B(_0575_));
 sg13g2_or2_1 _1372_ (.X(_0577_),
    .B(_0576_),
    .A(_0570_));
 sg13g2_o21ai_1 _1373_ (.B1(_0573_),
    .Y(_0032_),
    .A1(_0102_),
    .A2(_0577_));
 sg13g2_nand2_1 _1374_ (.Y(_0578_),
    .A(net113),
    .B(net224));
 sg13g2_xnor2_1 _1375_ (.Y(_0579_),
    .A(net266),
    .B(\hvsync_gen.vpos[0] ));
 sg13g2_o21ai_1 _1376_ (.B1(_0578_),
    .Y(_0033_),
    .A1(_0577_),
    .A2(_0579_));
 sg13g2_nor2_1 _1377_ (.A(_0159_),
    .B(net224),
    .Y(_0580_));
 sg13g2_o21ai_1 _1378_ (.B1(net293),
    .Y(_0581_),
    .A1(_0570_),
    .A2(_0575_));
 sg13g2_xnor2_1 _1379_ (.Y(_0582_),
    .A(net265),
    .B(_0580_));
 sg13g2_nor2_1 _1380_ (.A(_0581_),
    .B(_0582_),
    .Y(_0034_));
 sg13g2_a21oi_1 _1381_ (.A1(net265),
    .A2(_0580_),
    .Y(_0583_),
    .B1(net263));
 sg13g2_nor2_1 _1382_ (.A(_0299_),
    .B(net224),
    .Y(_0584_));
 sg13g2_nor3_1 _1383_ (.A(_0581_),
    .B(_0583_),
    .C(_0584_),
    .Y(_0035_));
 sg13g2_and2_1 _1384_ (.A(net261),
    .B(_0584_),
    .X(_0585_));
 sg13g2_nor2_1 _1385_ (.A(net261),
    .B(_0584_),
    .Y(_0586_));
 sg13g2_nor3_1 _1386_ (.A(_0581_),
    .B(_0585_),
    .C(_0586_),
    .Y(_0036_));
 sg13g2_nor2_1 _1387_ (.A(net259),
    .B(_0585_),
    .Y(_0587_));
 sg13g2_nor3_2 _1388_ (.A(_0151_),
    .B(_0299_),
    .C(net224),
    .Y(_0588_));
 sg13g2_nor3_1 _1389_ (.A(_0581_),
    .B(_0587_),
    .C(_0588_),
    .Y(_0037_));
 sg13g2_nand2_1 _1390_ (.Y(_0589_),
    .A(net257),
    .B(_0588_));
 sg13g2_xnor2_1 _1391_ (.Y(_0590_),
    .A(net257),
    .B(_0588_));
 sg13g2_nor2_1 _1392_ (.A(_0581_),
    .B(_0590_),
    .Y(_0038_));
 sg13g2_nand2_1 _1393_ (.Y(_0591_),
    .A(_0188_),
    .B(_0585_));
 sg13g2_a221oi_1 _1394_ (.B2(_0103_),
    .C1(_0581_),
    .B1(_0589_),
    .A1(_0188_),
    .Y(_0039_),
    .A2(_0585_));
 sg13g2_xnor2_1 _1395_ (.Y(_0592_),
    .A(_0106_),
    .B(_0591_));
 sg13g2_nor2_1 _1396_ (.A(_0581_),
    .B(_0592_),
    .Y(_0040_));
 sg13g2_nand2_1 _1397_ (.Y(_0593_),
    .A(net254),
    .B(net224));
 sg13g2_nor3_1 _1398_ (.A(_0021_),
    .B(_0190_),
    .C(_0299_),
    .Y(_0594_));
 sg13g2_xnor2_1 _1399_ (.Y(_0595_),
    .A(net254),
    .B(_0594_));
 sg13g2_o21ai_1 _1400_ (.B1(_0593_),
    .Y(_0041_),
    .A1(_0577_),
    .A2(_0595_));
 sg13g2_nand2b_2 _1401_ (.Y(_0596_),
    .B(\vga_image_generator.counter[27] ),
    .A_N(\vga_image_generator.counter[26] ));
 sg13g2_nor3_1 _1402_ (.A(\vga_image_generator.counter[24] ),
    .B(_0128_),
    .C(_0596_),
    .Y(_0597_));
 sg13g2_nor4_2 _1403_ (.A(_0117_),
    .B(\vga_image_generator.counter[20] ),
    .C(\vga_image_generator.counter[21] ),
    .Y(_0598_),
    .D(\vga_image_generator.counter[23] ));
 sg13g2_a21oi_1 _1404_ (.A1(_0597_),
    .A2(_0598_),
    .Y(_0599_),
    .B1(net109));
 sg13g2_nor2_1 _1405_ (.A(net283),
    .B(net110),
    .Y(_0042_));
 sg13g2_nor4_2 _1406_ (.A(_0117_),
    .B(\vga_image_generator.counter[20] ),
    .C(\vga_image_generator.counter[21] ),
    .Y(_0600_),
    .D(_0126_));
 sg13g2_nor3_2 _1407_ (.A(_0127_),
    .B(\vga_image_generator.counter[25] ),
    .C(_0596_),
    .Y(_0601_));
 sg13g2_a21oi_1 _1408_ (.A1(_0600_),
    .A2(_0601_),
    .Y(_0602_),
    .B1(net145));
 sg13g2_nor2_1 _1409_ (.A(net284),
    .B(net146),
    .Y(_0043_));
 sg13g2_nor4_2 _1410_ (.A(\vga_image_generator.counter[22] ),
    .B(\vga_image_generator.counter[20] ),
    .C(\vga_image_generator.counter[21] ),
    .Y(_0603_),
    .D(_0126_));
 sg13g2_a21oi_1 _1411_ (.A1(_0601_),
    .A2(_0603_),
    .Y(_0604_),
    .B1(net115));
 sg13g2_nor2_1 _1412_ (.A(net284),
    .B(net116),
    .Y(_0044_));
 sg13g2_a21oi_1 _1413_ (.A1(_0598_),
    .A2(_0601_),
    .Y(_0605_),
    .B1(net111));
 sg13g2_nor2_1 _1414_ (.A(net283),
    .B(net112),
    .Y(_0045_));
 sg13g2_nor4_2 _1415_ (.A(\vga_image_generator.counter[22] ),
    .B(\vga_image_generator.counter[20] ),
    .C(\vga_image_generator.counter[21] ),
    .Y(_0606_),
    .D(\vga_image_generator.counter[23] ));
 sg13g2_a21oi_1 _1416_ (.A1(_0601_),
    .A2(_0606_),
    .Y(_0607_),
    .B1(net150));
 sg13g2_nor2_1 _1417_ (.A(net284),
    .B(net151),
    .Y(_0046_));
 sg13g2_nor3_2 _1418_ (.A(\vga_image_generator.counter[24] ),
    .B(\vga_image_generator.counter[25] ),
    .C(_0596_),
    .Y(_0608_));
 sg13g2_a21oi_1 _1419_ (.A1(_0600_),
    .A2(_0608_),
    .Y(_0609_),
    .B1(net134));
 sg13g2_nor2_1 _1420_ (.A(net284),
    .B(net135),
    .Y(_0047_));
 sg13g2_a21oi_1 _1421_ (.A1(_0603_),
    .A2(_0608_),
    .Y(_0610_),
    .B1(net154));
 sg13g2_nor2_1 _1422_ (.A(net284),
    .B(net155),
    .Y(_0048_));
 sg13g2_a21oi_1 _1423_ (.A1(_0598_),
    .A2(_0608_),
    .Y(_0611_),
    .B1(net141));
 sg13g2_nor2_1 _1424_ (.A(net283),
    .B(net142),
    .Y(_0049_));
 sg13g2_a21oi_1 _1425_ (.A1(_0606_),
    .A2(_0608_),
    .Y(_0612_),
    .B1(net125));
 sg13g2_nor2_1 _1426_ (.A(net284),
    .B(net126),
    .Y(_0050_));
 sg13g2_nand2_1 _1427_ (.Y(_0613_),
    .A(\vga_image_generator.counter[25] ),
    .B(\vga_image_generator.counter[26] ));
 sg13g2_nand3_1 _1428_ (.B(\vga_image_generator.counter[25] ),
    .C(net184),
    .A(\vga_image_generator.counter[24] ),
    .Y(_0614_));
 sg13g2_nor2_2 _1429_ (.A(\vga_image_generator.counter[27] ),
    .B(_0614_),
    .Y(_0615_));
 sg13g2_a21oi_1 _1430_ (.A1(_0600_),
    .A2(_0615_),
    .Y(_0616_),
    .B1(net139));
 sg13g2_nor2_1 _1431_ (.A(net281),
    .B(net140),
    .Y(_0051_));
 sg13g2_a21oi_1 _1432_ (.A1(_0603_),
    .A2(_0615_),
    .Y(_0617_),
    .B1(net121));
 sg13g2_nor2_1 _1433_ (.A(net281),
    .B(net122),
    .Y(_0052_));
 sg13g2_a21oi_1 _1434_ (.A1(_0598_),
    .A2(_0615_),
    .Y(_0618_),
    .B1(net123));
 sg13g2_nor2_1 _1435_ (.A(net281),
    .B(net124),
    .Y(_0053_));
 sg13g2_a21oi_1 _1436_ (.A1(_0606_),
    .A2(_0615_),
    .Y(_0619_),
    .B1(net152));
 sg13g2_nor2_1 _1437_ (.A(net282),
    .B(net153),
    .Y(_0054_));
 sg13g2_nor3_2 _1438_ (.A(\vga_image_generator.counter[24] ),
    .B(\vga_image_generator.counter[27] ),
    .C(_0613_),
    .Y(_0620_));
 sg13g2_a21oi_1 _1439_ (.A1(_0600_),
    .A2(_0620_),
    .Y(_0621_),
    .B1(net143));
 sg13g2_nor2_1 _1440_ (.A(net281),
    .B(net144),
    .Y(_0055_));
 sg13g2_a21oi_1 _1441_ (.A1(_0603_),
    .A2(_0620_),
    .Y(_0622_),
    .B1(net132));
 sg13g2_nor2_1 _1442_ (.A(net282),
    .B(net133),
    .Y(_0056_));
 sg13g2_a21oi_1 _1443_ (.A1(_0598_),
    .A2(_0620_),
    .Y(_0623_),
    .B1(net107));
 sg13g2_nor2_1 _1444_ (.A(net281),
    .B(net108),
    .Y(_0057_));
 sg13g2_a21oi_1 _1445_ (.A1(_0606_),
    .A2(_0620_),
    .Y(_0624_),
    .B1(net117));
 sg13g2_nor2_1 _1446_ (.A(net282),
    .B(net118),
    .Y(_0058_));
 sg13g2_and2_1 _1447_ (.A(net293),
    .B(net100),
    .X(_0059_));
 sg13g2_o21ai_1 _1448_ (.B1(net293),
    .Y(_0625_),
    .A1(net166),
    .A2(\vga_image_generator.counter[0] ));
 sg13g2_a21oi_1 _1449_ (.A1(net166),
    .A2(\vga_image_generator.counter[0] ),
    .Y(_0060_),
    .B1(_0625_));
 sg13g2_a21oi_1 _1450_ (.A1(\vga_image_generator.counter[1] ),
    .A2(\vga_image_generator.counter[0] ),
    .Y(_0626_),
    .B1(net157));
 sg13g2_nand3_1 _1451_ (.B(\vga_image_generator.counter[0] ),
    .C(net157),
    .A(net166),
    .Y(_0627_));
 sg13g2_nand2_1 _1452_ (.Y(_0628_),
    .A(net293),
    .B(_0627_));
 sg13g2_nor2_1 _1453_ (.A(net158),
    .B(_0628_),
    .Y(_0061_));
 sg13g2_nand2b_1 _1454_ (.Y(_0629_),
    .B(_0627_),
    .A_N(net189));
 sg13g2_nand4_1 _1455_ (.B(\vga_image_generator.counter[0] ),
    .C(net157),
    .A(\vga_image_generator.counter[1] ),
    .Y(_0630_),
    .D(net189));
 sg13g2_and3_1 _1456_ (.X(_0062_),
    .A(net293),
    .B(net190),
    .C(_0630_));
 sg13g2_nor2_1 _1457_ (.A(_0120_),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_a21oi_1 _1458_ (.A1(_0120_),
    .A2(_0630_),
    .Y(_0632_),
    .B1(net284));
 sg13g2_nor2b_1 _1459_ (.A(_0631_),
    .B_N(net202),
    .Y(_0063_));
 sg13g2_nor2_1 _1460_ (.A(net163),
    .B(_0631_),
    .Y(_0633_));
 sg13g2_nor3_1 _1461_ (.A(_0120_),
    .B(_0121_),
    .C(_0630_),
    .Y(_0634_));
 sg13g2_nor3_1 _1462_ (.A(net284),
    .B(net164),
    .C(_0634_),
    .Y(_0064_));
 sg13g2_nor4_2 _1463_ (.A(_0120_),
    .B(_0121_),
    .C(_0122_),
    .Y(_0635_),
    .D(_0630_));
 sg13g2_o21ai_1 _1464_ (.B1(net293),
    .Y(_0636_),
    .A1(net175),
    .A2(_0634_));
 sg13g2_nor2_1 _1465_ (.A(_0635_),
    .B(net176),
    .Y(_0065_));
 sg13g2_nor2_1 _1466_ (.A(net173),
    .B(_0635_),
    .Y(_0637_));
 sg13g2_and2_1 _1467_ (.A(net173),
    .B(_0635_),
    .X(_0638_));
 sg13g2_nor3_1 _1468_ (.A(net283),
    .B(net174),
    .C(_0638_),
    .Y(_0066_));
 sg13g2_and2_1 _1469_ (.A(net178),
    .B(_0638_),
    .X(_0639_));
 sg13g2_o21ai_1 _1470_ (.B1(net291),
    .Y(_0640_),
    .A1(net178),
    .A2(_0638_));
 sg13g2_nor2_1 _1471_ (.A(_0639_),
    .B(_0640_),
    .Y(_0067_));
 sg13g2_or2_1 _1472_ (.X(_0641_),
    .B(_0639_),
    .A(net192));
 sg13g2_nand4_1 _1473_ (.B(net178),
    .C(net192),
    .A(net173),
    .Y(_0642_),
    .D(_0635_));
 sg13g2_and3_1 _1474_ (.X(_0068_),
    .A(net291),
    .B(_0641_),
    .C(_0642_));
 sg13g2_o21ai_1 _1475_ (.B1(net290),
    .Y(_0643_),
    .A1(_0123_),
    .A2(_0642_));
 sg13g2_a21oi_1 _1476_ (.A1(_0123_),
    .A2(_0642_),
    .Y(_0069_),
    .B1(_0643_));
 sg13g2_o21ai_1 _1477_ (.B1(_0124_),
    .Y(_0644_),
    .A1(_0123_),
    .A2(_0642_));
 sg13g2_nor3_1 _1478_ (.A(_0123_),
    .B(_0124_),
    .C(_0642_),
    .Y(_0645_));
 sg13g2_nand2_1 _1479_ (.Y(_0646_),
    .A(net290),
    .B(_0644_));
 sg13g2_nor2_1 _1480_ (.A(_0645_),
    .B(_0646_),
    .Y(_0070_));
 sg13g2_nor4_2 _1481_ (.A(_0123_),
    .B(_0124_),
    .C(_0125_),
    .Y(_0647_),
    .D(_0642_));
 sg13g2_o21ai_1 _1482_ (.B1(net290),
    .Y(_0648_),
    .A1(net170),
    .A2(_0645_));
 sg13g2_nor2_1 _1483_ (.A(_0647_),
    .B(net171),
    .Y(_0071_));
 sg13g2_xnor2_1 _1484_ (.Y(_0649_),
    .A(net179),
    .B(_0647_));
 sg13g2_nor2_1 _1485_ (.A(net283),
    .B(net180),
    .Y(_0072_));
 sg13g2_a21oi_1 _1486_ (.A1(\vga_image_generator.counter[13] ),
    .A2(_0647_),
    .Y(_0650_),
    .B1(net136));
 sg13g2_nand3_1 _1487_ (.B(net136),
    .C(_0647_),
    .A(\vga_image_generator.counter[13] ),
    .Y(_0651_));
 sg13g2_nand2_1 _1488_ (.Y(_0652_),
    .A(net290),
    .B(_0651_));
 sg13g2_nor2_1 _1489_ (.A(net137),
    .B(_0652_),
    .Y(_0073_));
 sg13g2_nor2b_1 _1490_ (.A(net160),
    .B_N(_0651_),
    .Y(_0653_));
 sg13g2_and4_2 _1491_ (.A(\vga_image_generator.counter[13] ),
    .B(net136),
    .C(net160),
    .D(_0647_),
    .X(_0654_));
 sg13g2_nor3_1 _1492_ (.A(net283),
    .B(net161),
    .C(_0654_),
    .Y(_0074_));
 sg13g2_o21ai_1 _1493_ (.B1(net290),
    .Y(_0655_),
    .A1(net148),
    .A2(_0654_));
 sg13g2_a21oi_1 _1494_ (.A1(net148),
    .A2(_0654_),
    .Y(_0075_),
    .B1(_0655_));
 sg13g2_a21oi_1 _1495_ (.A1(\vga_image_generator.counter[16] ),
    .A2(_0654_),
    .Y(_0656_),
    .B1(net130));
 sg13g2_and2_1 _1496_ (.A(net220),
    .B(net130),
    .X(_0657_));
 sg13g2_and2_1 _1497_ (.A(_0654_),
    .B(_0657_),
    .X(_0658_));
 sg13g2_nor3_1 _1498_ (.A(net283),
    .B(net131),
    .C(_0658_),
    .Y(_0076_));
 sg13g2_o21ai_1 _1499_ (.B1(net290),
    .Y(_0659_),
    .A1(net147),
    .A2(_0658_));
 sg13g2_a21oi_1 _1500_ (.A1(net147),
    .A2(_0658_),
    .Y(_0077_),
    .B1(_0659_));
 sg13g2_a21oi_1 _1501_ (.A1(\vga_image_generator.counter[18] ),
    .A2(_0658_),
    .Y(_0660_),
    .B1(net127));
 sg13g2_and4_1 _1502_ (.A(net147),
    .B(net127),
    .C(_0654_),
    .D(_0657_),
    .X(_0661_));
 sg13g2_nor3_1 _1503_ (.A(net281),
    .B(net128),
    .C(_0661_),
    .Y(_0078_));
 sg13g2_and2_1 _1504_ (.A(\vga_image_generator.counter[20] ),
    .B(_0661_),
    .X(_0662_));
 sg13g2_o21ai_1 _1505_ (.B1(net290),
    .Y(_0663_),
    .A1(net215),
    .A2(_0661_));
 sg13g2_nor2_1 _1506_ (.A(_0662_),
    .B(_0663_),
    .Y(_0079_));
 sg13g2_xnor2_1 _1507_ (.Y(_0664_),
    .A(net207),
    .B(_0662_));
 sg13g2_nor2_1 _1508_ (.A(net283),
    .B(_0664_),
    .Y(_0080_));
 sg13g2_a21oi_1 _1509_ (.A1(\vga_image_generator.counter[21] ),
    .A2(_0662_),
    .Y(_0665_),
    .B1(net186));
 sg13g2_nand4_1 _1510_ (.B(\vga_image_generator.counter[20] ),
    .C(\vga_image_generator.counter[21] ),
    .A(\vga_image_generator.counter[22] ),
    .Y(_0666_),
    .D(_0661_));
 sg13g2_nand2_1 _1511_ (.Y(_0667_),
    .A(net291),
    .B(_0666_));
 sg13g2_nor2_1 _1512_ (.A(net187),
    .B(_0667_),
    .Y(_0081_));
 sg13g2_o21ai_1 _1513_ (.B1(net290),
    .Y(_0668_),
    .A1(_0126_),
    .A2(_0666_));
 sg13g2_a21oi_1 _1514_ (.A1(_0126_),
    .A2(_0666_),
    .Y(_0082_),
    .B1(_0668_));
 sg13g2_o21ai_1 _1515_ (.B1(_0127_),
    .Y(_0669_),
    .A1(_0126_),
    .A2(_0666_));
 sg13g2_nor3_1 _1516_ (.A(_0126_),
    .B(_0127_),
    .C(_0666_),
    .Y(_0670_));
 sg13g2_nand2_1 _1517_ (.Y(_0671_),
    .A(net291),
    .B(_0669_));
 sg13g2_nor2_1 _1518_ (.A(_0670_),
    .B(_0671_),
    .Y(_0083_));
 sg13g2_nor4_1 _1519_ (.A(_0126_),
    .B(_0127_),
    .C(_0128_),
    .D(_0666_),
    .Y(_0672_));
 sg13g2_o21ai_1 _1520_ (.B1(net291),
    .Y(_0673_),
    .A1(net204),
    .A2(_0670_));
 sg13g2_nor2_1 _1521_ (.A(_0672_),
    .B(_0673_),
    .Y(_0084_));
 sg13g2_nor3_2 _1522_ (.A(_0126_),
    .B(_0614_),
    .C(_0666_),
    .Y(_0674_));
 sg13g2_o21ai_1 _1523_ (.B1(net291),
    .Y(_0675_),
    .A1(net184),
    .A2(_0672_));
 sg13g2_nor2_1 _1524_ (.A(_0674_),
    .B(_0675_),
    .Y(_0085_));
 sg13g2_o21ai_1 _1525_ (.B1(net291),
    .Y(_0676_),
    .A1(net188),
    .A2(_0674_));
 sg13g2_a21oi_1 _1526_ (.A1(net188),
    .A2(_0674_),
    .Y(_0086_),
    .B1(_0676_));
 sg13g2_and2_1 _1527_ (.A(net99),
    .B(_0571_),
    .X(_0087_));
 sg13g2_nor3_1 _1528_ (.A(net285),
    .B(_0139_),
    .C(_0177_),
    .Y(_0088_));
 sg13g2_xnor2_1 _1529_ (.Y(_0677_),
    .A(net252),
    .B(_0139_));
 sg13g2_nor2_1 _1530_ (.A(_0572_),
    .B(_0677_),
    .Y(_0089_));
 sg13g2_a21oi_1 _1531_ (.A1(net251),
    .A2(_0139_),
    .Y(_0678_),
    .B1(net249));
 sg13g2_nor3_1 _1532_ (.A(_0173_),
    .B(_0572_),
    .C(_0678_),
    .Y(_0090_));
 sg13g2_o21ai_1 _1533_ (.B1(net293),
    .Y(_0679_),
    .A1(net246),
    .A2(_0173_));
 sg13g2_nor2_1 _1534_ (.A(_0285_),
    .B(_0679_),
    .Y(_0091_));
 sg13g2_o21ai_1 _1535_ (.B1(net224),
    .Y(_0680_),
    .A1(net243),
    .A2(_0285_));
 sg13g2_a21oi_1 _1536_ (.A1(net243),
    .A2(_0285_),
    .Y(_0092_),
    .B1(_0680_));
 sg13g2_a21oi_1 _1537_ (.A1(_0173_),
    .A2(_0199_),
    .Y(_0681_),
    .B1(net242));
 sg13g2_nor2_2 _1538_ (.A(_0174_),
    .B(_0201_),
    .Y(_0682_));
 sg13g2_nor3_1 _1539_ (.A(_0572_),
    .B(_0681_),
    .C(_0682_),
    .Y(_0093_));
 sg13g2_or2_1 _1540_ (.X(_0683_),
    .B(_0682_),
    .A(net238));
 sg13g2_nand2_2 _1541_ (.Y(_0684_),
    .A(net238),
    .B(_0682_));
 sg13g2_and3_1 _1542_ (.X(_0094_),
    .A(net224),
    .B(_0683_),
    .C(_0684_));
 sg13g2_o21ai_1 _1543_ (.B1(net224),
    .Y(_0685_),
    .A1(_0109_),
    .A2(_0684_));
 sg13g2_a21oi_1 _1544_ (.A1(_0109_),
    .A2(_0684_),
    .Y(_0095_),
    .B1(_0685_));
 sg13g2_nor2_1 _1545_ (.A(_0018_),
    .B(_0684_),
    .Y(_0686_));
 sg13g2_xnor2_1 _1546_ (.Y(_0687_),
    .A(net168),
    .B(_0686_));
 sg13g2_nor2_1 _1547_ (.A(_0572_),
    .B(net169),
    .Y(_0096_));
 sg13g2_a21oi_1 _1548_ (.A1(_0597_),
    .A2(_0606_),
    .Y(_0688_),
    .B1(net119));
 sg13g2_nor2_1 _1549_ (.A(net282),
    .B(net120),
    .Y(_0097_));
 sg13g2_dfrbp_1 _1550_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net8),
    .D(_0027_),
    .Q_N(_0026_),
    .Q(\bnc_image_generator.counter[0] ));
 sg13g2_dfrbp_1 _1551_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net64),
    .D(_0028_),
    .Q_N(_0025_),
    .Q(\bnc_image_generator.counter[1] ));
 sg13g2_dfrbp_1 _1552_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net63),
    .D(_0029_),
    .Q_N(_0024_),
    .Q(\bnc_image_generator.counter[2] ));
 sg13g2_dfrbp_1 _1553_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net62),
    .D(_0030_),
    .Q_N(_0023_),
    .Q(\BNC1_out[0] ));
 sg13g2_dfrbp_1 _1554_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net19),
    .D(_0031_),
    .Q_N(_0750_),
    .Q(\bnc_image_generator.counter[4] ));
 sg13g2_dfrbp_1 _1555_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net61),
    .D(_0015_),
    .Q_N(_0749_),
    .Q(hsync));
 sg13g2_dfrbp_1 _1556_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net60),
    .D(net103),
    .Q_N(_0022_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _1557_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net58),
    .D(net114),
    .Q_N(_0748_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _1558_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net56),
    .D(_0034_),
    .Q_N(_0747_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _1559_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net54),
    .D(_0035_),
    .Q_N(_0746_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _1560_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net52),
    .D(_0036_),
    .Q_N(_0745_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _1561_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net50),
    .D(_0037_),
    .Q_N(_0744_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _1562_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net48),
    .D(_0038_),
    .Q_N(_0743_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _1563_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net46),
    .D(_0039_),
    .Q_N(_0742_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _1564_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net44),
    .D(_0040_),
    .Q_N(_0021_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _1565_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net76),
    .D(_0041_),
    .Q_N(_0751_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _1566_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net42),
    .D(net200),
    .Q_N(_0741_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 _1567_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net40),
    .D(_0042_),
    .Q_N(_0740_),
    .Q(\vga_image_generator.character_hold[17] ));
 sg13g2_dfrbp_1 _1568_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net38),
    .D(_0043_),
    .Q_N(_0739_),
    .Q(\vga_image_generator.character_hold[15] ));
 sg13g2_dfrbp_1 _1569_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net36),
    .D(_0044_),
    .Q_N(_0738_),
    .Q(\vga_image_generator.character_hold[14] ));
 sg13g2_dfrbp_1 _1570_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net34),
    .D(_0045_),
    .Q_N(_0737_),
    .Q(\vga_image_generator.character_hold[13] ));
 sg13g2_dfrbp_1 _1571_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net32),
    .D(_0046_),
    .Q_N(_0736_),
    .Q(\vga_image_generator.character_hold[12] ));
 sg13g2_dfrbp_1 _1572_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net30),
    .D(_0047_),
    .Q_N(_0735_),
    .Q(\vga_image_generator.character_hold[11] ));
 sg13g2_dfrbp_1 _1573_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net28),
    .D(_0048_),
    .Q_N(_0734_),
    .Q(\vga_image_generator.character_hold[10] ));
 sg13g2_dfrbp_1 _1574_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net26),
    .D(_0049_),
    .Q_N(_0733_),
    .Q(\vga_image_generator.character_hold[9] ));
 sg13g2_dfrbp_1 _1575_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net24),
    .D(_0050_),
    .Q_N(_0732_),
    .Q(\vga_image_generator.character_hold[8] ));
 sg13g2_dfrbp_1 _1576_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net22),
    .D(_0051_),
    .Q_N(_0731_),
    .Q(\vga_image_generator.character_hold[7] ));
 sg13g2_dfrbp_1 _1577_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net20),
    .D(_0052_),
    .Q_N(_0730_),
    .Q(\vga_image_generator.character_hold[6] ));
 sg13g2_dfrbp_1 _1578_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net17),
    .D(_0053_),
    .Q_N(_0729_),
    .Q(\vga_image_generator.character_hold[5] ));
 sg13g2_dfrbp_1 _1579_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net15),
    .D(_0054_),
    .Q_N(_0728_),
    .Q(\vga_image_generator.character_hold[4] ));
 sg13g2_dfrbp_1 _1580_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net13),
    .D(_0055_),
    .Q_N(_0727_),
    .Q(\vga_image_generator.character_hold[3] ));
 sg13g2_dfrbp_1 _1581_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net11),
    .D(_0056_),
    .Q_N(_0726_),
    .Q(\vga_image_generator.character_hold[2] ));
 sg13g2_dfrbp_1 _1582_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net9),
    .D(_0057_),
    .Q_N(_0725_),
    .Q(\vga_image_generator.character_hold[1] ));
 sg13g2_dfrbp_1 _1583_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net6),
    .D(_0058_),
    .Q_N(_0724_),
    .Q(\vga_image_generator.character_hold[0] ));
 sg13g2_dfrbp_1 _1584_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net4),
    .D(_0059_),
    .Q_N(_0020_),
    .Q(\vga_image_generator.counter[0] ));
 sg13g2_dfrbp_1 _1585_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net3),
    .D(net167),
    .Q_N(_0723_),
    .Q(\vga_image_generator.counter[1] ));
 sg13g2_dfrbp_1 _1586_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net75),
    .D(net159),
    .Q_N(_0722_),
    .Q(\vga_image_generator.counter[2] ));
 sg13g2_dfrbp_1 _1587_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net74),
    .D(net191),
    .Q_N(_0721_),
    .Q(\vga_image_generator.counter[3] ));
 sg13g2_dfrbp_1 _1588_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net73),
    .D(net203),
    .Q_N(_0720_),
    .Q(\vga_image_generator.counter[4] ));
 sg13g2_dfrbp_1 _1589_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net72),
    .D(net165),
    .Q_N(_0719_),
    .Q(\vga_image_generator.counter[5] ));
 sg13g2_dfrbp_1 _1590_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net71),
    .D(net177),
    .Q_N(_0718_),
    .Q(\vga_image_generator.counter[6] ));
 sg13g2_dfrbp_1 _1591_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net70),
    .D(_0066_),
    .Q_N(_0717_),
    .Q(\vga_image_generator.counter[7] ));
 sg13g2_dfrbp_1 _1592_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net69),
    .D(_0067_),
    .Q_N(_0716_),
    .Q(\vga_image_generator.counter[8] ));
 sg13g2_dfrbp_1 _1593_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net68),
    .D(_0068_),
    .Q_N(_0715_),
    .Q(\vga_image_generator.counter[9] ));
 sg13g2_dfrbp_1 _1594_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net67),
    .D(net183),
    .Q_N(_0714_),
    .Q(\vga_image_generator.counter[10] ));
 sg13g2_dfrbp_1 _1595_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net66),
    .D(_0070_),
    .Q_N(_0713_),
    .Q(\vga_image_generator.counter[11] ));
 sg13g2_dfrbp_1 _1596_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net65),
    .D(net172),
    .Q_N(_0712_),
    .Q(\vga_image_generator.counter[12] ));
 sg13g2_dfrbp_1 _1597_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net59),
    .D(_0072_),
    .Q_N(_0711_),
    .Q(\vga_image_generator.counter[13] ));
 sg13g2_dfrbp_1 _1598_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net57),
    .D(net138),
    .Q_N(_0710_),
    .Q(\vga_image_generator.counter[14] ));
 sg13g2_dfrbp_1 _1599_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net55),
    .D(net162),
    .Q_N(_0709_),
    .Q(\vga_image_generator.counter[15] ));
 sg13g2_dfrbp_1 _1600_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net53),
    .D(net149),
    .Q_N(_0708_),
    .Q(\vga_image_generator.counter[16] ));
 sg13g2_dfrbp_1 _1601_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net51),
    .D(_0076_),
    .Q_N(_0707_),
    .Q(\vga_image_generator.counter[17] ));
 sg13g2_dfrbp_1 _1602_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net49),
    .D(_0077_),
    .Q_N(_0706_),
    .Q(\vga_image_generator.counter[18] ));
 sg13g2_dfrbp_1 _1603_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net47),
    .D(net129),
    .Q_N(_0705_),
    .Q(\vga_image_generator.counter[19] ));
 sg13g2_dfrbp_1 _1604_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net45),
    .D(_0079_),
    .Q_N(_0704_),
    .Q(\vga_image_generator.counter[20] ));
 sg13g2_dfrbp_1 _1605_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net43),
    .D(_0080_),
    .Q_N(_0703_),
    .Q(\vga_image_generator.counter[21] ));
 sg13g2_dfrbp_1 _1606_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net41),
    .D(_0081_),
    .Q_N(_0702_),
    .Q(\vga_image_generator.counter[22] ));
 sg13g2_dfrbp_1 _1607_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net39),
    .D(_0082_),
    .Q_N(_0701_),
    .Q(\vga_image_generator.counter[23] ));
 sg13g2_dfrbp_1 _1608_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net37),
    .D(_0083_),
    .Q_N(_0700_),
    .Q(\vga_image_generator.counter[24] ));
 sg13g2_dfrbp_1 _1609_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net35),
    .D(_0084_),
    .Q_N(_0699_),
    .Q(\vga_image_generator.counter[25] ));
 sg13g2_dfrbp_1 _1610_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net33),
    .D(net185),
    .Q_N(_0698_),
    .Q(\vga_image_generator.counter[26] ));
 sg13g2_dfrbp_1 _1611_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net31),
    .D(_0086_),
    .Q_N(_0697_),
    .Q(\vga_image_generator.counter[27] ));
 sg13g2_dfrbp_1 _1612_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net29),
    .D(_0087_),
    .Q_N(_0019_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 _1613_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net27),
    .D(_0088_),
    .Q_N(_0696_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _1614_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net25),
    .D(_0089_),
    .Q_N(_0695_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _1615_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net23),
    .D(_0090_),
    .Q_N(_0694_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _1616_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net21),
    .D(_0091_),
    .Q_N(_0693_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _1617_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net18),
    .D(_0092_),
    .Q_N(_0692_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _1618_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net16),
    .D(_0093_),
    .Q_N(_0691_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _1619_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net14),
    .D(_0094_),
    .Q_N(_0690_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _1620_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net12),
    .D(_0095_),
    .Q_N(_0018_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _1621_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net10),
    .D(_0096_),
    .Q_N(_0017_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _1622_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net77),
    .D(_0097_),
    .Q_N(_0752_),
    .Q(\vga_image_generator.character_hold[16] ));
 sg13g2_dfrbp_1 _1623_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net78),
    .D(net196),
    .Q_N(_0753_),
    .Q(\BNC2Y_out[0] ));
 sg13g2_dfrbp_1 _1624_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net79),
    .D(_0009_),
    .Q_N(_0754_),
    .Q(\BNC2Y_out[4] ));
 sg13g2_dfrbp_1 _1625_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net80),
    .D(_0010_),
    .Q_N(_0755_),
    .Q(\BNC2Y_out[1] ));
 sg13g2_dfrbp_1 _1626_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net81),
    .D(_0011_),
    .Q_N(_0756_),
    .Q(\BNC2Y_out[5] ));
 sg13g2_dfrbp_1 _1627_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net82),
    .D(_0012_),
    .Q_N(_0757_),
    .Q(\BNC1_out[5] ));
 sg13g2_dfrbp_1 _1628_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net83),
    .D(_0013_),
    .Q_N(_0758_),
    .Q(\BNC1_out[1] ));
 sg13g2_dfrbp_1 _1629_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net84),
    .D(net106),
    .Q_N(_0759_),
    .Q(\BNC1_out[4] ));
 sg13g2_dfrbp_1 _1630_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net85),
    .D(_0000_),
    .Q_N(_0760_),
    .Q(\BNC2X_out[0] ));
 sg13g2_dfrbp_1 _1631_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net86),
    .D(_0001_),
    .Q_N(_0761_),
    .Q(\BNC2X_out[4] ));
 sg13g2_dfrbp_1 _1632_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net87),
    .D(_0002_),
    .Q_N(_0762_),
    .Q(\BNC2X_out[1] ));
 sg13g2_dfrbp_1 _1633_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net88),
    .D(_0003_),
    .Q_N(_0763_),
    .Q(\BNC2X_out[5] ));
 sg13g2_dfrbp_1 _1634_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net89),
    .D(_0004_),
    .Q_N(_0764_),
    .Q(\BNC1_out[7] ));
 sg13g2_dfrbp_1 _1635_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net90),
    .D(_0005_),
    .Q_N(_0765_),
    .Q(\BNC1_out[3] ));
 sg13g2_dfrbp_1 _1636_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net5),
    .D(_0006_),
    .Q_N(_0766_),
    .Q(\BNC1_out[6] ));
 sg13g2_dfrbp_1 _1637_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net7),
    .D(_0007_),
    .Q_N(_0689_),
    .Q(\BNC1_out[2] ));
 sg13g2_tiehi _1584__4 (.L_HI(net4));
 sg13g2_tiehi _1636__5 (.L_HI(net5));
 sg13g2_tiehi _1583__6 (.L_HI(net6));
 sg13g2_tiehi _1637__7 (.L_HI(net7));
 sg13g2_tiehi _1550__8 (.L_HI(net8));
 sg13g2_tiehi _1582__9 (.L_HI(net9));
 sg13g2_tiehi _1621__10 (.L_HI(net10));
 sg13g2_tiehi _1581__11 (.L_HI(net11));
 sg13g2_tiehi _1620__12 (.L_HI(net12));
 sg13g2_tiehi _1580__13 (.L_HI(net13));
 sg13g2_tiehi _1619__14 (.L_HI(net14));
 sg13g2_tiehi _1579__15 (.L_HI(net15));
 sg13g2_tiehi _1618__16 (.L_HI(net16));
 sg13g2_tiehi _1578__17 (.L_HI(net17));
 sg13g2_tiehi _1617__18 (.L_HI(net18));
 sg13g2_tiehi _1554__19 (.L_HI(net19));
 sg13g2_tiehi _1577__20 (.L_HI(net20));
 sg13g2_tiehi _1616__21 (.L_HI(net21));
 sg13g2_tiehi _1576__22 (.L_HI(net22));
 sg13g2_tiehi _1615__23 (.L_HI(net23));
 sg13g2_tiehi _1575__24 (.L_HI(net24));
 sg13g2_tiehi _1614__25 (.L_HI(net25));
 sg13g2_tiehi _1574__26 (.L_HI(net26));
 sg13g2_tiehi _1613__27 (.L_HI(net27));
 sg13g2_tiehi _1573__28 (.L_HI(net28));
 sg13g2_tiehi _1612__29 (.L_HI(net29));
 sg13g2_tiehi _1572__30 (.L_HI(net30));
 sg13g2_tiehi _1611__31 (.L_HI(net31));
 sg13g2_tiehi _1571__32 (.L_HI(net32));
 sg13g2_tiehi _1610__33 (.L_HI(net33));
 sg13g2_tiehi _1570__34 (.L_HI(net34));
 sg13g2_tiehi _1609__35 (.L_HI(net35));
 sg13g2_tiehi _1569__36 (.L_HI(net36));
 sg13g2_tiehi _1608__37 (.L_HI(net37));
 sg13g2_tiehi _1568__38 (.L_HI(net38));
 sg13g2_tiehi _1607__39 (.L_HI(net39));
 sg13g2_tiehi _1567__40 (.L_HI(net40));
 sg13g2_tiehi _1606__41 (.L_HI(net41));
 sg13g2_tiehi _1566__42 (.L_HI(net42));
 sg13g2_tiehi _1605__43 (.L_HI(net43));
 sg13g2_tiehi _1564__44 (.L_HI(net44));
 sg13g2_tiehi _1604__45 (.L_HI(net45));
 sg13g2_tiehi _1563__46 (.L_HI(net46));
 sg13g2_tiehi _1603__47 (.L_HI(net47));
 sg13g2_tiehi _1562__48 (.L_HI(net48));
 sg13g2_tiehi _1602__49 (.L_HI(net49));
 sg13g2_tiehi _1561__50 (.L_HI(net50));
 sg13g2_tiehi _1601__51 (.L_HI(net51));
 sg13g2_tiehi _1560__52 (.L_HI(net52));
 sg13g2_tiehi _1600__53 (.L_HI(net53));
 sg13g2_tiehi _1559__54 (.L_HI(net54));
 sg13g2_tiehi _1599__55 (.L_HI(net55));
 sg13g2_tiehi _1558__56 (.L_HI(net56));
 sg13g2_tiehi _1598__57 (.L_HI(net57));
 sg13g2_tiehi _1557__58 (.L_HI(net58));
 sg13g2_tiehi _1597__59 (.L_HI(net59));
 sg13g2_tiehi _1556__60 (.L_HI(net60));
 sg13g2_tiehi _1555__61 (.L_HI(net61));
 sg13g2_tiehi _1553__62 (.L_HI(net62));
 sg13g2_tiehi _1552__63 (.L_HI(net63));
 sg13g2_tiehi _1551__64 (.L_HI(net64));
 sg13g2_tiehi _1596__65 (.L_HI(net65));
 sg13g2_tiehi _1595__66 (.L_HI(net66));
 sg13g2_tiehi _1594__67 (.L_HI(net67));
 sg13g2_tiehi _1593__68 (.L_HI(net68));
 sg13g2_tiehi _1592__69 (.L_HI(net69));
 sg13g2_tiehi _1591__70 (.L_HI(net70));
 sg13g2_tiehi _1590__71 (.L_HI(net71));
 sg13g2_tiehi _1589__72 (.L_HI(net72));
 sg13g2_tiehi _1588__73 (.L_HI(net73));
 sg13g2_tiehi _1587__74 (.L_HI(net74));
 sg13g2_tiehi _1586__75 (.L_HI(net75));
 sg13g2_tiehi _1565__76 (.L_HI(net76));
 sg13g2_tiehi _1622__77 (.L_HI(net77));
 sg13g2_tiehi _1623__78 (.L_HI(net78));
 sg13g2_tiehi _1624__79 (.L_HI(net79));
 sg13g2_tiehi _1625__80 (.L_HI(net80));
 sg13g2_tiehi _1626__81 (.L_HI(net81));
 sg13g2_tiehi _1627__82 (.L_HI(net82));
 sg13g2_tiehi _1628__83 (.L_HI(net83));
 sg13g2_tiehi _1629__84 (.L_HI(net84));
 sg13g2_tiehi _1630__85 (.L_HI(net85));
 sg13g2_tiehi _1631__86 (.L_HI(net86));
 sg13g2_tiehi _1632__87 (.L_HI(net87));
 sg13g2_tiehi _1633__88 (.L_HI(net88));
 sg13g2_tiehi _1634__89 (.L_HI(net89));
 sg13g2_tiehi _1635__90 (.L_HI(net90));
 sg13g2_tiehi tt_um_cdc_test_91 (.L_HI(net91));
 sg13g2_tiehi tt_um_cdc_test_92 (.L_HI(net92));
 sg13g2_tiehi tt_um_cdc_test_93 (.L_HI(net93));
 sg13g2_tiehi tt_um_cdc_test_94 (.L_HI(net94));
 sg13g2_tiehi tt_um_cdc_test_95 (.L_HI(net95));
 sg13g2_tiehi tt_um_cdc_test_96 (.L_HI(net96));
 sg13g2_tiehi tt_um_cdc_test_97 (.L_HI(net97));
 sg13g2_tiehi tt_um_cdc_test_98 (.L_HI(net98));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_4 fanout224 (.X(net224),
    .A(_0571_));
 sg13g2_buf_2 fanout225 (.A(_0319_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_0311_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_0227_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_0213_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_0156_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_0119_),
    .X(net230));
 sg13g2_buf_1 fanout231 (.A(_0119_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(net233),
    .X(net232));
 sg13g2_buf_1 fanout233 (.A(_0017_),
    .X(net233));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(net168));
 sg13g2_buf_2 fanout235 (.A(net237),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(net237),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(\hvsync_gen.hpos[8] ),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(net219),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(\hvsync_gen.hpos[7] ),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net241),
    .X(net240));
 sg13g2_buf_1 fanout241 (.A(net242),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(net212),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(net205),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(net245),
    .X(net244));
 sg13g2_buf_4 fanout245 (.X(net245),
    .A(\hvsync_gen.hpos[5] ));
 sg13g2_buf_2 fanout246 (.A(net247),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(\hvsync_gen.hpos[4] ),
    .X(net247));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(net250));
 sg13g2_buf_2 fanout249 (.A(net250),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(\hvsync_gen.hpos[3] ),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(net214),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(net214),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(\hvsync_gen.hpos[1] ),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(net211),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(net210),
    .X(net255));
 sg13g2_buf_1 fanout256 (.A(\hvsync_gen.vpos[7] ),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(net198),
    .X(net257));
 sg13g2_buf_1 fanout258 (.A(net198),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(net209),
    .X(net259));
 sg13g2_buf_1 fanout260 (.A(\hvsync_gen.vpos[5] ),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(net206),
    .X(net261));
 sg13g2_buf_1 fanout262 (.A(\hvsync_gen.vpos[4] ),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(net264),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(\hvsync_gen.vpos[3] ),
    .X(net264));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(net216));
 sg13g2_buf_2 fanout266 (.A(net113),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(net268),
    .X(net267));
 sg13g2_buf_1 fanout268 (.A(net195),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(net195),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(net271),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(net274),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(net274),
    .X(net272));
 sg13g2_buf_1 fanout273 (.A(net274),
    .X(net273));
 sg13g2_buf_1 fanout274 (.A(net197),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(net277),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(net277),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(\bnc_image_generator.counter[2] ),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(net279),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(\bnc_image_generator.counter[1] ),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(\bnc_image_generator.counter[0] ),
    .X(net280));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(net285));
 sg13g2_buf_1 fanout282 (.A(net285),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(net285),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(net285),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_0129_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(net288),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(net288),
    .X(net287));
 sg13g2_buf_1 fanout288 (.A(ui_in[1]),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(net1),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(net292),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(net292),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(net294),
    .X(net292));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(net294));
 sg13g2_buf_2 fanout294 (.A(rst_n),
    .X(net294));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_tiehi _1585__3 (.L_HI(net3));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0019_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0020_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0026_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0022_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0032_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0023_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0531_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0014_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold9 (.A(\vga_image_generator.character_hold[1] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0623_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold11 (.A(\vga_image_generator.character_hold[17] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0599_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold13 (.A(\vga_image_generator.character_hold[13] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0605_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold15 (.A(\hvsync_gen.vpos[1] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0033_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold17 (.A(\vga_image_generator.character_hold[14] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0604_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold19 (.A(\vga_image_generator.character_hold[0] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0624_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold21 (.A(\vga_image_generator.character_hold[16] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0688_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold23 (.A(\vga_image_generator.character_hold[6] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0617_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold25 (.A(\vga_image_generator.character_hold[5] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0618_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold27 (.A(\vga_image_generator.character_hold[8] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0612_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold29 (.A(\vga_image_generator.counter[19] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0660_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0078_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold32 (.A(\vga_image_generator.counter[17] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0656_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold34 (.A(\vga_image_generator.character_hold[2] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0622_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold36 (.A(\vga_image_generator.character_hold[11] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0609_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold38 (.A(\vga_image_generator.counter[14] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0650_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0073_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold41 (.A(\vga_image_generator.character_hold[7] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0616_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold43 (.A(\vga_image_generator.character_hold[9] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0611_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold45 (.A(\vga_image_generator.character_hold[3] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0621_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold47 (.A(\vga_image_generator.character_hold[15] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0602_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold49 (.A(\vga_image_generator.counter[18] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold50 (.A(\vga_image_generator.counter[16] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0075_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold52 (.A(\vga_image_generator.character_hold[12] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0607_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold54 (.A(\vga_image_generator.character_hold[4] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0619_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold56 (.A(\vga_image_generator.character_hold[10] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0610_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold58 (.A(\bnc_image_generator.counter[1] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold59 (.A(\vga_image_generator.counter[2] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0626_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0061_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold62 (.A(\vga_image_generator.counter[15] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0653_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0074_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold65 (.A(\vga_image_generator.counter[5] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0633_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0064_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold68 (.A(\vga_image_generator.counter[1] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0060_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold70 (.A(\hvsync_gen.hpos[9] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0687_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold72 (.A(\vga_image_generator.counter[12] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0648_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0071_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold75 (.A(\vga_image_generator.counter[7] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0637_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold77 (.A(\vga_image_generator.counter[6] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0636_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0065_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold80 (.A(\vga_image_generator.counter[8] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold81 (.A(\vga_image_generator.counter[13] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0649_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0024_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold84 (.A(\vga_image_generator.counter[10] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0069_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold86 (.A(\vga_image_generator.counter[26] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0085_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold88 (.A(\vga_image_generator.counter[22] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0665_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold90 (.A(\vga_image_generator.counter[27] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold91 (.A(\vga_image_generator.counter[3] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0629_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0062_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold94 (.A(\vga_image_generator.counter[9] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold95 (.A(\vga_image_generator.counter[11] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold96 (.A(\vga_image_generator.counter[23] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold97 (.A(\bnc_image_generator.counter[4] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0008_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold99 (.A(\BNC1_out[0] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold100 (.A(\hvsync_gen.vpos[6] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0563_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0016_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold103 (.A(\vga_image_generator.counter[4] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0632_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0063_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold106 (.A(\vga_image_generator.counter[25] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold107 (.A(\hvsync_gen.hpos[5] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold108 (.A(\hvsync_gen.vpos[4] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold109 (.A(\vga_image_generator.counter[21] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0025_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold111 (.A(\hvsync_gen.vpos[5] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold112 (.A(\hvsync_gen.vpos[7] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold113 (.A(\hvsync_gen.vpos[9] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold114 (.A(\hvsync_gen.hpos[6] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold115 (.A(\bnc_image_generator.counter[0] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold116 (.A(\hvsync_gen.hpos[2] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold117 (.A(\vga_image_generator.counter[20] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold118 (.A(\hvsync_gen.vpos[2] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold119 (.A(\hvsync_gen.hpos[0] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold120 (.A(\vga_image_generator.counter[24] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold121 (.A(\hvsync_gen.hpos[7] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold122 (.A(\vga_image_generator.counter[16] ),
    .X(net220));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_fill_2 FILLER_9_70 ();
 sg13g2_decap_4 FILLER_9_89 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_4 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_4 FILLER_10_49 ();
 sg13g2_fill_2 FILLER_10_53 ();
 sg13g2_decap_8 FILLER_10_176 ();
 sg13g2_decap_8 FILLER_10_183 ();
 sg13g2_decap_8 FILLER_10_190 ();
 sg13g2_fill_2 FILLER_10_197 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_4 FILLER_10_291 ();
 sg13g2_fill_1 FILLER_10_295 ();
 sg13g2_decap_8 FILLER_10_300 ();
 sg13g2_decap_8 FILLER_10_307 ();
 sg13g2_decap_8 FILLER_10_314 ();
 sg13g2_decap_8 FILLER_10_321 ();
 sg13g2_decap_8 FILLER_10_328 ();
 sg13g2_decap_8 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_fill_1 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_190 ();
 sg13g2_fill_2 FILLER_11_197 ();
 sg13g2_decap_8 FILLER_11_242 ();
 sg13g2_decap_8 FILLER_11_249 ();
 sg13g2_decap_8 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_263 ();
 sg13g2_fill_1 FILLER_11_270 ();
 sg13g2_fill_2 FILLER_11_279 ();
 sg13g2_fill_1 FILLER_11_281 ();
 sg13g2_fill_2 FILLER_11_289 ();
 sg13g2_fill_1 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_320 ();
 sg13g2_decap_8 FILLER_11_327 ();
 sg13g2_decap_8 FILLER_11_334 ();
 sg13g2_decap_4 FILLER_11_341 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_4 FILLER_12_42 ();
 sg13g2_fill_1 FILLER_12_46 ();
 sg13g2_fill_2 FILLER_12_73 ();
 sg13g2_fill_2 FILLER_12_130 ();
 sg13g2_decap_8 FILLER_12_197 ();
 sg13g2_decap_4 FILLER_12_204 ();
 sg13g2_fill_1 FILLER_12_208 ();
 sg13g2_fill_2 FILLER_12_229 ();
 sg13g2_fill_2 FILLER_12_257 ();
 sg13g2_fill_2 FILLER_12_271 ();
 sg13g2_fill_1 FILLER_12_282 ();
 sg13g2_fill_1 FILLER_12_297 ();
 sg13g2_decap_4 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_369 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_fill_2 FILLER_13_132 ();
 sg13g2_fill_1 FILLER_13_138 ();
 sg13g2_fill_1 FILLER_13_165 ();
 sg13g2_fill_2 FILLER_13_207 ();
 sg13g2_fill_1 FILLER_13_209 ();
 sg13g2_fill_2 FILLER_13_236 ();
 sg13g2_fill_2 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_248 ();
 sg13g2_fill_1 FILLER_13_258 ();
 sg13g2_fill_1 FILLER_13_285 ();
 sg13g2_fill_1 FILLER_13_291 ();
 sg13g2_fill_1 FILLER_13_348 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_fill_1 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_76 ();
 sg13g2_fill_2 FILLER_14_115 ();
 sg13g2_fill_1 FILLER_14_121 ();
 sg13g2_fill_1 FILLER_14_185 ();
 sg13g2_fill_2 FILLER_14_216 ();
 sg13g2_fill_1 FILLER_14_230 ();
 sg13g2_fill_2 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_4 FILLER_15_42 ();
 sg13g2_fill_2 FILLER_15_46 ();
 sg13g2_fill_2 FILLER_15_122 ();
 sg13g2_fill_2 FILLER_15_180 ();
 sg13g2_fill_2 FILLER_15_190 ();
 sg13g2_fill_1 FILLER_15_271 ();
 sg13g2_fill_1 FILLER_15_286 ();
 sg13g2_fill_1 FILLER_15_317 ();
 sg13g2_fill_2 FILLER_15_344 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_4 FILLER_16_49 ();
 sg13g2_fill_1 FILLER_16_144 ();
 sg13g2_fill_2 FILLER_16_175 ();
 sg13g2_fill_1 FILLER_16_177 ();
 sg13g2_fill_1 FILLER_16_192 ();
 sg13g2_fill_1 FILLER_16_202 ();
 sg13g2_fill_2 FILLER_16_235 ();
 sg13g2_fill_1 FILLER_16_237 ();
 sg13g2_fill_2 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_259 ();
 sg13g2_decap_4 FILLER_16_313 ();
 sg13g2_fill_2 FILLER_16_329 ();
 sg13g2_fill_1 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_341 ();
 sg13g2_fill_1 FILLER_16_348 ();
 sg13g2_fill_2 FILLER_16_359 ();
 sg13g2_fill_1 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_4 FILLER_17_42 ();
 sg13g2_fill_1 FILLER_17_46 ();
 sg13g2_fill_1 FILLER_17_82 ();
 sg13g2_fill_2 FILLER_17_88 ();
 sg13g2_fill_2 FILLER_17_121 ();
 sg13g2_fill_1 FILLER_17_141 ();
 sg13g2_fill_2 FILLER_17_172 ();
 sg13g2_fill_1 FILLER_17_200 ();
 sg13g2_fill_2 FILLER_17_231 ();
 sg13g2_fill_2 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_fill_1 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_333 ();
 sg13g2_decap_8 FILLER_17_340 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_56 ();
 sg13g2_fill_1 FILLER_18_83 ();
 sg13g2_decap_4 FILLER_18_111 ();
 sg13g2_fill_2 FILLER_18_124 ();
 sg13g2_fill_1 FILLER_18_166 ();
 sg13g2_fill_2 FILLER_18_175 ();
 sg13g2_decap_4 FILLER_18_181 ();
 sg13g2_decap_4 FILLER_18_189 ();
 sg13g2_fill_2 FILLER_18_193 ();
 sg13g2_fill_2 FILLER_18_200 ();
 sg13g2_fill_1 FILLER_18_202 ();
 sg13g2_decap_4 FILLER_18_207 ();
 sg13g2_fill_1 FILLER_18_211 ();
 sg13g2_fill_2 FILLER_18_219 ();
 sg13g2_fill_2 FILLER_18_248 ();
 sg13g2_decap_4 FILLER_18_307 ();
 sg13g2_fill_2 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_327 ();
 sg13g2_fill_2 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_fill_2 FILLER_19_63 ();
 sg13g2_fill_2 FILLER_19_78 ();
 sg13g2_decap_8 FILLER_19_85 ();
 sg13g2_fill_2 FILLER_19_92 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_decap_8 FILLER_19_109 ();
 sg13g2_decap_8 FILLER_19_116 ();
 sg13g2_fill_2 FILLER_19_123 ();
 sg13g2_fill_1 FILLER_19_125 ();
 sg13g2_fill_1 FILLER_19_141 ();
 sg13g2_fill_2 FILLER_19_151 ();
 sg13g2_decap_4 FILLER_19_188 ();
 sg13g2_fill_1 FILLER_19_192 ();
 sg13g2_decap_4 FILLER_19_213 ();
 sg13g2_fill_1 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_fill_1 FILLER_19_275 ();
 sg13g2_fill_2 FILLER_19_298 ();
 sg13g2_fill_1 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_fill_1 FILLER_20_133 ();
 sg13g2_fill_1 FILLER_20_173 ();
 sg13g2_fill_2 FILLER_20_192 ();
 sg13g2_fill_1 FILLER_20_194 ();
 sg13g2_fill_2 FILLER_20_208 ();
 sg13g2_fill_1 FILLER_20_210 ();
 sg13g2_fill_2 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_238 ();
 sg13g2_fill_2 FILLER_20_248 ();
 sg13g2_fill_1 FILLER_20_250 ();
 sg13g2_fill_2 FILLER_20_266 ();
 sg13g2_fill_1 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_291 ();
 sg13g2_fill_2 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_302 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_fill_1 FILLER_20_325 ();
 sg13g2_fill_2 FILLER_20_349 ();
 sg13g2_fill_1 FILLER_20_351 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_fill_1 FILLER_20_366 ();
 sg13g2_decap_8 FILLER_20_379 ();
 sg13g2_decap_8 FILLER_20_386 ();
 sg13g2_decap_8 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_151 ();
 sg13g2_fill_1 FILLER_21_213 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_4 FILLER_21_231 ();
 sg13g2_decap_4 FILLER_21_239 ();
 sg13g2_fill_2 FILLER_21_243 ();
 sg13g2_decap_4 FILLER_21_249 ();
 sg13g2_decap_4 FILLER_21_279 ();
 sg13g2_fill_2 FILLER_21_308 ();
 sg13g2_fill_1 FILLER_21_310 ();
 sg13g2_fill_1 FILLER_21_321 ();
 sg13g2_decap_4 FILLER_21_339 ();
 sg13g2_fill_2 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_4 FILLER_22_119 ();
 sg13g2_fill_2 FILLER_22_149 ();
 sg13g2_fill_2 FILLER_22_174 ();
 sg13g2_fill_2 FILLER_22_185 ();
 sg13g2_fill_1 FILLER_22_204 ();
 sg13g2_fill_1 FILLER_22_219 ();
 sg13g2_fill_2 FILLER_22_230 ();
 sg13g2_decap_4 FILLER_22_246 ();
 sg13g2_fill_2 FILLER_22_257 ();
 sg13g2_fill_1 FILLER_22_259 ();
 sg13g2_fill_2 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_279 ();
 sg13g2_decap_8 FILLER_22_286 ();
 sg13g2_fill_1 FILLER_22_293 ();
 sg13g2_fill_2 FILLER_22_316 ();
 sg13g2_decap_4 FILLER_22_326 ();
 sg13g2_fill_2 FILLER_22_330 ();
 sg13g2_fill_1 FILLER_22_338 ();
 sg13g2_fill_2 FILLER_22_350 ();
 sg13g2_fill_2 FILLER_22_362 ();
 sg13g2_fill_1 FILLER_22_364 ();
 sg13g2_fill_2 FILLER_22_370 ();
 sg13g2_fill_1 FILLER_22_381 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_119 ();
 sg13g2_fill_2 FILLER_23_147 ();
 sg13g2_fill_1 FILLER_23_198 ();
 sg13g2_decap_8 FILLER_23_212 ();
 sg13g2_fill_2 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_221 ();
 sg13g2_fill_1 FILLER_23_226 ();
 sg13g2_fill_2 FILLER_23_232 ();
 sg13g2_fill_1 FILLER_23_234 ();
 sg13g2_fill_2 FILLER_23_246 ();
 sg13g2_decap_8 FILLER_23_265 ();
 sg13g2_decap_4 FILLER_23_272 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_decap_8 FILLER_23_293 ();
 sg13g2_fill_2 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_310 ();
 sg13g2_decap_4 FILLER_23_326 ();
 sg13g2_fill_2 FILLER_23_330 ();
 sg13g2_fill_1 FILLER_23_337 ();
 sg13g2_decap_4 FILLER_23_343 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_367 ();
 sg13g2_fill_2 FILLER_23_395 ();
 sg13g2_fill_1 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_fill_2 FILLER_24_119 ();
 sg13g2_fill_2 FILLER_24_146 ();
 sg13g2_fill_2 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_200 ();
 sg13g2_fill_2 FILLER_24_216 ();
 sg13g2_fill_1 FILLER_24_218 ();
 sg13g2_fill_2 FILLER_24_257 ();
 sg13g2_fill_1 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_272 ();
 sg13g2_fill_2 FILLER_24_279 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_fill_2 FILLER_24_314 ();
 sg13g2_fill_1 FILLER_24_316 ();
 sg13g2_fill_1 FILLER_24_335 ();
 sg13g2_fill_2 FILLER_24_341 ();
 sg13g2_fill_1 FILLER_24_343 ();
 sg13g2_fill_1 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_4 FILLER_25_119 ();
 sg13g2_fill_2 FILLER_25_123 ();
 sg13g2_fill_2 FILLER_25_155 ();
 sg13g2_fill_2 FILLER_25_192 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_fill_1 FILLER_25_221 ();
 sg13g2_fill_1 FILLER_25_228 ();
 sg13g2_fill_2 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_235 ();
 sg13g2_decap_8 FILLER_25_279 ();
 sg13g2_decap_4 FILLER_25_286 ();
 sg13g2_fill_1 FILLER_25_290 ();
 sg13g2_fill_2 FILLER_25_296 ();
 sg13g2_decap_4 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_317 ();
 sg13g2_fill_2 FILLER_25_326 ();
 sg13g2_fill_1 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_338 ();
 sg13g2_fill_1 FILLER_25_345 ();
 sg13g2_fill_1 FILLER_25_350 ();
 sg13g2_fill_1 FILLER_25_357 ();
 sg13g2_fill_2 FILLER_25_389 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_fill_2 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_111 ();
 sg13g2_decap_8 FILLER_26_118 ();
 sg13g2_decap_8 FILLER_26_125 ();
 sg13g2_decap_4 FILLER_26_132 ();
 sg13g2_fill_2 FILLER_26_153 ();
 sg13g2_fill_1 FILLER_26_155 ();
 sg13g2_fill_2 FILLER_26_183 ();
 sg13g2_fill_1 FILLER_26_185 ();
 sg13g2_fill_2 FILLER_26_201 ();
 sg13g2_fill_1 FILLER_26_203 ();
 sg13g2_fill_2 FILLER_26_260 ();
 sg13g2_fill_1 FILLER_26_262 ();
 sg13g2_decap_4 FILLER_26_267 ();
 sg13g2_decap_4 FILLER_26_275 ();
 sg13g2_decap_4 FILLER_26_284 ();
 sg13g2_fill_1 FILLER_26_293 ();
 sg13g2_decap_8 FILLER_26_309 ();
 sg13g2_fill_2 FILLER_26_316 ();
 sg13g2_fill_1 FILLER_26_346 ();
 sg13g2_decap_4 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_78 ();
 sg13g2_fill_2 FILLER_27_89 ();
 sg13g2_fill_2 FILLER_27_143 ();
 sg13g2_fill_1 FILLER_27_145 ();
 sg13g2_decap_4 FILLER_27_192 ();
 sg13g2_fill_2 FILLER_27_204 ();
 sg13g2_decap_4 FILLER_27_211 ();
 sg13g2_decap_4 FILLER_27_241 ();
 sg13g2_decap_4 FILLER_27_270 ();
 sg13g2_fill_2 FILLER_27_280 ();
 sg13g2_fill_1 FILLER_27_293 ();
 sg13g2_decap_4 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_321 ();
 sg13g2_fill_2 FILLER_27_327 ();
 sg13g2_fill_1 FILLER_27_329 ();
 sg13g2_fill_2 FILLER_27_358 ();
 sg13g2_fill_1 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_4 FILLER_28_42 ();
 sg13g2_decap_4 FILLER_28_117 ();
 sg13g2_fill_1 FILLER_28_138 ();
 sg13g2_decap_8 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_164 ();
 sg13g2_fill_2 FILLER_28_169 ();
 sg13g2_fill_2 FILLER_28_219 ();
 sg13g2_fill_1 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_4 FILLER_28_242 ();
 sg13g2_fill_1 FILLER_28_246 ();
 sg13g2_fill_2 FILLER_28_262 ();
 sg13g2_fill_1 FILLER_28_264 ();
 sg13g2_decap_4 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_287 ();
 sg13g2_fill_1 FILLER_28_323 ();
 sg13g2_fill_2 FILLER_28_362 ();
 sg13g2_fill_2 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_55 ();
 sg13g2_fill_2 FILLER_29_61 ();
 sg13g2_fill_1 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_118 ();
 sg13g2_fill_2 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_decap_4 FILLER_29_176 ();
 sg13g2_fill_2 FILLER_29_180 ();
 sg13g2_decap_8 FILLER_29_195 ();
 sg13g2_decap_8 FILLER_29_202 ();
 sg13g2_decap_4 FILLER_29_231 ();
 sg13g2_fill_1 FILLER_29_235 ();
 sg13g2_fill_1 FILLER_29_244 ();
 sg13g2_decap_4 FILLER_29_250 ();
 sg13g2_decap_4 FILLER_29_264 ();
 sg13g2_fill_2 FILLER_29_268 ();
 sg13g2_fill_2 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_276 ();
 sg13g2_fill_1 FILLER_29_286 ();
 sg13g2_fill_2 FILLER_29_310 ();
 sg13g2_decap_4 FILLER_29_329 ();
 sg13g2_fill_1 FILLER_29_333 ();
 sg13g2_fill_2 FILLER_29_345 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_376 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_4 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_46 ();
 sg13g2_fill_2 FILLER_30_64 ();
 sg13g2_fill_1 FILLER_30_66 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_fill_2 FILLER_30_104 ();
 sg13g2_fill_2 FILLER_30_130 ();
 sg13g2_fill_1 FILLER_30_132 ();
 sg13g2_decap_8 FILLER_30_200 ();
 sg13g2_decap_4 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_221 ();
 sg13g2_fill_2 FILLER_30_234 ();
 sg13g2_fill_1 FILLER_30_236 ();
 sg13g2_decap_8 FILLER_30_249 ();
 sg13g2_fill_2 FILLER_30_256 ();
 sg13g2_fill_1 FILLER_30_258 ();
 sg13g2_decap_4 FILLER_30_272 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_decap_4 FILLER_30_298 ();
 sg13g2_fill_2 FILLER_30_302 ();
 sg13g2_decap_8 FILLER_30_309 ();
 sg13g2_decap_8 FILLER_30_323 ();
 sg13g2_decap_8 FILLER_30_330 ();
 sg13g2_decap_8 FILLER_30_352 ();
 sg13g2_decap_4 FILLER_30_359 ();
 sg13g2_fill_1 FILLER_30_363 ();
 sg13g2_fill_2 FILLER_30_372 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_4 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_59 ();
 sg13g2_fill_1 FILLER_31_67 ();
 sg13g2_fill_2 FILLER_31_93 ();
 sg13g2_fill_1 FILLER_31_100 ();
 sg13g2_fill_2 FILLER_31_111 ();
 sg13g2_decap_4 FILLER_31_132 ();
 sg13g2_fill_2 FILLER_31_146 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_fill_2 FILLER_31_217 ();
 sg13g2_decap_4 FILLER_31_231 ();
 sg13g2_fill_2 FILLER_31_240 ();
 sg13g2_fill_2 FILLER_31_278 ();
 sg13g2_fill_1 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_348 ();
 sg13g2_decap_8 FILLER_31_354 ();
 sg13g2_decap_4 FILLER_31_365 ();
 sg13g2_fill_2 FILLER_31_369 ();
 sg13g2_decap_4 FILLER_31_376 ();
 sg13g2_fill_2 FILLER_31_380 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_4 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_46 ();
 sg13g2_decap_4 FILLER_32_72 ();
 sg13g2_fill_1 FILLER_32_90 ();
 sg13g2_fill_1 FILLER_32_108 ();
 sg13g2_fill_1 FILLER_32_113 ();
 sg13g2_fill_2 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_172 ();
 sg13g2_decap_4 FILLER_32_204 ();
 sg13g2_fill_2 FILLER_32_208 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_decap_4 FILLER_32_236 ();
 sg13g2_fill_2 FILLER_32_240 ();
 sg13g2_decap_8 FILLER_32_246 ();
 sg13g2_decap_8 FILLER_32_253 ();
 sg13g2_fill_2 FILLER_32_260 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_fill_1 FILLER_32_279 ();
 sg13g2_fill_1 FILLER_32_319 ();
 sg13g2_decap_4 FILLER_32_324 ();
 sg13g2_fill_1 FILLER_32_328 ();
 sg13g2_fill_2 FILLER_32_334 ();
 sg13g2_fill_2 FILLER_32_363 ();
 sg13g2_fill_1 FILLER_32_391 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_4 FILLER_33_35 ();
 sg13g2_fill_1 FILLER_33_66 ();
 sg13g2_fill_2 FILLER_33_76 ();
 sg13g2_fill_1 FILLER_33_78 ();
 sg13g2_fill_2 FILLER_33_85 ();
 sg13g2_fill_1 FILLER_33_87 ();
 sg13g2_fill_1 FILLER_33_111 ();
 sg13g2_fill_2 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_fill_1 FILLER_33_220 ();
 sg13g2_decap_8 FILLER_33_229 ();
 sg13g2_decap_4 FILLER_33_268 ();
 sg13g2_fill_2 FILLER_33_277 ();
 sg13g2_fill_1 FILLER_33_279 ();
 sg13g2_decap_8 FILLER_33_296 ();
 sg13g2_fill_2 FILLER_33_303 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_decap_4 FILLER_33_358 ();
 sg13g2_fill_1 FILLER_33_362 ();
 sg13g2_fill_1 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_4 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_61 ();
 sg13g2_fill_1 FILLER_34_83 ();
 sg13g2_fill_2 FILLER_34_115 ();
 sg13g2_fill_1 FILLER_34_128 ();
 sg13g2_fill_2 FILLER_34_150 ();
 sg13g2_decap_4 FILLER_34_190 ();
 sg13g2_decap_4 FILLER_34_199 ();
 sg13g2_fill_2 FILLER_34_203 ();
 sg13g2_fill_1 FILLER_34_214 ();
 sg13g2_decap_8 FILLER_34_233 ();
 sg13g2_fill_1 FILLER_34_240 ();
 sg13g2_decap_8 FILLER_34_253 ();
 sg13g2_fill_2 FILLER_34_260 ();
 sg13g2_fill_1 FILLER_34_262 ();
 sg13g2_fill_2 FILLER_34_268 ();
 sg13g2_fill_2 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_277 ();
 sg13g2_decap_4 FILLER_34_293 ();
 sg13g2_fill_2 FILLER_34_297 ();
 sg13g2_decap_4 FILLER_34_318 ();
 sg13g2_fill_1 FILLER_34_343 ();
 sg13g2_fill_2 FILLER_34_359 ();
 sg13g2_decap_4 FILLER_34_367 ();
 sg13g2_fill_1 FILLER_34_371 ();
 sg13g2_fill_2 FILLER_34_398 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_4 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_53 ();
 sg13g2_fill_2 FILLER_35_64 ();
 sg13g2_fill_1 FILLER_35_66 ();
 sg13g2_fill_2 FILLER_35_72 ();
 sg13g2_fill_1 FILLER_35_74 ();
 sg13g2_decap_8 FILLER_35_96 ();
 sg13g2_decap_8 FILLER_35_103 ();
 sg13g2_fill_2 FILLER_35_115 ();
 sg13g2_fill_1 FILLER_35_117 ();
 sg13g2_fill_2 FILLER_35_122 ();
 sg13g2_decap_8 FILLER_35_127 ();
 sg13g2_decap_8 FILLER_35_134 ();
 sg13g2_fill_1 FILLER_35_141 ();
 sg13g2_fill_2 FILLER_35_150 ();
 sg13g2_decap_8 FILLER_35_156 ();
 sg13g2_fill_1 FILLER_35_163 ();
 sg13g2_decap_4 FILLER_35_168 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_decap_4 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_203 ();
 sg13g2_fill_2 FILLER_35_218 ();
 sg13g2_decap_8 FILLER_35_225 ();
 sg13g2_decap_8 FILLER_35_232 ();
 sg13g2_fill_1 FILLER_35_254 ();
 sg13g2_fill_2 FILLER_35_260 ();
 sg13g2_fill_1 FILLER_35_273 ();
 sg13g2_fill_2 FILLER_35_294 ();
 sg13g2_decap_4 FILLER_35_304 ();
 sg13g2_fill_1 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_328 ();
 sg13g2_fill_2 FILLER_35_341 ();
 sg13g2_fill_1 FILLER_35_343 ();
 sg13g2_fill_2 FILLER_35_354 ();
 sg13g2_fill_1 FILLER_35_356 ();
 sg13g2_decap_4 FILLER_35_369 ();
 sg13g2_fill_2 FILLER_35_373 ();
 sg13g2_fill_2 FILLER_35_380 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_75 ();
 sg13g2_decap_4 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_163 ();
 sg13g2_fill_1 FILLER_36_170 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_fill_2 FILLER_36_182 ();
 sg13g2_decap_4 FILLER_36_188 ();
 sg13g2_decap_4 FILLER_36_196 ();
 sg13g2_fill_1 FILLER_36_200 ();
 sg13g2_decap_4 FILLER_36_229 ();
 sg13g2_fill_1 FILLER_36_233 ();
 sg13g2_decap_4 FILLER_36_279 ();
 sg13g2_fill_2 FILLER_36_315 ();
 sg13g2_fill_2 FILLER_36_330 ();
 sg13g2_fill_1 FILLER_36_332 ();
 sg13g2_fill_1 FILLER_36_342 ();
 sg13g2_fill_2 FILLER_36_395 ();
 sg13g2_fill_1 FILLER_36_397 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_fill_2 FILLER_37_56 ();
 sg13g2_fill_1 FILLER_37_58 ();
 sg13g2_fill_1 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_76 ();
 sg13g2_decap_8 FILLER_37_116 ();
 sg13g2_decap_8 FILLER_37_127 ();
 sg13g2_decap_4 FILLER_37_134 ();
 sg13g2_decap_4 FILLER_37_143 ();
 sg13g2_fill_1 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_156 ();
 sg13g2_decap_4 FILLER_37_176 ();
 sg13g2_fill_2 FILLER_37_180 ();
 sg13g2_fill_2 FILLER_37_186 ();
 sg13g2_fill_1 FILLER_37_197 ();
 sg13g2_fill_1 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_214 ();
 sg13g2_decap_8 FILLER_37_225 ();
 sg13g2_decap_8 FILLER_37_236 ();
 sg13g2_fill_2 FILLER_37_243 ();
 sg13g2_fill_2 FILLER_37_249 ();
 sg13g2_fill_2 FILLER_37_276 ();
 sg13g2_fill_1 FILLER_37_278 ();
 sg13g2_fill_2 FILLER_37_306 ();
 sg13g2_fill_1 FILLER_37_336 ();
 sg13g2_fill_2 FILLER_37_342 ();
 sg13g2_fill_1 FILLER_37_344 ();
 sg13g2_fill_2 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_384 ();
 sg13g2_fill_2 FILLER_37_391 ();
 sg13g2_fill_1 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_91 ();
 sg13g2_fill_2 FILLER_38_101 ();
 sg13g2_fill_2 FILLER_38_138 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_167 ();
 sg13g2_decap_4 FILLER_38_197 ();
 sg13g2_fill_1 FILLER_38_201 ();
 sg13g2_decap_4 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_214 ();
 sg13g2_decap_8 FILLER_38_247 ();
 sg13g2_decap_4 FILLER_38_254 ();
 sg13g2_fill_2 FILLER_38_284 ();
 sg13g2_decap_8 FILLER_38_316 ();
 sg13g2_fill_1 FILLER_38_323 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net91;
 assign uio_oe[1] = net92;
 assign uio_oe[2] = net93;
 assign uio_oe[3] = net94;
 assign uio_oe[4] = net95;
 assign uio_oe[5] = net96;
 assign uio_oe[6] = net97;
 assign uio_oe[7] = net98;
endmodule

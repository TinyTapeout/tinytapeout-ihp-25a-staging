module tt_um_wokwi_group_2 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire \proj_10.net10 ;
 wire \proj_10.net11 ;
 wire \proj_10.net12 ;
 wire \proj_10.net13 ;
 wire \proj_10.net14 ;
 wire \proj_10.net15 ;
 wire \proj_10.net16 ;
 wire \proj_10.net17 ;
 wire \proj_10.net23 ;
 wire \proj_10.net24 ;
 wire \proj_10.net25 ;
 wire \proj_10.net26 ;
 wire \proj_10.net27 ;
 wire \proj_10.net28 ;
 wire \proj_10.net29 ;
 wire \proj_10.net30 ;
 wire \proj_10.net31 ;
 wire \proj_10.net32 ;
 wire \proj_10.net33 ;
 wire \proj_10.net34 ;
 wire \proj_10.net35 ;
 wire \proj_10.net36 ;
 wire \proj_10.net37 ;
 wire \proj_10.net38 ;
 wire \proj_10.net39 ;
 wire \proj_10.net40 ;
 wire \proj_10.net41 ;
 wire \proj_10.net42 ;
 wire \proj_10.net43 ;
 wire \proj_10.net44 ;
 wire \proj_10.net45 ;
 wire \proj_10.net46 ;
 wire \proj_11.net10 ;
 wire \proj_11.net11 ;
 wire \proj_11.net12 ;
 wire \proj_11.net13 ;
 wire \proj_11.net19 ;
 wire \proj_11.net20 ;
 wire \proj_11.net21 ;
 wire \proj_11.net22 ;
 wire \proj_11.net23 ;
 wire \proj_11.net24 ;
 wire \proj_11.net25 ;
 wire \proj_11.net26 ;
 wire \proj_11.net27 ;
 wire \proj_11.net28 ;
 wire \proj_11.net29 ;
 wire \proj_11.net30 ;
 wire \proj_11.net9 ;
 wire \proj_12.net11 ;
 wire \proj_12.net12 ;
 wire \proj_12.net13 ;
 wire \proj_12.net14 ;
 wire \proj_12.net20 ;
 wire \proj_12.net21 ;
 wire \proj_12.net22 ;
 wire \proj_13.net10 ;
 wire \proj_13.net11 ;
 wire \proj_13.net12 ;
 wire \proj_13.net13 ;
 wire \proj_13.net14 ;
 wire \proj_13.net20 ;
 wire \proj_13.net21 ;
 wire \proj_13.net22 ;
 wire \proj_13.net23 ;
 wire \proj_13.net24 ;
 wire \proj_13.net9 ;
 wire \proj_14.net100 ;
 wire \proj_14.net102 ;
 wire \proj_14.net103 ;
 wire \proj_14.net105 ;
 wire \proj_14.net106 ;
 wire \proj_14.net108 ;
 wire \proj_14.net109 ;
 wire \proj_14.net11 ;
 wire \proj_14.net111 ;
 wire \proj_14.net112 ;
 wire \proj_14.net114 ;
 wire \proj_14.net116 ;
 wire \proj_14.net118 ;
 wire \proj_14.net119 ;
 wire \proj_14.net12 ;
 wire \proj_14.net121 ;
 wire \proj_14.net122 ;
 wire \proj_14.net124 ;
 wire \proj_14.net125 ;
 wire \proj_14.net127 ;
 wire \proj_14.net128 ;
 wire \proj_14.net130 ;
 wire \proj_14.net131 ;
 wire \proj_14.net133 ;
 wire \proj_14.net134 ;
 wire \proj_14.net136 ;
 wire \proj_14.net137 ;
 wire \proj_14.net139 ;
 wire \proj_14.net14 ;
 wire \proj_14.net140 ;
 wire \proj_14.net142 ;
 wire \proj_14.net143 ;
 wire \proj_14.net145 ;
 wire \proj_14.net146 ;
 wire \proj_14.net148 ;
 wire \proj_14.net149 ;
 wire \proj_14.net15 ;
 wire \proj_14.net151 ;
 wire \proj_14.net152 ;
 wire \proj_14.net154 ;
 wire \proj_14.net155 ;
 wire \proj_14.net157 ;
 wire \proj_14.net158 ;
 wire \proj_14.net160 ;
 wire \proj_14.net161 ;
 wire \proj_14.net163 ;
 wire \proj_14.net164 ;
 wire \proj_14.net166 ;
 wire \proj_14.net167 ;
 wire \proj_14.net169 ;
 wire \proj_14.net17 ;
 wire \proj_14.net170 ;
 wire \proj_14.net172 ;
 wire \proj_14.net173 ;
 wire \proj_14.net175 ;
 wire \proj_14.net176 ;
 wire \proj_14.net178 ;
 wire \proj_14.net179 ;
 wire \proj_14.net18 ;
 wire \proj_14.net181 ;
 wire \proj_14.net182 ;
 wire \proj_14.net184 ;
 wire \proj_14.net185 ;
 wire \proj_14.net187 ;
 wire \proj_14.net188 ;
 wire \proj_14.net190 ;
 wire \proj_14.net192 ;
 wire \proj_14.net194 ;
 wire \proj_14.net195 ;
 wire \proj_14.net197 ;
 wire \proj_14.net198 ;
 wire \proj_14.net20 ;
 wire \proj_14.net200 ;
 wire \proj_14.net201 ;
 wire \proj_14.net203 ;
 wire \proj_14.net204 ;
 wire \proj_14.net206 ;
 wire \proj_14.net207 ;
 wire \proj_14.net209 ;
 wire \proj_14.net21 ;
 wire \proj_14.net210 ;
 wire \proj_14.net212 ;
 wire \proj_14.net213 ;
 wire \proj_14.net215 ;
 wire \proj_14.net216 ;
 wire \proj_14.net218 ;
 wire \proj_14.net219 ;
 wire \proj_14.net221 ;
 wire \proj_14.net222 ;
 wire \proj_14.net224 ;
 wire \proj_14.net225 ;
 wire \proj_14.net227 ;
 wire \proj_14.net228 ;
 wire \proj_14.net23 ;
 wire \proj_14.net230 ;
 wire \proj_14.net231 ;
 wire \proj_14.net233 ;
 wire \proj_14.net234 ;
 wire \proj_14.net236 ;
 wire \proj_14.net237 ;
 wire \proj_14.net239 ;
 wire \proj_14.net24 ;
 wire \proj_14.net240 ;
 wire \proj_14.net242 ;
 wire \proj_14.net243 ;
 wire \proj_14.net245 ;
 wire \proj_14.net246 ;
 wire \proj_14.net248 ;
 wire \proj_14.net249 ;
 wire \proj_14.net251 ;
 wire \proj_14.net252 ;
 wire \proj_14.net254 ;
 wire \proj_14.net256 ;
 wire \proj_14.net258 ;
 wire \proj_14.net259 ;
 wire \proj_14.net26 ;
 wire \proj_14.net261 ;
 wire \proj_14.net262 ;
 wire \proj_14.net264 ;
 wire \proj_14.net265 ;
 wire \proj_14.net267 ;
 wire \proj_14.net268 ;
 wire \proj_14.net27 ;
 wire \proj_14.net270 ;
 wire \proj_14.net271 ;
 wire \proj_14.net273 ;
 wire \proj_14.net274 ;
 wire \proj_14.net276 ;
 wire \proj_14.net277 ;
 wire \proj_14.net279 ;
 wire \proj_14.net280 ;
 wire \proj_14.net282 ;
 wire \proj_14.net283 ;
 wire \proj_14.net285 ;
 wire \proj_14.net286 ;
 wire \proj_14.net288 ;
 wire \proj_14.net289 ;
 wire \proj_14.net29 ;
 wire \proj_14.net291 ;
 wire \proj_14.net292 ;
 wire \proj_14.net294 ;
 wire \proj_14.net295 ;
 wire \proj_14.net297 ;
 wire \proj_14.net298 ;
 wire \proj_14.net30 ;
 wire \proj_14.net300 ;
 wire \proj_14.net301 ;
 wire \proj_14.net303 ;
 wire \proj_14.net304 ;
 wire \proj_14.net306 ;
 wire \proj_14.net307 ;
 wire \proj_14.net309 ;
 wire \proj_14.net310 ;
 wire \proj_14.net312 ;
 wire \proj_14.net313 ;
 wire \proj_14.net315 ;
 wire \proj_14.net316 ;
 wire \proj_14.net318 ;
 wire \proj_14.net32 ;
 wire \proj_14.net320 ;
 wire \proj_14.net322 ;
 wire \proj_14.net323 ;
 wire \proj_14.net325 ;
 wire \proj_14.net326 ;
 wire \proj_14.net328 ;
 wire \proj_14.net329 ;
 wire \proj_14.net33 ;
 wire \proj_14.net332 ;
 wire \proj_14.net333 ;
 wire \proj_14.net335 ;
 wire \proj_14.net336 ;
 wire \proj_14.net338 ;
 wire \proj_14.net339 ;
 wire \proj_14.net341 ;
 wire \proj_14.net342 ;
 wire \proj_14.net344 ;
 wire \proj_14.net345 ;
 wire \proj_14.net347 ;
 wire \proj_14.net348 ;
 wire \proj_14.net35 ;
 wire \proj_14.net350 ;
 wire \proj_14.net351 ;
 wire \proj_14.net353 ;
 wire \proj_14.net354 ;
 wire \proj_14.net356 ;
 wire \proj_14.net357 ;
 wire \proj_14.net359 ;
 wire \proj_14.net36 ;
 wire \proj_14.net360 ;
 wire \proj_14.net362 ;
 wire \proj_14.net363 ;
 wire \proj_14.net365 ;
 wire \proj_14.net366 ;
 wire \proj_14.net368 ;
 wire \proj_14.net369 ;
 wire \proj_14.net371 ;
 wire \proj_14.net372 ;
 wire \proj_14.net374 ;
 wire \proj_14.net375 ;
 wire \proj_14.net377 ;
 wire \proj_14.net378 ;
 wire \proj_14.net38 ;
 wire \proj_14.net380 ;
 wire \proj_14.net381 ;
 wire \proj_14.net383 ;
 wire \proj_14.net385 ;
 wire \proj_14.net387 ;
 wire \proj_14.net388 ;
 wire \proj_14.net39 ;
 wire \proj_14.net390 ;
 wire \proj_14.net391 ;
 wire \proj_14.net393 ;
 wire \proj_14.net394 ;
 wire \proj_14.net396 ;
 wire \proj_14.net397 ;
 wire \proj_14.net399 ;
 wire \proj_14.net4 ;
 wire \proj_14.net400 ;
 wire \proj_14.net402 ;
 wire \proj_14.net403 ;
 wire \proj_14.net405 ;
 wire \proj_14.net406 ;
 wire \proj_14.net408 ;
 wire \proj_14.net409 ;
 wire \proj_14.net41 ;
 wire \proj_14.net411 ;
 wire \proj_14.net412 ;
 wire \proj_14.net414 ;
 wire \proj_14.net415 ;
 wire \proj_14.net417 ;
 wire \proj_14.net418 ;
 wire \proj_14.net42 ;
 wire \proj_14.net420 ;
 wire \proj_14.net421 ;
 wire \proj_14.net423 ;
 wire \proj_14.net424 ;
 wire \proj_14.net426 ;
 wire \proj_14.net427 ;
 wire \proj_14.net429 ;
 wire \proj_14.net430 ;
 wire \proj_14.net432 ;
 wire \proj_14.net433 ;
 wire \proj_14.net435 ;
 wire \proj_14.net436 ;
 wire \proj_14.net438 ;
 wire \proj_14.net439 ;
 wire \proj_14.net44 ;
 wire \proj_14.net441 ;
 wire \proj_14.net442 ;
 wire \proj_14.net444 ;
 wire \proj_14.net445 ;
 wire \proj_14.net447 ;
 wire \proj_14.net449 ;
 wire \proj_14.net45 ;
 wire \proj_14.net451 ;
 wire \proj_14.net452 ;
 wire \proj_14.net454 ;
 wire \proj_14.net455 ;
 wire \proj_14.net457 ;
 wire \proj_14.net458 ;
 wire \proj_14.net460 ;
 wire \proj_14.net461 ;
 wire \proj_14.net463 ;
 wire \proj_14.net464 ;
 wire \proj_14.net466 ;
 wire \proj_14.net467 ;
 wire \proj_14.net469 ;
 wire \proj_14.net47 ;
 wire \proj_14.net470 ;
 wire \proj_14.net472 ;
 wire \proj_14.net473 ;
 wire \proj_14.net475 ;
 wire \proj_14.net476 ;
 wire \proj_14.net478 ;
 wire \proj_14.net479 ;
 wire \proj_14.net48 ;
 wire \proj_14.net481 ;
 wire \proj_14.net482 ;
 wire \proj_14.net484 ;
 wire \proj_14.net485 ;
 wire \proj_14.net487 ;
 wire \proj_14.net488 ;
 wire \proj_14.net490 ;
 wire \proj_14.net491 ;
 wire \proj_14.net493 ;
 wire \proj_14.net494 ;
 wire \proj_14.net496 ;
 wire \proj_14.net497 ;
 wire \proj_14.net499 ;
 wire \proj_14.net50 ;
 wire \proj_14.net500 ;
 wire \proj_14.net502 ;
 wire \proj_14.net503 ;
 wire \proj_14.net505 ;
 wire \proj_14.net506 ;
 wire \proj_14.net508 ;
 wire \proj_14.net509 ;
 wire \proj_14.net51 ;
 wire \proj_14.net512 ;
 wire \proj_14.net514 ;
 wire \proj_14.net515 ;
 wire \proj_14.net517 ;
 wire \proj_14.net518 ;
 wire \proj_14.net520 ;
 wire \proj_14.net521 ;
 wire \proj_14.net53 ;
 wire \proj_14.net54 ;
 wire \proj_14.net56 ;
 wire \proj_14.net57 ;
 wire \proj_14.net59 ;
 wire \proj_14.net63 ;
 wire \proj_14.net64 ;
 wire \proj_14.net66 ;
 wire \proj_14.net67 ;
 wire \proj_14.net69 ;
 wire \proj_14.net70 ;
 wire \proj_14.net72 ;
 wire \proj_14.net73 ;
 wire \proj_14.net75 ;
 wire \proj_14.net76 ;
 wire \proj_14.net78 ;
 wire \proj_14.net79 ;
 wire \proj_14.net8 ;
 wire \proj_14.net81 ;
 wire \proj_14.net82 ;
 wire \proj_14.net84 ;
 wire \proj_14.net85 ;
 wire \proj_14.net87 ;
 wire \proj_14.net88 ;
 wire \proj_14.net9 ;
 wire \proj_14.net90 ;
 wire \proj_14.net91 ;
 wire \proj_14.net93 ;
 wire \proj_14.net94 ;
 wire \proj_14.net96 ;
 wire \proj_14.net97 ;
 wire \proj_14.net99 ;
 wire \proj_15.net10 ;
 wire \proj_15.net11 ;
 wire \proj_15.net12 ;
 wire \proj_15.net13 ;
 wire \proj_15.net14 ;
 wire \proj_15.net15 ;
 wire \proj_15.net16 ;
 wire \proj_15.net9 ;
 wire \proj__0.net10 ;
 wire \proj__0.net11 ;
 wire \proj__0.net3 ;
 wire \proj__0.net4 ;
 wire \proj__1.net10 ;
 wire \proj__1.net11 ;
 wire \proj__1.net9 ;
 wire \proj__2.net14 ;
 wire \proj__2.net3 ;
 wire \proj__2.net5 ;
 wire \proj__2.net6 ;
 wire \proj__2.net7 ;
 wire \proj__3.net10 ;
 wire \proj__3.net11 ;
 wire \proj__3.net12 ;
 wire \proj__3.net13 ;
 wire \proj__3.net3 ;
 wire \proj__3.net4 ;
 wire \proj__4.net10 ;
 wire \proj__4.net11 ;
 wire \proj__4.net12 ;
 wire \proj__4.net9 ;
 wire \proj__5.net8 ;
 wire \proj__5.net9 ;
 wire \proj__6.net3 ;
 wire \proj__6.net4 ;
 wire \proj__7.net3 ;
 wire \proj__8.net10 ;
 wire \proj__8.net11 ;
 wire \proj__8.net12 ;
 wire \proj__8.net18 ;
 wire \proj__8.net19 ;
 wire \proj__8.net20 ;
 wire \proj__8.net7 ;
 wire \proj__8.net8 ;
 wire \proj__8.net9 ;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net428;
 wire \proj_10.flop1/notq ;
 wire net429;
 wire \proj_10.flop10/notq ;
 wire net430;
 wire \proj_10.flop11/notq ;
 wire net431;
 wire \proj_10.flop12/notq ;
 wire net432;
 wire \proj_10.flop13/notq ;
 wire net433;
 wire \proj_10.flop14/notq ;
 wire net434;
 wire \proj_10.flop2/notq ;
 wire net435;
 wire \proj_10.flop3/notq ;
 wire net436;
 wire \proj_10.flop4/notq ;
 wire net437;
 wire \proj_10.flop5/notq ;
 wire net438;
 wire \proj_10.flop6/notq ;
 wire net439;
 wire \proj_10.flop7/notq ;
 wire net440;
 wire \proj_10.flop8/notq ;
 wire net441;
 wire \proj_10.flop9/notq ;
 wire net442;
 wire \proj_14.flop1/notq ;
 wire net443;
 wire \proj_14.flop10/notq ;
 wire net444;
 wire \proj_14.flop100/notq ;
 wire net445;
 wire \proj_14.flop101/notq ;
 wire net446;
 wire \proj_14.flop102/notq ;
 wire net447;
 wire \proj_14.flop103/notq ;
 wire net448;
 wire \proj_14.flop104/notq ;
 wire net449;
 wire \proj_14.flop105/notq ;
 wire net450;
 wire \proj_14.flop106/notq ;
 wire net451;
 wire \proj_14.flop107/notq ;
 wire net452;
 wire \proj_14.flop108/notq ;
 wire net453;
 wire \proj_14.flop109/notq ;
 wire net454;
 wire \proj_14.flop11/notq ;
 wire net455;
 wire \proj_14.flop110/notq ;
 wire net456;
 wire \proj_14.flop111/notq ;
 wire net457;
 wire \proj_14.flop112/notq ;
 wire net458;
 wire \proj_14.flop113/notq ;
 wire net459;
 wire \proj_14.flop114/notq ;
 wire net460;
 wire \proj_14.flop115/notq ;
 wire net461;
 wire \proj_14.flop116/notq ;
 wire net462;
 wire \proj_14.flop117/notq ;
 wire net463;
 wire \proj_14.flop118/notq ;
 wire net464;
 wire \proj_14.flop119/notq ;
 wire net465;
 wire \proj_14.flop12/notq ;
 wire net466;
 wire \proj_14.flop120/notq ;
 wire net467;
 wire \proj_14.flop121/notq ;
 wire net468;
 wire \proj_14.flop122/notq ;
 wire net469;
 wire \proj_14.flop123/notq ;
 wire net470;
 wire \proj_14.flop124/notq ;
 wire net471;
 wire \proj_14.flop125/notq ;
 wire net472;
 wire \proj_14.flop126/notq ;
 wire net473;
 wire \proj_14.flop127/notq ;
 wire net474;
 wire \proj_14.flop128/notq ;
 wire net475;
 wire \proj_14.flop129/notq ;
 wire net476;
 wire \proj_14.flop13/notq ;
 wire net477;
 wire \proj_14.flop130/notq ;
 wire net478;
 wire \proj_14.flop131/notq ;
 wire net479;
 wire \proj_14.flop132/notq ;
 wire net480;
 wire \proj_14.flop133/notq ;
 wire net481;
 wire \proj_14.flop134/notq ;
 wire net482;
 wire \proj_14.flop135/notq ;
 wire net483;
 wire \proj_14.flop136/notq ;
 wire net484;
 wire \proj_14.flop137/notq ;
 wire net485;
 wire \proj_14.flop138/notq ;
 wire net486;
 wire \proj_14.flop139/notq ;
 wire net487;
 wire \proj_14.flop14/notq ;
 wire net488;
 wire \proj_14.flop140/notq ;
 wire net489;
 wire \proj_14.flop141/notq ;
 wire net490;
 wire \proj_14.flop142/notq ;
 wire net491;
 wire \proj_14.flop143/notq ;
 wire net492;
 wire \proj_14.flop144/notq ;
 wire net493;
 wire \proj_14.flop145/notq ;
 wire net494;
 wire \proj_14.flop146/notq ;
 wire net495;
 wire \proj_14.flop147/notq ;
 wire net496;
 wire \proj_14.flop148/notq ;
 wire net497;
 wire \proj_14.flop149/notq ;
 wire net498;
 wire \proj_14.flop15/notq ;
 wire net499;
 wire \proj_14.flop150/notq ;
 wire net500;
 wire \proj_14.flop151/notq ;
 wire net501;
 wire \proj_14.flop152/notq ;
 wire net502;
 wire \proj_14.flop153/notq ;
 wire net503;
 wire \proj_14.flop154/notq ;
 wire net504;
 wire \proj_14.flop155/notq ;
 wire net505;
 wire \proj_14.flop156/notq ;
 wire net506;
 wire \proj_14.flop157/notq ;
 wire net507;
 wire \proj_14.flop158/notq ;
 wire net508;
 wire \proj_14.flop159/notq ;
 wire net509;
 wire \proj_14.flop16/notq ;
 wire net510;
 wire \proj_14.flop160/notq ;
 wire net511;
 wire \proj_14.flop161/notq ;
 wire net512;
 wire \proj_14.flop162/notq ;
 wire net513;
 wire \proj_14.flop163/notq ;
 wire net514;
 wire \proj_14.flop164/notq ;
 wire net515;
 wire \proj_14.flop165/notq ;
 wire net516;
 wire \proj_14.flop166/notq ;
 wire net517;
 wire \proj_14.flop167/notq ;
 wire net518;
 wire \proj_14.flop168/notq ;
 wire net519;
 wire \proj_14.flop17/notq ;
 wire net520;
 wire \proj_14.flop18/notq ;
 wire net521;
 wire \proj_14.flop19/notq ;
 wire net522;
 wire \proj_14.flop2/notq ;
 wire net523;
 wire \proj_14.flop20/notq ;
 wire net524;
 wire \proj_14.flop21/notq ;
 wire net525;
 wire \proj_14.flop22/notq ;
 wire net526;
 wire \proj_14.flop23/notq ;
 wire net527;
 wire \proj_14.flop24/notq ;
 wire net528;
 wire \proj_14.flop25/notq ;
 wire net529;
 wire \proj_14.flop26/notq ;
 wire net530;
 wire \proj_14.flop27/notq ;
 wire net531;
 wire \proj_14.flop28/notq ;
 wire net532;
 wire \proj_14.flop29/notq ;
 wire net533;
 wire \proj_14.flop3/notq ;
 wire net534;
 wire \proj_14.flop30/notq ;
 wire net535;
 wire \proj_14.flop31/notq ;
 wire net536;
 wire \proj_14.flop32/notq ;
 wire net537;
 wire \proj_14.flop33/notq ;
 wire net538;
 wire \proj_14.flop34/notq ;
 wire net539;
 wire \proj_14.flop35/notq ;
 wire net540;
 wire \proj_14.flop36/notq ;
 wire net541;
 wire \proj_14.flop37/notq ;
 wire net542;
 wire \proj_14.flop38/notq ;
 wire net543;
 wire \proj_14.flop39/notq ;
 wire net544;
 wire \proj_14.flop4/notq ;
 wire net545;
 wire \proj_14.flop40/notq ;
 wire net546;
 wire \proj_14.flop41/notq ;
 wire net547;
 wire \proj_14.flop42/notq ;
 wire net548;
 wire \proj_14.flop43/notq ;
 wire net549;
 wire \proj_14.flop44/notq ;
 wire net550;
 wire \proj_14.flop45/notq ;
 wire net551;
 wire \proj_14.flop46/notq ;
 wire net552;
 wire \proj_14.flop47/notq ;
 wire net553;
 wire \proj_14.flop48/notq ;
 wire net554;
 wire \proj_14.flop49/notq ;
 wire net555;
 wire \proj_14.flop5/notq ;
 wire net556;
 wire \proj_14.flop50/notq ;
 wire net557;
 wire \proj_14.flop51/notq ;
 wire net558;
 wire \proj_14.flop52/notq ;
 wire net559;
 wire \proj_14.flop53/notq ;
 wire net560;
 wire \proj_14.flop54/notq ;
 wire net561;
 wire \proj_14.flop55/notq ;
 wire net562;
 wire \proj_14.flop56/notq ;
 wire net563;
 wire \proj_14.flop57/notq ;
 wire net564;
 wire \proj_14.flop58/notq ;
 wire net565;
 wire \proj_14.flop59/notq ;
 wire net566;
 wire \proj_14.flop6/notq ;
 wire net567;
 wire \proj_14.flop60/notq ;
 wire net568;
 wire \proj_14.flop61/notq ;
 wire net569;
 wire \proj_14.flop62/notq ;
 wire net570;
 wire \proj_14.flop63/notq ;
 wire net571;
 wire \proj_14.flop64/notq ;
 wire net572;
 wire \proj_14.flop65/notq ;
 wire net573;
 wire \proj_14.flop66/notq ;
 wire net574;
 wire \proj_14.flop67/notq ;
 wire net575;
 wire \proj_14.flop68/notq ;
 wire net576;
 wire \proj_14.flop69/notq ;
 wire net577;
 wire \proj_14.flop7/notq ;
 wire net578;
 wire \proj_14.flop70/notq ;
 wire net579;
 wire \proj_14.flop71/notq ;
 wire net580;
 wire \proj_14.flop72/notq ;
 wire net581;
 wire \proj_14.flop73/notq ;
 wire net582;
 wire \proj_14.flop74/notq ;
 wire net583;
 wire \proj_14.flop75/notq ;
 wire net584;
 wire \proj_14.flop76/notq ;
 wire net585;
 wire \proj_14.flop77/notq ;
 wire net586;
 wire \proj_14.flop78/notq ;
 wire net587;
 wire \proj_14.flop79/notq ;
 wire net588;
 wire \proj_14.flop8/notq ;
 wire net589;
 wire \proj_14.flop80/notq ;
 wire net590;
 wire \proj_14.flop81/notq ;
 wire net591;
 wire \proj_14.flop82/notq ;
 wire net592;
 wire \proj_14.flop83/notq ;
 wire net593;
 wire \proj_14.flop84/notq ;
 wire net594;
 wire \proj_14.flop85/notq ;
 wire net595;
 wire \proj_14.flop86/notq ;
 wire net596;
 wire \proj_14.flop87/notq ;
 wire net597;
 wire \proj_14.flop88/notq ;
 wire net598;
 wire \proj_14.flop89/notq ;
 wire net599;
 wire \proj_14.flop9/notq ;
 wire net600;
 wire \proj_14.flop90/notq ;
 wire net601;
 wire \proj_14.flop91/notq ;
 wire net602;
 wire \proj_14.flop92/notq ;
 wire net603;
 wire \proj_14.flop93/notq ;
 wire net604;
 wire \proj_14.flop94/notq ;
 wire net605;
 wire \proj_14.flop95/notq ;
 wire net606;
 wire \proj_14.flop96/notq ;
 wire net607;
 wire \proj_14.flop97/notq ;
 wire net608;
 wire \proj_14.flop98/notq ;
 wire \proj_14.flop99/notq ;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;

 sg13g2_inv_1 _427_ (.Y(_050_),
    .A(net8));
 sg13g2_inv_1 _428_ (.Y(_051_),
    .A(\proj__0.net3 ));
 sg13g2_inv_1 _429_ (.Y(_052_),
    .A(\proj__0.net4 ));
 sg13g2_nor2_2 _430_ (.A(net11),
    .B(net10),
    .Y(_053_));
 sg13g2_nor2b_2 _431_ (.A(net8),
    .B_N(net9),
    .Y(_054_));
 sg13g2_and2_1 _432_ (.A(_053_),
    .B(_054_),
    .X(_055_));
 sg13g2_nand2_1 _433_ (.Y(_056_),
    .A(\proj__2.net3 ),
    .B(_055_));
 sg13g2_nor2b_2 _434_ (.A(net11),
    .B_N(net10),
    .Y(_057_));
 sg13g2_nand3_1 _435_ (.B(net177),
    .C(_057_),
    .A(net8),
    .Y(_058_));
 sg13g2_and2_1 _436_ (.A(net11),
    .B(net10),
    .X(_059_));
 sg13g2_nor2b_1 _437_ (.A(net9),
    .B_N(net8),
    .Y(_060_));
 sg13g2_and2_2 _438_ (.A(_059_),
    .B(_060_),
    .X(_061_));
 sg13g2_nand2_1 _439_ (.Y(_062_),
    .A(\proj_13.net9 ),
    .B(_061_));
 sg13g2_nor2_1 _440_ (.A(net8),
    .B(net9),
    .Y(_063_));
 sg13g2_nor2b_1 _441_ (.A(net10),
    .B_N(net11),
    .Y(_064_));
 sg13g2_and2_2 _442_ (.A(_063_),
    .B(_064_),
    .X(_065_));
 sg13g2_and2_2 _443_ (.A(_053_),
    .B(_060_),
    .X(_066_));
 sg13g2_a22oi_1 _444_ (.Y(_067_),
    .B1(_066_),
    .B2(\proj__1.net9 ),
    .A2(_065_),
    .A1(\proj__8.net7 ));
 sg13g2_and4_1 _445_ (.A(_056_),
    .B(_058_),
    .C(_062_),
    .D(_067_),
    .X(_068_));
 sg13g2_and2_1 _446_ (.A(_054_),
    .B(_059_),
    .X(_069_));
 sg13g2_and2_2 _447_ (.A(_054_),
    .B(_064_),
    .X(_070_));
 sg13g2_a22oi_1 _448_ (.Y(_071_),
    .B1(_070_),
    .B2(\proj_10.net10 ),
    .A2(_069_),
    .A1(net7));
 sg13g2_and2_1 _449_ (.A(net8),
    .B(net9),
    .X(_000_));
 sg13g2_and2_2 _450_ (.A(_064_),
    .B(_000_),
    .X(_001_));
 sg13g2_and2_2 _451_ (.A(_059_),
    .B(_063_),
    .X(_002_));
 sg13g2_a22oi_1 _452_ (.Y(_003_),
    .B1(_002_),
    .B2(\proj_12.net11 ),
    .A2(_001_),
    .A1(\proj_11.net9 ));
 sg13g2_and2_2 _453_ (.A(_059_),
    .B(_000_),
    .X(_004_));
 sg13g2_and2_1 _454_ (.A(_054_),
    .B(_057_),
    .X(_005_));
 sg13g2_a22oi_1 _455_ (.Y(_006_),
    .B1(_005_),
    .B2(\proj__6.net3 ),
    .A2(_004_),
    .A1(\proj_15.net9 ));
 sg13g2_and2_1 _456_ (.A(_053_),
    .B(_063_),
    .X(_007_));
 sg13g2_and2_2 _457_ (.A(_057_),
    .B(_063_),
    .X(_008_));
 sg13g2_a21oi_1 _458_ (.A1(\proj__4.net9 ),
    .A2(_008_),
    .Y(_009_),
    .B1(_007_));
 sg13g2_and4_1 _459_ (.A(_071_),
    .B(_003_),
    .C(_006_),
    .D(_009_),
    .X(_010_));
 sg13g2_a22oi_1 _460_ (.Y(uo_out[0]),
    .B1(_010_),
    .B2(_068_),
    .A2(_007_),
    .A1(_051_));
 sg13g2_a22oi_1 _461_ (.Y(_011_),
    .B1(_066_),
    .B2(\proj__1.net9 ),
    .A2(_053_),
    .A1(_050_));
 sg13g2_nand3_1 _462_ (.B(_057_),
    .C(_000_),
    .A(\proj__7.net3 ),
    .Y(_012_));
 sg13g2_nand2_1 _463_ (.Y(_013_),
    .A(\proj__6.net4 ),
    .B(_005_));
 sg13g2_and2_2 _464_ (.A(_057_),
    .B(_060_),
    .X(_014_));
 sg13g2_a22oi_1 _465_ (.Y(_015_),
    .B1(_014_),
    .B2(net176),
    .A2(_070_),
    .A1(\proj_10.net11 ));
 sg13g2_and4_1 _466_ (.A(_011_),
    .B(_012_),
    .C(_013_),
    .D(_015_),
    .X(_016_));
 sg13g2_a22oi_1 _467_ (.Y(_017_),
    .B1(_004_),
    .B2(\proj_15.net10 ),
    .A2(_069_),
    .A1(net163));
 sg13g2_a22oi_1 _468_ (.Y(_018_),
    .B1(_002_),
    .B2(\proj_12.net12 ),
    .A2(_001_),
    .A1(\proj_11.net10 ));
 sg13g2_and2_1 _469_ (.A(_053_),
    .B(_000_),
    .X(_019_));
 sg13g2_a22oi_1 _470_ (.Y(_020_),
    .B1(_019_),
    .B2(\proj__3.net3 ),
    .A2(_061_),
    .A1(\proj_13.net10 ));
 sg13g2_a22oi_1 _471_ (.Y(_021_),
    .B1(_008_),
    .B2(\proj__4.net10 ),
    .A2(_065_),
    .A1(\proj__8.net8 ));
 sg13g2_and4_1 _472_ (.A(_017_),
    .B(_018_),
    .C(_020_),
    .D(_021_),
    .X(_022_));
 sg13g2_a22oi_1 _473_ (.Y(uo_out[1]),
    .B1(_016_),
    .B2(_022_),
    .A2(_007_),
    .A1(_052_));
 sg13g2_a22oi_1 _474_ (.Y(_023_),
    .B1(_014_),
    .B2(net172),
    .A2(_066_),
    .A1(\proj__1.net10 ));
 sg13g2_a22oi_1 _475_ (.Y(_024_),
    .B1(_004_),
    .B2(\proj_15.net11 ),
    .A2(_070_),
    .A1(\proj_10.net12 ));
 sg13g2_a22oi_1 _476_ (.Y(_025_),
    .B1(_001_),
    .B2(\proj_11.net11 ),
    .A2(_065_),
    .A1(\proj__8.net8 ));
 sg13g2_a22oi_1 _477_ (.Y(_026_),
    .B1(_008_),
    .B2(\proj__4.net11 ),
    .A2(_002_),
    .A1(\proj_12.net13 ));
 sg13g2_and3_1 _478_ (.X(_027_),
    .A(_024_),
    .B(_025_),
    .C(_026_));
 sg13g2_a22oi_1 _479_ (.Y(_028_),
    .B1(_061_),
    .B2(\proj_13.net11 ),
    .A2(_055_),
    .A1(\proj__2.net5 ));
 sg13g2_nand3_1 _480_ (.B(_027_),
    .C(_028_),
    .A(_023_),
    .Y(uo_out[2]));
 sg13g2_nand2_1 _481_ (.Y(_029_),
    .A(\proj_13.net12 ),
    .B(_061_));
 sg13g2_a22oi_1 _482_ (.Y(_030_),
    .B1(_008_),
    .B2(\proj__4.net12 ),
    .A2(_002_),
    .A1(\proj_12.net14 ));
 sg13g2_a22oi_1 _483_ (.Y(_031_),
    .B1(_014_),
    .B2(\proj__5.net8 ),
    .A2(_070_),
    .A1(\proj_10.net13 ));
 sg13g2_and4_1 _484_ (.A(_056_),
    .B(_029_),
    .C(_030_),
    .D(_031_),
    .X(_032_));
 sg13g2_a22oi_1 _485_ (.Y(_033_),
    .B1(_001_),
    .B2(\proj_11.net12 ),
    .A2(_065_),
    .A1(\proj__8.net9 ));
 sg13g2_a22oi_1 _486_ (.Y(_034_),
    .B1(_004_),
    .B2(\proj_15.net12 ),
    .A2(_066_),
    .A1(\proj__1.net11 ));
 sg13g2_nand3_1 _487_ (.B(_033_),
    .C(_034_),
    .A(_032_),
    .Y(uo_out[3]));
 sg13g2_a22oi_1 _488_ (.Y(_035_),
    .B1(_004_),
    .B2(\proj_15.net13 ),
    .A2(_065_),
    .A1(\proj__8.net10 ));
 sg13g2_or2_2 _489_ (.X(_036_),
    .B(_008_),
    .A(_066_));
 sg13g2_a22oi_1 _490_ (.Y(_037_),
    .B1(_001_),
    .B2(\proj_11.net13 ),
    .A2(_070_),
    .A1(\proj_10.net14 ));
 sg13g2_a22oi_1 _491_ (.Y(_038_),
    .B1(_036_),
    .B2(net170),
    .A2(_014_),
    .A1(\proj__5.net8 ));
 sg13g2_nand4_1 _492_ (.B(_035_),
    .C(_037_),
    .A(_056_),
    .Y(uo_out[4]),
    .D(_038_));
 sg13g2_o21ai_1 _493_ (.B1(net169),
    .Y(_039_),
    .A1(_014_),
    .A2(_036_));
 sg13g2_a22oi_1 _494_ (.Y(_040_),
    .B1(_004_),
    .B2(\proj_15.net14 ),
    .A2(_065_),
    .A1(\proj__8.net11 ));
 sg13g2_a22oi_1 _495_ (.Y(_041_),
    .B1(_070_),
    .B2(\proj_10.net15 ),
    .A2(_055_),
    .A1(\proj__2.net6 ));
 sg13g2_a22oi_1 _496_ (.Y(_042_),
    .B1(_019_),
    .B2(\proj__3.net4 ),
    .A2(_061_),
    .A1(\proj_13.net13 ));
 sg13g2_nand4_1 _497_ (.B(_040_),
    .C(_041_),
    .A(_039_),
    .Y(uo_out[5]),
    .D(_042_));
 sg13g2_a22oi_1 _498_ (.Y(_043_),
    .B1(_036_),
    .B2(net151),
    .A2(_070_),
    .A1(\proj_10.net16 ));
 sg13g2_a22oi_1 _499_ (.Y(_044_),
    .B1(_004_),
    .B2(\proj_15.net15 ),
    .A2(_065_),
    .A1(\proj__8.net12 ));
 sg13g2_a22oi_1 _500_ (.Y(_045_),
    .B1(_014_),
    .B2(\proj__5.net9 ),
    .A2(_055_),
    .A1(\proj__2.net7 ));
 sg13g2_and2_1 _501_ (.A(_044_),
    .B(_045_),
    .X(_046_));
 sg13g2_nand3_1 _502_ (.B(_043_),
    .C(_046_),
    .A(_029_),
    .Y(uo_out[6]));
 sg13g2_a22oi_1 _503_ (.Y(_047_),
    .B1(_004_),
    .B2(\proj_15.net16 ),
    .A2(_061_),
    .A1(\proj_13.net14 ));
 sg13g2_nand2_1 _504_ (.Y(_048_),
    .A(\proj_14.net4 ),
    .B(_069_));
 sg13g2_a22oi_1 _505_ (.Y(_049_),
    .B1(_036_),
    .B2(net135),
    .A2(_070_),
    .A1(\proj_10.net17 ));
 sg13g2_nand3_1 _506_ (.B(_048_),
    .C(_049_),
    .A(_047_),
    .Y(uo_out[7]));
 sg13g2_tiehi \proj_14.mux100/_0__263  (.L_HI(net307));
 sg13g2_tiehi \proj_14.mux101/_0__264  (.L_HI(net308));
 sg13g2_tiehi \proj_14.mux102/_0__265  (.L_HI(net309));
 sg13g2_tiehi \proj_14.mux103/_0__266  (.L_HI(net310));
 sg13g2_tiehi \proj_14.mux104/_0__267  (.L_HI(net311));
 sg13g2_tiehi \proj_14.mux105/_0__268  (.L_HI(net312));
 sg13g2_tiehi \proj_14.mux106/_0__269  (.L_HI(net313));
 sg13g2_tiehi \proj_14.mux107/_0__270  (.L_HI(net314));
 sg13g2_tiehi \proj_14.mux108/_0__271  (.L_HI(net315));
 sg13g2_tiehi \proj_14.mux109/_0__272  (.L_HI(net316));
 sg13g2_tiehi \proj_14.mux11/_0__273  (.L_HI(net317));
 sg13g2_tiehi \proj_14.mux110/_0__274  (.L_HI(net318));
 sg13g2_tiehi \proj_14.mux112/_0__275  (.L_HI(net319));
 sg13g2_tiehi \proj_14.mux118/_0__276  (.L_HI(net320));
 sg13g2_tiehi \proj_14.mux120/_0__277  (.L_HI(net321));
 sg13g2_tiehi \proj_14.mux121/_0__278  (.L_HI(net322));
 sg13g2_tiehi \proj_14.mux122/_0__279  (.L_HI(net323));
 sg13g2_tiehi \proj_14.mux123/_0__280  (.L_HI(net324));
 sg13g2_tiehi \proj_14.mux124/_0__281  (.L_HI(net325));
 sg13g2_tiehi \proj_14.mux125/_0__282  (.L_HI(net326));
 sg13g2_tiehi \proj_14.mux126/_0__283  (.L_HI(net327));
 sg13g2_tiehi \proj_14.mux127/_0__284  (.L_HI(net328));
 sg13g2_tiehi \proj_14.mux128/_0__285  (.L_HI(net329));
 sg13g2_tiehi \proj_14.mux129/_0__286  (.L_HI(net330));
 sg13g2_tiehi \proj_14.mux13/_0__287  (.L_HI(net331));
 sg13g2_tiehi \proj_14.mux130/_0__288  (.L_HI(net332));
 sg13g2_tiehi \proj_14.mux131/_0__289  (.L_HI(net333));
 sg13g2_tiehi \proj_14.mux133/_0__290  (.L_HI(net334));
 sg13g2_tiehi \proj_14.mux136/_0__291  (.L_HI(net335));
 sg13g2_tiehi \proj_14.mux139/_0__292  (.L_HI(net336));
 sg13g2_tiehi \proj_14.mux141/_0__293  (.L_HI(net337));
 sg13g2_tiehi \proj_14.mux142/_0__294  (.L_HI(net338));
 sg13g2_tiehi \proj_14.mux143/_0__295  (.L_HI(net339));
 sg13g2_tiehi \proj_14.mux144/_0__296  (.L_HI(net340));
 sg13g2_tiehi \proj_14.mux145/_0__297  (.L_HI(net341));
 sg13g2_tiehi \proj_14.mux146/_0__298  (.L_HI(net342));
 sg13g2_tiehi \proj_14.mux147/_0__299  (.L_HI(net343));
 sg13g2_tiehi \proj_14.mux148/_0__300  (.L_HI(net344));
 sg13g2_tiehi \proj_14.mux149/_0__301  (.L_HI(net345));
 sg13g2_tiehi \proj_14.mux15/_0__302  (.L_HI(net346));
 sg13g2_tiehi \proj_14.mux150/_0__303  (.L_HI(net347));
 sg13g2_tiehi \proj_14.mux151/_0__304  (.L_HI(net348));
 sg13g2_tiehi \proj_14.mux152/_0__305  (.L_HI(net349));
 sg13g2_tiehi \proj_14.mux155/_0__306  (.L_HI(net350));
 sg13g2_tiehi \proj_14.mux157/_0__307  (.L_HI(net351));
 sg13g2_tiehi \proj_14.mux16/_0__308  (.L_HI(net352));
 sg13g2_tiehi \proj_14.mux162/_0__309  (.L_HI(net353));
 sg13g2_tiehi \proj_14.mux163/_0__310  (.L_HI(net354));
 sg13g2_tiehi \proj_14.mux164/_0__311  (.L_HI(net355));
 sg13g2_tiehi \proj_14.mux165/_0__312  (.L_HI(net356));
 sg13g2_tiehi \proj_14.mux166/_0__313  (.L_HI(net357));
 sg13g2_tiehi \proj_14.mux167/_0__314  (.L_HI(net358));
 sg13g2_tiehi \proj_14.mux168/_0__315  (.L_HI(net359));
 sg13g2_tiehi \proj_14.mux169/_0__316  (.L_HI(net360));
 sg13g2_tiehi \proj_14.mux17/_0__317  (.L_HI(net361));
 sg13g2_tiehi \proj_14.mux18/_0__318  (.L_HI(net362));
 sg13g2_tiehi \proj_14.mux19/_0__319  (.L_HI(net363));
 sg13g2_tiehi \proj_14.mux2/_0__320  (.L_HI(net364));
 sg13g2_tiehi \proj_14.mux20/_0__321  (.L_HI(net365));
 sg13g2_tiehi \proj_14.mux21/_0__322  (.L_HI(net366));
 sg13g2_tiehi \proj_14.mux22/_0__323  (.L_HI(net367));
 sg13g2_tiehi \proj_14.mux27/_0__324  (.L_HI(net368));
 sg13g2_tiehi \proj_14.mux3/_0__325  (.L_HI(net369));
 sg13g2_tiehi \proj_14.mux30/_0__326  (.L_HI(net370));
 sg13g2_tiehi \proj_14.mux32/_0__327  (.L_HI(net371));
 sg13g2_tiehi \proj_14.mux33/_0__328  (.L_HI(net372));
 sg13g2_tiehi \proj_14.mux34/_0__329  (.L_HI(net373));
 sg13g2_tiehi \proj_14.mux35/_0__330  (.L_HI(net374));
 sg13g2_tiehi \proj_14.mux36/_0__331  (.L_HI(net375));
 sg13g2_tiehi \proj_14.mux37/_0__332  (.L_HI(net376));
 sg13g2_tiehi \proj_14.mux38/_0__333  (.L_HI(net377));
 sg13g2_tiehi \proj_14.mux39/_0__334  (.L_HI(net378));
 sg13g2_tiehi \proj_14.mux4/_0__335  (.L_HI(net379));
 sg13g2_tiehi \proj_14.mux40/_0__336  (.L_HI(net380));
 sg13g2_tiehi \proj_14.mux41/_0__337  (.L_HI(net381));
 sg13g2_tiehi \proj_14.mux42/_0__338  (.L_HI(net382));
 sg13g2_tiehi \proj_14.mux43/_0__339  (.L_HI(net383));
 sg13g2_tiehi \proj_14.mux44/_0__340  (.L_HI(net384));
 sg13g2_tiehi \proj_14.mux45/_0__341  (.L_HI(net385));
 sg13g2_tiehi \proj_14.mux46/_0__342  (.L_HI(net386));
 sg13g2_tiehi \proj_14.mux47/_0__343  (.L_HI(net387));
 sg13g2_tiehi \proj_14.mux49/_0__344  (.L_HI(net388));
 sg13g2_tiehi \proj_14.mux5/_0__345  (.L_HI(net389));
 sg13g2_tiehi \proj_14.mux55/_0__346  (.L_HI(net390));
 sg13g2_tiehi \proj_14.mux57/_0__347  (.L_HI(net391));
 sg13g2_tiehi \proj_14.mux58/_0__348  (.L_HI(net392));
 sg13g2_tiehi \proj_14.mux59/_0__349  (.L_HI(net393));
 sg13g2_tiehi \proj_14.mux60/_0__350  (.L_HI(net394));
 sg13g2_tiehi \proj_14.mux61/_0__351  (.L_HI(net395));
 sg13g2_tiehi \proj_14.mux62/_0__352  (.L_HI(net396));
 sg13g2_tiehi \proj_14.mux63/_0__353  (.L_HI(net397));
 sg13g2_tiehi \proj_14.mux64/_0__354  (.L_HI(net398));
 sg13g2_tiehi \proj_14.mux65/_0__355  (.L_HI(net399));
 sg13g2_tiehi \proj_14.mux66/_0__356  (.L_HI(net400));
 sg13g2_tiehi \proj_14.mux67/_0__357  (.L_HI(net401));
 sg13g2_tiehi \proj_14.mux68/_0__358  (.L_HI(net402));
 sg13g2_tiehi \proj_14.mux7/_0__359  (.L_HI(net403));
 sg13g2_tiehi \proj_14.mux70/_0__360  (.L_HI(net404));
 sg13g2_tiehi \proj_14.mux71/_0__361  (.L_HI(net405));
 sg13g2_tiehi \proj_14.mux72/_0__362  (.L_HI(net406));
 sg13g2_tiehi \proj_14.mux73/_0__363  (.L_HI(net407));
 sg13g2_tiehi \proj_14.mux76/_0__364  (.L_HI(net408));
 sg13g2_tiehi \proj_14.mux78/_0__365  (.L_HI(net409));
 sg13g2_tiehi \proj_14.mux79/_0__366  (.L_HI(net410));
 sg13g2_tiehi \proj_14.mux8/_0__367  (.L_HI(net411));
 sg13g2_tiehi \proj_14.mux80/_0__368  (.L_HI(net412));
 sg13g2_tiehi \proj_14.mux81/_0__369  (.L_HI(net413));
 sg13g2_tiehi \proj_14.mux82/_0__370  (.L_HI(net414));
 sg13g2_tiehi \proj_14.mux83/_0__371  (.L_HI(net415));
 sg13g2_tiehi \proj_14.mux84/_0__372  (.L_HI(net416));
 sg13g2_tiehi \proj_14.mux85/_0__373  (.L_HI(net417));
 sg13g2_tiehi \proj_14.mux86/_0__374  (.L_HI(net418));
 sg13g2_tiehi \proj_14.mux87/_0__375  (.L_HI(net419));
 sg13g2_tiehi \proj_14.mux88/_0__376  (.L_HI(net420));
 sg13g2_tiehi \proj_14.mux89/_0__377  (.L_HI(net421));
 sg13g2_tiehi \proj_14.mux91/_0__378  (.L_HI(net422));
 sg13g2_tiehi \proj_14.mux92/_0__379  (.L_HI(net423));
 sg13g2_tiehi \proj_14.mux94/_0__380  (.L_HI(net424));
 sg13g2_tiehi \proj_14.mux97/_0__381  (.L_HI(net425));
 sg13g2_tiehi \proj_14.mux99/_0__382  (.L_HI(net426));
 sg13g2_tiehi \proj_10.flop1/_1__383  (.L_HI(net427));
 sg13g2_tielo \proj_10.flop10/_1__13  (.L_LO(net13));
 sg13g2_tielo \proj_10.flop11/_1__14  (.L_LO(net14));
 sg13g2_tielo \proj_10.flop12/_1__15  (.L_LO(net15));
 sg13g2_tielo \proj_10.flop13/_1__16  (.L_LO(net16));
 sg13g2_tielo \proj_10.flop14/_1__17  (.L_LO(net17));
 sg13g2_tielo \proj_10.flop2/_1__18  (.L_LO(net18));
 sg13g2_tielo \proj_10.flop3/_1__19  (.L_LO(net19));
 sg13g2_tielo \proj_10.flop4/_1__20  (.L_LO(net20));
 sg13g2_tielo \proj_10.flop5/_1__21  (.L_LO(net21));
 sg13g2_tielo \proj_10.flop6/_1__22  (.L_LO(net22));
 sg13g2_tielo \proj_10.flop7/_1__23  (.L_LO(net23));
 sg13g2_tielo \proj_10.flop8/_1__24  (.L_LO(net24));
 sg13g2_tielo \proj_10.flop9/_1__25  (.L_LO(net25));
 sg13g2_tielo \proj_10.xor1/_0__26  (.L_LO(net26));
 sg13g2_tielo \proj_10.xor1/_0__27  (.L_LO(net27));
 sg13g2_tielo \proj_12.nand1/_0__28  (.L_LO(net28));
 sg13g2_tielo \proj_12.nand1/_0__29  (.L_LO(net29));
 sg13g2_tielo \proj_14.flop1/_1__30  (.L_LO(net30));
 sg13g2_tielo \proj_14.flop10/_1__31  (.L_LO(net31));
 sg13g2_tielo \proj_14.flop100/_1__32  (.L_LO(net32));
 sg13g2_tielo \proj_14.flop101/_1__33  (.L_LO(net33));
 sg13g2_tielo \proj_14.flop102/_1__34  (.L_LO(net34));
 sg13g2_tielo \proj_14.flop103/_1__35  (.L_LO(net35));
 sg13g2_tielo \proj_14.flop104/_1__36  (.L_LO(net36));
 sg13g2_tielo \proj_14.flop105/_1__37  (.L_LO(net37));
 sg13g2_tielo \proj_14.flop106/_1__38  (.L_LO(net38));
 sg13g2_tielo \proj_14.flop107/_1__39  (.L_LO(net39));
 sg13g2_tielo \proj_14.flop108/_1__40  (.L_LO(net40));
 sg13g2_tielo \proj_14.flop109/_1__41  (.L_LO(net41));
 sg13g2_tielo \proj_14.flop11/_1__42  (.L_LO(net42));
 sg13g2_tielo \proj_14.flop110/_1__43  (.L_LO(net43));
 sg13g2_tielo \proj_14.flop111/_1__44  (.L_LO(net44));
 sg13g2_tielo \proj_14.flop112/_1__45  (.L_LO(net45));
 sg13g2_tielo \proj_14.flop113/_1__46  (.L_LO(net46));
 sg13g2_tielo \proj_14.flop114/_1__47  (.L_LO(net47));
 sg13g2_tielo \proj_14.flop115/_1__48  (.L_LO(net48));
 sg13g2_tielo \proj_14.flop116/_1__49  (.L_LO(net49));
 sg13g2_tielo \proj_14.flop117/_1__50  (.L_LO(net50));
 sg13g2_tielo \proj_14.flop118/_1__51  (.L_LO(net51));
 sg13g2_tielo \proj_14.flop119/_1__52  (.L_LO(net52));
 sg13g2_tielo \proj_14.flop12/_1__53  (.L_LO(net53));
 sg13g2_tielo \proj_14.flop120/_1__54  (.L_LO(net54));
 sg13g2_tielo \proj_14.flop121/_1__55  (.L_LO(net55));
 sg13g2_tielo \proj_14.flop122/_1__56  (.L_LO(net56));
 sg13g2_tielo \proj_14.flop123/_1__57  (.L_LO(net57));
 sg13g2_tielo \proj_14.flop124/_1__58  (.L_LO(net58));
 sg13g2_tielo \proj_14.flop125/_1__59  (.L_LO(net59));
 sg13g2_tielo \proj_14.flop126/_1__60  (.L_LO(net60));
 sg13g2_tielo \proj_14.flop127/_1__61  (.L_LO(net61));
 sg13g2_tielo \proj_14.flop128/_1__62  (.L_LO(net62));
 sg13g2_tielo \proj_14.flop129/_1__63  (.L_LO(net63));
 sg13g2_tielo \proj_14.flop13/_1__64  (.L_LO(net64));
 sg13g2_tielo \proj_14.flop130/_1__65  (.L_LO(net65));
 sg13g2_tielo \proj_14.flop131/_1__66  (.L_LO(net66));
 sg13g2_tielo \proj_14.flop132/_1__67  (.L_LO(net67));
 sg13g2_tielo \proj_14.flop133/_1__68  (.L_LO(net68));
 sg13g2_tielo \proj_14.flop134/_1__69  (.L_LO(net69));
 sg13g2_tielo \proj_14.flop135/_1__70  (.L_LO(net70));
 sg13g2_tielo \proj_14.flop136/_1__71  (.L_LO(net71));
 sg13g2_tielo \proj_14.flop137/_1__72  (.L_LO(net72));
 sg13g2_tielo \proj_14.flop138/_1__73  (.L_LO(net73));
 sg13g2_tielo \proj_14.flop139/_1__74  (.L_LO(net74));
 sg13g2_tielo \proj_14.flop14/_1__75  (.L_LO(net75));
 sg13g2_tielo \proj_14.flop140/_1__76  (.L_LO(net76));
 sg13g2_tielo \proj_14.flop141/_1__77  (.L_LO(net77));
 sg13g2_tielo \proj_14.flop142/_1__78  (.L_LO(net78));
 sg13g2_tielo \proj_14.flop143/_1__79  (.L_LO(net79));
 sg13g2_tielo \proj_14.flop144/_1__80  (.L_LO(net80));
 sg13g2_tielo \proj_14.flop145/_1__81  (.L_LO(net81));
 sg13g2_tielo \proj_14.flop146/_1__82  (.L_LO(net82));
 sg13g2_tielo \proj_14.flop147/_1__83  (.L_LO(net83));
 sg13g2_tielo \proj_14.flop148/_1__84  (.L_LO(net84));
 sg13g2_tielo \proj_14.flop149/_1__85  (.L_LO(net85));
 sg13g2_tielo \proj_14.flop15/_1__86  (.L_LO(net86));
 sg13g2_tielo \proj_14.flop150/_1__87  (.L_LO(net87));
 sg13g2_tielo \proj_14.flop151/_1__88  (.L_LO(net88));
 sg13g2_tielo \proj_14.flop152/_1__89  (.L_LO(net89));
 sg13g2_tielo \proj_14.flop153/_1__90  (.L_LO(net90));
 sg13g2_tielo \proj_14.flop154/_1__91  (.L_LO(net91));
 sg13g2_tielo \proj_14.flop155/_1__92  (.L_LO(net92));
 sg13g2_tielo \proj_14.flop156/_1__93  (.L_LO(net93));
 sg13g2_tielo \proj_14.flop157/_1__94  (.L_LO(net94));
 sg13g2_tielo \proj_14.flop158/_1__95  (.L_LO(net95));
 sg13g2_tielo \proj_14.flop159/_1__96  (.L_LO(net96));
 sg13g2_tielo \proj_14.flop16/_1__97  (.L_LO(net97));
 sg13g2_tielo \proj_14.flop160/_1__98  (.L_LO(net98));
 sg13g2_tielo \proj_14.flop161/_1__99  (.L_LO(net99));
 sg13g2_tielo \proj_14.flop162/_1__100  (.L_LO(net100));
 sg13g2_tielo \proj_14.flop163/_1__101  (.L_LO(net101));
 sg13g2_tielo \proj_14.flop164/_1__102  (.L_LO(net102));
 sg13g2_tielo \proj_14.flop165/_1__103  (.L_LO(net103));
 sg13g2_tielo \proj_14.flop166/_1__104  (.L_LO(net104));
 sg13g2_tielo \proj_14.flop167/_1__105  (.L_LO(net105));
 sg13g2_tielo \proj_14.flop168/_1__106  (.L_LO(net106));
 sg13g2_tielo \proj_14.flop17/_1__107  (.L_LO(net107));
 sg13g2_tielo \proj_14.flop18/_1__108  (.L_LO(net108));
 sg13g2_tielo \proj_14.flop19/_1__109  (.L_LO(net109));
 sg13g2_tielo \proj_14.flop2/_1__110  (.L_LO(net110));
 sg13g2_tielo \proj_14.flop20/_1__111  (.L_LO(net111));
 sg13g2_tielo \proj_14.flop21/_1__112  (.L_LO(net112));
 sg13g2_tielo \proj_14.flop22/_1__113  (.L_LO(net113));
 sg13g2_tielo \proj_14.flop23/_1__114  (.L_LO(net114));
 sg13g2_tielo \proj_14.flop24/_1__115  (.L_LO(net115));
 sg13g2_tielo \proj_14.flop25/_1__116  (.L_LO(net116));
 sg13g2_tielo \proj_14.flop26/_1__117  (.L_LO(net117));
 sg13g2_tielo \proj_14.flop27/_1__118  (.L_LO(net118));
 sg13g2_tielo \proj_14.flop28/_1__119  (.L_LO(net119));
 sg13g2_tielo \proj_14.flop29/_1__120  (.L_LO(net120));
 sg13g2_tielo \proj_14.flop3/_1__121  (.L_LO(net121));
 sg13g2_tielo \proj_14.flop30/_1__122  (.L_LO(net122));
 sg13g2_tielo \proj_14.flop31/_1__123  (.L_LO(net123));
 sg13g2_tielo \proj_14.flop32/_1__124  (.L_LO(net124));
 sg13g2_tielo \proj_14.flop33/_1__125  (.L_LO(net125));
 sg13g2_tielo \proj_14.flop34/_1__126  (.L_LO(net126));
 sg13g2_tielo \proj_14.flop35/_1__127  (.L_LO(net127));
 sg13g2_tielo \proj_14.flop36/_1__128  (.L_LO(net128));
 sg13g2_tielo \proj_14.flop37/_1__129  (.L_LO(net129));
 sg13g2_tielo \proj_14.flop38/_1__130  (.L_LO(net130));
 sg13g2_tielo \proj_14.flop39/_1__131  (.L_LO(net131));
 sg13g2_tielo \proj_14.flop4/_1__132  (.L_LO(net132));
 sg13g2_tielo \proj_14.flop40/_1__133  (.L_LO(net133));
 sg13g2_tielo \proj_14.flop41/_1__134  (.L_LO(net134));
 sg13g2_tielo \proj_14.flop42/_1__135  (.L_LO(net179));
 sg13g2_tielo \proj_14.flop43/_1__136  (.L_LO(net180));
 sg13g2_tielo \proj_14.flop44/_1__137  (.L_LO(net181));
 sg13g2_tielo \proj_14.flop45/_1__138  (.L_LO(net182));
 sg13g2_tielo \proj_14.flop46/_1__139  (.L_LO(net183));
 sg13g2_tielo \proj_14.flop47/_1__140  (.L_LO(net184));
 sg13g2_tielo \proj_14.flop48/_1__141  (.L_LO(net185));
 sg13g2_tielo \proj_14.flop49/_1__142  (.L_LO(net186));
 sg13g2_tielo \proj_14.flop5/_1__143  (.L_LO(net187));
 sg13g2_tielo \proj_14.flop50/_1__144  (.L_LO(net188));
 sg13g2_tielo \proj_14.flop51/_1__145  (.L_LO(net189));
 sg13g2_tielo \proj_14.flop52/_1__146  (.L_LO(net190));
 sg13g2_tielo \proj_14.flop53/_1__147  (.L_LO(net191));
 sg13g2_tielo \proj_14.flop54/_1__148  (.L_LO(net192));
 sg13g2_tielo \proj_14.flop55/_1__149  (.L_LO(net193));
 sg13g2_tielo \proj_14.flop56/_1__150  (.L_LO(net194));
 sg13g2_tielo \proj_14.flop57/_1__151  (.L_LO(net195));
 sg13g2_tielo \proj_14.flop58/_1__152  (.L_LO(net196));
 sg13g2_tielo \proj_14.flop59/_1__153  (.L_LO(net197));
 sg13g2_tielo \proj_14.flop6/_1__154  (.L_LO(net198));
 sg13g2_tielo \proj_14.flop60/_1__155  (.L_LO(net199));
 sg13g2_tielo \proj_14.flop61/_1__156  (.L_LO(net200));
 sg13g2_tielo \proj_14.flop62/_1__157  (.L_LO(net201));
 sg13g2_tielo \proj_14.flop63/_1__158  (.L_LO(net202));
 sg13g2_tielo \proj_14.flop64/_1__159  (.L_LO(net203));
 sg13g2_tielo \proj_14.flop65/_1__160  (.L_LO(net204));
 sg13g2_tielo \proj_14.flop66/_1__161  (.L_LO(net205));
 sg13g2_tielo \proj_14.flop67/_1__162  (.L_LO(net206));
 sg13g2_tielo \proj_14.flop68/_1__163  (.L_LO(net207));
 sg13g2_tielo \proj_14.flop69/_1__164  (.L_LO(net208));
 sg13g2_tielo \proj_14.flop7/_1__165  (.L_LO(net209));
 sg13g2_tielo \proj_14.flop70/_1__166  (.L_LO(net210));
 sg13g2_tielo \proj_14.flop71/_1__167  (.L_LO(net211));
 sg13g2_tielo \proj_14.flop72/_1__168  (.L_LO(net212));
 sg13g2_tielo \proj_14.flop73/_1__169  (.L_LO(net213));
 sg13g2_tielo \proj_14.flop74/_1__170  (.L_LO(net214));
 sg13g2_tielo \proj_14.flop75/_1__171  (.L_LO(net215));
 sg13g2_tielo \proj_14.flop76/_1__172  (.L_LO(net216));
 sg13g2_tielo \proj_14.flop77/_1__173  (.L_LO(net217));
 sg13g2_tielo \proj_14.flop78/_1__174  (.L_LO(net218));
 sg13g2_tielo \proj_14.flop79/_1__175  (.L_LO(net219));
 sg13g2_tielo \proj_14.flop8/_1__176  (.L_LO(net220));
 sg13g2_tielo \proj_14.flop80/_1__177  (.L_LO(net221));
 sg13g2_tielo \proj_14.flop81/_1__178  (.L_LO(net222));
 sg13g2_tielo \proj_14.flop82/_1__179  (.L_LO(net223));
 sg13g2_tielo \proj_14.flop83/_1__180  (.L_LO(net224));
 sg13g2_tielo \proj_14.flop84/_1__181  (.L_LO(net225));
 sg13g2_tielo \proj_14.flop85/_1__182  (.L_LO(net226));
 sg13g2_tielo \proj_14.flop86/_1__183  (.L_LO(net227));
 sg13g2_tielo \proj_14.flop87/_1__184  (.L_LO(net228));
 sg13g2_tielo \proj_14.flop88/_1__185  (.L_LO(net229));
 sg13g2_tielo \proj_14.flop89/_1__186  (.L_LO(net230));
 sg13g2_tielo \proj_14.flop9/_1__187  (.L_LO(net231));
 sg13g2_tielo \proj_14.flop90/_1__188  (.L_LO(net232));
 sg13g2_tielo \proj_14.flop91/_1__189  (.L_LO(net233));
 sg13g2_tielo \proj_14.flop92/_1__190  (.L_LO(net234));
 sg13g2_tielo \proj_14.flop93/_1__191  (.L_LO(net235));
 sg13g2_tielo \proj_14.flop94/_1__192  (.L_LO(net236));
 sg13g2_tielo \proj_14.flop95/_1__193  (.L_LO(net237));
 sg13g2_tielo \proj_14.flop96/_1__194  (.L_LO(net238));
 sg13g2_tielo \proj_14.flop97/_1__195  (.L_LO(net239));
 sg13g2_tielo \proj_14.flop98/_1__196  (.L_LO(net240));
 sg13g2_tielo \proj_14.flop99/_1__197  (.L_LO(net241));
 sg13g2_tielo \proj_14.mux10/_0__198  (.L_LO(net242));
 sg13g2_tielo \proj_14.mux111/_0__199  (.L_LO(net243));
 sg13g2_tielo \proj_14.mux113/_0__200  (.L_LO(net244));
 sg13g2_tielo \proj_14.mux114/_0__201  (.L_LO(net245));
 sg13g2_tielo \proj_14.mux115/_0__202  (.L_LO(net246));
 sg13g2_tielo \proj_14.mux116/_0__203  (.L_LO(net247));
 sg13g2_tielo \proj_14.mux117/_0__204  (.L_LO(net248));
 sg13g2_tielo \proj_14.mux119/_0__205  (.L_LO(net249));
 sg13g2_tielo \proj_14.mux12/_0__206  (.L_LO(net250));
 sg13g2_tielo \proj_14.mux132/_0__207  (.L_LO(net251));
 sg13g2_tielo \proj_14.mux134/_0__208  (.L_LO(net252));
 sg13g2_tielo \proj_14.mux135/_0__209  (.L_LO(net253));
 sg13g2_tielo \proj_14.mux137/_0__210  (.L_LO(net254));
 sg13g2_tielo \proj_14.mux138/_0__211  (.L_LO(net255));
 sg13g2_tielo \proj_14.mux14/_0__212  (.L_LO(net256));
 sg13g2_tielo \proj_14.mux140/_0__213  (.L_LO(net257));
 sg13g2_tielo \proj_14.mux153/_0__214  (.L_LO(net258));
 sg13g2_tielo \proj_14.mux154/_0__215  (.L_LO(net259));
 sg13g2_tielo \proj_14.mux156/_0__216  (.L_LO(net260));
 sg13g2_tielo \proj_14.mux158/_0__217  (.L_LO(net261));
 sg13g2_tielo \proj_14.mux159/_0__218  (.L_LO(net262));
 sg13g2_tielo \proj_14.mux160/_0__219  (.L_LO(net263));
 sg13g2_tielo \proj_14.mux161/_0__220  (.L_LO(net264));
 sg13g2_tielo \proj_14.mux23/_0__221  (.L_LO(net265));
 sg13g2_tielo \proj_14.mux24/_0__222  (.L_LO(net266));
 sg13g2_tielo \proj_14.mux25/_0__223  (.L_LO(net267));
 sg13g2_tielo \proj_14.mux26/_0__224  (.L_LO(net268));
 sg13g2_tielo \proj_14.mux28/_0__225  (.L_LO(net269));
 sg13g2_tielo \proj_14.mux29/_0__226  (.L_LO(net270));
 sg13g2_tielo \proj_14.mux31/_0__227  (.L_LO(net271));
 sg13g2_tielo \proj_14.mux48/_0__228  (.L_LO(net272));
 sg13g2_tielo \proj_14.mux50/_0__229  (.L_LO(net273));
 sg13g2_tielo \proj_14.mux51/_0__230  (.L_LO(net274));
 sg13g2_tielo \proj_14.mux52/_0__231  (.L_LO(net275));
 sg13g2_tielo \proj_14.mux53/_0__232  (.L_LO(net276));
 sg13g2_tielo \proj_14.mux54/_0__233  (.L_LO(net277));
 sg13g2_tielo \proj_14.mux56/_0__234  (.L_LO(net278));
 sg13g2_tielo \proj_14.mux6/_0__235  (.L_LO(net279));
 sg13g2_tielo \proj_14.mux69/_0__236  (.L_LO(net280));
 sg13g2_tielo \proj_14.mux74/_0__237  (.L_LO(net281));
 sg13g2_tielo \proj_14.mux75/_0__238  (.L_LO(net282));
 sg13g2_tielo \proj_14.mux77/_0__239  (.L_LO(net283));
 sg13g2_tielo \proj_14.mux9/_0__240  (.L_LO(net284));
 sg13g2_tielo \proj_14.mux90/_0__241  (.L_LO(net285));
 sg13g2_tielo \proj_14.mux93/_0__242  (.L_LO(net286));
 sg13g2_tielo \proj_14.mux95/_0__243  (.L_LO(net287));
 sg13g2_tielo \proj_14.mux96/_0__244  (.L_LO(net288));
 sg13g2_tielo \proj_14.mux98/_0__245  (.L_LO(net289));
 sg13g2_tielo tt_um_wokwi_group_2_246 (.L_LO(net290));
 sg13g2_tielo tt_um_wokwi_group_2_247 (.L_LO(net291));
 sg13g2_tielo tt_um_wokwi_group_2_248 (.L_LO(net292));
 sg13g2_tielo tt_um_wokwi_group_2_249 (.L_LO(net293));
 sg13g2_tielo tt_um_wokwi_group_2_250 (.L_LO(net294));
 sg13g2_tielo tt_um_wokwi_group_2_251 (.L_LO(net295));
 sg13g2_tielo tt_um_wokwi_group_2_252 (.L_LO(net296));
 sg13g2_tielo tt_um_wokwi_group_2_253 (.L_LO(net297));
 sg13g2_tielo tt_um_wokwi_group_2_254 (.L_LO(net298));
 sg13g2_tielo tt_um_wokwi_group_2_255 (.L_LO(net299));
 sg13g2_tielo tt_um_wokwi_group_2_256 (.L_LO(net300));
 sg13g2_tielo tt_um_wokwi_group_2_257 (.L_LO(net301));
 sg13g2_tielo tt_um_wokwi_group_2_258 (.L_LO(net302));
 sg13g2_tielo tt_um_wokwi_group_2_259 (.L_LO(net303));
 sg13g2_tielo tt_um_wokwi_group_2_260 (.L_LO(net304));
 sg13g2_tielo tt_um_wokwi_group_2_261 (.L_LO(net305));
 sg13g2_tiehi \proj_14.mux1/_0__262  (.L_HI(net306));
 sg13g2_and2_1 \proj_10.and1/_0_  (.A(\proj_10.net37 ),
    .B(\proj_10.net28 ),
    .X(\proj_10.net41 ));
 sg13g2_and2_1 \proj_10.and10/_0_  (.A(\proj_10.net41 ),
    .B(\proj_10.net38 ),
    .X(\proj_10.net44 ));
 sg13g2_and2_1 \proj_10.and11/_0_  (.A(\proj_10.net45 ),
    .B(\proj_10.net43 ),
    .X(\proj_10.net46 ));
 sg13g2_and2_1 \proj_10.and2/_0_  (.A(\proj_10.net24 ),
    .B(\proj_10.net23 ),
    .X(\proj_10.net25 ));
 sg13g2_and2_1 \proj_10.and3/_0_  (.A(\proj_10.net27 ),
    .B(\proj_10.net26 ),
    .X(\proj_10.net28 ));
 sg13g2_and2_1 \proj_10.and4/_0_  (.A(\proj_10.net26 ),
    .B(\proj_10.net29 ),
    .X(\proj_10.net30 ));
 sg13g2_and2_1 \proj_10.and5/_0_  (.A(\proj_10.net31 ),
    .B(\proj_10.net23 ),
    .X(\proj_10.net32 ));
 sg13g2_and2_1 \proj_10.and6/_0_  (.A(\proj_10.net33 ),
    .B(\proj_10.net25 ),
    .X(\proj_10.net26 ));
 sg13g2_and2_1 \proj_10.and7/_0_  (.A(\proj_10.net34 ),
    .B(\proj_10.net25 ),
    .X(\proj_10.net35 ));
 sg13g2_and2_1 \proj_10.and8/_0_  (.A(\proj_10.net28 ),
    .B(\proj_10.net36 ),
    .X(\proj_10.net42 ));
 sg13g2_and2_1 \proj_10.and9/_0_  (.A(\proj_10.net41 ),
    .B(\proj_10.net39 ),
    .X(\proj_10.net43 ));
 sg13g2_dfrbp_1 \proj_10.flop1/_1_  (.CLK(net12),
    .RESET_B(net427),
    .D(net1),
    .Q_N(\proj_10.flop1/notq ),
    .Q(\proj_10.net40 ));
 sg13g2_tiehi \proj_10.flop10/_1__384  (.L_HI(net428));
 sg13g2_dfrbp_1 \proj_10.flop10/_1_  (.CLK(net13),
    .RESET_B(net428),
    .D(net169),
    .Q_N(\proj_10.flop10/notq ),
    .Q(\proj_10.net38 ));
 sg13g2_tiehi \proj_10.flop11/_1__385  (.L_HI(net429));
 sg13g2_dfrbp_1 \proj_10.flop11/_1_  (.CLK(net14),
    .RESET_B(net429),
    .D(net170),
    .Q_N(\proj_10.flop11/notq ),
    .Q(\proj_10.net36 ));
 sg13g2_tiehi \proj_10.flop12/_1__386  (.L_HI(net430));
 sg13g2_dfrbp_1 \proj_10.flop12/_1_  (.CLK(net15),
    .RESET_B(net430),
    .D(\proj_10.net46 ),
    .Q_N(\proj_10.flop12/notq ),
    .Q(\proj_10.net16 ));
 sg13g2_tiehi \proj_10.flop13/_1__387  (.L_HI(net431));
 sg13g2_dfrbp_1 \proj_10.flop13/_1_  (.CLK(net16),
    .RESET_B(net431),
    .D(\proj_10.net44 ),
    .Q_N(\proj_10.flop13/notq ),
    .Q(\proj_10.net15 ));
 sg13g2_tiehi \proj_10.flop14/_1__388  (.L_HI(net432));
 sg13g2_dfrbp_1 \proj_10.flop14/_1_  (.CLK(net17),
    .RESET_B(net432),
    .D(\proj_10.net42 ),
    .Q_N(\proj_10.flop14/notq ),
    .Q(\proj_10.net14 ));
 sg13g2_tiehi \proj_10.flop2/_1__389  (.L_HI(net433));
 sg13g2_dfrbp_1 \proj_10.flop2/_1_  (.CLK(net18),
    .RESET_B(net433),
    .D(net171),
    .Q_N(\proj_10.flop2/notq ),
    .Q(\proj_10.net29 ));
 sg13g2_tiehi \proj_10.flop3/_1__390  (.L_HI(net434));
 sg13g2_dfrbp_1 \proj_10.flop3/_1_  (.CLK(net19),
    .RESET_B(net434),
    .D(net173),
    .Q_N(\proj_10.flop3/notq ),
    .Q(\proj_10.net34 ));
 sg13g2_tiehi \proj_10.flop4/_1__391  (.L_HI(net435));
 sg13g2_dfrbp_1 \proj_10.flop4/_1_  (.CLK(net20),
    .RESET_B(net435),
    .D(net175),
    .Q_N(\proj_10.flop4/notq ),
    .Q(\proj_10.net31 ));
 sg13g2_tiehi \proj_10.flop5/_1__392  (.L_HI(net436));
 sg13g2_dfrbp_1 \proj_10.flop5/_1_  (.CLK(net21),
    .RESET_B(net436),
    .D(\proj_10.net30 ),
    .Q_N(\proj_10.flop5/notq ),
    .Q(\proj_10.net13 ));
 sg13g2_tiehi \proj_10.flop6/_1__393  (.L_HI(net437));
 sg13g2_dfrbp_1 \proj_10.flop6/_1_  (.CLK(net22),
    .RESET_B(net437),
    .D(\proj_10.net35 ),
    .Q_N(\proj_10.flop6/notq ),
    .Q(\proj_10.net12 ));
 sg13g2_tiehi \proj_10.flop7/_1__394  (.L_HI(net438));
 sg13g2_dfrbp_1 \proj_10.flop7/_1_  (.CLK(net23),
    .RESET_B(net438),
    .D(\proj_10.net32 ),
    .Q_N(\proj_10.flop7/notq ),
    .Q(\proj_10.net11 ));
 sg13g2_tiehi \proj_10.flop8/_1__395  (.L_HI(net439));
 sg13g2_dfrbp_1 \proj_10.flop8/_1_  (.CLK(net24),
    .RESET_B(net439),
    .D(\proj_10.net40 ),
    .Q_N(\proj_10.flop8/notq ),
    .Q(\proj_10.net10 ));
 sg13g2_tiehi \proj_10.flop9/_1__396  (.L_HI(net440));
 sg13g2_dfrbp_1 \proj_10.flop9/_1_  (.CLK(net25),
    .RESET_B(net440),
    .D(net151),
    .Q_N(\proj_10.flop9/notq ),
    .Q(\proj_10.net45 ));
 sg13g2_tiehi \proj_14.flop1/_1__397  (.L_HI(net441));
 sg13g2_inv_1 \proj_10.not1/_0_  (.Y(\proj_10.net24 ),
    .A(\proj_10.net31 ));
 sg13g2_inv_1 \proj_10.not2/_0_  (.Y(\proj_10.net27 ),
    .A(\proj_10.net29 ));
 sg13g2_inv_1 \proj_10.not3/_0_  (.Y(\proj_10.net37 ),
    .A(\proj_10.net36 ));
 sg13g2_inv_1 \proj_10.not5/_0_  (.Y(\proj_10.net39 ),
    .A(\proj_10.net38 ));
 sg13g2_inv_1 \proj_10.not6/_0_  (.Y(\proj_10.net23 ),
    .A(\proj_10.net40 ));
 sg13g2_inv_1 \proj_10.not7/_0_  (.Y(\proj_10.net33 ),
    .A(\proj_10.net34 ));
 sg13g2_xor2_1 \proj_10.xor1/_0_  (.B(net26),
    .A(net27),
    .X(\proj_10.net17 ));
 sg13g2_and2_1 \proj_11.and1/_0_  (.A(net5),
    .B(net177),
    .X(\proj_11.net19 ));
 sg13g2_and2_1 \proj_11.and2/_0_  (.A(\proj_11.net20 ),
    .B(\proj_11.net19 ),
    .X(\proj_11.net21 ));
 sg13g2_and2_1 \proj_11.and3/_0_  (.A(net6),
    .B(net174),
    .X(\proj_11.net22 ));
 sg13g2_and2_1 \proj_11.and4/_0_  (.A(net163),
    .B(net173),
    .X(\proj_11.net24 ));
 sg13g2_and2_1 \proj_11.and5/_0_  (.A(\proj_11.net25 ),
    .B(\proj_11.net23 ),
    .X(\proj_11.net26 ));
 sg13g2_and2_1 \proj_11.and6/_0_  (.A(net135),
    .B(net171),
    .X(\proj_11.net28 ));
 sg13g2_and2_1 \proj_11.and7/_0_  (.A(\proj_11.net29 ),
    .B(\proj_11.net27 ),
    .X(\proj_11.net30 ));
 sg13g2_or2_1 \proj_11.or1/_0_  (.X(\proj_11.net23 ),
    .B(\proj_11.net21 ),
    .A(\proj_11.net22 ));
 sg13g2_or2_1 \proj_11.or2/_0_  (.X(\proj_11.net27 ),
    .B(\proj_11.net26 ),
    .A(\proj_11.net24 ));
 sg13g2_or2_1 \proj_11.or3/_0_  (.X(\proj_11.net13 ),
    .B(\proj_11.net30 ),
    .A(\proj_11.net28 ));
 sg13g2_xor2_1 \proj_11.xor1/_0_  (.B(net178),
    .A(net5),
    .X(\proj_11.net9 ));
 sg13g2_xor2_1 \proj_11.xor2/_0_  (.B(net174),
    .A(net169),
    .X(\proj_11.net20 ));
 sg13g2_xor2_1 \proj_11.xor3/_0_  (.B(\proj_11.net20 ),
    .A(\proj_11.net19 ),
    .X(\proj_11.net10 ));
 sg13g2_xor2_1 \proj_11.xor4/_0_  (.B(\proj_11.net25 ),
    .A(\proj_11.net23 ),
    .X(\proj_11.net11 ));
 sg13g2_xor2_1 \proj_11.xor5/_0_  (.B(net173),
    .A(net163),
    .X(\proj_11.net25 ));
 sg13g2_xor2_1 \proj_11.xor6/_0_  (.B(net171),
    .A(net135),
    .X(\proj_11.net29 ));
 sg13g2_xor2_1 \proj_11.xor7/_0_  (.B(\proj_11.net29 ),
    .A(\proj_11.net27 ),
    .X(\proj_11.net12 ));
 sg13g2_and2_1 \proj_12.and1/_0_  (.A(net178),
    .B(net176),
    .X(\proj_12.net21 ));
 sg13g2_and2_1 \proj_12.and2/_0_  (.A(net170),
    .B(net4),
    .X(\proj_12.net12 ));
 sg13g2_mux2_1 \proj_12.mux1/_0_  (.A0(\proj_12.net21 ),
    .A1(\proj_12.net20 ),
    .S(net3),
    .X(\proj_12.net22 ));
 sg13g2_nand2_1 \proj_12.nand1/_0_  (.Y(\proj_12.net20 ),
    .A(net29),
    .B(net28));
 sg13g2_nand2_1 \proj_12.nand2/_0_  (.Y(\proj_12.net13 ),
    .A(net163),
    .B(net6));
 sg13g2_inv_1 \proj_12.not1/_0_  (.Y(\proj_12.net11 ),
    .A(\proj_12.net22 ));
 sg13g2_xor2_1 \proj_12.xor1/_0_  (.B(net135),
    .A(net168),
    .X(\proj_12.net14 ));
 sg13g2_and2_1 \proj_13.and1/_0_  (.A(net172),
    .B(net135),
    .X(\proj_13.net13 ));
 sg13g2_and2_1 \proj_13.and2/_0_  (.A(\proj_13.net14 ),
    .B(\proj_13.net23 ),
    .X(\proj_13.net10 ));
 sg13g2_and2_1 \proj_13.and3/_0_  (.A(\proj_13.net24 ),
    .B(\proj_13.net22 ),
    .X(\proj_13.net11 ));
 sg13g2_and2_1 \proj_13.and4/_0_  (.A(net163),
    .B(net170),
    .X(\proj_13.net14 ));
 sg13g2_nand2_1 \proj_13.nand1/_0_  (.Y(\proj_13.net9 ),
    .A(net175),
    .B(\proj_13.net21 ));
 sg13g2_nand2_1 \proj_13.nand2/_0_  (.Y(\proj_13.net21 ),
    .A(\proj_13.net13 ),
    .B(\proj_13.net20 ));
 sg13g2_inv_1 \proj_13.not1/_0_  (.Y(\proj_13.net20 ),
    .A(net177));
 sg13g2_inv_1 \proj_13.not2/_0_  (.Y(\proj_13.net24 ),
    .A(net172));
 sg13g2_or2_1 \proj_13.or1/_0_  (.X(\proj_13.net22 ),
    .B(\proj_13.net14 ),
    .A(\proj_13.net12 ));
 sg13g2_or2_1 \proj_13.or2/_0_  (.X(\proj_13.net23 ),
    .B(net4),
    .A(net6));
 sg13g2_xor2_1 \proj_13.xor1/_0_  (.B(net174),
    .A(net172),
    .X(\proj_13.net12 ));
 sg13g2_dfrbp_1 \proj_14.flop1/_1_  (.CLK(net30),
    .RESET_B(net441),
    .D(\proj_14.net8 ),
    .Q_N(\proj_14.flop1/notq ),
    .Q(\proj_14.net9 ));
 sg13g2_tiehi \proj_14.flop10/_1__398  (.L_HI(net442));
 sg13g2_dfrbp_1 \proj_14.flop10/_1_  (.CLK(net31),
    .RESET_B(net442),
    .D(\proj_14.net33 ),
    .Q_N(\proj_14.flop10/notq ),
    .Q(\proj_14.net32 ));
 sg13g2_tiehi \proj_14.flop100/_1__399  (.L_HI(net443));
 sg13g2_dfrbp_1 \proj_14.flop100/_1_  (.CLK(net32),
    .RESET_B(net443),
    .D(\proj_14.net313 ),
    .Q_N(\proj_14.flop100/notq ),
    .Q(\proj_14.net312 ));
 sg13g2_tiehi \proj_14.flop101/_1__400  (.L_HI(net444));
 sg13g2_dfrbp_1 \proj_14.flop101/_1_  (.CLK(net33),
    .RESET_B(net444),
    .D(\proj_14.net316 ),
    .Q_N(\proj_14.flop101/notq ),
    .Q(\proj_14.net315 ));
 sg13g2_tiehi \proj_14.flop102/_1__401  (.L_HI(net445));
 sg13g2_dfrbp_1 \proj_14.flop102/_1_  (.CLK(net34),
    .RESET_B(net445),
    .D(\proj_14.net320 ),
    .Q_N(\proj_14.flop102/notq ),
    .Q(\proj_14.net254 ));
 sg13g2_tiehi \proj_14.flop103/_1__402  (.L_HI(net446));
 sg13g2_dfrbp_1 \proj_14.flop103/_1_  (.CLK(net35),
    .RESET_B(net446),
    .D(\proj_14.net323 ),
    .Q_N(\proj_14.flop103/notq ),
    .Q(\proj_14.net322 ));
 sg13g2_tiehi \proj_14.flop104/_1__403  (.L_HI(net447));
 sg13g2_dfrbp_1 \proj_14.flop104/_1_  (.CLK(net36),
    .RESET_B(net447),
    .D(\proj_14.net326 ),
    .Q_N(\proj_14.flop104/notq ),
    .Q(\proj_14.net325 ));
 sg13g2_tiehi \proj_14.flop105/_1__404  (.L_HI(net448));
 sg13g2_dfrbp_1 \proj_14.flop105/_1_  (.CLK(net37),
    .RESET_B(net448),
    .D(\proj_14.net329 ),
    .Q_N(\proj_14.flop105/notq ),
    .Q(\proj_14.net328 ));
 sg13g2_tiehi \proj_14.flop106/_1__405  (.L_HI(net449));
 sg13g2_dfrbp_1 \proj_14.flop106/_1_  (.CLK(net38),
    .RESET_B(net449),
    .D(\proj_14.net332 ),
    .Q_N(\proj_14.flop106/notq ),
    .Q(\proj_14.net333 ));
 sg13g2_tiehi \proj_14.flop107/_1__406  (.L_HI(net450));
 sg13g2_dfrbp_1 \proj_14.flop107/_1_  (.CLK(net39),
    .RESET_B(net450),
    .D(\proj_14.net336 ),
    .Q_N(\proj_14.flop107/notq ),
    .Q(\proj_14.net335 ));
 sg13g2_tiehi \proj_14.flop108/_1__407  (.L_HI(net451));
 sg13g2_dfrbp_1 \proj_14.flop108/_1_  (.CLK(net40),
    .RESET_B(net451),
    .D(\proj_14.net339 ),
    .Q_N(\proj_14.flop108/notq ),
    .Q(\proj_14.net338 ));
 sg13g2_tiehi \proj_14.flop109/_1__408  (.L_HI(net452));
 sg13g2_dfrbp_1 \proj_14.flop109/_1_  (.CLK(net41),
    .RESET_B(net452),
    .D(\proj_14.net342 ),
    .Q_N(\proj_14.flop109/notq ),
    .Q(\proj_14.net341 ));
 sg13g2_tiehi \proj_14.flop11/_1__409  (.L_HI(net453));
 sg13g2_dfrbp_1 \proj_14.flop11/_1_  (.CLK(net42),
    .RESET_B(net453),
    .D(\proj_14.net36 ),
    .Q_N(\proj_14.flop11/notq ),
    .Q(\proj_14.net35 ));
 sg13g2_tiehi \proj_14.flop110/_1__410  (.L_HI(net454));
 sg13g2_dfrbp_1 \proj_14.flop110/_1_  (.CLK(net43),
    .RESET_B(net454),
    .D(\proj_14.net345 ),
    .Q_N(\proj_14.flop110/notq ),
    .Q(\proj_14.net344 ));
 sg13g2_tiehi \proj_14.flop111/_1__411  (.L_HI(net455));
 sg13g2_dfrbp_1 \proj_14.flop111/_1_  (.CLK(net44),
    .RESET_B(net455),
    .D(\proj_14.net348 ),
    .Q_N(\proj_14.flop111/notq ),
    .Q(\proj_14.net347 ));
 sg13g2_tiehi \proj_14.flop112/_1__412  (.L_HI(net456));
 sg13g2_dfrbp_1 \proj_14.flop112/_1_  (.CLK(net45),
    .RESET_B(net456),
    .D(\proj_14.net351 ),
    .Q_N(\proj_14.flop112/notq ),
    .Q(\proj_14.net350 ));
 sg13g2_tiehi \proj_14.flop113/_1__413  (.L_HI(net457));
 sg13g2_dfrbp_1 \proj_14.flop113/_1_  (.CLK(net46),
    .RESET_B(net457),
    .D(\proj_14.net354 ),
    .Q_N(\proj_14.flop113/notq ),
    .Q(\proj_14.net353 ));
 sg13g2_tiehi \proj_14.flop114/_1__414  (.L_HI(net458));
 sg13g2_dfrbp_1 \proj_14.flop114/_1_  (.CLK(net47),
    .RESET_B(net458),
    .D(\proj_14.net357 ),
    .Q_N(\proj_14.flop114/notq ),
    .Q(\proj_14.net356 ));
 sg13g2_tiehi \proj_14.flop115/_1__415  (.L_HI(net459));
 sg13g2_dfrbp_1 \proj_14.flop115/_1_  (.CLK(net48),
    .RESET_B(net459),
    .D(\proj_14.net360 ),
    .Q_N(\proj_14.flop115/notq ),
    .Q(\proj_14.net359 ));
 sg13g2_tiehi \proj_14.flop116/_1__416  (.L_HI(net460));
 sg13g2_dfrbp_1 \proj_14.flop116/_1_  (.CLK(net49),
    .RESET_B(net460),
    .D(\proj_14.net363 ),
    .Q_N(\proj_14.flop116/notq ),
    .Q(\proj_14.net362 ));
 sg13g2_tiehi \proj_14.flop117/_1__417  (.L_HI(net461));
 sg13g2_dfrbp_1 \proj_14.flop117/_1_  (.CLK(net50),
    .RESET_B(net461),
    .D(\proj_14.net366 ),
    .Q_N(\proj_14.flop117/notq ),
    .Q(\proj_14.net365 ));
 sg13g2_tiehi \proj_14.flop118/_1__418  (.L_HI(net462));
 sg13g2_dfrbp_1 \proj_14.flop118/_1_  (.CLK(net51),
    .RESET_B(net462),
    .D(\proj_14.net369 ),
    .Q_N(\proj_14.flop118/notq ),
    .Q(\proj_14.net368 ));
 sg13g2_tiehi \proj_14.flop119/_1__419  (.L_HI(net463));
 sg13g2_dfrbp_1 \proj_14.flop119/_1_  (.CLK(net52),
    .RESET_B(net463),
    .D(\proj_14.net372 ),
    .Q_N(\proj_14.flop119/notq ),
    .Q(\proj_14.net371 ));
 sg13g2_tiehi \proj_14.flop12/_1__420  (.L_HI(net464));
 sg13g2_dfrbp_1 \proj_14.flop12/_1_  (.CLK(net53),
    .RESET_B(net464),
    .D(\proj_14.net39 ),
    .Q_N(\proj_14.flop12/notq ),
    .Q(\proj_14.net38 ));
 sg13g2_tiehi \proj_14.flop120/_1__421  (.L_HI(net465));
 sg13g2_dfrbp_1 \proj_14.flop120/_1_  (.CLK(net54),
    .RESET_B(net465),
    .D(\proj_14.net375 ),
    .Q_N(\proj_14.flop120/notq ),
    .Q(\proj_14.net374 ));
 sg13g2_tiehi \proj_14.flop121/_1__422  (.L_HI(net466));
 sg13g2_dfrbp_1 \proj_14.flop121/_1_  (.CLK(net55),
    .RESET_B(net466),
    .D(\proj_14.net378 ),
    .Q_N(\proj_14.flop121/notq ),
    .Q(\proj_14.net377 ));
 sg13g2_tiehi \proj_14.flop122/_1__423  (.L_HI(net467));
 sg13g2_dfrbp_1 \proj_14.flop122/_1_  (.CLK(net56),
    .RESET_B(net467),
    .D(\proj_14.net381 ),
    .Q_N(\proj_14.flop122/notq ),
    .Q(\proj_14.net380 ));
 sg13g2_tiehi \proj_14.flop123/_1__424  (.L_HI(net468));
 sg13g2_dfrbp_1 \proj_14.flop123/_1_  (.CLK(net57),
    .RESET_B(net468),
    .D(\proj_14.net385 ),
    .Q_N(\proj_14.flop123/notq ),
    .Q(\proj_14.net318 ));
 sg13g2_tiehi \proj_14.flop124/_1__425  (.L_HI(net469));
 sg13g2_dfrbp_1 \proj_14.flop124/_1_  (.CLK(net58),
    .RESET_B(net469),
    .D(\proj_14.net388 ),
    .Q_N(\proj_14.flop124/notq ),
    .Q(\proj_14.net387 ));
 sg13g2_tiehi \proj_14.flop125/_1__426  (.L_HI(net470));
 sg13g2_dfrbp_1 \proj_14.flop125/_1_  (.CLK(net59),
    .RESET_B(net470),
    .D(\proj_14.net391 ),
    .Q_N(\proj_14.flop125/notq ),
    .Q(\proj_14.net390 ));
 sg13g2_tiehi \proj_14.flop126/_1__427  (.L_HI(net471));
 sg13g2_dfrbp_1 \proj_14.flop126/_1_  (.CLK(net60),
    .RESET_B(net471),
    .D(\proj_14.net394 ),
    .Q_N(\proj_14.flop126/notq ),
    .Q(\proj_14.net393 ));
 sg13g2_tiehi \proj_14.flop127/_1__428  (.L_HI(net472));
 sg13g2_dfrbp_1 \proj_14.flop127/_1_  (.CLK(net61),
    .RESET_B(net472),
    .D(\proj_14.net396 ),
    .Q_N(\proj_14.flop127/notq ),
    .Q(\proj_14.net397 ));
 sg13g2_tiehi \proj_14.flop128/_1__429  (.L_HI(net473));
 sg13g2_dfrbp_1 \proj_14.flop128/_1_  (.CLK(net62),
    .RESET_B(net473),
    .D(\proj_14.net400 ),
    .Q_N(\proj_14.flop128/notq ),
    .Q(\proj_14.net399 ));
 sg13g2_tiehi \proj_14.flop129/_1__430  (.L_HI(net474));
 sg13g2_dfrbp_1 \proj_14.flop129/_1_  (.CLK(net63),
    .RESET_B(net474),
    .D(\proj_14.net403 ),
    .Q_N(\proj_14.flop129/notq ),
    .Q(\proj_14.net402 ));
 sg13g2_tiehi \proj_14.flop13/_1__431  (.L_HI(net475));
 sg13g2_dfrbp_1 \proj_14.flop13/_1_  (.CLK(net64),
    .RESET_B(net475),
    .D(\proj_14.net42 ),
    .Q_N(\proj_14.flop13/notq ),
    .Q(\proj_14.net41 ));
 sg13g2_tiehi \proj_14.flop130/_1__432  (.L_HI(net476));
 sg13g2_dfrbp_1 \proj_14.flop130/_1_  (.CLK(net65),
    .RESET_B(net476),
    .D(\proj_14.net406 ),
    .Q_N(\proj_14.flop130/notq ),
    .Q(\proj_14.net405 ));
 sg13g2_tiehi \proj_14.flop131/_1__433  (.L_HI(net477));
 sg13g2_dfrbp_1 \proj_14.flop131/_1_  (.CLK(net66),
    .RESET_B(net477),
    .D(\proj_14.net409 ),
    .Q_N(\proj_14.flop131/notq ),
    .Q(\proj_14.net408 ));
 sg13g2_tiehi \proj_14.flop132/_1__434  (.L_HI(net478));
 sg13g2_dfrbp_1 \proj_14.flop132/_1_  (.CLK(net67),
    .RESET_B(net478),
    .D(\proj_14.net412 ),
    .Q_N(\proj_14.flop132/notq ),
    .Q(\proj_14.net411 ));
 sg13g2_tiehi \proj_14.flop133/_1__435  (.L_HI(net479));
 sg13g2_dfrbp_1 \proj_14.flop133/_1_  (.CLK(net68),
    .RESET_B(net479),
    .D(\proj_14.net415 ),
    .Q_N(\proj_14.flop133/notq ),
    .Q(\proj_14.net414 ));
 sg13g2_tiehi \proj_14.flop134/_1__436  (.L_HI(net480));
 sg13g2_dfrbp_1 \proj_14.flop134/_1_  (.CLK(net69),
    .RESET_B(net480),
    .D(\proj_14.net418 ),
    .Q_N(\proj_14.flop134/notq ),
    .Q(\proj_14.net417 ));
 sg13g2_tiehi \proj_14.flop135/_1__437  (.L_HI(net481));
 sg13g2_dfrbp_1 \proj_14.flop135/_1_  (.CLK(net70),
    .RESET_B(net481),
    .D(\proj_14.net421 ),
    .Q_N(\proj_14.flop135/notq ),
    .Q(\proj_14.net420 ));
 sg13g2_tiehi \proj_14.flop136/_1__438  (.L_HI(net482));
 sg13g2_dfrbp_1 \proj_14.flop136/_1_  (.CLK(net71),
    .RESET_B(net482),
    .D(\proj_14.net424 ),
    .Q_N(\proj_14.flop136/notq ),
    .Q(\proj_14.net423 ));
 sg13g2_tiehi \proj_14.flop137/_1__439  (.L_HI(net483));
 sg13g2_dfrbp_1 \proj_14.flop137/_1_  (.CLK(net72),
    .RESET_B(net483),
    .D(\proj_14.net427 ),
    .Q_N(\proj_14.flop137/notq ),
    .Q(\proj_14.net426 ));
 sg13g2_tiehi \proj_14.flop138/_1__440  (.L_HI(net484));
 sg13g2_dfrbp_1 \proj_14.flop138/_1_  (.CLK(net73),
    .RESET_B(net484),
    .D(\proj_14.net430 ),
    .Q_N(\proj_14.flop138/notq ),
    .Q(\proj_14.net429 ));
 sg13g2_tiehi \proj_14.flop139/_1__441  (.L_HI(net485));
 sg13g2_dfrbp_1 \proj_14.flop139/_1_  (.CLK(net74),
    .RESET_B(net485),
    .D(\proj_14.net433 ),
    .Q_N(\proj_14.flop139/notq ),
    .Q(\proj_14.net432 ));
 sg13g2_tiehi \proj_14.flop14/_1__442  (.L_HI(net486));
 sg13g2_dfrbp_1 \proj_14.flop14/_1_  (.CLK(net75),
    .RESET_B(net486),
    .D(\proj_14.net45 ),
    .Q_N(\proj_14.flop14/notq ),
    .Q(\proj_14.net44 ));
 sg13g2_tiehi \proj_14.flop140/_1__443  (.L_HI(net487));
 sg13g2_dfrbp_1 \proj_14.flop140/_1_  (.CLK(net76),
    .RESET_B(net487),
    .D(\proj_14.net436 ),
    .Q_N(\proj_14.flop140/notq ),
    .Q(\proj_14.net435 ));
 sg13g2_tiehi \proj_14.flop141/_1__444  (.L_HI(net488));
 sg13g2_dfrbp_1 \proj_14.flop141/_1_  (.CLK(net77),
    .RESET_B(net488),
    .D(\proj_14.net439 ),
    .Q_N(\proj_14.flop141/notq ),
    .Q(\proj_14.net438 ));
 sg13g2_tiehi \proj_14.flop142/_1__445  (.L_HI(net489));
 sg13g2_dfrbp_1 \proj_14.flop142/_1_  (.CLK(net78),
    .RESET_B(net489),
    .D(\proj_14.net442 ),
    .Q_N(\proj_14.flop142/notq ),
    .Q(\proj_14.net441 ));
 sg13g2_tiehi \proj_14.flop143/_1__446  (.L_HI(net490));
 sg13g2_dfrbp_1 \proj_14.flop143/_1_  (.CLK(net79),
    .RESET_B(net490),
    .D(\proj_14.net445 ),
    .Q_N(\proj_14.flop143/notq ),
    .Q(\proj_14.net444 ));
 sg13g2_tiehi \proj_14.flop144/_1__447  (.L_HI(net491));
 sg13g2_dfrbp_1 \proj_14.flop144/_1_  (.CLK(net80),
    .RESET_B(net491),
    .D(\proj_14.net449 ),
    .Q_N(\proj_14.flop144/notq ),
    .Q(\proj_14.net383 ));
 sg13g2_tiehi \proj_14.flop145/_1__448  (.L_HI(net492));
 sg13g2_dfrbp_1 \proj_14.flop145/_1_  (.CLK(net81),
    .RESET_B(net492),
    .D(\proj_14.net452 ),
    .Q_N(\proj_14.flop145/notq ),
    .Q(\proj_14.net451 ));
 sg13g2_tiehi \proj_14.flop146/_1__449  (.L_HI(net493));
 sg13g2_dfrbp_1 \proj_14.flop146/_1_  (.CLK(net82),
    .RESET_B(net493),
    .D(\proj_14.net455 ),
    .Q_N(\proj_14.flop146/notq ),
    .Q(\proj_14.net454 ));
 sg13g2_tiehi \proj_14.flop147/_1__450  (.L_HI(net494));
 sg13g2_dfrbp_1 \proj_14.flop147/_1_  (.CLK(net83),
    .RESET_B(net494),
    .D(\proj_14.net458 ),
    .Q_N(\proj_14.flop147/notq ),
    .Q(\proj_14.net457 ));
 sg13g2_tiehi \proj_14.flop148/_1__451  (.L_HI(net495));
 sg13g2_dfrbp_1 \proj_14.flop148/_1_  (.CLK(net84),
    .RESET_B(net495),
    .D(\proj_14.net460 ),
    .Q_N(\proj_14.flop148/notq ),
    .Q(\proj_14.net461 ));
 sg13g2_tiehi \proj_14.flop149/_1__452  (.L_HI(net496));
 sg13g2_dfrbp_1 \proj_14.flop149/_1_  (.CLK(net85),
    .RESET_B(net496),
    .D(\proj_14.net464 ),
    .Q_N(\proj_14.flop149/notq ),
    .Q(\proj_14.net463 ));
 sg13g2_tiehi \proj_14.flop15/_1__453  (.L_HI(net497));
 sg13g2_dfrbp_1 \proj_14.flop15/_1_  (.CLK(net86),
    .RESET_B(net497),
    .D(\proj_14.net48 ),
    .Q_N(\proj_14.flop15/notq ),
    .Q(\proj_14.net47 ));
 sg13g2_tiehi \proj_14.flop150/_1__454  (.L_HI(net498));
 sg13g2_dfrbp_1 \proj_14.flop150/_1_  (.CLK(net87),
    .RESET_B(net498),
    .D(\proj_14.net467 ),
    .Q_N(\proj_14.flop150/notq ),
    .Q(\proj_14.net466 ));
 sg13g2_tiehi \proj_14.flop151/_1__455  (.L_HI(net499));
 sg13g2_dfrbp_1 \proj_14.flop151/_1_  (.CLK(net88),
    .RESET_B(net499),
    .D(\proj_14.net470 ),
    .Q_N(\proj_14.flop151/notq ),
    .Q(\proj_14.net469 ));
 sg13g2_tiehi \proj_14.flop152/_1__456  (.L_HI(net500));
 sg13g2_dfrbp_1 \proj_14.flop152/_1_  (.CLK(net89),
    .RESET_B(net500),
    .D(\proj_14.net473 ),
    .Q_N(\proj_14.flop152/notq ),
    .Q(\proj_14.net472 ));
 sg13g2_tiehi \proj_14.flop153/_1__457  (.L_HI(net501));
 sg13g2_dfrbp_1 \proj_14.flop153/_1_  (.CLK(net90),
    .RESET_B(net501),
    .D(\proj_14.net476 ),
    .Q_N(\proj_14.flop153/notq ),
    .Q(\proj_14.net475 ));
 sg13g2_tiehi \proj_14.flop154/_1__458  (.L_HI(net502));
 sg13g2_dfrbp_1 \proj_14.flop154/_1_  (.CLK(net91),
    .RESET_B(net502),
    .D(\proj_14.net479 ),
    .Q_N(\proj_14.flop154/notq ),
    .Q(\proj_14.net478 ));
 sg13g2_tiehi \proj_14.flop155/_1__459  (.L_HI(net503));
 sg13g2_dfrbp_1 \proj_14.flop155/_1_  (.CLK(net92),
    .RESET_B(net503),
    .D(\proj_14.net482 ),
    .Q_N(\proj_14.flop155/notq ),
    .Q(\proj_14.net481 ));
 sg13g2_tiehi \proj_14.flop156/_1__460  (.L_HI(net504));
 sg13g2_dfrbp_1 \proj_14.flop156/_1_  (.CLK(net93),
    .RESET_B(net504),
    .D(\proj_14.net485 ),
    .Q_N(\proj_14.flop156/notq ),
    .Q(\proj_14.net484 ));
 sg13g2_tiehi \proj_14.flop157/_1__461  (.L_HI(net505));
 sg13g2_dfrbp_1 \proj_14.flop157/_1_  (.CLK(net94),
    .RESET_B(net505),
    .D(\proj_14.net488 ),
    .Q_N(\proj_14.flop157/notq ),
    .Q(\proj_14.net487 ));
 sg13g2_tiehi \proj_14.flop158/_1__462  (.L_HI(net506));
 sg13g2_dfrbp_1 \proj_14.flop158/_1_  (.CLK(net95),
    .RESET_B(net506),
    .D(\proj_14.net491 ),
    .Q_N(\proj_14.flop158/notq ),
    .Q(\proj_14.net490 ));
 sg13g2_tiehi \proj_14.flop159/_1__463  (.L_HI(net507));
 sg13g2_dfrbp_1 \proj_14.flop159/_1_  (.CLK(net96),
    .RESET_B(net507),
    .D(\proj_14.net494 ),
    .Q_N(\proj_14.flop159/notq ),
    .Q(\proj_14.net493 ));
 sg13g2_tiehi \proj_14.flop16/_1__464  (.L_HI(net508));
 sg13g2_dfrbp_1 \proj_14.flop16/_1_  (.CLK(net97),
    .RESET_B(net508),
    .D(\proj_14.net51 ),
    .Q_N(\proj_14.flop16/notq ),
    .Q(\proj_14.net50 ));
 sg13g2_tiehi \proj_14.flop160/_1__465  (.L_HI(net509));
 sg13g2_dfrbp_1 \proj_14.flop160/_1_  (.CLK(net98),
    .RESET_B(net509),
    .D(\proj_14.net497 ),
    .Q_N(\proj_14.flop160/notq ),
    .Q(\proj_14.net496 ));
 sg13g2_tiehi \proj_14.flop161/_1__466  (.L_HI(net510));
 sg13g2_dfrbp_1 \proj_14.flop161/_1_  (.CLK(net99),
    .RESET_B(net510),
    .D(\proj_14.net500 ),
    .Q_N(\proj_14.flop161/notq ),
    .Q(\proj_14.net499 ));
 sg13g2_tiehi \proj_14.flop162/_1__467  (.L_HI(net511));
 sg13g2_dfrbp_1 \proj_14.flop162/_1_  (.CLK(net100),
    .RESET_B(net511),
    .D(\proj_14.net503 ),
    .Q_N(\proj_14.flop162/notq ),
    .Q(\proj_14.net502 ));
 sg13g2_tiehi \proj_14.flop163/_1__468  (.L_HI(net512));
 sg13g2_dfrbp_1 \proj_14.flop163/_1_  (.CLK(net101),
    .RESET_B(net512),
    .D(\proj_14.net506 ),
    .Q_N(\proj_14.flop163/notq ),
    .Q(\proj_14.net505 ));
 sg13g2_tiehi \proj_14.flop164/_1__469  (.L_HI(net513));
 sg13g2_dfrbp_1 \proj_14.flop164/_1_  (.CLK(net102),
    .RESET_B(net513),
    .D(\proj_14.net509 ),
    .Q_N(\proj_14.flop164/notq ),
    .Q(\proj_14.net508 ));
 sg13g2_tiehi \proj_14.flop165/_1__470  (.L_HI(net514));
 sg13g2_dfrbp_1 \proj_14.flop165/_1_  (.CLK(net103),
    .RESET_B(net514),
    .D(\proj_14.net512 ),
    .Q_N(\proj_14.flop165/notq ),
    .Q(\proj_14.net447 ));
 sg13g2_tiehi \proj_14.flop166/_1__471  (.L_HI(net515));
 sg13g2_dfrbp_1 \proj_14.flop166/_1_  (.CLK(net104),
    .RESET_B(net515),
    .D(\proj_14.net515 ),
    .Q_N(\proj_14.flop166/notq ),
    .Q(\proj_14.net514 ));
 sg13g2_tiehi \proj_14.flop167/_1__472  (.L_HI(net516));
 sg13g2_dfrbp_1 \proj_14.flop167/_1_  (.CLK(net105),
    .RESET_B(net516),
    .D(\proj_14.net518 ),
    .Q_N(\proj_14.flop167/notq ),
    .Q(\proj_14.net517 ));
 sg13g2_tiehi \proj_14.flop168/_1__473  (.L_HI(net517));
 sg13g2_dfrbp_1 \proj_14.flop168/_1_  (.CLK(net106),
    .RESET_B(net517),
    .D(\proj_14.net521 ),
    .Q_N(\proj_14.flop168/notq ),
    .Q(\proj_14.net520 ));
 sg13g2_tiehi \proj_14.flop17/_1__474  (.L_HI(net518));
 sg13g2_dfrbp_1 \proj_14.flop17/_1_  (.CLK(net107),
    .RESET_B(net518),
    .D(\proj_14.net54 ),
    .Q_N(\proj_14.flop17/notq ),
    .Q(\proj_14.net53 ));
 sg13g2_tiehi \proj_14.flop18/_1__475  (.L_HI(net519));
 sg13g2_dfrbp_1 \proj_14.flop18/_1_  (.CLK(net108),
    .RESET_B(net519),
    .D(\proj_14.net57 ),
    .Q_N(\proj_14.flop18/notq ),
    .Q(\proj_14.net56 ));
 sg13g2_tiehi \proj_14.flop19/_1__476  (.L_HI(net520));
 sg13g2_dfrbp_1 \proj_14.flop19/_1_  (.CLK(net109),
    .RESET_B(net520),
    .D(\proj_14.net67 ),
    .Q_N(\proj_14.flop19/notq ),
    .Q(\proj_14.net66 ));
 sg13g2_tiehi \proj_14.flop2/_1__477  (.L_HI(net521));
 sg13g2_dfrbp_1 \proj_14.flop2/_1_  (.CLK(net110),
    .RESET_B(net521),
    .D(\proj_14.net63 ),
    .Q_N(\proj_14.flop2/notq ),
    .Q(\proj_14.net64 ));
 sg13g2_tiehi \proj_14.flop20/_1__478  (.L_HI(net522));
 sg13g2_dfrbp_1 \proj_14.flop20/_1_  (.CLK(net111),
    .RESET_B(net522),
    .D(\proj_14.net70 ),
    .Q_N(\proj_14.flop20/notq ),
    .Q(\proj_14.net69 ));
 sg13g2_tiehi \proj_14.flop21/_1__479  (.L_HI(net523));
 sg13g2_dfrbp_1 \proj_14.flop21/_1_  (.CLK(net112),
    .RESET_B(net523),
    .D(\proj_14.net73 ),
    .Q_N(\proj_14.flop21/notq ),
    .Q(\proj_14.net72 ));
 sg13g2_tiehi \proj_14.flop22/_1__480  (.L_HI(net524));
 sg13g2_dfrbp_1 \proj_14.flop22/_1_  (.CLK(net113),
    .RESET_B(net524),
    .D(\proj_14.net76 ),
    .Q_N(\proj_14.flop22/notq ),
    .Q(\proj_14.net75 ));
 sg13g2_tiehi \proj_14.flop23/_1__481  (.L_HI(net525));
 sg13g2_dfrbp_1 \proj_14.flop23/_1_  (.CLK(net114),
    .RESET_B(net525),
    .D(\proj_14.net79 ),
    .Q_N(\proj_14.flop23/notq ),
    .Q(\proj_14.net78 ));
 sg13g2_tiehi \proj_14.flop24/_1__482  (.L_HI(net526));
 sg13g2_dfrbp_1 \proj_14.flop24/_1_  (.CLK(net115),
    .RESET_B(net526),
    .D(\proj_14.net82 ),
    .Q_N(\proj_14.flop24/notq ),
    .Q(\proj_14.net81 ));
 sg13g2_tiehi \proj_14.flop25/_1__483  (.L_HI(net527));
 sg13g2_dfrbp_1 \proj_14.flop25/_1_  (.CLK(net116),
    .RESET_B(net527),
    .D(\proj_14.net85 ),
    .Q_N(\proj_14.flop25/notq ),
    .Q(\proj_14.net84 ));
 sg13g2_tiehi \proj_14.flop26/_1__484  (.L_HI(net528));
 sg13g2_dfrbp_1 \proj_14.flop26/_1_  (.CLK(net117),
    .RESET_B(net528),
    .D(\proj_14.net88 ),
    .Q_N(\proj_14.flop26/notq ),
    .Q(\proj_14.net87 ));
 sg13g2_tiehi \proj_14.flop27/_1__485  (.L_HI(net529));
 sg13g2_dfrbp_1 \proj_14.flop27/_1_  (.CLK(net118),
    .RESET_B(net529),
    .D(\proj_14.net91 ),
    .Q_N(\proj_14.flop27/notq ),
    .Q(\proj_14.net90 ));
 sg13g2_tiehi \proj_14.flop28/_1__486  (.L_HI(net530));
 sg13g2_dfrbp_1 \proj_14.flop28/_1_  (.CLK(net119),
    .RESET_B(net530),
    .D(\proj_14.net94 ),
    .Q_N(\proj_14.flop28/notq ),
    .Q(\proj_14.net93 ));
 sg13g2_tiehi \proj_14.flop29/_1__487  (.L_HI(net531));
 sg13g2_dfrbp_1 \proj_14.flop29/_1_  (.CLK(net120),
    .RESET_B(net531),
    .D(\proj_14.net97 ),
    .Q_N(\proj_14.flop29/notq ),
    .Q(\proj_14.net96 ));
 sg13g2_tiehi \proj_14.flop3/_1__488  (.L_HI(net532));
 sg13g2_dfrbp_1 \proj_14.flop3/_1_  (.CLK(net121),
    .RESET_B(net532),
    .D(\proj_14.net12 ),
    .Q_N(\proj_14.flop3/notq ),
    .Q(\proj_14.net11 ));
 sg13g2_tiehi \proj_14.flop30/_1__489  (.L_HI(net533));
 sg13g2_dfrbp_1 \proj_14.flop30/_1_  (.CLK(net122),
    .RESET_B(net533),
    .D(\proj_14.net100 ),
    .Q_N(\proj_14.flop30/notq ),
    .Q(\proj_14.net99 ));
 sg13g2_tiehi \proj_14.flop31/_1__490  (.L_HI(net534));
 sg13g2_dfrbp_1 \proj_14.flop31/_1_  (.CLK(net123),
    .RESET_B(net534),
    .D(\proj_14.net103 ),
    .Q_N(\proj_14.flop31/notq ),
    .Q(\proj_14.net102 ));
 sg13g2_tiehi \proj_14.flop32/_1__491  (.L_HI(net535));
 sg13g2_dfrbp_1 \proj_14.flop32/_1_  (.CLK(net124),
    .RESET_B(net535),
    .D(\proj_14.net106 ),
    .Q_N(\proj_14.flop32/notq ),
    .Q(\proj_14.net105 ));
 sg13g2_tiehi \proj_14.flop33/_1__492  (.L_HI(net536));
 sg13g2_dfrbp_1 \proj_14.flop33/_1_  (.CLK(net125),
    .RESET_B(net536),
    .D(\proj_14.net109 ),
    .Q_N(\proj_14.flop33/notq ),
    .Q(\proj_14.net108 ));
 sg13g2_tiehi \proj_14.flop34/_1__493  (.L_HI(net537));
 sg13g2_dfrbp_1 \proj_14.flop34/_1_  (.CLK(net126),
    .RESET_B(net537),
    .D(\proj_14.net112 ),
    .Q_N(\proj_14.flop34/notq ),
    .Q(\proj_14.net111 ));
 sg13g2_tiehi \proj_14.flop35/_1__494  (.L_HI(net538));
 sg13g2_dfrbp_1 \proj_14.flop35/_1_  (.CLK(net127),
    .RESET_B(net538),
    .D(\proj_14.net116 ),
    .Q_N(\proj_14.flop35/notq ),
    .Q(\proj_14.net59 ));
 sg13g2_tiehi \proj_14.flop36/_1__495  (.L_HI(net539));
 sg13g2_dfrbp_1 \proj_14.flop36/_1_  (.CLK(net128),
    .RESET_B(net539),
    .D(\proj_14.net119 ),
    .Q_N(\proj_14.flop36/notq ),
    .Q(\proj_14.net118 ));
 sg13g2_tiehi \proj_14.flop37/_1__496  (.L_HI(net540));
 sg13g2_dfrbp_1 \proj_14.flop37/_1_  (.CLK(net129),
    .RESET_B(net540),
    .D(\proj_14.net122 ),
    .Q_N(\proj_14.flop37/notq ),
    .Q(\proj_14.net121 ));
 sg13g2_tiehi \proj_14.flop38/_1__497  (.L_HI(net541));
 sg13g2_dfrbp_1 \proj_14.flop38/_1_  (.CLK(net130),
    .RESET_B(net541),
    .D(\proj_14.net125 ),
    .Q_N(\proj_14.flop38/notq ),
    .Q(\proj_14.net124 ));
 sg13g2_tiehi \proj_14.flop39/_1__498  (.L_HI(net542));
 sg13g2_dfrbp_1 \proj_14.flop39/_1_  (.CLK(net131),
    .RESET_B(net542),
    .D(\proj_14.net127 ),
    .Q_N(\proj_14.flop39/notq ),
    .Q(\proj_14.net128 ));
 sg13g2_tiehi \proj_14.flop4/_1__499  (.L_HI(net543));
 sg13g2_dfrbp_1 \proj_14.flop4/_1_  (.CLK(net132),
    .RESET_B(net543),
    .D(\proj_14.net15 ),
    .Q_N(\proj_14.flop4/notq ),
    .Q(\proj_14.net14 ));
 sg13g2_tiehi \proj_14.flop40/_1__500  (.L_HI(net544));
 sg13g2_dfrbp_1 \proj_14.flop40/_1_  (.CLK(net133),
    .RESET_B(net544),
    .D(\proj_14.net131 ),
    .Q_N(\proj_14.flop40/notq ),
    .Q(\proj_14.net130 ));
 sg13g2_tiehi \proj_14.flop41/_1__501  (.L_HI(net545));
 sg13g2_dfrbp_1 \proj_14.flop41/_1_  (.CLK(net134),
    .RESET_B(net545),
    .D(\proj_14.net134 ),
    .Q_N(\proj_14.flop41/notq ),
    .Q(\proj_14.net133 ));
 sg13g2_tiehi \proj_14.flop42/_1__502  (.L_HI(net546));
 sg13g2_dfrbp_1 \proj_14.flop42/_1_  (.CLK(net179),
    .RESET_B(net546),
    .D(\proj_14.net137 ),
    .Q_N(\proj_14.flop42/notq ),
    .Q(\proj_14.net136 ));
 sg13g2_tiehi \proj_14.flop43/_1__503  (.L_HI(net547));
 sg13g2_dfrbp_1 \proj_14.flop43/_1_  (.CLK(net180),
    .RESET_B(net547),
    .D(\proj_14.net139 ),
    .Q_N(\proj_14.flop43/notq ),
    .Q(\proj_14.net140 ));
 sg13g2_tiehi \proj_14.flop44/_1__504  (.L_HI(net548));
 sg13g2_dfrbp_1 \proj_14.flop44/_1_  (.CLK(net181),
    .RESET_B(net548),
    .D(\proj_14.net143 ),
    .Q_N(\proj_14.flop44/notq ),
    .Q(\proj_14.net142 ));
 sg13g2_tiehi \proj_14.flop45/_1__505  (.L_HI(net549));
 sg13g2_dfrbp_1 \proj_14.flop45/_1_  (.CLK(net182),
    .RESET_B(net549),
    .D(\proj_14.net146 ),
    .Q_N(\proj_14.flop45/notq ),
    .Q(\proj_14.net145 ));
 sg13g2_tiehi \proj_14.flop46/_1__506  (.L_HI(net550));
 sg13g2_dfrbp_1 \proj_14.flop46/_1_  (.CLK(net183),
    .RESET_B(net550),
    .D(\proj_14.net149 ),
    .Q_N(\proj_14.flop46/notq ),
    .Q(\proj_14.net148 ));
 sg13g2_tiehi \proj_14.flop47/_1__507  (.L_HI(net551));
 sg13g2_dfrbp_1 \proj_14.flop47/_1_  (.CLK(net184),
    .RESET_B(net551),
    .D(\proj_14.net152 ),
    .Q_N(\proj_14.flop47/notq ),
    .Q(\proj_14.net151 ));
 sg13g2_tiehi \proj_14.flop48/_1__508  (.L_HI(net552));
 sg13g2_dfrbp_1 \proj_14.flop48/_1_  (.CLK(net185),
    .RESET_B(net552),
    .D(\proj_14.net155 ),
    .Q_N(\proj_14.flop48/notq ),
    .Q(\proj_14.net154 ));
 sg13g2_tiehi \proj_14.flop49/_1__509  (.L_HI(net553));
 sg13g2_dfrbp_1 \proj_14.flop49/_1_  (.CLK(net186),
    .RESET_B(net553),
    .D(\proj_14.net158 ),
    .Q_N(\proj_14.flop49/notq ),
    .Q(\proj_14.net157 ));
 sg13g2_tiehi \proj_14.flop5/_1__510  (.L_HI(net554));
 sg13g2_dfrbp_1 \proj_14.flop5/_1_  (.CLK(net187),
    .RESET_B(net554),
    .D(\proj_14.net18 ),
    .Q_N(\proj_14.flop5/notq ),
    .Q(\proj_14.net17 ));
 sg13g2_tiehi \proj_14.flop50/_1__511  (.L_HI(net555));
 sg13g2_dfrbp_1 \proj_14.flop50/_1_  (.CLK(net188),
    .RESET_B(net555),
    .D(\proj_14.net161 ),
    .Q_N(\proj_14.flop50/notq ),
    .Q(\proj_14.net160 ));
 sg13g2_tiehi \proj_14.flop51/_1__512  (.L_HI(net556));
 sg13g2_dfrbp_1 \proj_14.flop51/_1_  (.CLK(net189),
    .RESET_B(net556),
    .D(\proj_14.net164 ),
    .Q_N(\proj_14.flop51/notq ),
    .Q(\proj_14.net163 ));
 sg13g2_tiehi \proj_14.flop52/_1__513  (.L_HI(net557));
 sg13g2_dfrbp_1 \proj_14.flop52/_1_  (.CLK(net190),
    .RESET_B(net557),
    .D(\proj_14.net167 ),
    .Q_N(\proj_14.flop52/notq ),
    .Q(\proj_14.net166 ));
 sg13g2_tiehi \proj_14.flop53/_1__514  (.L_HI(net558));
 sg13g2_dfrbp_1 \proj_14.flop53/_1_  (.CLK(net191),
    .RESET_B(net558),
    .D(\proj_14.net170 ),
    .Q_N(\proj_14.flop53/notq ),
    .Q(\proj_14.net169 ));
 sg13g2_tiehi \proj_14.flop54/_1__515  (.L_HI(net559));
 sg13g2_dfrbp_1 \proj_14.flop54/_1_  (.CLK(net192),
    .RESET_B(net559),
    .D(\proj_14.net173 ),
    .Q_N(\proj_14.flop54/notq ),
    .Q(\proj_14.net172 ));
 sg13g2_tiehi \proj_14.flop55/_1__516  (.L_HI(net560));
 sg13g2_dfrbp_1 \proj_14.flop55/_1_  (.CLK(net193),
    .RESET_B(net560),
    .D(\proj_14.net176 ),
    .Q_N(\proj_14.flop55/notq ),
    .Q(\proj_14.net175 ));
 sg13g2_tiehi \proj_14.flop56/_1__517  (.L_HI(net561));
 sg13g2_dfrbp_1 \proj_14.flop56/_1_  (.CLK(net194),
    .RESET_B(net561),
    .D(\proj_14.net179 ),
    .Q_N(\proj_14.flop56/notq ),
    .Q(\proj_14.net178 ));
 sg13g2_tiehi \proj_14.flop57/_1__518  (.L_HI(net562));
 sg13g2_dfrbp_1 \proj_14.flop57/_1_  (.CLK(net195),
    .RESET_B(net562),
    .D(\proj_14.net182 ),
    .Q_N(\proj_14.flop57/notq ),
    .Q(\proj_14.net181 ));
 sg13g2_tiehi \proj_14.flop58/_1__519  (.L_HI(net563));
 sg13g2_dfrbp_1 \proj_14.flop58/_1_  (.CLK(net196),
    .RESET_B(net563),
    .D(\proj_14.net185 ),
    .Q_N(\proj_14.flop58/notq ),
    .Q(\proj_14.net184 ));
 sg13g2_tiehi \proj_14.flop59/_1__520  (.L_HI(net564));
 sg13g2_dfrbp_1 \proj_14.flop59/_1_  (.CLK(net197),
    .RESET_B(net564),
    .D(\proj_14.net188 ),
    .Q_N(\proj_14.flop59/notq ),
    .Q(\proj_14.net187 ));
 sg13g2_tiehi \proj_14.flop6/_1__521  (.L_HI(net565));
 sg13g2_dfrbp_1 \proj_14.flop6/_1_  (.CLK(net198),
    .RESET_B(net565),
    .D(\proj_14.net21 ),
    .Q_N(\proj_14.flop6/notq ),
    .Q(\proj_14.net20 ));
 sg13g2_tiehi \proj_14.flop60/_1__522  (.L_HI(net566));
 sg13g2_dfrbp_1 \proj_14.flop60/_1_  (.CLK(net199),
    .RESET_B(net566),
    .D(\proj_14.net192 ),
    .Q_N(\proj_14.flop60/notq ),
    .Q(\proj_14.net114 ));
 sg13g2_tiehi \proj_14.flop61/_1__523  (.L_HI(net567));
 sg13g2_dfrbp_1 \proj_14.flop61/_1_  (.CLK(net200),
    .RESET_B(net567),
    .D(\proj_14.net195 ),
    .Q_N(\proj_14.flop61/notq ),
    .Q(\proj_14.net194 ));
 sg13g2_tiehi \proj_14.flop62/_1__524  (.L_HI(net568));
 sg13g2_dfrbp_1 \proj_14.flop62/_1_  (.CLK(net201),
    .RESET_B(net568),
    .D(\proj_14.net198 ),
    .Q_N(\proj_14.flop62/notq ),
    .Q(\proj_14.net197 ));
 sg13g2_tiehi \proj_14.flop63/_1__525  (.L_HI(net569));
 sg13g2_dfrbp_1 \proj_14.flop63/_1_  (.CLK(net202),
    .RESET_B(net569),
    .D(\proj_14.net201 ),
    .Q_N(\proj_14.flop63/notq ),
    .Q(\proj_14.net200 ));
 sg13g2_tiehi \proj_14.flop64/_1__526  (.L_HI(net570));
 sg13g2_dfrbp_1 \proj_14.flop64/_1_  (.CLK(net203),
    .RESET_B(net570),
    .D(\proj_14.net203 ),
    .Q_N(\proj_14.flop64/notq ),
    .Q(\proj_14.net204 ));
 sg13g2_tiehi \proj_14.flop65/_1__527  (.L_HI(net571));
 sg13g2_dfrbp_1 \proj_14.flop65/_1_  (.CLK(net204),
    .RESET_B(net571),
    .D(\proj_14.net207 ),
    .Q_N(\proj_14.flop65/notq ),
    .Q(\proj_14.net206 ));
 sg13g2_tiehi \proj_14.flop66/_1__528  (.L_HI(net572));
 sg13g2_dfrbp_1 \proj_14.flop66/_1_  (.CLK(net205),
    .RESET_B(net572),
    .D(\proj_14.net210 ),
    .Q_N(\proj_14.flop66/notq ),
    .Q(\proj_14.net209 ));
 sg13g2_tiehi \proj_14.flop67/_1__529  (.L_HI(net573));
 sg13g2_dfrbp_1 \proj_14.flop67/_1_  (.CLK(net206),
    .RESET_B(net573),
    .D(\proj_14.net213 ),
    .Q_N(\proj_14.flop67/notq ),
    .Q(\proj_14.net212 ));
 sg13g2_tiehi \proj_14.flop68/_1__530  (.L_HI(net574));
 sg13g2_dfrbp_1 \proj_14.flop68/_1_  (.CLK(net207),
    .RESET_B(net574),
    .D(\proj_14.net216 ),
    .Q_N(\proj_14.flop68/notq ),
    .Q(\proj_14.net215 ));
 sg13g2_tiehi \proj_14.flop69/_1__531  (.L_HI(net575));
 sg13g2_dfrbp_1 \proj_14.flop69/_1_  (.CLK(net208),
    .RESET_B(net575),
    .D(\proj_14.net219 ),
    .Q_N(\proj_14.flop69/notq ),
    .Q(\proj_14.net218 ));
 sg13g2_tiehi \proj_14.flop7/_1__532  (.L_HI(net576));
 sg13g2_dfrbp_1 \proj_14.flop7/_1_  (.CLK(net209),
    .RESET_B(net576),
    .D(\proj_14.net24 ),
    .Q_N(\proj_14.flop7/notq ),
    .Q(\proj_14.net23 ));
 sg13g2_tiehi \proj_14.flop70/_1__533  (.L_HI(net577));
 sg13g2_dfrbp_1 \proj_14.flop70/_1_  (.CLK(net210),
    .RESET_B(net577),
    .D(\proj_14.net222 ),
    .Q_N(\proj_14.flop70/notq ),
    .Q(\proj_14.net221 ));
 sg13g2_tiehi \proj_14.flop71/_1__534  (.L_HI(net578));
 sg13g2_dfrbp_1 \proj_14.flop71/_1_  (.CLK(net211),
    .RESET_B(net578),
    .D(\proj_14.net225 ),
    .Q_N(\proj_14.flop71/notq ),
    .Q(\proj_14.net224 ));
 sg13g2_tiehi \proj_14.flop72/_1__535  (.L_HI(net579));
 sg13g2_dfrbp_1 \proj_14.flop72/_1_  (.CLK(net212),
    .RESET_B(net579),
    .D(\proj_14.net228 ),
    .Q_N(\proj_14.flop72/notq ),
    .Q(\proj_14.net227 ));
 sg13g2_tiehi \proj_14.flop73/_1__536  (.L_HI(net580));
 sg13g2_dfrbp_1 \proj_14.flop73/_1_  (.CLK(net213),
    .RESET_B(net580),
    .D(\proj_14.net231 ),
    .Q_N(\proj_14.flop73/notq ),
    .Q(\proj_14.net230 ));
 sg13g2_tiehi \proj_14.flop74/_1__537  (.L_HI(net581));
 sg13g2_dfrbp_1 \proj_14.flop74/_1_  (.CLK(net214),
    .RESET_B(net581),
    .D(\proj_14.net234 ),
    .Q_N(\proj_14.flop74/notq ),
    .Q(\proj_14.net233 ));
 sg13g2_tiehi \proj_14.flop75/_1__538  (.L_HI(net582));
 sg13g2_dfrbp_1 \proj_14.flop75/_1_  (.CLK(net215),
    .RESET_B(net582),
    .D(\proj_14.net237 ),
    .Q_N(\proj_14.flop75/notq ),
    .Q(\proj_14.net236 ));
 sg13g2_tiehi \proj_14.flop76/_1__539  (.L_HI(net583));
 sg13g2_dfrbp_1 \proj_14.flop76/_1_  (.CLK(net216),
    .RESET_B(net583),
    .D(\proj_14.net240 ),
    .Q_N(\proj_14.flop76/notq ),
    .Q(\proj_14.net239 ));
 sg13g2_tiehi \proj_14.flop77/_1__540  (.L_HI(net584));
 sg13g2_dfrbp_1 \proj_14.flop77/_1_  (.CLK(net217),
    .RESET_B(net584),
    .D(\proj_14.net243 ),
    .Q_N(\proj_14.flop77/notq ),
    .Q(\proj_14.net242 ));
 sg13g2_tiehi \proj_14.flop78/_1__541  (.L_HI(net585));
 sg13g2_dfrbp_1 \proj_14.flop78/_1_  (.CLK(net218),
    .RESET_B(net585),
    .D(\proj_14.net246 ),
    .Q_N(\proj_14.flop78/notq ),
    .Q(\proj_14.net245 ));
 sg13g2_tiehi \proj_14.flop79/_1__542  (.L_HI(net586));
 sg13g2_dfrbp_1 \proj_14.flop79/_1_  (.CLK(net219),
    .RESET_B(net586),
    .D(\proj_14.net249 ),
    .Q_N(\proj_14.flop79/notq ),
    .Q(\proj_14.net248 ));
 sg13g2_tiehi \proj_14.flop8/_1__543  (.L_HI(net587));
 sg13g2_dfrbp_1 \proj_14.flop8/_1_  (.CLK(net220),
    .RESET_B(net587),
    .D(\proj_14.net27 ),
    .Q_N(\proj_14.flop8/notq ),
    .Q(\proj_14.net26 ));
 sg13g2_tiehi \proj_14.flop80/_1__544  (.L_HI(net588));
 sg13g2_dfrbp_1 \proj_14.flop80/_1_  (.CLK(net221),
    .RESET_B(net588),
    .D(\proj_14.net252 ),
    .Q_N(\proj_14.flop80/notq ),
    .Q(\proj_14.net251 ));
 sg13g2_tiehi \proj_14.flop81/_1__545  (.L_HI(net589));
 sg13g2_dfrbp_1 \proj_14.flop81/_1_  (.CLK(net222),
    .RESET_B(net589),
    .D(\proj_14.net256 ),
    .Q_N(\proj_14.flop81/notq ),
    .Q(\proj_14.net190 ));
 sg13g2_tiehi \proj_14.flop82/_1__546  (.L_HI(net590));
 sg13g2_dfrbp_1 \proj_14.flop82/_1_  (.CLK(net223),
    .RESET_B(net590),
    .D(\proj_14.net259 ),
    .Q_N(\proj_14.flop82/notq ),
    .Q(\proj_14.net258 ));
 sg13g2_tiehi \proj_14.flop83/_1__547  (.L_HI(net591));
 sg13g2_dfrbp_1 \proj_14.flop83/_1_  (.CLK(net224),
    .RESET_B(net591),
    .D(\proj_14.net262 ),
    .Q_N(\proj_14.flop83/notq ),
    .Q(\proj_14.net261 ));
 sg13g2_tiehi \proj_14.flop84/_1__548  (.L_HI(net592));
 sg13g2_dfrbp_1 \proj_14.flop84/_1_  (.CLK(net225),
    .RESET_B(net592),
    .D(\proj_14.net265 ),
    .Q_N(\proj_14.flop84/notq ),
    .Q(\proj_14.net264 ));
 sg13g2_tiehi \proj_14.flop85/_1__549  (.L_HI(net593));
 sg13g2_dfrbp_1 \proj_14.flop85/_1_  (.CLK(net226),
    .RESET_B(net593),
    .D(\proj_14.net267 ),
    .Q_N(\proj_14.flop85/notq ),
    .Q(\proj_14.net268 ));
 sg13g2_tiehi \proj_14.flop86/_1__550  (.L_HI(net594));
 sg13g2_dfrbp_1 \proj_14.flop86/_1_  (.CLK(net227),
    .RESET_B(net594),
    .D(\proj_14.net271 ),
    .Q_N(\proj_14.flop86/notq ),
    .Q(\proj_14.net270 ));
 sg13g2_tiehi \proj_14.flop87/_1__551  (.L_HI(net595));
 sg13g2_dfrbp_1 \proj_14.flop87/_1_  (.CLK(net228),
    .RESET_B(net595),
    .D(\proj_14.net274 ),
    .Q_N(\proj_14.flop87/notq ),
    .Q(\proj_14.net273 ));
 sg13g2_tiehi \proj_14.flop88/_1__552  (.L_HI(net596));
 sg13g2_dfrbp_1 \proj_14.flop88/_1_  (.CLK(net229),
    .RESET_B(net596),
    .D(\proj_14.net277 ),
    .Q_N(\proj_14.flop88/notq ),
    .Q(\proj_14.net276 ));
 sg13g2_tiehi \proj_14.flop89/_1__553  (.L_HI(net597));
 sg13g2_dfrbp_1 \proj_14.flop89/_1_  (.CLK(net230),
    .RESET_B(net597),
    .D(\proj_14.net280 ),
    .Q_N(\proj_14.flop89/notq ),
    .Q(\proj_14.net279 ));
 sg13g2_tiehi \proj_14.flop9/_1__554  (.L_HI(net598));
 sg13g2_dfrbp_1 \proj_14.flop9/_1_  (.CLK(net231),
    .RESET_B(net598),
    .D(\proj_14.net30 ),
    .Q_N(\proj_14.flop9/notq ),
    .Q(\proj_14.net29 ));
 sg13g2_tiehi \proj_14.flop90/_1__555  (.L_HI(net599));
 sg13g2_dfrbp_1 \proj_14.flop90/_1_  (.CLK(net232),
    .RESET_B(net599),
    .D(\proj_14.net283 ),
    .Q_N(\proj_14.flop90/notq ),
    .Q(\proj_14.net282 ));
 sg13g2_tiehi \proj_14.flop91/_1__556  (.L_HI(net600));
 sg13g2_dfrbp_1 \proj_14.flop91/_1_  (.CLK(net233),
    .RESET_B(net600),
    .D(\proj_14.net286 ),
    .Q_N(\proj_14.flop91/notq ),
    .Q(\proj_14.net285 ));
 sg13g2_tiehi \proj_14.flop92/_1__557  (.L_HI(net601));
 sg13g2_dfrbp_1 \proj_14.flop92/_1_  (.CLK(net234),
    .RESET_B(net601),
    .D(\proj_14.net289 ),
    .Q_N(\proj_14.flop92/notq ),
    .Q(\proj_14.net288 ));
 sg13g2_tiehi \proj_14.flop93/_1__558  (.L_HI(net602));
 sg13g2_dfrbp_1 \proj_14.flop93/_1_  (.CLK(net235),
    .RESET_B(net602),
    .D(\proj_14.net292 ),
    .Q_N(\proj_14.flop93/notq ),
    .Q(\proj_14.net291 ));
 sg13g2_tiehi \proj_14.flop94/_1__559  (.L_HI(net603));
 sg13g2_dfrbp_1 \proj_14.flop94/_1_  (.CLK(net236),
    .RESET_B(net603),
    .D(\proj_14.net295 ),
    .Q_N(\proj_14.flop94/notq ),
    .Q(\proj_14.net294 ));
 sg13g2_tiehi \proj_14.flop95/_1__560  (.L_HI(net604));
 sg13g2_dfrbp_1 \proj_14.flop95/_1_  (.CLK(net237),
    .RESET_B(net604),
    .D(\proj_14.net298 ),
    .Q_N(\proj_14.flop95/notq ),
    .Q(\proj_14.net297 ));
 sg13g2_tiehi \proj_14.flop96/_1__561  (.L_HI(net605));
 sg13g2_dfrbp_1 \proj_14.flop96/_1_  (.CLK(net238),
    .RESET_B(net605),
    .D(\proj_14.net301 ),
    .Q_N(\proj_14.flop96/notq ),
    .Q(\proj_14.net300 ));
 sg13g2_tiehi \proj_14.flop97/_1__562  (.L_HI(net606));
 sg13g2_dfrbp_1 \proj_14.flop97/_1_  (.CLK(net239),
    .RESET_B(net606),
    .D(\proj_14.net304 ),
    .Q_N(\proj_14.flop97/notq ),
    .Q(\proj_14.net303 ));
 sg13g2_tiehi \proj_14.flop98/_1__563  (.L_HI(net607));
 sg13g2_dfrbp_1 \proj_14.flop98/_1_  (.CLK(net240),
    .RESET_B(net607),
    .D(\proj_14.net307 ),
    .Q_N(\proj_14.flop98/notq ),
    .Q(\proj_14.net306 ));
 sg13g2_tiehi \proj_14.flop99/_1__564  (.L_HI(net608));
 sg13g2_dfrbp_1 \proj_14.flop99/_1_  (.CLK(net241),
    .RESET_B(net608),
    .D(\proj_14.net310 ),
    .Q_N(\proj_14.flop99/notq ),
    .Q(\proj_14.net309 ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_mux2_1 \proj_14.mux1/_0_  (.A0(net306),
    .A1(\proj_14.net11 ),
    .S(net149),
    .X(\proj_14.net8 ));
 sg13g2_mux2_1 \proj_14.mux10/_0_  (.A0(net242),
    .A1(\proj_14.net35 ),
    .S(net145),
    .X(\proj_14.net33 ));
 sg13g2_mux2_1 \proj_14.mux100/_0_  (.A0(net307),
    .A1(\proj_14.net312 ),
    .S(net136),
    .X(\proj_14.net310 ));
 sg13g2_mux2_1 \proj_14.mux101/_0_  (.A0(net308),
    .A1(\proj_14.net315 ),
    .S(net136),
    .X(\proj_14.net313 ));
 sg13g2_mux2_1 \proj_14.mux102/_0_  (.A0(net309),
    .A1(\proj_14.net318 ),
    .S(net136),
    .X(\proj_14.net316 ));
 sg13g2_mux2_1 \proj_14.mux103/_0_  (.A0(net310),
    .A1(\proj_14.net322 ),
    .S(net158),
    .X(\proj_14.net320 ));
 sg13g2_mux2_1 \proj_14.mux104/_0_  (.A0(net311),
    .A1(\proj_14.net325 ),
    .S(net158),
    .X(\proj_14.net323 ));
 sg13g2_mux2_1 \proj_14.mux105/_0_  (.A0(net312),
    .A1(\proj_14.net328 ),
    .S(net158),
    .X(\proj_14.net326 ));
 sg13g2_mux2_1 \proj_14.mux106/_0_  (.A0(net313),
    .A1(\proj_14.net268 ),
    .S(net158),
    .X(\proj_14.net329 ));
 sg13g2_mux2_1 \proj_14.mux107/_0_  (.A0(net314),
    .A1(\proj_14.net335 ),
    .S(net138),
    .X(\proj_14.net332 ));
 sg13g2_mux2_1 \proj_14.mux108/_0_  (.A0(net315),
    .A1(\proj_14.net338 ),
    .S(net138),
    .X(\proj_14.net336 ));
 sg13g2_mux2_1 \proj_14.mux109/_0_  (.A0(net316),
    .A1(\proj_14.net341 ),
    .S(net138),
    .X(\proj_14.net339 ));
 sg13g2_mux2_1 \proj_14.mux11/_0_  (.A0(net317),
    .A1(\proj_14.net38 ),
    .S(net145),
    .X(\proj_14.net36 ));
 sg13g2_mux2_1 \proj_14.mux110/_0_  (.A0(net318),
    .A1(\proj_14.net344 ),
    .S(net139),
    .X(\proj_14.net342 ));
 sg13g2_mux2_1 \proj_14.mux111/_0_  (.A0(net243),
    .A1(\proj_14.net347 ),
    .S(net143),
    .X(\proj_14.net345 ));
 sg13g2_mux2_1 \proj_14.mux112/_0_  (.A0(net319),
    .A1(\proj_14.net350 ),
    .S(net143),
    .X(\proj_14.net348 ));
 sg13g2_mux2_1 \proj_14.mux113/_0_  (.A0(net244),
    .A1(\proj_14.net353 ),
    .S(net143),
    .X(\proj_14.net351 ));
 sg13g2_mux2_1 \proj_14.mux114/_0_  (.A0(net245),
    .A1(\proj_14.net356 ),
    .S(net144),
    .X(\proj_14.net354 ));
 sg13g2_mux2_1 \proj_14.mux115/_0_  (.A0(net246),
    .A1(\proj_14.net359 ),
    .S(net144),
    .X(\proj_14.net357 ));
 sg13g2_mux2_1 \proj_14.mux116/_0_  (.A0(net247),
    .A1(\proj_14.net362 ),
    .S(net155),
    .X(\proj_14.net360 ));
 sg13g2_mux2_1 \proj_14.mux117/_0_  (.A0(net248),
    .A1(\proj_14.net365 ),
    .S(net155),
    .X(\proj_14.net363 ));
 sg13g2_mux2_1 \proj_14.mux118/_0_  (.A0(net320),
    .A1(\proj_14.net368 ),
    .S(net162),
    .X(\proj_14.net366 ));
 sg13g2_mux2_1 \proj_14.mux119/_0_  (.A0(net249),
    .A1(\proj_14.net371 ),
    .S(net162),
    .X(\proj_14.net369 ));
 sg13g2_mux2_1 \proj_14.mux12/_0_  (.A0(net250),
    .A1(\proj_14.net41 ),
    .S(net148),
    .X(\proj_14.net39 ));
 sg13g2_mux2_1 \proj_14.mux120/_0_  (.A0(net321),
    .A1(\proj_14.net374 ),
    .S(net163),
    .X(\proj_14.net372 ));
 sg13g2_mux2_1 \proj_14.mux121/_0_  (.A0(net322),
    .A1(\proj_14.net377 ),
    .S(net162),
    .X(\proj_14.net375 ));
 sg13g2_mux2_1 \proj_14.mux122/_0_  (.A0(net323),
    .A1(\proj_14.net380 ),
    .S(net164),
    .X(\proj_14.net378 ));
 sg13g2_mux2_1 \proj_14.mux123/_0_  (.A0(net324),
    .A1(\proj_14.net383 ),
    .S(net164),
    .X(\proj_14.net381 ));
 sg13g2_mux2_1 \proj_14.mux124/_0_  (.A0(net325),
    .A1(\proj_14.net387 ),
    .S(net136),
    .X(\proj_14.net385 ));
 sg13g2_mux2_1 \proj_14.mux125/_0_  (.A0(net326),
    .A1(\proj_14.net390 ),
    .S(net136),
    .X(\proj_14.net388 ));
 sg13g2_mux2_1 \proj_14.mux126/_0_  (.A0(net327),
    .A1(\proj_14.net393 ),
    .S(net138),
    .X(\proj_14.net391 ));
 sg13g2_mux2_1 \proj_14.mux127/_0_  (.A0(net328),
    .A1(\proj_14.net333 ),
    .S(net138),
    .X(\proj_14.net394 ));
 sg13g2_mux2_1 \proj_14.mux128/_0_  (.A0(net329),
    .A1(\proj_14.net399 ),
    .S(net160),
    .X(\proj_14.net396 ));
 sg13g2_mux2_1 \proj_14.mux129/_0_  (.A0(net330),
    .A1(\proj_14.net402 ),
    .S(net160),
    .X(\proj_14.net400 ));
 sg13g2_mux2_1 \proj_14.mux13/_0_  (.A0(net331),
    .A1(\proj_14.net44 ),
    .S(net148),
    .X(\proj_14.net42 ));
 sg13g2_mux2_1 \proj_14.mux130/_0_  (.A0(net332),
    .A1(\proj_14.net405 ),
    .S(net159),
    .X(\proj_14.net403 ));
 sg13g2_mux2_1 \proj_14.mux131/_0_  (.A0(net333),
    .A1(\proj_14.net408 ),
    .S(net159),
    .X(\proj_14.net406 ));
 sg13g2_mux2_1 \proj_14.mux132/_0_  (.A0(net251),
    .A1(\proj_14.net411 ),
    .S(net155),
    .X(\proj_14.net409 ));
 sg13g2_mux2_1 \proj_14.mux133/_0_  (.A0(net334),
    .A1(\proj_14.net414 ),
    .S(net155),
    .X(\proj_14.net412 ));
 sg13g2_mux2_1 \proj_14.mux134/_0_  (.A0(net252),
    .A1(\proj_14.net417 ),
    .S(net155),
    .X(\proj_14.net415 ));
 sg13g2_mux2_1 \proj_14.mux135/_0_  (.A0(net253),
    .A1(\proj_14.net420 ),
    .S(net153),
    .X(\proj_14.net418 ));
 sg13g2_mux2_1 \proj_14.mux136/_0_  (.A0(net335),
    .A1(\proj_14.net423 ),
    .S(net153),
    .X(\proj_14.net421 ));
 sg13g2_mux2_1 \proj_14.mux137/_0_  (.A0(net254),
    .A1(\proj_14.net426 ),
    .S(net142),
    .X(\proj_14.net424 ));
 sg13g2_mux2_1 \proj_14.mux138/_0_  (.A0(net255),
    .A1(\proj_14.net429 ),
    .S(net142),
    .X(\proj_14.net427 ));
 sg13g2_mux2_1 \proj_14.mux139/_0_  (.A0(net336),
    .A1(\proj_14.net432 ),
    .S(net143),
    .X(\proj_14.net430 ));
 sg13g2_mux2_1 \proj_14.mux14/_0_  (.A0(net256),
    .A1(\proj_14.net47 ),
    .S(net148),
    .X(\proj_14.net45 ));
 sg13g2_mux2_1 \proj_14.mux140/_0_  (.A0(net257),
    .A1(\proj_14.net435 ),
    .S(net143),
    .X(\proj_14.net433 ));
 sg13g2_mux2_1 \proj_14.mux141/_0_  (.A0(net337),
    .A1(\proj_14.net438 ),
    .S(net138),
    .X(\proj_14.net436 ));
 sg13g2_mux2_1 \proj_14.mux142/_0_  (.A0(net338),
    .A1(\proj_14.net441 ),
    .S(net137),
    .X(\proj_14.net439 ));
 sg13g2_mux2_1 \proj_14.mux143/_0_  (.A0(net339),
    .A1(\proj_14.net444 ),
    .S(net138),
    .X(\proj_14.net442 ));
 sg13g2_mux2_1 \proj_14.mux144/_0_  (.A0(net340),
    .A1(\proj_14.net447 ),
    .S(net139),
    .X(\proj_14.net445 ));
 sg13g2_mux2_1 \proj_14.mux145/_0_  (.A0(net341),
    .A1(\proj_14.net451 ),
    .S(net159),
    .X(\proj_14.net449 ));
 sg13g2_mux2_1 \proj_14.mux146/_0_  (.A0(net342),
    .A1(\proj_14.net454 ),
    .S(net160),
    .X(\proj_14.net452 ));
 sg13g2_mux2_1 \proj_14.mux147/_0_  (.A0(net343),
    .A1(\proj_14.net457 ),
    .S(net160),
    .X(\proj_14.net455 ));
 sg13g2_mux2_1 \proj_14.mux148/_0_  (.A0(net344),
    .A1(\proj_14.net397 ),
    .S(net159),
    .X(\proj_14.net458 ));
 sg13g2_mux2_1 \proj_14.mux149/_0_  (.A0(net345),
    .A1(\proj_14.net463 ),
    .S(net145),
    .X(\proj_14.net460 ));
 sg13g2_mux2_1 \proj_14.mux15/_0_  (.A0(net346),
    .A1(\proj_14.net50 ),
    .S(net145),
    .X(\proj_14.net48 ));
 sg13g2_mux2_1 \proj_14.mux150/_0_  (.A0(net347),
    .A1(\proj_14.net466 ),
    .S(net145),
    .X(\proj_14.net464 ));
 sg13g2_mux2_1 \proj_14.mux151/_0_  (.A0(net348),
    .A1(\proj_14.net469 ),
    .S(net145),
    .X(\proj_14.net467 ));
 sg13g2_mux2_1 \proj_14.mux152/_0_  (.A0(net349),
    .A1(\proj_14.net472 ),
    .S(net145),
    .X(\proj_14.net470 ));
 sg13g2_mux2_1 \proj_14.mux153/_0_  (.A0(net258),
    .A1(\proj_14.net475 ),
    .S(net145),
    .X(\proj_14.net473 ));
 sg13g2_mux2_1 \proj_14.mux154/_0_  (.A0(net259),
    .A1(\proj_14.net478 ),
    .S(net146),
    .X(\proj_14.net476 ));
 sg13g2_mux2_1 \proj_14.mux155/_0_  (.A0(net350),
    .A1(\proj_14.net481 ),
    .S(net146),
    .X(\proj_14.net479 ));
 sg13g2_mux2_1 \proj_14.mux156/_0_  (.A0(net260),
    .A1(\proj_14.net484 ),
    .S(net146),
    .X(\proj_14.net482 ));
 sg13g2_mux2_1 \proj_14.mux157/_0_  (.A0(net351),
    .A1(\proj_14.net487 ),
    .S(net146),
    .X(\proj_14.net485 ));
 sg13g2_mux2_1 \proj_14.mux158/_0_  (.A0(net261),
    .A1(\proj_14.net490 ),
    .S(net146),
    .X(\proj_14.net488 ));
 sg13g2_mux2_1 \proj_14.mux159/_0_  (.A0(net262),
    .A1(\proj_14.net493 ),
    .S(net146),
    .X(\proj_14.net491 ));
 sg13g2_mux2_1 \proj_14.mux16/_0_  (.A0(net352),
    .A1(\proj_14.net53 ),
    .S(net143),
    .X(\proj_14.net51 ));
 sg13g2_mux2_1 \proj_14.mux160/_0_  (.A0(net263),
    .A1(\proj_14.net496 ),
    .S(net146),
    .X(\proj_14.net494 ));
 sg13g2_mux2_1 \proj_14.mux161/_0_  (.A0(net264),
    .A1(\proj_14.net499 ),
    .S(net146),
    .X(\proj_14.net497 ));
 sg13g2_mux2_1 \proj_14.mux162/_0_  (.A0(net353),
    .A1(\proj_14.net502 ),
    .S(net147),
    .X(\proj_14.net500 ));
 sg13g2_mux2_1 \proj_14.mux163/_0_  (.A0(net354),
    .A1(\proj_14.net505 ),
    .S(net147),
    .X(\proj_14.net503 ));
 sg13g2_mux2_1 \proj_14.mux164/_0_  (.A0(net355),
    .A1(\proj_14.net508 ),
    .S(net147),
    .X(\proj_14.net506 ));
 sg13g2_mux2_1 \proj_14.mux165/_0_  (.A0(net356),
    .A1(\proj_14.net4 ),
    .S(net147),
    .X(\proj_14.net509 ));
 sg13g2_mux2_1 \proj_14.mux166/_0_  (.A0(net357),
    .A1(\proj_14.net514 ),
    .S(net139),
    .X(\proj_14.net512 ));
 sg13g2_mux2_1 \proj_14.mux167/_0_  (.A0(net358),
    .A1(\proj_14.net517 ),
    .S(net139),
    .X(\proj_14.net515 ));
 sg13g2_mux2_1 \proj_14.mux168/_0_  (.A0(net359),
    .A1(\proj_14.net520 ),
    .S(net139),
    .X(\proj_14.net518 ));
 sg13g2_mux2_1 \proj_14.mux169/_0_  (.A0(net360),
    .A1(\proj_14.net461 ),
    .S(net138),
    .X(\proj_14.net521 ));
 sg13g2_mux2_1 \proj_14.mux17/_0_  (.A0(net361),
    .A1(\proj_14.net56 ),
    .S(net149),
    .X(\proj_14.net54 ));
 sg13g2_mux2_1 \proj_14.mux18/_0_  (.A0(net362),
    .A1(\proj_14.net59 ),
    .S(net150),
    .X(\proj_14.net57 ));
 sg13g2_mux2_1 \proj_14.mux19/_0_  (.A0(net363),
    .A1(\proj_14.net66 ),
    .S(net162),
    .X(\proj_14.net63 ));
 sg13g2_mux2_1 \proj_14.mux2/_0_  (.A0(net364),
    .A1(\proj_14.net128 ),
    .S(net135),
    .X(\proj_14.net4 ));
 sg13g2_mux2_1 \proj_14.mux20/_0_  (.A0(net365),
    .A1(\proj_14.net69 ),
    .S(net163),
    .X(\proj_14.net67 ));
 sg13g2_mux2_1 \proj_14.mux21/_0_  (.A0(net366),
    .A1(\proj_14.net72 ),
    .S(net162),
    .X(\proj_14.net70 ));
 sg13g2_mux2_1 \proj_14.mux22/_0_  (.A0(net367),
    .A1(\proj_14.net75 ),
    .S(net164),
    .X(\proj_14.net73 ));
 sg13g2_mux2_1 \proj_14.mux23/_0_  (.A0(net265),
    .A1(\proj_14.net78 ),
    .S(net164),
    .X(\proj_14.net76 ));
 sg13g2_mux2_1 \proj_14.mux24/_0_  (.A0(net266),
    .A1(\proj_14.net81 ),
    .S(net164),
    .X(\proj_14.net79 ));
 sg13g2_mux2_1 \proj_14.mux25/_0_  (.A0(net267),
    .A1(\proj_14.net84 ),
    .S(net164),
    .X(\proj_14.net82 ));
 sg13g2_mux2_1 \proj_14.mux26/_0_  (.A0(net268),
    .A1(\proj_14.net87 ),
    .S(net164),
    .X(\proj_14.net85 ));
 sg13g2_mux2_1 \proj_14.mux27/_0_  (.A0(net368),
    .A1(\proj_14.net90 ),
    .S(net166),
    .X(\proj_14.net88 ));
 sg13g2_mux2_1 \proj_14.mux28/_0_  (.A0(net269),
    .A1(\proj_14.net93 ),
    .S(net166),
    .X(\proj_14.net91 ));
 sg13g2_mux2_1 \proj_14.mux29/_0_  (.A0(net270),
    .A1(\proj_14.net96 ),
    .S(net166),
    .X(\proj_14.net94 ));
 sg13g2_mux2_1 \proj_14.mux3/_0_  (.A0(net369),
    .A1(\proj_14.net14 ),
    .S(net149),
    .X(\proj_14.net12 ));
 sg13g2_mux2_1 \proj_14.mux30/_0_  (.A0(net370),
    .A1(\proj_14.net99 ),
    .S(net166),
    .X(\proj_14.net97 ));
 sg13g2_mux2_1 \proj_14.mux31/_0_  (.A0(net271),
    .A1(\proj_14.net102 ),
    .S(net167),
    .X(\proj_14.net100 ));
 sg13g2_mux2_1 \proj_14.mux32/_0_  (.A0(net371),
    .A1(\proj_14.net105 ),
    .S(net166),
    .X(\proj_14.net103 ));
 sg13g2_mux2_1 \proj_14.mux33/_0_  (.A0(net372),
    .A1(\proj_14.net108 ),
    .S(net167),
    .X(\proj_14.net106 ));
 sg13g2_mux2_1 \proj_14.mux34/_0_  (.A0(net373),
    .A1(\proj_14.net111 ),
    .S(net166),
    .X(\proj_14.net109 ));
 sg13g2_mux2_1 \proj_14.mux35/_0_  (.A0(net374),
    .A1(\proj_14.net114 ),
    .S(net166),
    .X(\proj_14.net112 ));
 sg13g2_mux2_1 \proj_14.mux36/_0_  (.A0(net375),
    .A1(\proj_14.net118 ),
    .S(net150),
    .X(\proj_14.net116 ));
 sg13g2_mux2_1 \proj_14.mux37/_0_  (.A0(net376),
    .A1(\proj_14.net121 ),
    .S(net162),
    .X(\proj_14.net119 ));
 sg13g2_mux2_1 \proj_14.mux38/_0_  (.A0(net377),
    .A1(\proj_14.net124 ),
    .S(net162),
    .X(\proj_14.net122 ));
 sg13g2_mux2_1 \proj_14.mux39/_0_  (.A0(net378),
    .A1(\proj_14.net64 ),
    .S(net162),
    .X(\proj_14.net125 ));
 sg13g2_mux2_1 \proj_14.mux4/_0_  (.A0(net379),
    .A1(\proj_14.net17 ),
    .S(net149),
    .X(\proj_14.net15 ));
 sg13g2_mux2_1 \proj_14.mux40/_0_  (.A0(net380),
    .A1(\proj_14.net130 ),
    .S(net150),
    .X(\proj_14.net127 ));
 sg13g2_mux2_1 \proj_14.mux41/_0_  (.A0(net381),
    .A1(\proj_14.net133 ),
    .S(net149),
    .X(\proj_14.net131 ));
 sg13g2_mux2_1 \proj_14.mux42/_0_  (.A0(net382),
    .A1(\proj_14.net136 ),
    .S(net150),
    .X(\proj_14.net134 ));
 sg13g2_mux2_1 \proj_14.mux43/_0_  (.A0(net383),
    .A1(\proj_14.net9 ),
    .S(net149),
    .X(\proj_14.net137 ));
 sg13g2_mux2_1 \proj_14.mux44/_0_  (.A0(net384),
    .A1(\proj_14.net142 ),
    .S(net165),
    .X(\proj_14.net139 ));
 sg13g2_mux2_1 \proj_14.mux45/_0_  (.A0(net385),
    .A1(\proj_14.net145 ),
    .S(net164),
    .X(\proj_14.net143 ));
 sg13g2_mux2_1 \proj_14.mux46/_0_  (.A0(net386),
    .A1(\proj_14.net148 ),
    .S(net159),
    .X(\proj_14.net146 ));
 sg13g2_mux2_1 \proj_14.mux47/_0_  (.A0(net387),
    .A1(\proj_14.net151 ),
    .S(net159),
    .X(\proj_14.net149 ));
 sg13g2_mux2_1 \proj_14.mux48/_0_  (.A0(net272),
    .A1(\proj_14.net154 ),
    .S(net159),
    .X(\proj_14.net152 ));
 sg13g2_mux2_1 \proj_14.mux49/_0_  (.A0(net388),
    .A1(\proj_14.net157 ),
    .S(net159),
    .X(\proj_14.net155 ));
 sg13g2_mux2_1 \proj_14.mux5/_0_  (.A0(net389),
    .A1(\proj_14.net20 ),
    .S(net149),
    .X(\proj_14.net18 ));
 sg13g2_mux2_1 \proj_14.mux50/_0_  (.A0(net273),
    .A1(\proj_14.net160 ),
    .S(net156),
    .X(\proj_14.net158 ));
 sg13g2_mux2_1 \proj_14.mux51/_0_  (.A0(net274),
    .A1(\proj_14.net163 ),
    .S(net156),
    .X(\proj_14.net161 ));
 sg13g2_mux2_1 \proj_14.mux52/_0_  (.A0(net275),
    .A1(\proj_14.net166 ),
    .S(net156),
    .X(\proj_14.net164 ));
 sg13g2_mux2_1 \proj_14.mux53/_0_  (.A0(net276),
    .A1(\proj_14.net169 ),
    .S(net155),
    .X(\proj_14.net167 ));
 sg13g2_mux2_1 \proj_14.mux54/_0_  (.A0(net277),
    .A1(\proj_14.net172 ),
    .S(net155),
    .X(\proj_14.net170 ));
 sg13g2_mux2_1 \proj_14.mux55/_0_  (.A0(net390),
    .A1(\proj_14.net175 ),
    .S(net155),
    .X(\proj_14.net173 ));
 sg13g2_mux2_1 \proj_14.mux56/_0_  (.A0(net278),
    .A1(\proj_14.net178 ),
    .S(net143),
    .X(\proj_14.net176 ));
 sg13g2_mux2_1 \proj_14.mux57/_0_  (.A0(net391),
    .A1(\proj_14.net181 ),
    .S(net144),
    .X(\proj_14.net179 ));
 sg13g2_mux2_1 \proj_14.mux58/_0_  (.A0(net392),
    .A1(\proj_14.net184 ),
    .S(net143),
    .X(\proj_14.net182 ));
 sg13g2_mux2_1 \proj_14.mux59/_0_  (.A0(net393),
    .A1(\proj_14.net187 ),
    .S(net141),
    .X(\proj_14.net185 ));
 sg13g2_mux2_1 \proj_14.mux6/_0_  (.A0(net279),
    .A1(\proj_14.net23 ),
    .S(net149),
    .X(\proj_14.net21 ));
 sg13g2_mux2_1 \proj_14.mux60/_0_  (.A0(net394),
    .A1(\proj_14.net190 ),
    .S(net141),
    .X(\proj_14.net188 ));
 sg13g2_mux2_1 \proj_14.mux61/_0_  (.A0(net395),
    .A1(\proj_14.net194 ),
    .S(net166),
    .X(\proj_14.net192 ));
 sg13g2_mux2_1 \proj_14.mux62/_0_  (.A0(net396),
    .A1(\proj_14.net197 ),
    .S(net165),
    .X(\proj_14.net195 ));
 sg13g2_mux2_1 \proj_14.mux63/_0_  (.A0(net397),
    .A1(\proj_14.net200 ),
    .S(net165),
    .X(\proj_14.net198 ));
 sg13g2_mux2_1 \proj_14.mux64/_0_  (.A0(net398),
    .A1(\proj_14.net140 ),
    .S(net165),
    .X(\proj_14.net201 ));
 sg13g2_mux2_1 \proj_14.mux65/_0_  (.A0(net399),
    .A1(\proj_14.net206 ),
    .S(net142),
    .X(\proj_14.net203 ));
 sg13g2_mux2_1 \proj_14.mux66/_0_  (.A0(net400),
    .A1(\proj_14.net209 ),
    .S(net153),
    .X(\proj_14.net207 ));
 sg13g2_mux2_1 \proj_14.mux67/_0_  (.A0(net401),
    .A1(\proj_14.net212 ),
    .S(net153),
    .X(\proj_14.net210 ));
 sg13g2_mux2_1 \proj_14.mux68/_0_  (.A0(net402),
    .A1(\proj_14.net215 ),
    .S(net153),
    .X(\proj_14.net213 ));
 sg13g2_mux2_1 \proj_14.mux69/_0_  (.A0(net280),
    .A1(\proj_14.net218 ),
    .S(net154),
    .X(\proj_14.net216 ));
 sg13g2_mux2_1 \proj_14.mux7/_0_  (.A0(net403),
    .A1(\proj_14.net26 ),
    .S(net151),
    .X(\proj_14.net24 ));
 sg13g2_mux2_1 \proj_14.mux70/_0_  (.A0(net404),
    .A1(\proj_14.net221 ),
    .S(net154),
    .X(\proj_14.net219 ));
 sg13g2_mux2_1 \proj_14.mux71/_0_  (.A0(net405),
    .A1(\proj_14.net224 ),
    .S(net158),
    .X(\proj_14.net222 ));
 sg13g2_mux2_1 \proj_14.mux72/_0_  (.A0(net406),
    .A1(\proj_14.net227 ),
    .S(net158),
    .X(\proj_14.net225 ));
 sg13g2_mux2_1 \proj_14.mux73/_0_  (.A0(net407),
    .A1(\proj_14.net230 ),
    .S(net158),
    .X(\proj_14.net228 ));
 sg13g2_mux2_1 \proj_14.mux74/_0_  (.A0(net281),
    .A1(\proj_14.net233 ),
    .S(net157),
    .X(\proj_14.net231 ));
 sg13g2_mux2_1 \proj_14.mux75/_0_  (.A0(net282),
    .A1(\proj_14.net236 ),
    .S(net157),
    .X(\proj_14.net234 ));
 sg13g2_mux2_1 \proj_14.mux76/_0_  (.A0(net408),
    .A1(\proj_14.net239 ),
    .S(net157),
    .X(\proj_14.net237 ));
 sg13g2_mux2_1 \proj_14.mux77/_0_  (.A0(net283),
    .A1(\proj_14.net242 ),
    .S(net157),
    .X(\proj_14.net240 ));
 sg13g2_mux2_1 \proj_14.mux78/_0_  (.A0(net409),
    .A1(\proj_14.net245 ),
    .S(net157),
    .X(\proj_14.net243 ));
 sg13g2_mux2_1 \proj_14.mux79/_0_  (.A0(net410),
    .A1(\proj_14.net248 ),
    .S(net157),
    .X(\proj_14.net246 ));
 sg13g2_mux2_1 \proj_14.mux8/_0_  (.A0(net411),
    .A1(\proj_14.net29 ),
    .S(net147),
    .X(\proj_14.net27 ));
 sg13g2_mux2_1 \proj_14.mux80/_0_  (.A0(net412),
    .A1(\proj_14.net251 ),
    .S(net157),
    .X(\proj_14.net249 ));
 sg13g2_mux2_1 \proj_14.mux81/_0_  (.A0(net413),
    .A1(\proj_14.net254 ),
    .S(net157),
    .X(\proj_14.net252 ));
 sg13g2_mux2_1 \proj_14.mux82/_0_  (.A0(net414),
    .A1(\proj_14.net258 ),
    .S(net137),
    .X(\proj_14.net256 ));
 sg13g2_mux2_1 \proj_14.mux83/_0_  (.A0(net415),
    .A1(\proj_14.net261 ),
    .S(net137),
    .X(\proj_14.net259 ));
 sg13g2_mux2_1 \proj_14.mux84/_0_  (.A0(net416),
    .A1(\proj_14.net264 ),
    .S(net141),
    .X(\proj_14.net262 ));
 sg13g2_mux2_1 \proj_14.mux85/_0_  (.A0(net417),
    .A1(\proj_14.net204 ),
    .S(net142),
    .X(\proj_14.net265 ));
 sg13g2_mux2_1 \proj_14.mux86/_0_  (.A0(net418),
    .A1(\proj_14.net270 ),
    .S(net154),
    .X(\proj_14.net267 ));
 sg13g2_mux2_1 \proj_14.mux87/_0_  (.A0(net419),
    .A1(\proj_14.net273 ),
    .S(net153),
    .X(\proj_14.net271 ));
 sg13g2_mux2_1 \proj_14.mux88/_0_  (.A0(net420),
    .A1(\proj_14.net276 ),
    .S(net154),
    .X(\proj_14.net274 ));
 sg13g2_mux2_1 \proj_14.mux89/_0_  (.A0(net421),
    .A1(\proj_14.net279 ),
    .S(net153),
    .X(\proj_14.net277 ));
 sg13g2_mux2_1 \proj_14.mux9/_0_  (.A0(net284),
    .A1(\proj_14.net32 ),
    .S(net147),
    .X(\proj_14.net30 ));
 sg13g2_mux2_1 \proj_14.mux90/_0_  (.A0(net285),
    .A1(\proj_14.net282 ),
    .S(net153),
    .X(\proj_14.net280 ));
 sg13g2_mux2_1 \proj_14.mux91/_0_  (.A0(net422),
    .A1(\proj_14.net285 ),
    .S(net141),
    .X(\proj_14.net283 ));
 sg13g2_mux2_1 \proj_14.mux92/_0_  (.A0(net423),
    .A1(\proj_14.net288 ),
    .S(net141),
    .X(\proj_14.net286 ));
 sg13g2_mux2_1 \proj_14.mux93/_0_  (.A0(net286),
    .A1(\proj_14.net291 ),
    .S(net141),
    .X(\proj_14.net289 ));
 sg13g2_mux2_1 \proj_14.mux94/_0_  (.A0(net424),
    .A1(\proj_14.net294 ),
    .S(net141),
    .X(\proj_14.net292 ));
 sg13g2_mux2_1 \proj_14.mux95/_0_  (.A0(net287),
    .A1(\proj_14.net297 ),
    .S(net141),
    .X(\proj_14.net295 ));
 sg13g2_mux2_1 \proj_14.mux96/_0_  (.A0(net288),
    .A1(\proj_14.net300 ),
    .S(net136),
    .X(\proj_14.net298 ));
 sg13g2_mux2_1 \proj_14.mux97/_0_  (.A0(net425),
    .A1(\proj_14.net303 ),
    .S(net136),
    .X(\proj_14.net301 ));
 sg13g2_mux2_1 \proj_14.mux98/_0_  (.A0(net289),
    .A1(\proj_14.net306 ),
    .S(net137),
    .X(\proj_14.net304 ));
 sg13g2_mux2_1 \proj_14.mux99/_0_  (.A0(net426),
    .A1(\proj_14.net309 ),
    .S(net136),
    .X(\proj_14.net307 ));
 sg13g2_and2_1 \proj_15.and1/_0_  (.A(net173),
    .B(net175),
    .X(\proj_15.net10 ));
 sg13g2_and2_1 \proj_15.and2/_0_  (.A(net172),
    .B(net174),
    .X(\proj_15.net14 ));
 sg13g2_nand2_1 \proj_15.nand1/_0_  (.Y(\proj_15.net11 ),
    .A(net170),
    .B(net171));
 sg13g2_inv_1 \proj_15.not1/_0_  (.Y(\proj_15.net9 ),
    .A(net178));
 sg13g2_or2_1 \proj_15.or1/_0_  (.X(\proj_15.net13 ),
    .B(net135),
    .A(net177));
 sg13g2_or2_1 \proj_15.or2/_0_  (.X(\proj_15.net15 ),
    .B(net171),
    .A(net170));
 sg13g2_xor2_1 \proj_15.xor1/_0_  (.B(net169),
    .A(net151),
    .X(\proj_15.net12 ));
 sg13g2_xor2_1 \proj_15.xor2/_0_  (.B(net169),
    .A(net151),
    .X(\proj_15.net16 ));
 sg13g2_inv_1 \proj__0.not1/_0_  (.Y(\proj__0.net4 ),
    .A(\proj__0.net11 ));
 sg13g2_inv_1 \proj__0.not2/_0_  (.Y(\proj__0.net3 ),
    .A(\proj__0.net10 ));
 sg13g2_or2_1 \proj__0.or1/_0_  (.X(\proj__0.net10 ),
    .B(net178),
    .A(\proj__0.net4 ));
 sg13g2_or2_1 \proj__0.or2/_0_  (.X(\proj__0.net11 ),
    .B(\proj__0.net3 ),
    .A(net175));
 sg13g2_nand2_1 \proj__1.nand1/_0_  (.Y(\proj__1.net9 ),
    .A(net175),
    .B(net177));
 sg13g2_inv_1 \proj__1.not3/_0_  (.Y(\proj__1.net10 ),
    .A(net172));
 sg13g2_inv_1 \proj__1.not4/_0_  (.Y(\proj__1.net11 ),
    .A(net171));
 sg13g2_and2_1 \proj__2.and1/_0_  (.A(net174),
    .B(net177),
    .X(\proj__2.net7 ));
 sg13g2_and2_1 \proj__2.and2/_0_  (.A(\proj__2.net3 ),
    .B(\proj__2.net5 ),
    .X(\proj__2.net6 ));
 sg13g2_inv_1 \proj__2.not1/_0_  (.Y(\proj__2.net3 ),
    .A(\proj__2.net14 ));
 sg13g2_inv_1 \proj__2.not2/_0_  (.Y(\proj__2.net5 ),
    .A(\proj__2.net7 ));
 sg13g2_xor2_1 \proj__2.xor1/_0_  (.B(net177),
    .A(net174),
    .X(\proj__2.net14 ));
 sg13g2_and2_1 \proj__3.and1/_0_  (.A(net2),
    .B(\proj__3.net10 ),
    .X(\proj__3.net11 ));
 sg13g2_and2_1 \proj__3.and2/_0_  (.A(net174),
    .B(net169),
    .X(\proj__3.net4 ));
 sg13g2_and2_1 \proj__3.and3/_0_  (.A(\proj__3.net12 ),
    .B(net169),
    .X(\proj__3.net13 ));
 sg13g2_and2_1 \proj__3.and4/_0_  (.A(\proj__3.net13 ),
    .B(\proj__3.net11 ),
    .X(\proj__3.net3 ));
 sg13g2_inv_1 \proj__3.not1/_0_  (.Y(\proj__3.net10 ),
    .A(net169));
 sg13g2_inv_1 \proj__3.not2/_0_  (.Y(\proj__3.net12 ),
    .A(net176));
 sg13g2_inv_1 \proj__4.not1/_0_  (.Y(\proj__4.net9 ),
    .A(net1));
 sg13g2_inv_1 \proj__4.not2/_0_  (.Y(\proj__4.net10 ),
    .A(net175));
 sg13g2_inv_1 \proj__4.not3/_0_  (.Y(\proj__4.net11 ),
    .A(net172));
 sg13g2_inv_1 \proj__4.not4/_0_  (.Y(\proj__4.net12 ),
    .A(net171));
 sg13g2_inv_1 \proj__5.not1/_0_  (.Y(\proj__5.net9 ),
    .A(net168));
 sg13g2_or2_1 \proj__5.or1/_0_  (.X(\proj__5.net8 ),
    .B(net171),
    .A(net170));
 sg13g2_and2_1 \proj__6.and2/_0_  (.A(net176),
    .B(net178),
    .X(\proj__6.net4 ));
 sg13g2_xor2_1 \proj__6.xor1/_0_  (.B(net178),
    .A(net176),
    .X(\proj__6.net3 ));
 sg13g2_xor2_1 \proj__7.xor1/_0_  (.B(net178),
    .A(net176),
    .X(\proj__7.net3 ));
 sg13g2_and2_1 \proj__8.and1/_0_  (.A(net172),
    .B(net174),
    .X(\proj__8.net18 ));
 sg13g2_and2_1 \proj__8.and2/_0_  (.A(net177),
    .B(\proj__8.net19 ),
    .X(\proj__8.net20 ));
 sg13g2_inv_1 \proj__8.not1/_0_  (.Y(\proj__8.net8 ),
    .A(\proj__8.net18 ));
 sg13g2_inv_1 \proj__8.not2/_0_  (.Y(\proj__8.net19 ),
    .A(\proj__8.net18 ));
 sg13g2_or2_1 \proj__8.or1/_0_  (.X(\proj__8.net12 ),
    .B(\proj__8.net18 ),
    .A(net170));
 sg13g2_or2_1 \proj__8.or2/_0_  (.X(\proj__8.net11 ),
    .B(\proj__8.net20 ),
    .A(\proj__8.net12 ));
 sg13g2_or2_1 \proj__8.or3/_0_  (.X(\proj__8.net7 ),
    .B(\proj__8.net20 ),
    .A(net135));
 sg13g2_or2_1 \proj__8.or4/_0_  (.X(\proj__8.net10 ),
    .B(net168),
    .A(\proj__8.net20 ));
 sg13g2_or2_1 \proj__8.or5/_0_  (.X(\proj__8.net9 ),
    .B(\proj__8.net10 ),
    .A(\proj__8.net20 ));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(net7));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(net140));
 sg13g2_buf_2 fanout137 (.A(net140),
    .X(net137));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(net140));
 sg13g2_buf_2 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(net152),
    .X(net140));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(net144));
 sg13g2_buf_2 fanout142 (.A(net144),
    .X(net142));
 sg13g2_buf_4 fanout143 (.X(net143),
    .A(net144));
 sg13g2_buf_2 fanout144 (.A(net152),
    .X(net144));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(net148));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(net148));
 sg13g2_buf_2 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(net152),
    .X(net148));
 sg13g2_buf_4 fanout149 (.X(net149),
    .A(net151));
 sg13g2_buf_2 fanout150 (.A(net151),
    .X(net150));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(net152));
 sg13g2_buf_2 fanout152 (.A(ui_in[6]),
    .X(net152));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(net156));
 sg13g2_buf_2 fanout154 (.A(net156),
    .X(net154));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(net156));
 sg13g2_buf_2 fanout156 (.A(net161),
    .X(net156));
 sg13g2_buf_4 fanout157 (.X(net157),
    .A(net158));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(net161));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(net161));
 sg13g2_buf_2 fanout160 (.A(net161),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(ui_in[6]),
    .X(net161));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(net163));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(net168));
 sg13g2_buf_4 fanout164 (.X(net164),
    .A(net167));
 sg13g2_buf_2 fanout165 (.A(net167),
    .X(net165));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(net167));
 sg13g2_buf_2 fanout167 (.A(net168),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(ui_in[6]),
    .X(net168));
 sg13g2_buf_4 fanout169 (.X(net169),
    .A(net6));
 sg13g2_buf_2 fanout170 (.A(net5),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(net4),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(net173),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(net3),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(net176),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(net2),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(net178),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(net1),
    .X(net178));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[0]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[3]),
    .X(net11));
 sg13g2_tielo \proj_10.flop1/_1__12  (.L_LO(net12));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_4 FILLER_2_70 ();
 sg13g2_fill_1 FILLER_2_74 ();
 sg13g2_fill_2 FILLER_2_79 ();
 sg13g2_decap_4 FILLER_2_85 ();
 sg13g2_fill_1 FILLER_2_89 ();
 sg13g2_decap_8 FILLER_2_100 ();
 sg13g2_decap_8 FILLER_2_107 ();
 sg13g2_decap_8 FILLER_2_114 ();
 sg13g2_decap_8 FILLER_2_121 ();
 sg13g2_decap_8 FILLER_2_128 ();
 sg13g2_decap_8 FILLER_2_135 ();
 sg13g2_decap_8 FILLER_2_142 ();
 sg13g2_decap_8 FILLER_2_149 ();
 sg13g2_decap_8 FILLER_2_156 ();
 sg13g2_decap_8 FILLER_2_163 ();
 sg13g2_decap_8 FILLER_2_170 ();
 sg13g2_decap_8 FILLER_2_177 ();
 sg13g2_decap_8 FILLER_2_184 ();
 sg13g2_decap_8 FILLER_2_191 ();
 sg13g2_decap_8 FILLER_2_198 ();
 sg13g2_decap_8 FILLER_2_205 ();
 sg13g2_decap_8 FILLER_2_212 ();
 sg13g2_decap_8 FILLER_2_219 ();
 sg13g2_decap_8 FILLER_2_226 ();
 sg13g2_decap_8 FILLER_2_233 ();
 sg13g2_decap_8 FILLER_2_240 ();
 sg13g2_decap_8 FILLER_2_247 ();
 sg13g2_decap_8 FILLER_2_254 ();
 sg13g2_decap_8 FILLER_2_261 ();
 sg13g2_decap_8 FILLER_2_268 ();
 sg13g2_decap_8 FILLER_2_275 ();
 sg13g2_decap_8 FILLER_2_282 ();
 sg13g2_decap_8 FILLER_2_289 ();
 sg13g2_decap_8 FILLER_2_296 ();
 sg13g2_decap_8 FILLER_2_303 ();
 sg13g2_decap_8 FILLER_2_310 ();
 sg13g2_decap_8 FILLER_2_317 ();
 sg13g2_decap_8 FILLER_2_324 ();
 sg13g2_decap_8 FILLER_2_331 ();
 sg13g2_decap_8 FILLER_2_338 ();
 sg13g2_decap_8 FILLER_2_345 ();
 sg13g2_decap_8 FILLER_2_352 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_373 ();
 sg13g2_decap_8 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_fill_1 FILLER_3_31 ();
 sg13g2_fill_2 FILLER_3_36 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_4 FILLER_3_56 ();
 sg13g2_fill_2 FILLER_3_100 ();
 sg13g2_decap_4 FILLER_3_132 ();
 sg13g2_fill_1 FILLER_3_136 ();
 sg13g2_fill_2 FILLER_3_141 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_fill_1 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_165 ();
 sg13g2_decap_8 FILLER_3_172 ();
 sg13g2_decap_8 FILLER_3_179 ();
 sg13g2_decap_8 FILLER_3_186 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_8 FILLER_3_207 ();
 sg13g2_decap_8 FILLER_3_214 ();
 sg13g2_decap_8 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_8 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_fill_2 FILLER_3_347 ();
 sg13g2_fill_2 FILLER_3_363 ();
 sg13g2_decap_8 FILLER_3_369 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_fill_1 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_27 ();
 sg13g2_fill_2 FILLER_4_68 ();
 sg13g2_decap_4 FILLER_4_74 ();
 sg13g2_fill_1 FILLER_4_78 ();
 sg13g2_fill_1 FILLER_4_83 ();
 sg13g2_fill_2 FILLER_4_110 ();
 sg13g2_fill_1 FILLER_4_112 ();
 sg13g2_decap_4 FILLER_4_117 ();
 sg13g2_fill_2 FILLER_4_121 ();
 sg13g2_fill_1 FILLER_4_163 ();
 sg13g2_decap_8 FILLER_4_190 ();
 sg13g2_decap_8 FILLER_4_197 ();
 sg13g2_decap_8 FILLER_4_204 ();
 sg13g2_decap_8 FILLER_4_211 ();
 sg13g2_decap_8 FILLER_4_218 ();
 sg13g2_decap_8 FILLER_4_225 ();
 sg13g2_decap_8 FILLER_4_232 ();
 sg13g2_decap_8 FILLER_4_239 ();
 sg13g2_decap_8 FILLER_4_246 ();
 sg13g2_decap_8 FILLER_4_253 ();
 sg13g2_decap_8 FILLER_4_260 ();
 sg13g2_decap_8 FILLER_4_267 ();
 sg13g2_decap_8 FILLER_4_274 ();
 sg13g2_decap_8 FILLER_4_281 ();
 sg13g2_decap_8 FILLER_4_288 ();
 sg13g2_decap_8 FILLER_4_295 ();
 sg13g2_decap_8 FILLER_4_302 ();
 sg13g2_decap_4 FILLER_4_309 ();
 sg13g2_fill_2 FILLER_4_313 ();
 sg13g2_fill_2 FILLER_4_351 ();
 sg13g2_fill_1 FILLER_4_353 ();
 sg13g2_fill_2 FILLER_4_380 ();
 sg13g2_fill_1 FILLER_4_382 ();
 sg13g2_decap_4 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_4 ();
 sg13g2_fill_2 FILLER_5_10 ();
 sg13g2_decap_8 FILLER_5_16 ();
 sg13g2_fill_2 FILLER_5_23 ();
 sg13g2_fill_1 FILLER_5_25 ();
 sg13g2_decap_8 FILLER_5_34 ();
 sg13g2_fill_2 FILLER_5_41 ();
 sg13g2_fill_1 FILLER_5_43 ();
 sg13g2_fill_1 FILLER_5_88 ();
 sg13g2_fill_2 FILLER_5_93 ();
 sg13g2_decap_8 FILLER_5_99 ();
 sg13g2_fill_1 FILLER_5_106 ();
 sg13g2_fill_2 FILLER_5_115 ();
 sg13g2_fill_2 FILLER_5_121 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_fill_2 FILLER_5_140 ();
 sg13g2_fill_2 FILLER_5_146 ();
 sg13g2_decap_8 FILLER_5_152 ();
 sg13g2_decap_8 FILLER_5_159 ();
 sg13g2_fill_2 FILLER_5_166 ();
 sg13g2_fill_2 FILLER_5_172 ();
 sg13g2_fill_2 FILLER_5_178 ();
 sg13g2_decap_8 FILLER_5_194 ();
 sg13g2_decap_8 FILLER_5_201 ();
 sg13g2_decap_8 FILLER_5_208 ();
 sg13g2_decap_8 FILLER_5_215 ();
 sg13g2_decap_8 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_229 ();
 sg13g2_decap_8 FILLER_5_236 ();
 sg13g2_decap_8 FILLER_5_243 ();
 sg13g2_decap_8 FILLER_5_250 ();
 sg13g2_decap_8 FILLER_5_257 ();
 sg13g2_decap_8 FILLER_5_264 ();
 sg13g2_decap_8 FILLER_5_271 ();
 sg13g2_decap_8 FILLER_5_278 ();
 sg13g2_decap_4 FILLER_5_285 ();
 sg13g2_fill_2 FILLER_5_289 ();
 sg13g2_fill_2 FILLER_5_317 ();
 sg13g2_fill_2 FILLER_5_323 ();
 sg13g2_decap_4 FILLER_5_329 ();
 sg13g2_fill_1 FILLER_5_333 ();
 sg13g2_fill_2 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_fill_1 FILLER_5_372 ();
 sg13g2_decap_4 FILLER_5_405 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_4 ();
 sg13g2_decap_4 FILLER_6_42 ();
 sg13g2_fill_2 FILLER_6_56 ();
 sg13g2_fill_1 FILLER_6_58 ();
 sg13g2_decap_8 FILLER_6_69 ();
 sg13g2_decap_4 FILLER_6_76 ();
 sg13g2_fill_1 FILLER_6_80 ();
 sg13g2_decap_4 FILLER_6_133 ();
 sg13g2_fill_2 FILLER_6_163 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_4 FILLER_6_182 ();
 sg13g2_fill_1 FILLER_6_186 ();
 sg13g2_fill_1 FILLER_6_217 ();
 sg13g2_decap_4 FILLER_6_222 ();
 sg13g2_fill_2 FILLER_6_226 ();
 sg13g2_fill_2 FILLER_6_242 ();
 sg13g2_fill_1 FILLER_6_248 ();
 sg13g2_fill_2 FILLER_6_259 ();
 sg13g2_fill_1 FILLER_6_261 ();
 sg13g2_decap_4 FILLER_6_272 ();
 sg13g2_fill_1 FILLER_6_276 ();
 sg13g2_decap_8 FILLER_6_281 ();
 sg13g2_decap_8 FILLER_6_288 ();
 sg13g2_fill_1 FILLER_6_295 ();
 sg13g2_fill_2 FILLER_6_300 ();
 sg13g2_decap_4 FILLER_6_306 ();
 sg13g2_fill_1 FILLER_6_310 ();
 sg13g2_fill_1 FILLER_6_325 ();
 sg13g2_decap_8 FILLER_6_330 ();
 sg13g2_decap_8 FILLER_6_337 ();
 sg13g2_decap_8 FILLER_6_344 ();
 sg13g2_fill_1 FILLER_6_351 ();
 sg13g2_decap_4 FILLER_6_378 ();
 sg13g2_fill_1 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_7 ();
 sg13g2_fill_1 FILLER_7_9 ();
 sg13g2_fill_2 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_20 ();
 sg13g2_decap_4 FILLER_7_27 ();
 sg13g2_fill_2 FILLER_7_57 ();
 sg13g2_fill_1 FILLER_7_59 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_fill_2 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_132 ();
 sg13g2_decap_8 FILLER_7_139 ();
 sg13g2_fill_2 FILLER_7_146 ();
 sg13g2_fill_1 FILLER_7_148 ();
 sg13g2_fill_1 FILLER_7_163 ();
 sg13g2_fill_2 FILLER_7_168 ();
 sg13g2_fill_2 FILLER_7_196 ();
 sg13g2_decap_4 FILLER_7_202 ();
 sg13g2_fill_1 FILLER_7_206 ();
 sg13g2_fill_2 FILLER_7_263 ();
 sg13g2_fill_1 FILLER_7_265 ();
 sg13g2_decap_4 FILLER_7_344 ();
 sg13g2_fill_1 FILLER_7_348 ();
 sg13g2_fill_2 FILLER_7_371 ();
 sg13g2_fill_2 FILLER_7_385 ();
 sg13g2_fill_1 FILLER_7_387 ();
 sg13g2_fill_2 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_398 ();
 sg13g2_decap_4 FILLER_7_405 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_4 FILLER_8_46 ();
 sg13g2_fill_1 FILLER_8_50 ();
 sg13g2_decap_8 FILLER_8_55 ();
 sg13g2_decap_8 FILLER_8_62 ();
 sg13g2_fill_2 FILLER_8_73 ();
 sg13g2_decap_8 FILLER_8_79 ();
 sg13g2_fill_1 FILLER_8_86 ();
 sg13g2_decap_4 FILLER_8_91 ();
 sg13g2_fill_2 FILLER_8_95 ();
 sg13g2_fill_2 FILLER_8_101 ();
 sg13g2_decap_4 FILLER_8_107 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_4 FILLER_8_154 ();
 sg13g2_fill_1 FILLER_8_158 ();
 sg13g2_fill_2 FILLER_8_195 ();
 sg13g2_fill_2 FILLER_8_201 ();
 sg13g2_decap_8 FILLER_8_207 ();
 sg13g2_fill_1 FILLER_8_214 ();
 sg13g2_decap_8 FILLER_8_225 ();
 sg13g2_fill_1 FILLER_8_232 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_8 FILLER_8_254 ();
 sg13g2_decap_4 FILLER_8_261 ();
 sg13g2_fill_2 FILLER_8_265 ();
 sg13g2_decap_8 FILLER_8_275 ();
 sg13g2_decap_8 FILLER_8_282 ();
 sg13g2_fill_2 FILLER_8_289 ();
 sg13g2_fill_2 FILLER_8_295 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_fill_1 FILLER_8_315 ();
 sg13g2_fill_2 FILLER_8_356 ();
 sg13g2_decap_4 FILLER_8_368 ();
 sg13g2_fill_1 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_11 ();
 sg13g2_fill_2 FILLER_9_38 ();
 sg13g2_decap_4 FILLER_9_76 ();
 sg13g2_fill_2 FILLER_9_80 ();
 sg13g2_fill_1 FILLER_9_118 ();
 sg13g2_fill_1 FILLER_9_123 ();
 sg13g2_fill_2 FILLER_9_146 ();
 sg13g2_fill_1 FILLER_9_148 ();
 sg13g2_decap_8 FILLER_9_172 ();
 sg13g2_decap_4 FILLER_9_179 ();
 sg13g2_fill_2 FILLER_9_183 ();
 sg13g2_fill_2 FILLER_9_189 ();
 sg13g2_fill_1 FILLER_9_191 ();
 sg13g2_decap_4 FILLER_9_218 ();
 sg13g2_fill_1 FILLER_9_222 ();
 sg13g2_decap_4 FILLER_9_249 ();
 sg13g2_fill_2 FILLER_9_253 ();
 sg13g2_fill_2 FILLER_9_281 ();
 sg13g2_decap_4 FILLER_9_293 ();
 sg13g2_fill_2 FILLER_9_297 ();
 sg13g2_decap_4 FILLER_9_325 ();
 sg13g2_fill_2 FILLER_9_333 ();
 sg13g2_fill_2 FILLER_9_339 ();
 sg13g2_fill_2 FILLER_9_345 ();
 sg13g2_fill_2 FILLER_9_357 ();
 sg13g2_fill_1 FILLER_9_359 ();
 sg13g2_fill_2 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_374 ();
 sg13g2_fill_2 FILLER_9_381 ();
 sg13g2_fill_1 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_14 ();
 sg13g2_fill_1 FILLER_10_16 ();
 sg13g2_fill_2 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_27 ();
 sg13g2_fill_2 FILLER_10_34 ();
 sg13g2_fill_1 FILLER_10_36 ();
 sg13g2_decap_4 FILLER_10_41 ();
 sg13g2_fill_2 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_55 ();
 sg13g2_fill_2 FILLER_10_62 ();
 sg13g2_decap_8 FILLER_10_68 ();
 sg13g2_decap_4 FILLER_10_75 ();
 sg13g2_fill_1 FILLER_10_79 ();
 sg13g2_decap_8 FILLER_10_93 ();
 sg13g2_decap_8 FILLER_10_100 ();
 sg13g2_fill_2 FILLER_10_133 ();
 sg13g2_fill_2 FILLER_10_161 ();
 sg13g2_fill_1 FILLER_10_163 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_4 FILLER_10_214 ();
 sg13g2_fill_2 FILLER_10_218 ();
 sg13g2_decap_4 FILLER_10_224 ();
 sg13g2_fill_2 FILLER_10_232 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_4 FILLER_10_245 ();
 sg13g2_decap_4 FILLER_10_253 ();
 sg13g2_fill_2 FILLER_10_257 ();
 sg13g2_fill_2 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_269 ();
 sg13g2_fill_1 FILLER_10_294 ();
 sg13g2_decap_4 FILLER_10_317 ();
 sg13g2_fill_1 FILLER_10_321 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_fill_2 FILLER_10_381 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_4 ();
 sg13g2_fill_2 FILLER_11_9 ();
 sg13g2_fill_1 FILLER_11_15 ();
 sg13g2_decap_4 FILLER_11_36 ();
 sg13g2_fill_2 FILLER_11_44 ();
 sg13g2_fill_2 FILLER_11_116 ();
 sg13g2_decap_4 FILLER_11_122 ();
 sg13g2_fill_2 FILLER_11_126 ();
 sg13g2_fill_2 FILLER_11_138 ();
 sg13g2_fill_2 FILLER_11_144 ();
 sg13g2_decap_8 FILLER_11_150 ();
 sg13g2_decap_4 FILLER_11_157 ();
 sg13g2_fill_1 FILLER_11_161 ();
 sg13g2_fill_2 FILLER_11_166 ();
 sg13g2_fill_1 FILLER_11_168 ();
 sg13g2_fill_2 FILLER_11_173 ();
 sg13g2_decap_8 FILLER_11_179 ();
 sg13g2_decap_4 FILLER_11_226 ();
 sg13g2_fill_2 FILLER_11_240 ();
 sg13g2_fill_1 FILLER_11_242 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_fill_2 FILLER_11_280 ();
 sg13g2_decap_4 FILLER_11_291 ();
 sg13g2_fill_2 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_decap_4 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_4 FILLER_11_347 ();
 sg13g2_fill_1 FILLER_11_351 ();
 sg13g2_decap_8 FILLER_11_356 ();
 sg13g2_decap_8 FILLER_11_363 ();
 sg13g2_fill_1 FILLER_11_370 ();
 sg13g2_fill_2 FILLER_11_385 ();
 sg13g2_fill_1 FILLER_11_387 ();
 sg13g2_fill_2 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_4 FILLER_12_30 ();
 sg13g2_fill_1 FILLER_12_34 ();
 sg13g2_fill_1 FILLER_12_69 ();
 sg13g2_fill_2 FILLER_12_88 ();
 sg13g2_fill_1 FILLER_12_90 ();
 sg13g2_fill_2 FILLER_12_95 ();
 sg13g2_fill_2 FILLER_12_101 ();
 sg13g2_fill_1 FILLER_12_103 ();
 sg13g2_fill_2 FILLER_12_118 ();
 sg13g2_decap_4 FILLER_12_124 ();
 sg13g2_fill_1 FILLER_12_128 ();
 sg13g2_fill_2 FILLER_12_147 ();
 sg13g2_decap_4 FILLER_12_153 ();
 sg13g2_fill_2 FILLER_12_157 ();
 sg13g2_fill_2 FILLER_12_169 ();
 sg13g2_fill_1 FILLER_12_171 ();
 sg13g2_fill_2 FILLER_12_176 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_4 FILLER_12_189 ();
 sg13g2_fill_1 FILLER_12_193 ();
 sg13g2_fill_2 FILLER_12_198 ();
 sg13g2_decap_4 FILLER_12_204 ();
 sg13g2_fill_2 FILLER_12_208 ();
 sg13g2_decap_8 FILLER_12_240 ();
 sg13g2_fill_1 FILLER_12_247 ();
 sg13g2_fill_1 FILLER_12_274 ();
 sg13g2_fill_2 FILLER_12_301 ();
 sg13g2_fill_2 FILLER_12_329 ();
 sg13g2_fill_2 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_15 ();
 sg13g2_fill_1 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_36 ();
 sg13g2_decap_4 FILLER_13_43 ();
 sg13g2_decap_8 FILLER_13_51 ();
 sg13g2_decap_8 FILLER_13_68 ();
 sg13g2_fill_2 FILLER_13_75 ();
 sg13g2_decap_8 FILLER_13_85 ();
 sg13g2_decap_4 FILLER_13_92 ();
 sg13g2_fill_2 FILLER_13_136 ();
 sg13g2_fill_2 FILLER_13_164 ();
 sg13g2_fill_1 FILLER_13_166 ();
 sg13g2_fill_2 FILLER_13_203 ();
 sg13g2_fill_1 FILLER_13_205 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_fill_2 FILLER_13_217 ();
 sg13g2_fill_2 FILLER_13_223 ();
 sg13g2_decap_4 FILLER_13_229 ();
 sg13g2_fill_1 FILLER_13_233 ();
 sg13g2_fill_2 FILLER_13_242 ();
 sg13g2_decap_4 FILLER_13_248 ();
 sg13g2_decap_8 FILLER_13_262 ();
 sg13g2_decap_8 FILLER_13_269 ();
 sg13g2_fill_2 FILLER_13_276 ();
 sg13g2_fill_1 FILLER_13_278 ();
 sg13g2_decap_8 FILLER_13_293 ();
 sg13g2_decap_8 FILLER_13_318 ();
 sg13g2_fill_2 FILLER_13_325 ();
 sg13g2_decap_4 FILLER_13_331 ();
 sg13g2_fill_2 FILLER_13_339 ();
 sg13g2_decap_8 FILLER_13_345 ();
 sg13g2_fill_1 FILLER_13_352 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_33 ();
 sg13g2_fill_2 FILLER_14_40 ();
 sg13g2_decap_4 FILLER_14_72 ();
 sg13g2_fill_2 FILLER_14_76 ();
 sg13g2_decap_4 FILLER_14_104 ();
 sg13g2_fill_2 FILLER_14_108 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_fill_2 FILLER_14_162 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_4 FILLER_14_182 ();
 sg13g2_fill_1 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_decap_4 FILLER_14_228 ();
 sg13g2_fill_1 FILLER_14_232 ();
 sg13g2_fill_1 FILLER_14_285 ();
 sg13g2_fill_2 FILLER_14_312 ();
 sg13g2_decap_4 FILLER_14_340 ();
 sg13g2_fill_1 FILLER_14_344 ();
 sg13g2_decap_4 FILLER_14_353 ();
 sg13g2_fill_2 FILLER_14_357 ();
 sg13g2_fill_2 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_28 ();
 sg13g2_fill_1 FILLER_15_30 ();
 sg13g2_decap_8 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_46 ();
 sg13g2_decap_8 FILLER_15_61 ();
 sg13g2_decap_8 FILLER_15_68 ();
 sg13g2_fill_2 FILLER_15_75 ();
 sg13g2_fill_1 FILLER_15_77 ();
 sg13g2_decap_4 FILLER_15_96 ();
 sg13g2_decap_8 FILLER_15_114 ();
 sg13g2_decap_8 FILLER_15_121 ();
 sg13g2_fill_2 FILLER_15_199 ();
 sg13g2_decap_4 FILLER_15_205 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_4 FILLER_15_252 ();
 sg13g2_decap_4 FILLER_15_260 ();
 sg13g2_fill_2 FILLER_15_268 ();
 sg13g2_decap_8 FILLER_15_274 ();
 sg13g2_fill_2 FILLER_15_281 ();
 sg13g2_decap_4 FILLER_15_287 ();
 sg13g2_fill_2 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_fill_1 FILLER_15_308 ();
 sg13g2_decap_4 FILLER_15_313 ();
 sg13g2_fill_2 FILLER_15_317 ();
 sg13g2_fill_2 FILLER_15_323 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_fill_1 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_decap_4 FILLER_15_348 ();
 sg13g2_fill_2 FILLER_15_352 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_11 ();
 sg13g2_decap_4 FILLER_16_17 ();
 sg13g2_fill_2 FILLER_16_67 ();
 sg13g2_decap_4 FILLER_16_73 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_4 FILLER_16_105 ();
 sg13g2_fill_2 FILLER_16_113 ();
 sg13g2_fill_2 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_125 ();
 sg13g2_fill_1 FILLER_16_132 ();
 sg13g2_fill_2 FILLER_16_137 ();
 sg13g2_decap_8 FILLER_16_143 ();
 sg13g2_decap_8 FILLER_16_150 ();
 sg13g2_fill_2 FILLER_16_157 ();
 sg13g2_fill_1 FILLER_16_159 ();
 sg13g2_fill_2 FILLER_16_178 ();
 sg13g2_decap_4 FILLER_16_184 ();
 sg13g2_fill_2 FILLER_16_188 ();
 sg13g2_fill_2 FILLER_16_216 ();
 sg13g2_fill_1 FILLER_16_218 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_fill_2 FILLER_16_228 ();
 sg13g2_fill_2 FILLER_16_234 ();
 sg13g2_fill_2 FILLER_16_250 ();
 sg13g2_decap_4 FILLER_16_256 ();
 sg13g2_fill_1 FILLER_16_260 ();
 sg13g2_fill_2 FILLER_16_279 ();
 sg13g2_fill_1 FILLER_16_285 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_fill_2 FILLER_16_348 ();
 sg13g2_fill_2 FILLER_16_354 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_fill_2 FILLER_16_391 ();
 sg13g2_fill_1 FILLER_16_393 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_fill_1 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_40 ();
 sg13g2_decap_8 FILLER_17_46 ();
 sg13g2_fill_1 FILLER_17_53 ();
 sg13g2_fill_2 FILLER_17_84 ();
 sg13g2_fill_1 FILLER_17_86 ();
 sg13g2_fill_2 FILLER_17_91 ();
 sg13g2_fill_1 FILLER_17_93 ();
 sg13g2_decap_4 FILLER_17_98 ();
 sg13g2_fill_1 FILLER_17_102 ();
 sg13g2_fill_2 FILLER_17_117 ();
 sg13g2_fill_2 FILLER_17_123 ();
 sg13g2_fill_2 FILLER_17_129 ();
 sg13g2_fill_1 FILLER_17_131 ();
 sg13g2_fill_2 FILLER_17_142 ();
 sg13g2_fill_2 FILLER_17_148 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_fill_1 FILLER_17_165 ();
 sg13g2_fill_2 FILLER_17_170 ();
 sg13g2_fill_1 FILLER_17_176 ();
 sg13g2_decap_8 FILLER_17_191 ();
 sg13g2_decap_4 FILLER_17_198 ();
 sg13g2_fill_1 FILLER_17_202 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_213 ();
 sg13g2_decap_8 FILLER_17_229 ();
 sg13g2_fill_1 FILLER_17_236 ();
 sg13g2_fill_2 FILLER_17_267 ();
 sg13g2_fill_1 FILLER_17_269 ();
 sg13g2_fill_2 FILLER_17_310 ();
 sg13g2_fill_1 FILLER_17_312 ();
 sg13g2_fill_2 FILLER_17_317 ();
 sg13g2_fill_2 FILLER_17_323 ();
 sg13g2_fill_1 FILLER_17_325 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_4 FILLER_17_384 ();
 sg13g2_fill_2 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_4 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_53 ();
 sg13g2_fill_2 FILLER_18_64 ();
 sg13g2_fill_1 FILLER_18_66 ();
 sg13g2_fill_2 FILLER_18_71 ();
 sg13g2_fill_2 FILLER_18_165 ();
 sg13g2_fill_1 FILLER_18_197 ();
 sg13g2_decap_4 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_246 ();
 sg13g2_decap_8 FILLER_18_253 ();
 sg13g2_fill_2 FILLER_18_260 ();
 sg13g2_decap_8 FILLER_18_276 ();
 sg13g2_decap_8 FILLER_18_283 ();
 sg13g2_decap_4 FILLER_18_290 ();
 sg13g2_decap_8 FILLER_18_324 ();
 sg13g2_decap_4 FILLER_18_331 ();
 sg13g2_fill_1 FILLER_18_335 ();
 sg13g2_decap_4 FILLER_18_344 ();
 sg13g2_fill_2 FILLER_18_353 ();
 sg13g2_fill_2 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_4 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_32 ();
 sg13g2_fill_2 FILLER_19_60 ();
 sg13g2_decap_8 FILLER_19_88 ();
 sg13g2_decap_4 FILLER_19_95 ();
 sg13g2_fill_1 FILLER_19_99 ();
 sg13g2_decap_4 FILLER_19_104 ();
 sg13g2_decap_8 FILLER_19_118 ();
 sg13g2_decap_8 FILLER_19_125 ();
 sg13g2_decap_4 FILLER_19_132 ();
 sg13g2_fill_1 FILLER_19_136 ();
 sg13g2_decap_8 FILLER_19_141 ();
 sg13g2_decap_8 FILLER_19_148 ();
 sg13g2_decap_4 FILLER_19_155 ();
 sg13g2_fill_1 FILLER_19_159 ();
 sg13g2_decap_8 FILLER_19_164 ();
 sg13g2_decap_8 FILLER_19_171 ();
 sg13g2_fill_2 FILLER_19_178 ();
 sg13g2_fill_1 FILLER_19_180 ();
 sg13g2_decap_8 FILLER_19_191 ();
 sg13g2_decap_8 FILLER_19_198 ();
 sg13g2_decap_8 FILLER_19_220 ();
 sg13g2_fill_2 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_259 ();
 sg13g2_fill_2 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_303 ();
 sg13g2_fill_2 FILLER_19_308 ();
 sg13g2_decap_4 FILLER_19_318 ();
 sg13g2_fill_1 FILLER_19_322 ();
 sg13g2_fill_1 FILLER_19_333 ();
 sg13g2_fill_2 FILLER_19_338 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_4 FILLER_19_351 ();
 sg13g2_fill_1 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_fill_2 FILLER_20_56 ();
 sg13g2_fill_2 FILLER_20_62 ();
 sg13g2_fill_1 FILLER_20_64 ();
 sg13g2_fill_2 FILLER_20_117 ();
 sg13g2_fill_1 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_fill_2 FILLER_20_189 ();
 sg13g2_fill_2 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_227 ();
 sg13g2_fill_1 FILLER_20_234 ();
 sg13g2_decap_8 FILLER_20_239 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_decap_8 FILLER_20_253 ();
 sg13g2_decap_8 FILLER_20_260 ();
 sg13g2_fill_2 FILLER_20_267 ();
 sg13g2_fill_2 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_279 ();
 sg13g2_decap_4 FILLER_20_286 ();
 sg13g2_fill_2 FILLER_20_290 ();
 sg13g2_fill_2 FILLER_20_296 ();
 sg13g2_fill_1 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_decap_4 FILLER_20_379 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_4 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_18 ();
 sg13g2_fill_2 FILLER_21_49 ();
 sg13g2_fill_1 FILLER_21_51 ();
 sg13g2_fill_2 FILLER_21_62 ();
 sg13g2_fill_1 FILLER_21_64 ();
 sg13g2_decap_4 FILLER_21_69 ();
 sg13g2_fill_2 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_83 ();
 sg13g2_decap_4 FILLER_21_90 ();
 sg13g2_fill_1 FILLER_21_94 ();
 sg13g2_fill_2 FILLER_21_99 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_4 FILLER_21_116 ();
 sg13g2_fill_2 FILLER_21_120 ();
 sg13g2_fill_2 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_146 ();
 sg13g2_fill_1 FILLER_21_185 ();
 sg13g2_decap_4 FILLER_21_190 ();
 sg13g2_fill_2 FILLER_21_194 ();
 sg13g2_fill_2 FILLER_21_200 ();
 sg13g2_decap_4 FILLER_21_206 ();
 sg13g2_fill_2 FILLER_21_210 ();
 sg13g2_fill_1 FILLER_21_248 ();
 sg13g2_decap_8 FILLER_21_267 ();
 sg13g2_fill_1 FILLER_21_274 ();
 sg13g2_fill_2 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_317 ();
 sg13g2_decap_8 FILLER_21_324 ();
 sg13g2_decap_8 FILLER_21_331 ();
 sg13g2_decap_8 FILLER_21_338 ();
 sg13g2_decap_4 FILLER_21_345 ();
 sg13g2_fill_1 FILLER_21_349 ();
 sg13g2_decap_4 FILLER_21_380 ();
 sg13g2_fill_2 FILLER_21_392 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_4 ();
 sg13g2_fill_2 FILLER_22_9 ();
 sg13g2_fill_2 FILLER_22_15 ();
 sg13g2_fill_1 FILLER_22_17 ();
 sg13g2_fill_2 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_34 ();
 sg13g2_decap_8 FILLER_22_41 ();
 sg13g2_fill_2 FILLER_22_48 ();
 sg13g2_decap_4 FILLER_22_80 ();
 sg13g2_fill_2 FILLER_22_84 ();
 sg13g2_fill_2 FILLER_22_90 ();
 sg13g2_decap_4 FILLER_22_96 ();
 sg13g2_fill_2 FILLER_22_100 ();
 sg13g2_fill_2 FILLER_22_132 ();
 sg13g2_fill_2 FILLER_22_160 ();
 sg13g2_fill_1 FILLER_22_192 ();
 sg13g2_fill_2 FILLER_22_197 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_4 FILLER_22_210 ();
 sg13g2_fill_1 FILLER_22_214 ();
 sg13g2_fill_1 FILLER_22_225 ();
 sg13g2_decap_4 FILLER_22_230 ();
 sg13g2_fill_2 FILLER_22_234 ();
 sg13g2_fill_2 FILLER_22_250 ();
 sg13g2_decap_8 FILLER_22_296 ();
 sg13g2_decap_4 FILLER_22_339 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_decap_4 FILLER_22_354 ();
 sg13g2_fill_1 FILLER_22_358 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_fill_2 FILLER_22_383 ();
 sg13g2_fill_2 FILLER_22_389 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_fill_1 FILLER_23_34 ();
 sg13g2_fill_2 FILLER_23_53 ();
 sg13g2_fill_2 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_65 ();
 sg13g2_decap_4 FILLER_23_76 ();
 sg13g2_fill_1 FILLER_23_80 ();
 sg13g2_decap_4 FILLER_23_125 ();
 sg13g2_fill_2 FILLER_23_129 ();
 sg13g2_decap_4 FILLER_23_135 ();
 sg13g2_fill_2 FILLER_23_143 ();
 sg13g2_decap_4 FILLER_23_149 ();
 sg13g2_fill_1 FILLER_23_157 ();
 sg13g2_decap_4 FILLER_23_162 ();
 sg13g2_fill_1 FILLER_23_166 ();
 sg13g2_fill_2 FILLER_23_171 ();
 sg13g2_fill_1 FILLER_23_177 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_261 ();
 sg13g2_fill_2 FILLER_23_268 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_decap_4 FILLER_23_275 ();
 sg13g2_fill_2 FILLER_23_283 ();
 sg13g2_decap_8 FILLER_23_289 ();
 sg13g2_decap_8 FILLER_23_296 ();
 sg13g2_fill_2 FILLER_23_303 ();
 sg13g2_fill_1 FILLER_23_305 ();
 sg13g2_fill_2 FILLER_23_310 ();
 sg13g2_decap_8 FILLER_23_316 ();
 sg13g2_decap_4 FILLER_23_323 ();
 sg13g2_fill_1 FILLER_23_327 ();
 sg13g2_fill_2 FILLER_23_368 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_21 ();
 sg13g2_fill_2 FILLER_24_30 ();
 sg13g2_decap_8 FILLER_24_36 ();
 sg13g2_fill_2 FILLER_24_43 ();
 sg13g2_decap_4 FILLER_24_75 ();
 sg13g2_fill_2 FILLER_24_79 ();
 sg13g2_decap_4 FILLER_24_86 ();
 sg13g2_decap_8 FILLER_24_94 ();
 sg13g2_decap_4 FILLER_24_101 ();
 sg13g2_fill_1 FILLER_24_115 ();
 sg13g2_decap_8 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_127 ();
 sg13g2_decap_8 FILLER_24_138 ();
 sg13g2_fill_2 FILLER_24_145 ();
 sg13g2_fill_1 FILLER_24_147 ();
 sg13g2_fill_2 FILLER_24_158 ();
 sg13g2_fill_2 FILLER_24_164 ();
 sg13g2_decap_8 FILLER_24_170 ();
 sg13g2_decap_4 FILLER_24_177 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_fill_2 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_236 ();
 sg13g2_decap_8 FILLER_24_243 ();
 sg13g2_fill_1 FILLER_24_300 ();
 sg13g2_decap_4 FILLER_24_327 ();
 sg13g2_fill_1 FILLER_24_331 ();
 sg13g2_fill_1 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_fill_2 FILLER_24_348 ();
 sg13g2_fill_2 FILLER_24_354 ();
 sg13g2_fill_2 FILLER_24_360 ();
 sg13g2_fill_1 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_4 FILLER_24_381 ();
 sg13g2_fill_2 FILLER_24_385 ();
 sg13g2_fill_2 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_47 ();
 sg13g2_decap_4 FILLER_25_54 ();
 sg13g2_fill_1 FILLER_25_58 ();
 sg13g2_decap_8 FILLER_25_73 ();
 sg13g2_decap_4 FILLER_25_80 ();
 sg13g2_fill_1 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_145 ();
 sg13g2_fill_2 FILLER_25_152 ();
 sg13g2_fill_1 FILLER_25_154 ();
 sg13g2_fill_2 FILLER_25_191 ();
 sg13g2_fill_1 FILLER_25_193 ();
 sg13g2_decap_4 FILLER_25_220 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_fill_2 FILLER_25_229 ();
 sg13g2_fill_1 FILLER_25_231 ();
 sg13g2_fill_1 FILLER_25_236 ();
 sg13g2_decap_4 FILLER_25_247 ();
 sg13g2_fill_1 FILLER_25_281 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_fill_2 FILLER_25_315 ();
 sg13g2_decap_4 FILLER_25_377 ();
 sg13g2_fill_1 FILLER_25_381 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_4 ();
 sg13g2_fill_2 FILLER_26_10 ();
 sg13g2_decap_8 FILLER_26_16 ();
 sg13g2_decap_8 FILLER_26_23 ();
 sg13g2_fill_1 FILLER_26_30 ();
 sg13g2_decap_8 FILLER_26_41 ();
 sg13g2_decap_4 FILLER_26_48 ();
 sg13g2_decap_4 FILLER_26_90 ();
 sg13g2_fill_2 FILLER_26_94 ();
 sg13g2_decap_8 FILLER_26_100 ();
 sg13g2_fill_2 FILLER_26_107 ();
 sg13g2_decap_8 FILLER_26_113 ();
 sg13g2_fill_2 FILLER_26_120 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_4 FILLER_26_137 ();
 sg13g2_fill_1 FILLER_26_145 ();
 sg13g2_decap_8 FILLER_26_160 ();
 sg13g2_decap_4 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_171 ();
 sg13g2_fill_2 FILLER_26_177 ();
 sg13g2_fill_1 FILLER_26_179 ();
 sg13g2_decap_8 FILLER_26_188 ();
 sg13g2_decap_4 FILLER_26_195 ();
 sg13g2_fill_2 FILLER_26_203 ();
 sg13g2_fill_2 FILLER_26_209 ();
 sg13g2_decap_8 FILLER_26_251 ();
 sg13g2_fill_2 FILLER_26_258 ();
 sg13g2_fill_2 FILLER_26_264 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_fill_2 FILLER_26_284 ();
 sg13g2_fill_1 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_291 ();
 sg13g2_decap_4 FILLER_26_297 ();
 sg13g2_decap_8 FILLER_26_331 ();
 sg13g2_fill_2 FILLER_26_342 ();
 sg13g2_fill_1 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_decap_4 FILLER_26_356 ();
 sg13g2_fill_2 FILLER_26_360 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_27 ();
 sg13g2_decap_4 FILLER_27_59 ();
 sg13g2_fill_2 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_69 ();
 sg13g2_decap_4 FILLER_27_75 ();
 sg13g2_fill_1 FILLER_27_79 ();
 sg13g2_decap_8 FILLER_27_116 ();
 sg13g2_fill_2 FILLER_27_123 ();
 sg13g2_fill_1 FILLER_27_125 ();
 sg13g2_decap_4 FILLER_27_162 ();
 sg13g2_fill_2 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_194 ();
 sg13g2_decap_8 FILLER_27_199 ();
 sg13g2_decap_4 FILLER_27_206 ();
 sg13g2_fill_1 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_223 ();
 sg13g2_decap_8 FILLER_27_230 ();
 sg13g2_decap_4 FILLER_27_237 ();
 sg13g2_fill_2 FILLER_27_241 ();
 sg13g2_decap_4 FILLER_27_255 ();
 sg13g2_fill_2 FILLER_27_259 ();
 sg13g2_decap_4 FILLER_27_287 ();
 sg13g2_fill_2 FILLER_27_291 ();
 sg13g2_decap_8 FILLER_27_298 ();
 sg13g2_fill_1 FILLER_27_305 ();
 sg13g2_fill_2 FILLER_27_310 ();
 sg13g2_decap_4 FILLER_27_316 ();
 sg13g2_fill_1 FILLER_27_320 ();
 sg13g2_decap_4 FILLER_27_357 ();
 sg13g2_fill_2 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_14 ();
 sg13g2_decap_4 FILLER_28_32 ();
 sg13g2_fill_2 FILLER_28_36 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_48 ();
 sg13g2_decap_8 FILLER_28_86 ();
 sg13g2_fill_2 FILLER_28_93 ();
 sg13g2_fill_2 FILLER_28_99 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_fill_2 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_144 ();
 sg13g2_fill_1 FILLER_28_146 ();
 sg13g2_decap_4 FILLER_28_151 ();
 sg13g2_fill_2 FILLER_28_159 ();
 sg13g2_decap_8 FILLER_28_165 ();
 sg13g2_fill_2 FILLER_28_172 ();
 sg13g2_fill_2 FILLER_28_177 ();
 sg13g2_fill_1 FILLER_28_179 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_fill_2 FILLER_28_217 ();
 sg13g2_fill_1 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_236 ();
 sg13g2_fill_1 FILLER_28_238 ();
 sg13g2_fill_2 FILLER_28_277 ();
 sg13g2_fill_1 FILLER_28_314 ();
 sg13g2_decap_8 FILLER_28_319 ();
 sg13g2_fill_2 FILLER_28_330 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_fill_2 FILLER_28_343 ();
 sg13g2_fill_1 FILLER_28_345 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_26 ();
 sg13g2_decap_4 FILLER_29_33 ();
 sg13g2_fill_1 FILLER_29_37 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_4 FILLER_29_60 ();
 sg13g2_fill_2 FILLER_29_123 ();
 sg13g2_fill_2 FILLER_29_129 ();
 sg13g2_fill_2 FILLER_29_135 ();
 sg13g2_decap_8 FILLER_29_141 ();
 sg13g2_fill_2 FILLER_29_148 ();
 sg13g2_fill_2 FILLER_29_176 ();
 sg13g2_fill_2 FILLER_29_188 ();
 sg13g2_fill_1 FILLER_29_190 ();
 sg13g2_decap_8 FILLER_29_199 ();
 sg13g2_decap_4 FILLER_29_206 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_fill_1 FILLER_29_219 ();
 sg13g2_decap_8 FILLER_29_240 ();
 sg13g2_decap_8 FILLER_29_258 ();
 sg13g2_decap_4 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_283 ();
 sg13g2_fill_2 FILLER_29_288 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_299 ();
 sg13g2_fill_1 FILLER_29_303 ();
 sg13g2_decap_8 FILLER_29_338 ();
 sg13g2_fill_1 FILLER_29_349 ();
 sg13g2_fill_2 FILLER_29_364 ();
 sg13g2_fill_1 FILLER_29_366 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_fill_1 FILLER_29_378 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_fill_1 FILLER_30_9 ();
 sg13g2_fill_1 FILLER_30_50 ();
 sg13g2_fill_2 FILLER_30_55 ();
 sg13g2_fill_1 FILLER_30_57 ();
 sg13g2_decap_8 FILLER_30_66 ();
 sg13g2_decap_4 FILLER_30_73 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_fill_2 FILLER_30_96 ();
 sg13g2_decap_8 FILLER_30_102 ();
 sg13g2_fill_2 FILLER_30_109 ();
 sg13g2_decap_4 FILLER_30_115 ();
 sg13g2_fill_2 FILLER_30_123 ();
 sg13g2_fill_1 FILLER_30_125 ();
 sg13g2_decap_8 FILLER_30_155 ();
 sg13g2_decap_8 FILLER_30_162 ();
 sg13g2_decap_8 FILLER_30_169 ();
 sg13g2_fill_2 FILLER_30_186 ();
 sg13g2_fill_2 FILLER_30_206 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_decap_8 FILLER_30_244 ();
 sg13g2_decap_4 FILLER_30_251 ();
 sg13g2_fill_1 FILLER_30_255 ();
 sg13g2_fill_2 FILLER_30_262 ();
 sg13g2_fill_1 FILLER_30_264 ();
 sg13g2_decap_4 FILLER_30_279 ();
 sg13g2_fill_1 FILLER_30_294 ();
 sg13g2_decap_4 FILLER_30_300 ();
 sg13g2_fill_2 FILLER_30_304 ();
 sg13g2_fill_2 FILLER_30_332 ();
 sg13g2_fill_1 FILLER_30_334 ();
 sg13g2_fill_2 FILLER_30_370 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_14 ();
 sg13g2_fill_1 FILLER_31_18 ();
 sg13g2_fill_2 FILLER_31_23 ();
 sg13g2_decap_8 FILLER_31_29 ();
 sg13g2_fill_1 FILLER_31_36 ();
 sg13g2_decap_8 FILLER_31_73 ();
 sg13g2_fill_2 FILLER_31_80 ();
 sg13g2_fill_1 FILLER_31_118 ();
 sg13g2_fill_2 FILLER_31_123 ();
 sg13g2_decap_8 FILLER_31_129 ();
 sg13g2_decap_8 FILLER_31_136 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_fill_2 FILLER_31_187 ();
 sg13g2_fill_2 FILLER_31_194 ();
 sg13g2_fill_2 FILLER_31_213 ();
 sg13g2_decap_8 FILLER_31_228 ();
 sg13g2_decap_4 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_291 ();
 sg13g2_decap_8 FILLER_31_298 ();
 sg13g2_decap_4 FILLER_31_305 ();
 sg13g2_fill_1 FILLER_31_309 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_decap_8 FILLER_31_320 ();
 sg13g2_decap_8 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_341 ();
 sg13g2_decap_4 FILLER_31_347 ();
 sg13g2_fill_2 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_361 ();
 sg13g2_decap_4 FILLER_31_368 ();
 sg13g2_fill_2 FILLER_31_372 ();
 sg13g2_decap_8 FILLER_31_396 ();
 sg13g2_decap_4 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_4 FILLER_32_35 ();
 sg13g2_decap_4 FILLER_32_53 ();
 sg13g2_decap_4 FILLER_32_61 ();
 sg13g2_fill_1 FILLER_32_65 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_4 FILLER_32_77 ();
 sg13g2_fill_1 FILLER_32_81 ();
 sg13g2_fill_1 FILLER_32_86 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_decap_4 FILLER_32_97 ();
 sg13g2_fill_1 FILLER_32_101 ();
 sg13g2_decap_4 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_110 ();
 sg13g2_decap_8 FILLER_32_141 ();
 sg13g2_fill_2 FILLER_32_157 ();
 sg13g2_decap_8 FILLER_32_163 ();
 sg13g2_decap_4 FILLER_32_170 ();
 sg13g2_fill_1 FILLER_32_174 ();
 sg13g2_fill_2 FILLER_32_184 ();
 sg13g2_fill_1 FILLER_32_191 ();
 sg13g2_decap_4 FILLER_32_200 ();
 sg13g2_fill_1 FILLER_32_204 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_fill_1 FILLER_32_218 ();
 sg13g2_fill_1 FILLER_32_224 ();
 sg13g2_decap_4 FILLER_32_233 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_decap_4 FILLER_32_277 ();
 sg13g2_fill_2 FILLER_32_281 ();
 sg13g2_fill_1 FILLER_32_300 ();
 sg13g2_decap_4 FILLER_32_309 ();
 sg13g2_decap_8 FILLER_32_367 ();
 sg13g2_decap_4 FILLER_32_374 ();
 sg13g2_fill_1 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_4 FILLER_33_35 ();
 sg13g2_fill_2 FILLER_33_39 ();
 sg13g2_decap_8 FILLER_33_117 ();
 sg13g2_decap_4 FILLER_33_124 ();
 sg13g2_fill_2 FILLER_33_132 ();
 sg13g2_decap_8 FILLER_33_138 ();
 sg13g2_fill_1 FILLER_33_145 ();
 sg13g2_decap_8 FILLER_33_172 ();
 sg13g2_decap_4 FILLER_33_179 ();
 sg13g2_decap_4 FILLER_33_194 ();
 sg13g2_fill_1 FILLER_33_198 ();
 sg13g2_fill_2 FILLER_33_216 ();
 sg13g2_decap_8 FILLER_33_236 ();
 sg13g2_fill_1 FILLER_33_254 ();
 sg13g2_decap_4 FILLER_33_273 ();
 sg13g2_fill_2 FILLER_33_296 ();
 sg13g2_decap_8 FILLER_33_311 ();
 sg13g2_decap_8 FILLER_33_318 ();
 sg13g2_fill_2 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_335 ();
 sg13g2_decap_8 FILLER_33_342 ();
 sg13g2_decap_4 FILLER_33_349 ();
 sg13g2_fill_1 FILLER_33_353 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_fill_1 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_59 ();
 sg13g2_decap_8 FILLER_34_64 ();
 sg13g2_decap_8 FILLER_34_71 ();
 sg13g2_decap_4 FILLER_34_92 ();
 sg13g2_fill_2 FILLER_34_96 ();
 sg13g2_fill_2 FILLER_34_155 ();
 sg13g2_fill_2 FILLER_34_165 ();
 sg13g2_fill_1 FILLER_34_167 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_fill_1 FILLER_34_187 ();
 sg13g2_fill_1 FILLER_34_194 ();
 sg13g2_decap_8 FILLER_34_209 ();
 sg13g2_decap_8 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_239 ();
 sg13g2_fill_2 FILLER_34_248 ();
 sg13g2_decap_8 FILLER_34_254 ();
 sg13g2_decap_8 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_284 ();
 sg13g2_decap_4 FILLER_34_293 ();
 sg13g2_fill_1 FILLER_34_297 ();
 sg13g2_decap_4 FILLER_34_303 ();
 sg13g2_fill_2 FILLER_34_343 ();
 sg13g2_fill_1 FILLER_34_345 ();
 sg13g2_fill_2 FILLER_34_356 ();
 sg13g2_fill_2 FILLER_34_362 ();
 sg13g2_decap_4 FILLER_34_372 ();
 sg13g2_fill_1 FILLER_34_376 ();
 sg13g2_fill_1 FILLER_34_381 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_18 ();
 sg13g2_fill_2 FILLER_35_24 ();
 sg13g2_decap_8 FILLER_35_48 ();
 sg13g2_fill_1 FILLER_35_69 ();
 sg13g2_decap_8 FILLER_35_74 ();
 sg13g2_decap_4 FILLER_35_81 ();
 sg13g2_fill_2 FILLER_35_89 ();
 sg13g2_decap_8 FILLER_35_95 ();
 sg13g2_decap_4 FILLER_35_102 ();
 sg13g2_fill_1 FILLER_35_106 ();
 sg13g2_fill_2 FILLER_35_111 ();
 sg13g2_fill_1 FILLER_35_113 ();
 sg13g2_decap_8 FILLER_35_118 ();
 sg13g2_decap_4 FILLER_35_125 ();
 sg13g2_fill_1 FILLER_35_129 ();
 sg13g2_fill_2 FILLER_35_134 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_fill_2 FILLER_35_157 ();
 sg13g2_fill_2 FILLER_35_175 ();
 sg13g2_decap_4 FILLER_35_196 ();
 sg13g2_fill_2 FILLER_35_208 ();
 sg13g2_fill_2 FILLER_35_227 ();
 sg13g2_decap_4 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_260 ();
 sg13g2_decap_4 FILLER_35_301 ();
 sg13g2_fill_1 FILLER_35_305 ();
 sg13g2_fill_2 FILLER_35_324 ();
 sg13g2_fill_1 FILLER_35_330 ();
 sg13g2_decap_8 FILLER_35_335 ();
 sg13g2_decap_4 FILLER_35_342 ();
 sg13g2_fill_1 FILLER_35_386 ();
 sg13g2_fill_2 FILLER_35_391 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_52 ();
 sg13g2_fill_1 FILLER_36_54 ();
 sg13g2_decap_8 FILLER_36_85 ();
 sg13g2_decap_8 FILLER_36_92 ();
 sg13g2_decap_8 FILLER_36_99 ();
 sg13g2_decap_8 FILLER_36_106 ();
 sg13g2_decap_8 FILLER_36_113 ();
 sg13g2_decap_4 FILLER_36_120 ();
 sg13g2_fill_1 FILLER_36_124 ();
 sg13g2_fill_1 FILLER_36_151 ();
 sg13g2_fill_2 FILLER_36_166 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_fill_1 FILLER_36_182 ();
 sg13g2_fill_2 FILLER_36_203 ();
 sg13g2_decap_4 FILLER_36_209 ();
 sg13g2_fill_1 FILLER_36_216 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_4 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_258 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_decap_4 FILLER_36_277 ();
 sg13g2_decap_8 FILLER_36_298 ();
 sg13g2_decap_4 FILLER_36_305 ();
 sg13g2_fill_2 FILLER_36_309 ();
 sg13g2_decap_4 FILLER_36_315 ();
 sg13g2_fill_2 FILLER_36_319 ();
 sg13g2_decap_4 FILLER_36_351 ();
 sg13g2_fill_1 FILLER_36_359 ();
 sg13g2_decap_4 FILLER_36_370 ();
 sg13g2_fill_1 FILLER_36_374 ();
 sg13g2_fill_2 FILLER_36_379 ();
 sg13g2_fill_1 FILLER_36_381 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_4 FILLER_37_21 ();
 sg13g2_fill_2 FILLER_37_25 ();
 sg13g2_fill_1 FILLER_37_57 ();
 sg13g2_decap_8 FILLER_37_72 ();
 sg13g2_decap_8 FILLER_37_79 ();
 sg13g2_decap_8 FILLER_37_86 ();
 sg13g2_decap_8 FILLER_37_93 ();
 sg13g2_decap_8 FILLER_37_100 ();
 sg13g2_decap_8 FILLER_37_107 ();
 sg13g2_decap_8 FILLER_37_114 ();
 sg13g2_decap_8 FILLER_37_121 ();
 sg13g2_fill_1 FILLER_37_128 ();
 sg13g2_fill_2 FILLER_37_155 ();
 sg13g2_fill_1 FILLER_37_183 ();
 sg13g2_decap_8 FILLER_37_188 ();
 sg13g2_decap_4 FILLER_37_195 ();
 sg13g2_fill_1 FILLER_37_238 ();
 sg13g2_fill_2 FILLER_37_285 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_fill_1 FILLER_37_338 ();
 sg13g2_fill_2 FILLER_37_365 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_4 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_36 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_8 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_206 ();
 sg13g2_fill_2 FILLER_38_213 ();
 sg13g2_fill_1 FILLER_38_223 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_4 FILLER_38_236 ();
 sg13g2_fill_2 FILLER_38_240 ();
 sg13g2_decap_8 FILLER_38_251 ();
 sg13g2_decap_8 FILLER_38_258 ();
 sg13g2_fill_2 FILLER_38_265 ();
 sg13g2_fill_1 FILLER_38_278 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_decap_4 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 assign uio_oe[0] = net290;
 assign uio_oe[1] = net291;
 assign uio_oe[2] = net292;
 assign uio_oe[3] = net293;
 assign uio_oe[4] = net294;
 assign uio_oe[5] = net295;
 assign uio_oe[6] = net296;
 assign uio_oe[7] = net297;
 assign uio_out[0] = net298;
 assign uio_out[1] = net299;
 assign uio_out[2] = net300;
 assign uio_out[3] = net301;
 assign uio_out[4] = net302;
 assign uio_out[5] = net303;
 assign uio_out[6] = net304;
 assign uio_out[7] = net305;
endmodule
